magic
tech sky130A
magscale 1 2
timestamp 1542649553
<< checkpaint >>
rect -12658 -11586 596582 715522
<< viali >>
rect 478943 431409 478977 431443
rect 485831 431409 485865 431443
rect 478581 410397 478615 410431
rect 485111 410397 485145 410431
rect 479474 389453 479508 389487
rect 490610 389453 490644 389487
rect 477091 356813 477125 356847
rect 480143 356813 480177 356847
rect 482075 340833 482109 340867
rect 475442 340357 475476 340391
rect 478759 340357 478793 340391
rect 478939 320365 478973 320399
rect 485827 320365 485861 320399
rect 478580 305405 478614 305439
rect 485110 305405 485144 305439
rect 490610 285957 490644 285991
rect 479474 285821 479508 285855
rect 477101 265829 477135 265863
rect 208685 69853 208719 69887
<< metal1 >>
rect 470234 451485 470854 451491
rect 470234 451177 470262 451485
rect 470826 451177 470854 451485
rect 470234 451171 470854 451177
rect 471330 450644 471336 450696
rect 471388 450684 471394 450696
rect 471388 450656 471652 450684
rect 471388 450644 471394 450656
rect 468994 450399 469614 450405
rect 468994 450091 469022 450399
rect 469586 450091 469614 450399
rect 468994 450085 469614 450091
rect 475378 449436 475384 449488
rect 475436 449436 475442 449488
rect 478690 449436 478696 449488
rect 478748 449436 478754 449488
rect 482002 449436 482008 449488
rect 482060 449436 482066 449488
rect 485314 449436 485320 449488
rect 485372 449436 485378 449488
rect 488644 449392 488672 449462
rect 491938 449392 491944 449404
rect 488644 449364 491944 449392
rect 491938 449352 491944 449364
rect 491996 449352 492002 449404
rect 470234 449314 470854 449320
rect 470234 449006 470262 449314
rect 470826 449006 470854 449314
rect 470234 449000 470854 449006
rect 478690 446224 478696 446276
rect 478748 446264 478754 446276
rect 478748 446236 480254 446264
rect 478748 446224 478754 446236
rect 480226 445924 480254 446236
rect 515398 445924 515404 445936
rect 480226 445896 515404 445924
rect 515398 445884 515404 445896
rect 515456 445884 515462 445936
rect 482002 445816 482008 445868
rect 482060 445856 482066 445868
rect 520918 445856 520924 445868
rect 482060 445828 520924 445856
rect 482060 445816 482066 445828
rect 520918 445816 520924 445828
rect 520976 445816 520982 445868
rect 485314 445748 485320 445800
rect 485372 445788 485378 445800
rect 523678 445788 523684 445800
rect 485372 445760 523684 445788
rect 485372 445748 485378 445760
rect 523678 445748 523684 445760
rect 523736 445748 523742 445800
rect 475378 445680 475384 445732
rect 475436 445720 475442 445732
rect 535454 445720 535460 445732
rect 475436 445692 535460 445720
rect 475436 445680 475442 445692
rect 535454 445680 535460 445692
rect 535512 445680 535518 445732
rect 490558 442960 490564 443012
rect 490616 443000 490622 443012
rect 535454 443000 535460 443012
rect 490616 442972 535460 443000
rect 490616 442960 490622 442972
rect 535454 442960 535460 442972
rect 535512 442960 535518 443012
rect 493318 441600 493324 441652
rect 493376 441640 493382 441652
rect 535454 441640 535460 441652
rect 493376 441612 535460 441640
rect 493376 441600 493382 441612
rect 535454 441600 535460 441612
rect 535512 441600 535518 441652
rect 494698 440240 494704 440292
rect 494756 440280 494762 440292
rect 535454 440280 535460 440292
rect 494756 440252 535460 440280
rect 494756 440240 494762 440252
rect 535454 440240 535460 440252
rect 535512 440240 535518 440292
rect 496078 438880 496084 438932
rect 496136 438920 496142 438932
rect 535454 438920 535460 438932
rect 496136 438892 535460 438920
rect 496136 438880 496142 438892
rect 535454 438880 535460 438892
rect 535512 438880 535518 438932
rect 497458 437452 497464 437504
rect 497516 437492 497522 437504
rect 535454 437492 535460 437504
rect 497516 437464 535460 437492
rect 497516 437452 497522 437464
rect 535454 437452 535460 437464
rect 535512 437452 535518 437504
rect 498838 436092 498844 436144
rect 498896 436132 498902 436144
rect 535454 436132 535460 436144
rect 498896 436104 535460 436132
rect 498896 436092 498902 436104
rect 535454 436092 535460 436104
rect 535512 436092 535518 436144
rect 500218 434732 500224 434784
rect 500276 434772 500282 434784
rect 535454 434772 535460 434784
rect 500276 434744 535460 434772
rect 500276 434732 500282 434744
rect 535454 434732 535460 434744
rect 535512 434732 535518 434784
rect 501598 433304 501604 433356
rect 501656 433344 501662 433356
rect 535454 433344 535460 433356
rect 501656 433316 535460 433344
rect 501656 433304 501662 433316
rect 535454 433304 535460 433316
rect 535512 433304 535518 433356
rect 470234 433086 470854 433092
rect 470234 432778 470262 433086
rect 470826 432778 470854 433086
rect 470234 432772 470854 432778
rect 471612 432290 471664 432296
rect 471612 432232 471664 432238
rect 468994 431999 469614 432005
rect 468994 431691 469022 431999
rect 469586 431691 469614 431999
rect 502978 431944 502984 431996
rect 503036 431984 503042 431996
rect 535454 431984 535460 431996
rect 503036 431956 535460 431984
rect 503036 431944 503042 431956
rect 535454 431944 535460 431956
rect 535512 431944 535518 431996
rect 468994 431685 469614 431691
rect 478966 431449 478972 431452
rect 478931 431443 478972 431449
rect 478931 431409 478943 431443
rect 478931 431403 478972 431409
rect 478966 431400 478972 431403
rect 479024 431400 479030 431452
rect 485774 431400 485780 431452
rect 485832 431449 485838 431452
rect 485832 431443 485877 431449
rect 485865 431409 485877 431443
rect 485832 431403 485877 431409
rect 485832 431400 485838 431403
rect 475470 431035 475476 431087
rect 475528 431035 475534 431087
rect 482370 431035 482376 431087
rect 482428 431035 482434 431087
rect 489302 431047 489592 431075
rect 489564 431032 489592 431047
rect 492030 431032 492036 431044
rect 489564 431004 492036 431032
rect 492030 430992 492036 431004
rect 492088 430992 492094 431044
rect 470234 430914 470854 430920
rect 470234 430606 470262 430914
rect 470826 430606 470854 430914
rect 470234 430600 470854 430606
rect 475470 429088 475476 429140
rect 475528 429128 475534 429140
rect 490558 429128 490564 429140
rect 475528 429100 490564 429128
rect 475528 429088 475534 429100
rect 490558 429088 490564 429100
rect 490616 429088 490622 429140
rect 482370 427796 482376 427848
rect 482428 427836 482434 427848
rect 522298 427836 522304 427848
rect 482428 427808 522304 427836
rect 482428 427796 482434 427808
rect 522298 427796 522304 427808
rect 522356 427796 522362 427848
rect 470234 412086 470854 412092
rect 470234 411778 470262 412086
rect 470826 411778 470854 412086
rect 470234 411772 470854 411778
rect 471238 411204 471244 411256
rect 471296 411244 471302 411256
rect 471624 411244 471652 411263
rect 471296 411216 471652 411244
rect 473722 411232 473728 411284
rect 473780 411232 473786 411284
rect 471296 411204 471302 411216
rect 468994 411000 469614 411006
rect 468994 410692 469022 411000
rect 469586 410692 469614 411000
rect 468994 410686 469614 410692
rect 477788 410440 478478 410457
rect 477788 410428 478420 410440
rect 478414 410388 478420 410428
rect 478472 410388 478478 410440
rect 478598 410437 478604 410440
rect 478569 410431 478604 410437
rect 478569 410397 478581 410431
rect 478569 410391 478604 410397
rect 478598 410388 478604 410391
rect 478656 410388 478662 410440
rect 485130 410437 485136 410440
rect 485099 410431 485136 410437
rect 485099 410397 485111 410431
rect 485099 410391 485136 410397
rect 485130 410388 485136 410391
rect 485188 410388 485194 410440
rect 475286 410036 475292 410088
rect 475344 410036 475350 410088
rect 481818 410036 481824 410088
rect 481876 410036 481882 410088
rect 488382 410048 488672 410076
rect 488644 410020 488672 410048
rect 490742 410020 490748 410032
rect 488644 409992 490748 410020
rect 490742 409980 490748 409992
rect 490800 409980 490806 410032
rect 470234 409914 470854 409920
rect 470234 409606 470262 409914
rect 470826 409606 470854 409914
rect 515398 409776 515404 409828
rect 515456 409816 515462 409828
rect 535454 409816 535460 409828
rect 515456 409788 535460 409816
rect 515456 409776 515462 409788
rect 535454 409776 535460 409788
rect 535512 409776 535518 409828
rect 470234 409600 470854 409606
rect 475286 408416 475292 408468
rect 475344 408456 475350 408468
rect 493318 408456 493324 408468
rect 475344 408428 493324 408456
rect 475344 408416 475350 408428
rect 493318 408416 493324 408428
rect 493376 408416 493382 408468
rect 478598 407056 478604 407108
rect 478656 407096 478662 407108
rect 535454 407096 535460 407108
rect 478656 407068 535460 407096
rect 478656 407056 478662 407068
rect 535454 407056 535460 407068
rect 535512 407056 535518 407108
rect 515398 404336 515404 404388
rect 515456 404376 515462 404388
rect 535454 404376 535460 404388
rect 515456 404348 535460 404376
rect 515456 404336 515462 404348
rect 535454 404336 535460 404348
rect 535512 404336 535518 404388
rect 516778 402976 516784 403028
rect 516836 403016 516842 403028
rect 535454 403016 535460 403028
rect 516836 402988 535460 403016
rect 516836 402976 516842 402988
rect 535454 402976 535460 402988
rect 535512 402976 535518 403028
rect 518158 398828 518164 398880
rect 518216 398868 518222 398880
rect 535454 398868 535460 398880
rect 518216 398840 535460 398868
rect 518216 398828 518222 398840
rect 535454 398828 535460 398840
rect 535512 398828 535518 398880
rect 519538 396040 519544 396092
rect 519596 396080 519602 396092
rect 535454 396080 535460 396092
rect 519596 396052 535460 396080
rect 519596 396040 519602 396052
rect 535454 396040 535460 396052
rect 535512 396040 535518 396092
rect 470234 391087 470854 391093
rect 470234 390779 470262 391087
rect 470826 390779 470854 391087
rect 470234 390773 470854 390779
rect 471238 390260 471244 390312
rect 471296 390300 471302 390312
rect 471296 390272 471652 390300
rect 471296 390260 471302 390272
rect 471624 390096 471652 390272
rect 471698 390096 471704 390108
rect 471624 390068 471704 390096
rect 471698 390056 471704 390068
rect 471756 390056 471762 390108
rect 468994 390004 469614 390010
rect 468994 389696 469022 390004
rect 469586 389696 469614 390004
rect 468994 389690 469614 389696
rect 479426 389444 479432 389496
rect 479484 389493 479490 389496
rect 479484 389487 479520 389493
rect 479508 389453 479520 389487
rect 479484 389447 479520 389453
rect 490598 389487 490656 389493
rect 490598 389453 490610 389487
rect 490644 389484 490656 389487
rect 493318 389484 493324 389496
rect 490644 389456 493324 389484
rect 490644 389453 490656 389456
rect 490598 389447 490656 389453
rect 479484 389444 479490 389447
rect 493318 389444 493324 389456
rect 493376 389444 493382 389496
rect 475746 389036 475752 389088
rect 475804 389036 475810 389088
rect 483198 389036 483204 389088
rect 483256 389036 483262 389088
rect 486878 389036 486884 389088
rect 486936 389036 486942 389088
rect 470234 388914 470854 388920
rect 470234 388606 470262 388914
rect 470826 388606 470854 388914
rect 470234 388600 470854 388606
rect 475746 387744 475752 387796
rect 475804 387744 475810 387796
rect 479426 387744 479432 387796
rect 479484 387784 479490 387796
rect 515398 387784 515404 387796
rect 479484 387756 515404 387784
rect 479484 387744 479490 387756
rect 515398 387744 515404 387756
rect 515456 387744 515462 387796
rect 475764 387716 475792 387744
rect 494698 387716 494704 387728
rect 475764 387688 494704 387716
rect 494698 387676 494704 387688
rect 494756 387676 494762 387728
rect 483198 386384 483204 386436
rect 483256 386424 483262 386436
rect 484302 386424 484308 386436
rect 483256 386396 484308 386424
rect 483256 386384 483262 386396
rect 484302 386384 484308 386396
rect 484360 386384 484366 386436
rect 520918 373940 520924 373992
rect 520976 373980 520982 373992
rect 535454 373980 535460 373992
rect 520976 373952 535460 373980
rect 520976 373940 520982 373952
rect 535454 373940 535460 373952
rect 535512 373940 535518 373992
rect 522298 372512 522304 372564
rect 522356 372552 522362 372564
rect 535454 372552 535460 372564
rect 522356 372524 535460 372552
rect 522356 372512 522362 372524
rect 535454 372512 535460 372524
rect 535512 372512 535518 372564
rect 484302 369792 484308 369844
rect 484360 369832 484366 369844
rect 535454 369832 535460 369844
rect 484360 369804 535460 369832
rect 484360 369792 484366 369804
rect 535454 369792 535460 369804
rect 535512 369792 535518 369844
rect 520918 367072 520924 367124
rect 520976 367112 520982 367124
rect 535454 367112 535460 367124
rect 520976 367084 535460 367112
rect 520976 367072 520982 367084
rect 535454 367072 535460 367084
rect 535512 367072 535518 367124
rect 515398 365712 515404 365764
rect 515456 365752 515462 365764
rect 535454 365752 535460 365764
rect 515456 365724 535460 365752
rect 515456 365712 515462 365724
rect 535454 365712 535460 365724
rect 535512 365712 535518 365764
rect 522298 361564 522304 361616
rect 522356 361604 522362 361616
rect 535454 361604 535460 361616
rect 522356 361576 535460 361604
rect 522356 361564 522362 361576
rect 535454 361564 535460 361576
rect 535512 361564 535518 361616
rect 470234 358487 470854 358493
rect 470234 358179 470262 358487
rect 470826 358179 470854 358487
rect 470234 358173 470854 358179
rect 471698 357552 471704 357604
rect 471756 357592 471762 357604
rect 473648 357592 473676 357664
rect 475102 357620 475108 357672
rect 475160 357620 475166 357672
rect 478874 357631 478880 357683
rect 478932 357631 478938 357683
rect 481818 357631 481824 357683
rect 481876 357631 481882 357683
rect 484946 357631 484952 357683
rect 485004 357631 485010 357683
rect 471756 357564 473676 357592
rect 471756 357552 471762 357564
rect 468994 357401 469614 357407
rect 468994 357093 469022 357401
rect 469586 357093 469614 357401
rect 468994 357087 469614 357093
rect 477034 356804 477040 356856
rect 477092 356853 477098 356856
rect 480162 356853 480168 356856
rect 477092 356847 477137 356853
rect 477125 356813 477137 356847
rect 477092 356807 477137 356813
rect 480131 356847 480168 356853
rect 480131 356813 480143 356847
rect 480131 356807 480168 356813
rect 477092 356804 477098 356807
rect 480162 356804 480168 356807
rect 480220 356804 480226 356856
rect 483198 356435 483204 356487
rect 483256 356435 483262 356487
rect 486234 356435 486240 356487
rect 486292 356435 486298 356487
rect 489288 356436 489316 356461
rect 492122 356436 492128 356448
rect 489288 356408 492128 356436
rect 492122 356396 492128 356408
rect 492180 356396 492186 356448
rect 470234 356314 470854 356320
rect 470234 356006 470262 356314
rect 470826 356006 470854 356314
rect 470234 356000 470854 356006
rect 483198 354628 483204 354680
rect 483256 354668 483262 354680
rect 520918 354668 520924 354680
rect 483256 354640 520924 354668
rect 483256 354628 483262 354640
rect 520918 354628 520924 354640
rect 520976 354628 520982 354680
rect 480162 354560 480168 354612
rect 480220 354600 480226 354612
rect 516778 354600 516784 354612
rect 480220 354572 516784 354600
rect 480220 354560 480226 354572
rect 516778 354560 516784 354572
rect 516836 354560 516842 354612
rect 477126 354492 477132 354544
rect 477184 354532 477190 354544
rect 496078 354532 496084 354544
rect 477184 354504 496084 354532
rect 477184 354492 477190 354504
rect 496078 354492 496084 354504
rect 496136 354492 496142 354544
rect 486234 353608 486240 353660
rect 486292 353648 486298 353660
rect 486292 353620 489914 353648
rect 486292 353608 486298 353620
rect 489886 353308 489914 353620
rect 525058 353308 525064 353320
rect 489886 353280 525064 353308
rect 525058 353268 525064 353280
rect 525116 353268 525122 353320
rect 470234 342486 470854 342492
rect 470234 342178 470262 342486
rect 470826 342178 470854 342486
rect 470234 342172 470854 342178
rect 471698 341776 471704 341828
rect 471756 341776 471762 341828
rect 471238 341708 471244 341760
rect 471296 341748 471302 341760
rect 471716 341748 471744 341776
rect 471296 341720 471744 341748
rect 471296 341708 471302 341720
rect 471716 341663 471744 341720
rect 468994 341399 469614 341405
rect 468994 341091 469022 341399
rect 469586 341091 469614 341399
rect 468994 341085 469614 341091
rect 482094 340873 482100 340876
rect 482063 340867 482100 340873
rect 474642 340803 474648 340855
rect 474700 340803 474706 340855
rect 482063 340833 482075 340867
rect 482063 340827 482100 340833
rect 482094 340824 482100 340827
rect 482152 340824 482158 340876
rect 485590 340478 485596 340490
rect 485438 340450 485596 340478
rect 485590 340438 485596 340450
rect 485648 340438 485654 340490
rect 475470 340397 475476 340400
rect 475430 340391 475476 340397
rect 475430 340357 475442 340391
rect 475430 340351 475476 340357
rect 475470 340348 475476 340351
rect 475528 340348 475534 340400
rect 478782 340397 478788 340400
rect 478747 340391 478788 340397
rect 478747 340357 478759 340391
rect 478747 340351 478788 340357
rect 478782 340348 478788 340351
rect 478840 340348 478846 340400
rect 488736 340388 488764 340464
rect 492214 340388 492220 340400
rect 488736 340360 492220 340388
rect 492214 340348 492220 340360
rect 492272 340348 492278 340400
rect 470234 340314 470854 340320
rect 470234 340006 470262 340314
rect 470826 340006 470854 340314
rect 470234 340000 470854 340006
rect 475470 339396 475476 339448
rect 475528 339396 475534 339448
rect 478782 339396 478788 339448
rect 478840 339436 478846 339448
rect 536374 339436 536380 339448
rect 478840 339408 536380 339436
rect 478840 339396 478846 339408
rect 536374 339396 536380 339408
rect 536432 339396 536438 339448
rect 475488 339300 475516 339396
rect 482094 339328 482100 339380
rect 482152 339368 482158 339380
rect 515398 339368 515404 339380
rect 482152 339340 515404 339368
rect 482152 339328 482158 339340
rect 515398 339328 515404 339340
rect 515456 339328 515462 339380
rect 497458 339300 497464 339312
rect 475488 339272 497464 339300
rect 497458 339260 497464 339272
rect 497516 339260 497522 339312
rect 523678 338036 523684 338088
rect 523736 338076 523742 338088
rect 535454 338076 535460 338088
rect 523736 338048 535460 338076
rect 523736 338036 523742 338048
rect 535454 338036 535460 338048
rect 535512 338036 535518 338088
rect 525058 332528 525064 332580
rect 525116 332568 525122 332580
rect 535454 332568 535460 332580
rect 525116 332540 535460 332568
rect 525116 332528 525122 332540
rect 535454 332528 535460 332540
rect 535512 332528 535518 332580
rect 485682 331168 485688 331220
rect 485740 331208 485746 331220
rect 535454 331208 535460 331220
rect 485740 331180 535460 331208
rect 485740 331168 485746 331180
rect 535454 331168 535460 331180
rect 535512 331168 535518 331220
rect 523678 325660 523684 325712
rect 523736 325700 523742 325712
rect 535454 325700 535460 325712
rect 523736 325672 535460 325700
rect 523736 325660 523742 325672
rect 535454 325660 535460 325672
rect 535512 325660 535518 325712
rect 470234 322486 470854 322492
rect 470234 322178 470262 322486
rect 470826 322178 470854 322486
rect 470234 322172 470854 322178
rect 471238 321580 471244 321632
rect 471296 321620 471302 321632
rect 471624 321620 471652 321663
rect 471296 321592 471652 321620
rect 471296 321580 471302 321592
rect 468994 321399 469614 321405
rect 468994 321091 469022 321399
rect 469586 321091 469614 321399
rect 468994 321085 469614 321091
rect 475470 320435 475476 320487
rect 475528 320435 475534 320487
rect 482370 320424 482376 320476
rect 482428 320424 482434 320476
rect 478927 320399 478985 320405
rect 478927 320365 478939 320399
rect 478973 320396 478985 320399
rect 479058 320396 479064 320408
rect 478973 320368 479064 320396
rect 478973 320365 478985 320368
rect 478927 320359 478985 320365
rect 479058 320356 479064 320368
rect 479116 320356 479122 320408
rect 485815 320399 485873 320405
rect 485815 320365 485827 320399
rect 485861 320396 485873 320399
rect 485958 320396 485964 320408
rect 485861 320368 485964 320396
rect 485861 320365 485873 320368
rect 485815 320359 485873 320365
rect 485958 320356 485964 320368
rect 486016 320356 486022 320408
rect 489288 320396 489316 320461
rect 492306 320396 492312 320408
rect 489288 320368 492312 320396
rect 492306 320356 492312 320368
rect 492364 320356 492370 320408
rect 470234 320314 470854 320320
rect 470234 320006 470262 320314
rect 470826 320006 470854 320314
rect 470234 320000 470854 320006
rect 475470 318724 475476 318776
rect 475528 318724 475534 318776
rect 479058 318724 479064 318776
rect 479116 318764 479122 318776
rect 536282 318764 536288 318776
rect 479116 318736 536288 318764
rect 479116 318724 479122 318736
rect 536282 318724 536288 318736
rect 536340 318724 536346 318776
rect 475488 318560 475516 318724
rect 482370 318656 482376 318708
rect 482428 318696 482434 318708
rect 536558 318696 536564 318708
rect 482428 318668 536564 318696
rect 482428 318656 482434 318668
rect 536558 318656 536564 318668
rect 536616 318656 536622 318708
rect 485958 318588 485964 318640
rect 486016 318628 486022 318640
rect 536006 318628 536012 318640
rect 486016 318600 536012 318628
rect 486016 318588 486022 318600
rect 536006 318588 536012 318600
rect 536064 318588 536070 318640
rect 498838 318560 498844 318572
rect 475488 318532 498844 318560
rect 498838 318520 498844 318532
rect 498896 318520 498902 318572
rect 470234 307086 470854 307092
rect 470234 306778 470262 307086
rect 470826 306778 470854 307086
rect 470234 306772 470854 306778
rect 471238 306280 471244 306332
rect 471296 306320 471302 306332
rect 471296 306292 471652 306320
rect 471296 306280 471302 306292
rect 471624 306264 471652 306292
rect 473722 306232 473728 306284
rect 473780 306232 473786 306284
rect 468994 306001 469614 306007
rect 468994 305693 469022 306001
rect 469586 305693 469614 306001
rect 468994 305687 469614 305693
rect 478598 305445 478604 305448
rect 478568 305439 478604 305445
rect 478568 305405 478580 305439
rect 478568 305399 478604 305405
rect 478598 305396 478604 305399
rect 478656 305396 478662 305448
rect 485130 305445 485136 305448
rect 485098 305439 485136 305445
rect 485098 305405 485110 305439
rect 485098 305399 485136 305405
rect 485130 305396 485136 305399
rect 485188 305396 485194 305448
rect 475286 305036 475292 305088
rect 475344 305036 475350 305088
rect 481818 305036 481824 305088
rect 481876 305036 481882 305088
rect 488382 305048 488672 305076
rect 488644 305028 488672 305048
rect 490558 305028 490564 305040
rect 488644 305000 490564 305028
rect 490558 304988 490564 305000
rect 490616 304988 490622 305040
rect 470234 304914 470854 304920
rect 470234 304606 470262 304914
rect 470826 304606 470854 304914
rect 470234 304600 470854 304606
rect 485056 303640 485268 303668
rect 475286 303560 475292 303612
rect 475344 303560 475350 303612
rect 478598 303560 478604 303612
rect 478656 303600 478662 303612
rect 478656 303572 480254 303600
rect 478656 303560 478662 303572
rect 475304 303396 475332 303560
rect 480226 303464 480254 303572
rect 481818 303560 481824 303612
rect 481876 303600 481882 303612
rect 485056 303600 485084 303640
rect 481876 303572 485084 303600
rect 481876 303560 481882 303572
rect 485130 303560 485136 303612
rect 485188 303560 485194 303612
rect 485240 303600 485268 303640
rect 536466 303600 536472 303612
rect 485240 303572 536472 303600
rect 536466 303560 536472 303572
rect 536524 303560 536530 303612
rect 485148 303532 485176 303560
rect 536650 303532 536656 303544
rect 485148 303504 536656 303532
rect 536650 303492 536656 303504
rect 536708 303492 536714 303544
rect 518158 303464 518164 303476
rect 480226 303436 518164 303464
rect 518158 303424 518164 303436
rect 518216 303424 518222 303476
rect 500218 303396 500224 303408
rect 475304 303368 500224 303396
rect 500218 303356 500224 303368
rect 500276 303356 500282 303408
rect 491938 300772 491944 300824
rect 491996 300812 492002 300824
rect 535454 300812 535460 300824
rect 491996 300784 535460 300812
rect 491996 300772 492002 300784
rect 535454 300772 535460 300784
rect 535512 300772 535518 300824
rect 492030 299412 492036 299464
rect 492088 299452 492094 299464
rect 535454 299452 535460 299464
rect 492088 299424 535460 299452
rect 492088 299412 492094 299424
rect 535454 299412 535460 299424
rect 535512 299412 535518 299464
rect 490742 298052 490748 298104
rect 490800 298092 490806 298104
rect 535454 298092 535460 298104
rect 490800 298064 535460 298092
rect 490800 298052 490806 298064
rect 535454 298052 535460 298064
rect 535512 298052 535518 298104
rect 492122 296624 492128 296676
rect 492180 296664 492186 296676
rect 535546 296664 535552 296676
rect 492180 296636 535552 296664
rect 492180 296624 492186 296636
rect 535546 296624 535552 296636
rect 535604 296624 535610 296676
rect 493318 296556 493324 296608
rect 493376 296596 493382 296608
rect 535454 296596 535460 296608
rect 493376 296568 535460 296596
rect 493376 296556 493382 296568
rect 535454 296556 535460 296568
rect 535512 296556 535518 296608
rect 492214 295264 492220 295316
rect 492272 295304 492278 295316
rect 535454 295304 535460 295316
rect 492272 295276 535460 295304
rect 492272 295264 492278 295276
rect 535454 295264 535460 295276
rect 535512 295264 535518 295316
rect 492306 293904 492312 293956
rect 492364 293944 492370 293956
rect 535546 293944 535552 293956
rect 492364 293916 535552 293944
rect 492364 293904 492370 293916
rect 535546 293904 535552 293916
rect 535604 293904 535610 293956
rect 490558 292476 490564 292528
rect 490616 292516 490622 292528
rect 535454 292516 535460 292528
rect 490616 292488 535460 292516
rect 490616 292476 490622 292488
rect 535454 292476 535460 292488
rect 535512 292476 535518 292528
rect 492950 289824 492956 289876
rect 493008 289864 493014 289876
rect 535454 289864 535460 289876
rect 493008 289836 535460 289864
rect 493008 289824 493014 289836
rect 535454 289824 535460 289836
rect 535512 289824 535518 289876
rect 491938 288396 491944 288448
rect 491996 288436 492002 288448
rect 535454 288436 535460 288448
rect 491996 288408 535460 288436
rect 491996 288396 492002 288408
rect 535454 288396 535460 288408
rect 535512 288396 535518 288448
rect 470234 287487 470854 287493
rect 470234 287179 470262 287487
rect 470826 287179 470854 287487
rect 470234 287173 470854 287179
rect 488632 286680 488684 286686
rect 471238 286628 471244 286680
rect 471296 286668 471302 286680
rect 471296 286640 471652 286668
rect 471296 286628 471302 286640
rect 471624 286532 471652 286640
rect 488632 286622 488684 286628
rect 471698 286532 471704 286544
rect 471624 286504 471704 286532
rect 471698 286492 471704 286504
rect 471756 286492 471762 286544
rect 468994 286402 469614 286408
rect 468994 286094 469022 286402
rect 469586 286094 469614 286402
rect 468994 286088 469614 286094
rect 490598 285991 490656 285997
rect 490598 285957 490610 285991
rect 490644 285988 490656 285991
rect 490644 285960 490880 285988
rect 490644 285957 490656 285960
rect 490598 285951 490656 285957
rect 479426 285812 479432 285864
rect 479484 285861 479490 285864
rect 479484 285855 479520 285861
rect 479508 285821 479520 285855
rect 479484 285815 479520 285821
rect 479484 285812 479490 285815
rect 490852 285648 490880 285960
rect 492950 285648 492956 285660
rect 490852 285620 492956 285648
rect 492950 285608 492956 285620
rect 493008 285608 493014 285660
rect 475746 285436 475752 285488
rect 475804 285436 475810 285488
rect 483198 285436 483204 285488
rect 483256 285436 483262 285488
rect 486878 285436 486884 285488
rect 486936 285436 486942 285488
rect 470234 285314 470854 285320
rect 470234 285006 470262 285314
rect 470826 285006 470854 285314
rect 470234 285000 470854 285006
rect 475746 284248 475752 284300
rect 475804 284248 475810 284300
rect 479426 284248 479432 284300
rect 479484 284288 479490 284300
rect 536098 284288 536104 284300
rect 479484 284260 536104 284288
rect 479484 284248 479490 284260
rect 536098 284248 536104 284260
rect 536156 284248 536162 284300
rect 475764 284084 475792 284248
rect 483198 284180 483204 284232
rect 483256 284180 483262 284232
rect 522298 284220 522304 284232
rect 485746 284192 522304 284220
rect 483216 284152 483244 284180
rect 485746 284152 485774 284192
rect 522298 284180 522304 284192
rect 522356 284180 522362 284232
rect 483216 284124 485774 284152
rect 486878 284112 486884 284164
rect 486936 284152 486942 284164
rect 523678 284152 523684 284164
rect 486936 284124 523684 284152
rect 486936 284112 486942 284124
rect 523678 284112 523684 284124
rect 523736 284112 523742 284164
rect 501598 284084 501604 284096
rect 475764 284056 501604 284084
rect 501598 284044 501604 284056
rect 501656 284044 501662 284096
rect 471698 270444 471704 270496
rect 471756 270484 471762 270496
rect 473722 270484 473728 270496
rect 471756 270456 473728 270484
rect 471756 270444 471762 270456
rect 473722 270444 473728 270456
rect 473780 270444 473786 270496
rect 470234 267487 470854 267493
rect 470234 267179 470262 267487
rect 470826 267179 470854 267487
rect 470234 267173 470854 267179
rect 473648 266540 473676 266664
rect 473722 266540 473728 266552
rect 473648 266512 473728 266540
rect 473722 266500 473728 266512
rect 473780 266500 473786 266552
rect 468994 266401 469614 266407
rect 468994 266093 469022 266401
rect 469586 266093 469614 266401
rect 468994 266087 469614 266093
rect 491938 265996 491944 266008
rect 489288 265968 491944 265996
rect 477126 265869 477132 265872
rect 477089 265863 477132 265869
rect 477089 265829 477101 265863
rect 477089 265823 477132 265829
rect 477126 265820 477132 265823
rect 477184 265820 477190 265872
rect 489288 265731 489316 265968
rect 491938 265956 491944 265968
rect 491996 265956 492002 266008
rect 480162 265435 480168 265487
rect 480220 265435 480226 265487
rect 483198 265435 483204 265487
rect 483256 265435 483262 265487
rect 486234 265435 486240 265487
rect 486292 265435 486298 265487
rect 470234 265314 470854 265320
rect 470234 265006 470262 265314
rect 470826 265006 470854 265314
rect 470234 265000 470854 265006
rect 494716 263588 494928 263616
rect 477126 263508 477132 263560
rect 477184 263508 477190 263560
rect 480162 263508 480168 263560
rect 480220 263548 480226 263560
rect 480220 263508 480254 263548
rect 483198 263508 483204 263560
rect 483256 263508 483262 263560
rect 486234 263508 486240 263560
rect 486292 263548 486298 263560
rect 494716 263548 494744 263588
rect 486292 263520 494744 263548
rect 494900 263548 494928 263588
rect 494900 263520 495020 263548
rect 486292 263508 486298 263520
rect 477144 263344 477172 263508
rect 480226 263412 480254 263508
rect 483216 263480 483244 263508
rect 494790 263480 494796 263492
rect 483216 263452 494796 263480
rect 494790 263440 494796 263452
rect 494848 263440 494854 263492
rect 494992 263480 495020 263520
rect 495066 263508 495072 263560
rect 495124 263548 495130 263560
rect 536190 263548 536196 263560
rect 495124 263520 536196 263548
rect 495124 263508 495130 263520
rect 536190 263508 536196 263520
rect 536248 263508 536254 263560
rect 536374 263480 536380 263492
rect 494992 263452 536380 263480
rect 536374 263440 536380 263452
rect 536432 263440 536438 263492
rect 519538 263412 519544 263424
rect 480226 263384 519544 263412
rect 519538 263372 519544 263384
rect 519596 263372 519602 263424
rect 502978 263344 502984 263356
rect 477144 263316 502984 263344
rect 502978 263304 502984 263316
rect 503036 263304 503042 263356
rect 473722 206932 473728 206984
rect 473780 206972 473786 206984
rect 580166 206972 580172 206984
rect 473780 206944 580172 206972
rect 473780 206932 473786 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 208673 69887 208731 69893
rect 208673 69853 208685 69887
rect 208719 69884 208731 69887
rect 536098 69884 536104 69896
rect 208719 69856 536104 69884
rect 208719 69853 208731 69856
rect 208673 69847 208731 69853
rect 536098 69844 536104 69856
rect 536156 69844 536162 69896
<< via1 >>
rect 470262 451177 470826 451485
rect 471336 450644 471388 450696
rect 469022 450091 469586 450399
rect 475384 449436 475436 449488
rect 478696 449436 478748 449488
rect 482008 449436 482060 449488
rect 485320 449436 485372 449488
rect 491944 449352 491996 449404
rect 470262 449006 470826 449314
rect 478696 446224 478748 446276
rect 515404 445884 515456 445936
rect 482008 445816 482060 445868
rect 520924 445816 520976 445868
rect 485320 445748 485372 445800
rect 523684 445748 523736 445800
rect 475384 445680 475436 445732
rect 535460 445680 535512 445732
rect 490564 442960 490616 443012
rect 535460 442960 535512 443012
rect 493324 441600 493376 441652
rect 535460 441600 535512 441652
rect 494704 440240 494756 440292
rect 535460 440240 535512 440292
rect 496084 438880 496136 438932
rect 535460 438880 535512 438932
rect 497464 437452 497516 437504
rect 535460 437452 535512 437504
rect 498844 436092 498896 436144
rect 535460 436092 535512 436144
rect 500224 434732 500276 434784
rect 535460 434732 535512 434784
rect 501604 433304 501656 433356
rect 535460 433304 535512 433356
rect 470262 432778 470826 433086
rect 471612 432238 471664 432290
rect 469022 431691 469586 431999
rect 502984 431944 503036 431996
rect 535460 431944 535512 431996
rect 478972 431443 479024 431452
rect 478972 431409 478977 431443
rect 478977 431409 479024 431443
rect 478972 431400 479024 431409
rect 485780 431443 485832 431452
rect 485780 431409 485831 431443
rect 485831 431409 485832 431443
rect 485780 431400 485832 431409
rect 475476 431035 475528 431087
rect 482376 431035 482428 431087
rect 492036 430992 492088 431044
rect 470262 430606 470826 430914
rect 475476 429088 475528 429140
rect 490564 429088 490616 429140
rect 482376 427796 482428 427848
rect 522304 427796 522356 427848
rect 470262 411778 470826 412086
rect 471244 411204 471296 411256
rect 473728 411232 473780 411284
rect 469022 410692 469586 411000
rect 478420 410388 478472 410440
rect 478604 410431 478656 410440
rect 478604 410397 478615 410431
rect 478615 410397 478656 410431
rect 478604 410388 478656 410397
rect 485136 410431 485188 410440
rect 485136 410397 485145 410431
rect 485145 410397 485188 410431
rect 485136 410388 485188 410397
rect 475292 410036 475344 410088
rect 481824 410036 481876 410088
rect 490748 409980 490800 410032
rect 470262 409606 470826 409914
rect 515404 409776 515456 409828
rect 535460 409776 535512 409828
rect 475292 408416 475344 408468
rect 493324 408416 493376 408468
rect 478604 407056 478656 407108
rect 535460 407056 535512 407108
rect 515404 404336 515456 404388
rect 535460 404336 535512 404388
rect 516784 402976 516836 403028
rect 535460 402976 535512 403028
rect 518164 398828 518216 398880
rect 535460 398828 535512 398880
rect 519544 396040 519596 396092
rect 535460 396040 535512 396092
rect 470262 390779 470826 391087
rect 471244 390260 471296 390312
rect 471704 390056 471756 390108
rect 469022 389696 469586 390004
rect 479432 389487 479484 389496
rect 479432 389453 479474 389487
rect 479474 389453 479484 389487
rect 479432 389444 479484 389453
rect 493324 389444 493376 389496
rect 475752 389036 475804 389088
rect 483204 389036 483256 389088
rect 486884 389036 486936 389088
rect 470262 388606 470826 388914
rect 475752 387744 475804 387796
rect 479432 387744 479484 387796
rect 515404 387744 515456 387796
rect 494704 387676 494756 387728
rect 483204 386384 483256 386436
rect 484308 386384 484360 386436
rect 520924 373940 520976 373992
rect 535460 373940 535512 373992
rect 522304 372512 522356 372564
rect 535460 372512 535512 372564
rect 484308 369792 484360 369844
rect 535460 369792 535512 369844
rect 520924 367072 520976 367124
rect 535460 367072 535512 367124
rect 515404 365712 515456 365764
rect 535460 365712 535512 365764
rect 522304 361564 522356 361616
rect 535460 361564 535512 361616
rect 470262 358179 470826 358487
rect 471704 357552 471756 357604
rect 475108 357620 475160 357672
rect 478880 357631 478932 357683
rect 481824 357631 481876 357683
rect 484952 357631 485004 357683
rect 469022 357093 469586 357401
rect 477040 356847 477092 356856
rect 477040 356813 477091 356847
rect 477091 356813 477092 356847
rect 477040 356804 477092 356813
rect 480168 356847 480220 356856
rect 480168 356813 480177 356847
rect 480177 356813 480220 356847
rect 480168 356804 480220 356813
rect 483204 356435 483256 356487
rect 486240 356435 486292 356487
rect 492128 356396 492180 356448
rect 470262 356006 470826 356314
rect 483204 354628 483256 354680
rect 520924 354628 520976 354680
rect 480168 354560 480220 354612
rect 516784 354560 516836 354612
rect 477132 354492 477184 354544
rect 496084 354492 496136 354544
rect 486240 353608 486292 353660
rect 525064 353268 525116 353320
rect 470262 342178 470826 342486
rect 471704 341776 471756 341828
rect 471244 341708 471296 341760
rect 469022 341091 469586 341399
rect 482100 340867 482152 340876
rect 474648 340803 474700 340855
rect 482100 340833 482109 340867
rect 482109 340833 482152 340867
rect 482100 340824 482152 340833
rect 485596 340438 485648 340490
rect 475476 340348 475528 340400
rect 478788 340391 478840 340400
rect 478788 340357 478793 340391
rect 478793 340357 478840 340391
rect 478788 340348 478840 340357
rect 492220 340348 492272 340400
rect 470262 340006 470826 340314
rect 475476 339396 475528 339448
rect 478788 339396 478840 339448
rect 536380 339396 536432 339448
rect 482100 339328 482152 339380
rect 515404 339328 515456 339380
rect 497464 339260 497516 339312
rect 523684 338036 523736 338088
rect 535460 338036 535512 338088
rect 525064 332528 525116 332580
rect 535460 332528 535512 332580
rect 485688 331168 485740 331220
rect 535460 331168 535512 331220
rect 523684 325660 523736 325712
rect 535460 325660 535512 325712
rect 470262 322178 470826 322486
rect 471244 321580 471296 321632
rect 469022 321091 469586 321399
rect 475476 320435 475528 320487
rect 482376 320424 482428 320476
rect 479064 320356 479116 320408
rect 485964 320356 486016 320408
rect 492312 320356 492364 320408
rect 470262 320006 470826 320314
rect 475476 318724 475528 318776
rect 479064 318724 479116 318776
rect 536288 318724 536340 318776
rect 482376 318656 482428 318708
rect 536564 318656 536616 318708
rect 485964 318588 486016 318640
rect 536012 318588 536064 318640
rect 498844 318520 498896 318572
rect 470262 306778 470826 307086
rect 471244 306280 471296 306332
rect 473728 306232 473780 306284
rect 469022 305693 469586 306001
rect 478604 305439 478656 305448
rect 478604 305405 478614 305439
rect 478614 305405 478656 305439
rect 478604 305396 478656 305405
rect 485136 305439 485188 305448
rect 485136 305405 485144 305439
rect 485144 305405 485188 305439
rect 485136 305396 485188 305405
rect 475292 305036 475344 305088
rect 481824 305036 481876 305088
rect 490564 304988 490616 305040
rect 470262 304606 470826 304914
rect 475292 303560 475344 303612
rect 478604 303560 478656 303612
rect 481824 303560 481876 303612
rect 485136 303560 485188 303612
rect 536472 303560 536524 303612
rect 536656 303492 536708 303544
rect 518164 303424 518216 303476
rect 500224 303356 500276 303408
rect 491944 300772 491996 300824
rect 535460 300772 535512 300824
rect 492036 299412 492088 299464
rect 535460 299412 535512 299464
rect 490748 298052 490800 298104
rect 535460 298052 535512 298104
rect 492128 296624 492180 296676
rect 535552 296624 535604 296676
rect 493324 296556 493376 296608
rect 535460 296556 535512 296608
rect 492220 295264 492272 295316
rect 535460 295264 535512 295316
rect 492312 293904 492364 293956
rect 535552 293904 535604 293956
rect 490564 292476 490616 292528
rect 535460 292476 535512 292528
rect 492956 289824 493008 289876
rect 535460 289824 535512 289876
rect 491944 288396 491996 288448
rect 535460 288396 535512 288448
rect 470262 287179 470826 287487
rect 471244 286628 471296 286680
rect 488632 286628 488684 286680
rect 471704 286492 471756 286544
rect 469022 286094 469586 286402
rect 479432 285855 479484 285864
rect 479432 285821 479474 285855
rect 479474 285821 479484 285855
rect 479432 285812 479484 285821
rect 492956 285608 493008 285660
rect 475752 285436 475804 285488
rect 483204 285436 483256 285488
rect 486884 285436 486936 285488
rect 470262 285006 470826 285314
rect 475752 284248 475804 284300
rect 479432 284248 479484 284300
rect 536104 284248 536156 284300
rect 483204 284180 483256 284232
rect 522304 284180 522356 284232
rect 486884 284112 486936 284164
rect 523684 284112 523736 284164
rect 501604 284044 501656 284096
rect 471704 270444 471756 270496
rect 473728 270444 473780 270496
rect 470262 267179 470826 267487
rect 473728 266500 473780 266552
rect 469022 266093 469586 266401
rect 477132 265863 477184 265872
rect 477132 265829 477135 265863
rect 477135 265829 477184 265863
rect 477132 265820 477184 265829
rect 491944 265956 491996 266008
rect 480168 265435 480220 265487
rect 483204 265435 483256 265487
rect 486240 265435 486292 265487
rect 470262 265006 470826 265314
rect 477132 263508 477184 263560
rect 480168 263508 480220 263560
rect 483204 263508 483256 263560
rect 486240 263508 486292 263560
rect 494796 263440 494848 263492
rect 495072 263508 495124 263560
rect 536196 263508 536248 263560
rect 536380 263440 536432 263492
rect 519544 263372 519596 263424
rect 502984 263304 503036 263356
rect 473728 206932 473780 206984
rect 580172 206932 580224 206984
rect 536104 69844 536156 69896
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 470262 451485 470826 451491
rect 470262 451171 470826 451177
rect 471256 450758 471376 450786
rect 469022 450399 469586 450405
rect 469022 450085 469586 450091
rect 470262 449314 470826 449320
rect 470262 449000 470826 449006
rect 470262 433086 470826 433092
rect 470262 432772 470826 432778
rect 471256 432290 471284 450758
rect 471348 450702 471376 450758
rect 471336 450696 471388 450702
rect 471336 450638 471388 450644
rect 474108 450350 474554 450378
rect 474108 449721 474136 450350
rect 477843 450256 477899 450265
rect 477843 450191 477899 450200
rect 481160 450256 481216 450265
rect 481160 450191 481216 450200
rect 484477 450256 484533 450265
rect 484477 450191 484533 450200
rect 487793 450256 487849 450265
rect 487793 450191 487849 450200
rect 474094 449712 474150 449721
rect 474094 449647 474150 449656
rect 475384 449488 475436 449494
rect 475384 449430 475436 449436
rect 478696 449488 478748 449494
rect 478696 449430 478748 449436
rect 482008 449488 482060 449494
rect 482008 449430 482060 449436
rect 485320 449488 485372 449494
rect 485320 449430 485372 449436
rect 475396 445738 475424 449430
rect 478708 446282 478736 449430
rect 478696 446276 478748 446282
rect 478696 446218 478748 446224
rect 482020 445874 482048 449430
rect 482008 445868 482060 445874
rect 482008 445810 482060 445816
rect 485332 445806 485360 449430
rect 491944 449404 491996 449410
rect 491944 449346 491996 449352
rect 485320 445800 485372 445806
rect 485320 445742 485372 445748
rect 475384 445732 475436 445738
rect 475384 445674 475436 445680
rect 490564 443012 490616 443018
rect 490564 442954 490616 442960
rect 483570 432304 483626 432313
rect 471612 432290 471664 432296
rect 471256 432262 471612 432290
rect 469022 431999 469586 432005
rect 469022 431685 469586 431691
rect 470262 430914 470826 430920
rect 470262 430600 470826 430606
rect 470262 412086 470826 412092
rect 470262 411772 470826 411778
rect 471256 411262 471284 432262
rect 483143 432262 483570 432290
rect 483570 432239 483626 432248
rect 471612 432232 471664 432238
rect 481270 432168 481326 432177
rect 481326 432126 481573 432154
rect 481270 432103 481326 432112
rect 474292 431990 474685 432018
rect 488092 431990 488461 432018
rect 474292 431905 474320 431990
rect 488092 431905 488120 431990
rect 474278 431896 474334 431905
rect 474278 431831 474334 431840
rect 488078 431896 488134 431905
rect 488078 431831 488134 431840
rect 478102 431624 478158 431633
rect 478102 431559 478158 431568
rect 478972 431452 479024 431458
rect 478972 431394 479024 431400
rect 485780 431452 485832 431458
rect 485780 431394 485832 431400
rect 475476 431087 475528 431093
rect 475476 431029 475528 431035
rect 475488 429146 475516 431029
rect 475476 429140 475528 429146
rect 475476 429082 475528 429088
rect 478984 427961 479012 431394
rect 482376 431087 482428 431093
rect 482376 431029 482428 431035
rect 478970 427952 479026 427961
rect 478970 427887 479026 427896
rect 482388 427854 482416 431029
rect 485792 427961 485820 431394
rect 490576 429146 490604 442954
rect 490564 429140 490616 429146
rect 490564 429082 490616 429088
rect 485778 427952 485834 427961
rect 485778 427887 485834 427896
rect 482376 427848 482428 427854
rect 482376 427790 482428 427796
rect 473728 411284 473780 411290
rect 471244 411256 471296 411262
rect 473728 411226 473780 411232
rect 471244 411198 471296 411204
rect 469022 411000 469586 411006
rect 469022 410686 469586 410692
rect 470262 409914 470826 409920
rect 470262 409600 470826 409606
rect 470262 391087 470826 391093
rect 470262 390773 470826 390779
rect 471256 390318 471284 411198
rect 473740 410961 473768 411226
rect 473726 410952 473782 410961
rect 473726 410887 473782 410896
rect 478420 410440 478472 410446
rect 478420 410382 478472 410388
rect 478604 410440 478656 410446
rect 478604 410382 478656 410388
rect 478432 410145 478460 410382
rect 478418 410136 478474 410145
rect 475292 410088 475344 410094
rect 478418 410071 478474 410080
rect 475292 410030 475344 410036
rect 475304 408474 475332 410030
rect 475292 408468 475344 408474
rect 475292 408410 475344 408416
rect 478616 407114 478644 410382
rect 481019 410258 481047 410516
rect 484136 410502 484298 410530
rect 484136 410417 484164 410502
rect 485136 410440 485188 410446
rect 484122 410408 484178 410417
rect 485136 410382 485188 410388
rect 484122 410343 484178 410352
rect 481019 410230 481128 410258
rect 481100 410122 481128 410230
rect 481362 410136 481418 410145
rect 481100 410094 481362 410122
rect 481362 410071 481418 410080
rect 481824 410088 481876 410094
rect 481824 410030 481876 410036
rect 481836 407153 481864 410030
rect 485148 407153 485176 410382
rect 487549 410258 487577 410516
rect 487549 410230 487660 410258
rect 487632 410122 487660 410230
rect 487802 410136 487858 410145
rect 487632 410094 487802 410122
rect 487802 410071 487858 410080
rect 490748 410032 490800 410038
rect 490748 409974 490800 409980
rect 481822 407144 481878 407153
rect 478604 407108 478656 407114
rect 481822 407079 481878 407088
rect 485134 407144 485190 407153
rect 485134 407079 485190 407088
rect 478604 407050 478656 407056
rect 471244 390312 471296 390318
rect 471244 390254 471296 390260
rect 488552 390238 488658 390266
rect 488552 390153 488580 390238
rect 488538 390144 488594 390153
rect 471704 390108 471756 390114
rect 488538 390079 488594 390088
rect 471704 390050 471756 390056
rect 469022 390004 469586 390010
rect 469022 389690 469586 389696
rect 470262 388914 470826 388920
rect 470262 388600 470826 388606
rect 470262 358487 470826 358493
rect 470262 358173 470826 358179
rect 471716 357610 471744 390050
rect 479432 389496 479484 389502
rect 479432 389438 479484 389444
rect 482098 389464 482154 389473
rect 474936 389337 474964 389436
rect 478648 389337 478676 389436
rect 474922 389328 474978 389337
rect 474922 389263 474978 389272
rect 478634 389328 478690 389337
rect 478634 389263 478690 389272
rect 475752 389088 475804 389094
rect 475752 389030 475804 389036
rect 475764 387802 475792 389030
rect 479444 387802 479472 389438
rect 482154 389422 482374 389450
rect 482098 389399 482154 389408
rect 483204 389088 483256 389094
rect 483204 389030 483256 389036
rect 486884 389088 486936 389094
rect 486884 389030 486936 389036
rect 475752 387796 475804 387802
rect 475752 387738 475804 387744
rect 479432 387796 479484 387802
rect 479432 387738 479484 387744
rect 483216 386442 483244 389030
rect 486896 386481 486924 389030
rect 486882 386472 486938 386481
rect 483204 386436 483256 386442
rect 483204 386378 483256 386384
rect 484308 386436 484360 386442
rect 486882 386407 486938 386416
rect 484308 386378 484360 386384
rect 484320 369850 484348 386378
rect 484308 369844 484360 369850
rect 484308 369786 484360 369792
rect 478878 358048 478934 358057
rect 478878 357983 478934 357992
rect 481822 358048 481878 358057
rect 481822 357983 481878 357992
rect 484950 358048 485006 358057
rect 484950 357983 485006 357992
rect 488354 358048 488410 358057
rect 488354 357983 488410 357992
rect 478892 357689 478920 357983
rect 481836 357689 481864 357983
rect 484964 357689 484992 357983
rect 478880 357683 478932 357689
rect 475108 357672 475160 357678
rect 478880 357625 478932 357631
rect 481824 357683 481876 357689
rect 481824 357625 481876 357631
rect 484952 357683 485004 357689
rect 484952 357625 485004 357631
rect 475108 357614 475160 357620
rect 471704 357604 471756 357610
rect 471704 357546 471756 357552
rect 469022 357401 469586 357407
rect 469022 357087 469586 357093
rect 470262 356314 470826 356320
rect 470262 356000 470826 356006
rect 471716 354674 471744 357546
rect 475014 357504 475070 357513
rect 475120 357490 475148 357614
rect 475070 357462 475148 357490
rect 488368 357490 488396 357983
rect 488368 357462 488487 357490
rect 475014 357439 475070 357448
rect 477040 356856 477092 356862
rect 477040 356798 477092 356804
rect 480168 356856 480220 356862
rect 480168 356798 480220 356804
rect 477052 354674 477080 356798
rect 471716 354646 471928 354674
rect 477052 354646 477172 354674
rect 471900 345014 471928 354646
rect 477144 354550 477172 354646
rect 480180 354618 480208 356798
rect 483204 356487 483256 356493
rect 483204 356429 483256 356435
rect 486240 356487 486292 356493
rect 486240 356429 486292 356435
rect 483216 354686 483244 356429
rect 483204 354680 483256 354686
rect 483204 354622 483256 354628
rect 480168 354612 480220 354618
rect 480168 354554 480220 354560
rect 477132 354544 477184 354550
rect 477132 354486 477184 354492
rect 486252 353666 486280 356429
rect 486240 353660 486292 353666
rect 486240 353602 486292 353608
rect 471716 344986 471928 345014
rect 470262 342486 470826 342492
rect 470262 342172 470826 342178
rect 471716 341834 471744 344986
rect 471704 341828 471756 341834
rect 471704 341770 471756 341776
rect 471244 341760 471296 341766
rect 471244 341702 471296 341708
rect 469022 341399 469586 341405
rect 469022 341085 469586 341091
rect 470262 340314 470826 340320
rect 470262 340000 470826 340006
rect 470262 322486 470826 322492
rect 470262 322172 470826 322178
rect 471256 321638 471284 341702
rect 484504 341414 484577 341442
rect 484504 341306 484532 341414
rect 484412 341278 484532 341306
rect 484412 341057 484440 341278
rect 484398 341048 484454 341057
rect 477906 340992 477915 341048
rect 477971 340992 477980 341048
rect 481223 340992 481232 341048
rect 481288 340992 481297 341048
rect 487885 340992 487894 341048
rect 487950 340992 487959 341048
rect 484398 340983 484454 340992
rect 482100 340876 482152 340882
rect 474648 340855 474700 340861
rect 482100 340818 482152 340824
rect 474648 340797 474700 340803
rect 474554 340504 474610 340513
rect 474660 340490 474688 340797
rect 474610 340462 474688 340490
rect 474554 340439 474610 340448
rect 475476 340400 475528 340406
rect 475476 340342 475528 340348
rect 478788 340400 478840 340406
rect 478788 340342 478840 340348
rect 475488 339454 475516 340342
rect 478800 339454 478828 340342
rect 475476 339448 475528 339454
rect 475476 339390 475528 339396
rect 478788 339448 478840 339454
rect 478788 339390 478840 339396
rect 482112 339386 482140 340818
rect 485596 340490 485648 340496
rect 485596 340432 485648 340438
rect 482100 339380 482152 339386
rect 482100 339322 482152 339328
rect 485608 335354 485636 340432
rect 485608 335326 485728 335354
rect 485700 331226 485728 335326
rect 485688 331220 485740 331226
rect 485688 331162 485740 331168
rect 471244 321632 471296 321638
rect 471244 321574 471296 321580
rect 469022 321399 469586 321405
rect 469022 321085 469586 321091
rect 470262 320314 470826 320320
rect 470262 320000 470826 320006
rect 470262 307086 470826 307092
rect 470262 306772 470826 306778
rect 471256 306338 471284 321574
rect 474278 321328 474334 321337
rect 484582 321328 484638 321337
rect 474334 321286 474680 321314
rect 474278 321263 474334 321272
rect 484638 321286 485012 321314
rect 484582 321263 484638 321272
rect 488170 321056 488226 321065
rect 478125 321014 478184 321042
rect 478156 320929 478184 321014
rect 481560 320929 481588 321042
rect 488226 321014 488456 321042
rect 488170 320991 488226 321000
rect 478142 320920 478198 320929
rect 478142 320855 478198 320864
rect 481546 320920 481602 320929
rect 481546 320855 481602 320864
rect 475476 320487 475528 320493
rect 475476 320429 475528 320435
rect 482376 320476 482428 320482
rect 475488 318782 475516 320429
rect 482376 320418 482428 320424
rect 479064 320408 479116 320414
rect 479064 320350 479116 320356
rect 479076 318782 479104 320350
rect 475476 318776 475528 318782
rect 475476 318718 475528 318724
rect 479064 318776 479116 318782
rect 479064 318718 479116 318724
rect 482388 318714 482416 320418
rect 485964 320408 486016 320414
rect 485964 320350 486016 320356
rect 482376 318708 482428 318714
rect 482376 318650 482428 318656
rect 485976 318646 486004 320350
rect 485964 318640 486016 318646
rect 485964 318582 486016 318588
rect 471244 306332 471296 306338
rect 471244 306274 471296 306280
rect 473728 306284 473780 306290
rect 469022 306001 469586 306007
rect 469022 305687 469586 305693
rect 470262 304914 470826 304920
rect 470262 304600 470826 304606
rect 470262 287487 470826 287493
rect 470262 287173 470826 287179
rect 471256 286686 471284 306274
rect 473728 306226 473780 306232
rect 473740 305969 473768 306226
rect 487525 306176 487534 306232
rect 487590 306176 487599 306232
rect 481004 306096 481060 306105
rect 481004 306031 481060 306040
rect 473726 305960 473782 305969
rect 473726 305895 473782 305904
rect 477739 305688 477795 305697
rect 477739 305623 477795 305632
rect 484122 305552 484178 305561
rect 484178 305510 484297 305538
rect 484122 305487 484178 305496
rect 478604 305448 478656 305454
rect 478604 305390 478656 305396
rect 485136 305448 485188 305454
rect 485136 305390 485188 305396
rect 475292 305088 475344 305094
rect 475292 305030 475344 305036
rect 475304 303618 475332 305030
rect 478616 303618 478644 305390
rect 481824 305088 481876 305094
rect 481824 305030 481876 305036
rect 481836 303618 481864 305030
rect 485148 303618 485176 305390
rect 490564 305040 490616 305046
rect 490564 304982 490616 304988
rect 475292 303612 475344 303618
rect 475292 303554 475344 303560
rect 478604 303612 478656 303618
rect 478604 303554 478656 303560
rect 481824 303612 481876 303618
rect 481824 303554 481876 303560
rect 485136 303612 485188 303618
rect 485136 303554 485188 303560
rect 490576 292534 490604 304982
rect 490760 298110 490788 409974
rect 491956 300830 491984 449346
rect 515404 445936 515456 445942
rect 515404 445878 515456 445884
rect 493324 441652 493376 441658
rect 493324 441594 493376 441600
rect 492036 431044 492088 431050
rect 492036 430986 492088 430992
rect 491944 300824 491996 300830
rect 491944 300766 491996 300772
rect 492048 299470 492076 430986
rect 493336 408474 493364 441594
rect 494704 440292 494756 440298
rect 494704 440234 494756 440240
rect 493324 408468 493376 408474
rect 493324 408410 493376 408416
rect 493324 389496 493376 389502
rect 493324 389438 493376 389444
rect 492128 356448 492180 356454
rect 492128 356390 492180 356396
rect 492036 299464 492088 299470
rect 492036 299406 492088 299412
rect 490748 298104 490800 298110
rect 490748 298046 490800 298052
rect 492140 296682 492168 356390
rect 492220 340400 492272 340406
rect 492220 340342 492272 340348
rect 492128 296676 492180 296682
rect 492128 296618 492180 296624
rect 492232 295322 492260 340342
rect 492312 320408 492364 320414
rect 492312 320350 492364 320356
rect 492220 295316 492272 295322
rect 492220 295258 492272 295264
rect 492324 293962 492352 320350
rect 493336 296614 493364 389438
rect 494716 387734 494744 440234
rect 496084 438932 496136 438938
rect 496084 438874 496136 438880
rect 494704 387728 494756 387734
rect 494704 387670 494756 387676
rect 496096 354550 496124 438874
rect 497464 437504 497516 437510
rect 497464 437446 497516 437452
rect 496084 354544 496136 354550
rect 496084 354486 496136 354492
rect 497476 339318 497504 437446
rect 498844 436144 498896 436150
rect 498844 436086 498896 436092
rect 497464 339312 497516 339318
rect 497464 339254 497516 339260
rect 498856 318578 498884 436086
rect 500224 434784 500276 434790
rect 500224 434726 500276 434732
rect 498844 318572 498896 318578
rect 498844 318514 498896 318520
rect 500236 303414 500264 434726
rect 501604 433356 501656 433362
rect 501604 433298 501656 433304
rect 500224 303408 500276 303414
rect 500224 303350 500276 303356
rect 493324 296608 493376 296614
rect 493324 296550 493376 296556
rect 492312 293956 492364 293962
rect 492312 293898 492364 293904
rect 490564 292528 490616 292534
rect 490564 292470 490616 292476
rect 492956 289876 493008 289882
rect 492956 289818 493008 289824
rect 491944 288448 491996 288454
rect 491944 288390 491996 288396
rect 478633 286920 478689 286929
rect 478633 286855 478689 286864
rect 471244 286680 471296 286686
rect 471244 286622 471296 286628
rect 474912 286592 474921 286648
rect 474977 286592 474986 286648
rect 478647 286620 478675 286855
rect 488632 286680 488684 286686
rect 488630 286648 488632 286657
rect 488684 286648 488686 286657
rect 488630 286583 488686 286592
rect 471704 286544 471756 286550
rect 471704 286486 471756 286492
rect 469022 286402 469586 286408
rect 469022 286088 469586 286094
rect 470262 285314 470826 285320
rect 470262 285000 470826 285006
rect 471716 270502 471744 286486
rect 479432 285864 479484 285870
rect 485870 285832 485926 285841
rect 479432 285806 479484 285812
rect 475752 285488 475804 285494
rect 475752 285430 475804 285436
rect 475764 284306 475792 285430
rect 479444 284306 479472 285806
rect 482336 285776 482345 285832
rect 482401 285776 482410 285832
rect 485926 285790 486085 285818
rect 485870 285767 485926 285776
rect 483204 285488 483256 285494
rect 483204 285430 483256 285436
rect 486884 285488 486936 285494
rect 486884 285430 486936 285436
rect 475752 284300 475804 284306
rect 475752 284242 475804 284248
rect 479432 284300 479484 284306
rect 479432 284242 479484 284248
rect 483216 284238 483244 285430
rect 483204 284232 483256 284238
rect 483204 284174 483256 284180
rect 486896 284170 486924 285430
rect 486884 284164 486936 284170
rect 486884 284106 486936 284112
rect 471704 270496 471756 270502
rect 471704 270438 471756 270444
rect 473728 270496 473780 270502
rect 473728 270438 473780 270444
rect 470262 267487 470826 267493
rect 470262 267173 470826 267179
rect 473740 266558 473768 270438
rect 473728 266552 473780 266558
rect 473728 266494 473780 266500
rect 469022 266401 469586 266407
rect 469022 266087 469586 266093
rect 470262 265314 470826 265320
rect 470262 265000 470826 265006
rect 473740 206990 473768 266494
rect 491956 266014 491984 288390
rect 492968 285666 492996 289818
rect 492956 285660 493008 285666
rect 492956 285602 493008 285608
rect 501616 284102 501644 433298
rect 502984 431996 503036 432002
rect 502984 431938 503036 431944
rect 501604 284096 501656 284102
rect 501604 284038 501656 284044
rect 491944 266008 491996 266014
rect 479062 265976 479118 265985
rect 479118 265948 479341 265962
rect 491944 265950 491996 265956
rect 479118 265934 479355 265948
rect 479062 265911 479118 265920
rect 477132 265872 477184 265878
rect 477132 265814 477184 265820
rect 476275 265690 476303 265812
rect 476275 265662 476344 265690
rect 476316 265010 476344 265662
rect 476486 265024 476542 265033
rect 476316 264982 476486 265010
rect 476486 264959 476542 264968
rect 477144 263566 477172 265814
rect 479327 265690 479355 265934
rect 482379 265690 482407 265812
rect 485431 265690 485459 265812
rect 479327 265662 479380 265690
rect 482379 265662 482416 265690
rect 485431 265662 485728 265690
rect 479352 265010 479380 265662
rect 480168 265487 480220 265493
rect 480168 265429 480220 265435
rect 479522 265024 479578 265033
rect 479352 264982 479522 265010
rect 479522 264959 479578 264968
rect 480180 263566 480208 265429
rect 482388 265010 482416 265662
rect 483204 265487 483256 265493
rect 483204 265429 483256 265435
rect 482834 265024 482890 265033
rect 482388 264982 482834 265010
rect 482834 264959 482890 264968
rect 483216 263566 483244 265429
rect 485700 265033 485728 265662
rect 488483 265554 488511 265812
rect 488722 265568 488778 265577
rect 488483 265526 488722 265554
rect 488722 265503 488778 265512
rect 486240 265487 486292 265493
rect 486240 265429 486292 265435
rect 485686 265024 485742 265033
rect 485686 264959 485742 264968
rect 486252 263566 486280 265429
rect 477132 263560 477184 263566
rect 477132 263502 477184 263508
rect 480168 263560 480220 263566
rect 480168 263502 480220 263508
rect 483204 263560 483256 263566
rect 483204 263502 483256 263508
rect 486240 263560 486292 263566
rect 495072 263560 495124 263566
rect 486240 263502 486292 263508
rect 494808 263508 495072 263514
rect 494808 263502 495124 263508
rect 494808 263498 495112 263502
rect 494796 263492 495112 263498
rect 494848 263486 495112 263492
rect 494796 263434 494848 263440
rect 502996 263362 503024 431938
rect 515416 409834 515444 445878
rect 520924 445868 520976 445874
rect 520924 445810 520976 445816
rect 515404 409828 515456 409834
rect 515404 409770 515456 409776
rect 515404 404388 515456 404394
rect 515404 404330 515456 404336
rect 515416 387802 515444 404330
rect 516784 403028 516836 403034
rect 516784 402970 516836 402976
rect 515404 387796 515456 387802
rect 515404 387738 515456 387744
rect 515404 365764 515456 365770
rect 515404 365706 515456 365712
rect 515416 339386 515444 365706
rect 516796 354618 516824 402970
rect 518164 398880 518216 398886
rect 518164 398822 518216 398828
rect 516784 354612 516836 354618
rect 516784 354554 516836 354560
rect 515404 339380 515456 339386
rect 515404 339322 515456 339328
rect 518176 303482 518204 398822
rect 519544 396092 519596 396098
rect 519544 396034 519596 396040
rect 518164 303476 518216 303482
rect 518164 303418 518216 303424
rect 519556 263430 519584 396034
rect 520936 373998 520964 445810
rect 523684 445800 523736 445806
rect 523684 445742 523736 445748
rect 522304 427848 522356 427854
rect 522304 427790 522356 427796
rect 520924 373992 520976 373998
rect 520924 373934 520976 373940
rect 522316 372570 522344 427790
rect 522304 372564 522356 372570
rect 522304 372506 522356 372512
rect 520924 367124 520976 367130
rect 520924 367066 520976 367072
rect 520936 354686 520964 367066
rect 522304 361616 522356 361622
rect 522304 361558 522356 361564
rect 520924 354680 520976 354686
rect 520924 354622 520976 354628
rect 522316 284238 522344 361558
rect 523696 338094 523724 445742
rect 535460 445732 535512 445738
rect 535460 445674 535512 445680
rect 535472 444825 535500 445674
rect 538692 445182 539258 445210
rect 546710 445182 547368 445210
rect 535458 444816 535514 444825
rect 535458 444751 535514 444760
rect 535458 443456 535514 443465
rect 535458 443391 535514 443400
rect 535472 443018 535500 443391
rect 535460 443012 535512 443018
rect 535460 442954 535512 442960
rect 535458 442096 535514 442105
rect 535458 442031 535514 442040
rect 535472 441658 535500 442031
rect 535460 441652 535512 441658
rect 535460 441594 535512 441600
rect 535458 440736 535514 440745
rect 535458 440671 535514 440680
rect 535472 440298 535500 440671
rect 535460 440292 535512 440298
rect 535460 440234 535512 440240
rect 535458 439376 535514 439385
rect 535458 439311 535514 439320
rect 535472 438938 535500 439311
rect 535460 438932 535512 438938
rect 535460 438874 535512 438880
rect 535458 438016 535514 438025
rect 535458 437951 535514 437960
rect 535472 437510 535500 437951
rect 535460 437504 535512 437510
rect 535460 437446 535512 437452
rect 535458 436656 535514 436665
rect 535458 436591 535514 436600
rect 535472 436150 535500 436591
rect 535460 436144 535512 436150
rect 535460 436086 535512 436092
rect 535458 435296 535514 435305
rect 535458 435231 535514 435240
rect 535472 434790 535500 435231
rect 535460 434784 535512 434790
rect 535460 434726 535512 434732
rect 535458 433936 535514 433945
rect 535458 433871 535514 433880
rect 535472 433362 535500 433871
rect 535460 433356 535512 433362
rect 535460 433298 535512 433304
rect 535458 432576 535514 432585
rect 535458 432511 535514 432520
rect 535472 432002 535500 432511
rect 535460 431996 535512 432002
rect 535460 431938 535512 431944
rect 536746 424416 536802 424425
rect 536746 424351 536802 424360
rect 535460 409828 535512 409834
rect 535460 409770 535512 409776
rect 535472 409329 535500 409770
rect 535458 409320 535514 409329
rect 535458 409255 535514 409264
rect 535460 407108 535512 407114
rect 535460 407050 535512 407056
rect 535472 406609 535500 407050
rect 535458 406600 535514 406609
rect 535458 406535 535514 406544
rect 535458 404560 535514 404569
rect 535458 404495 535514 404504
rect 535472 404394 535500 404495
rect 535460 404388 535512 404394
rect 535460 404330 535512 404336
rect 535458 403200 535514 403209
rect 535458 403135 535514 403144
rect 535472 403034 535500 403135
rect 535460 403028 535512 403034
rect 535460 402970 535512 402976
rect 536378 401704 536434 401713
rect 536378 401639 536434 401648
rect 536286 400344 536342 400353
rect 536286 400279 536342 400288
rect 535458 399120 535514 399129
rect 535458 399055 535514 399064
rect 535472 398886 535500 399055
rect 535460 398880 535512 398886
rect 535460 398822 535512 398828
rect 536102 397488 536158 397497
rect 536102 397423 536158 397432
rect 535458 396400 535514 396409
rect 535458 396335 535514 396344
rect 535472 396098 535500 396335
rect 535460 396092 535512 396098
rect 535460 396034 535512 396040
rect 535460 373992 535512 373998
rect 535460 373934 535512 373940
rect 535472 372881 535500 373934
rect 535458 372872 535514 372881
rect 535458 372807 535514 372816
rect 535460 372564 535512 372570
rect 535460 372506 535512 372512
rect 535472 371521 535500 372506
rect 535458 371512 535514 371521
rect 535458 371447 535514 371456
rect 535460 369844 535512 369850
rect 535460 369786 535512 369792
rect 535472 368801 535500 369786
rect 535458 368792 535514 368801
rect 535458 368727 535514 368736
rect 535458 367432 535514 367441
rect 535458 367367 535514 367376
rect 535472 367130 535500 367367
rect 535460 367124 535512 367130
rect 535460 367066 535512 367072
rect 535458 366072 535514 366081
rect 535458 366007 535514 366016
rect 535472 365770 535500 366007
rect 535460 365764 535512 365770
rect 535460 365706 535512 365712
rect 535458 361992 535514 362001
rect 535458 361927 535514 361936
rect 535472 361622 535500 361927
rect 535460 361616 535512 361622
rect 535460 361558 535512 361564
rect 525064 353320 525116 353326
rect 525064 353262 525116 353268
rect 523684 338088 523736 338094
rect 523684 338030 523736 338036
rect 525076 332586 525104 353262
rect 535460 338088 535512 338094
rect 535460 338030 535512 338036
rect 535472 336841 535500 338030
rect 535458 336832 535514 336841
rect 535458 336767 535514 336776
rect 525064 332580 525116 332586
rect 525064 332522 525116 332528
rect 535460 332580 535512 332586
rect 535460 332522 535512 332528
rect 535472 331401 535500 332522
rect 535458 331392 535514 331401
rect 535458 331327 535514 331336
rect 535460 331220 535512 331226
rect 535460 331162 535512 331168
rect 535472 330041 535500 331162
rect 535458 330032 535514 330041
rect 535458 329967 535514 329976
rect 536010 328672 536066 328681
rect 536010 328607 536066 328616
rect 535458 325952 535514 325961
rect 535458 325887 535514 325896
rect 535472 325718 535500 325887
rect 523684 325712 523736 325718
rect 523684 325654 523736 325660
rect 535460 325712 535512 325718
rect 535460 325654 535512 325660
rect 522304 284232 522356 284238
rect 522304 284174 522356 284180
rect 523696 284170 523724 325654
rect 536024 318646 536052 328607
rect 536012 318640 536064 318646
rect 536012 318582 536064 318588
rect 535460 300824 535512 300830
rect 535458 300792 535460 300801
rect 535512 300792 535514 300801
rect 535458 300727 535514 300736
rect 535460 299464 535512 299470
rect 535458 299432 535460 299441
rect 535512 299432 535514 299441
rect 535458 299367 535514 299376
rect 535460 298104 535512 298110
rect 535458 298072 535460 298081
rect 535512 298072 535514 298081
rect 535458 298007 535514 298016
rect 535458 296712 535514 296721
rect 535458 296647 535514 296656
rect 535552 296676 535604 296682
rect 535472 296614 535500 296647
rect 535552 296618 535604 296624
rect 535460 296608 535512 296614
rect 535460 296550 535512 296556
rect 535564 295361 535592 296618
rect 535550 295352 535606 295361
rect 535460 295316 535512 295322
rect 535550 295287 535606 295296
rect 535460 295258 535512 295264
rect 535472 294001 535500 295258
rect 535458 293992 535514 294001
rect 535458 293927 535514 293936
rect 535552 293956 535604 293962
rect 535552 293898 535604 293904
rect 535564 292641 535592 293898
rect 535550 292632 535606 292641
rect 535550 292567 535606 292576
rect 535460 292528 535512 292534
rect 535460 292470 535512 292476
rect 535472 291281 535500 292470
rect 535458 291272 535514 291281
rect 535458 291207 535514 291216
rect 535458 289912 535514 289921
rect 535458 289847 535460 289856
rect 535512 289847 535514 289856
rect 535460 289818 535512 289824
rect 535458 288552 535514 288561
rect 535458 288487 535514 288496
rect 535472 288454 535500 288487
rect 535460 288448 535512 288454
rect 535460 288390 535512 288396
rect 536116 284306 536144 397423
rect 536194 360632 536250 360641
rect 536194 360567 536250 360576
rect 536104 284300 536156 284306
rect 536104 284242 536156 284248
rect 523684 284164 523736 284170
rect 523684 284106 523736 284112
rect 536102 280392 536158 280401
rect 536102 280327 536158 280336
rect 519544 263424 519596 263430
rect 519544 263366 519596 263372
rect 502984 263356 503036 263362
rect 502984 263298 503036 263304
rect 473728 206984 473780 206990
rect 473728 206926 473780 206932
rect 536116 69902 536144 280327
rect 536208 263566 536236 360567
rect 536300 318782 536328 400279
rect 536392 339454 536420 401639
rect 536760 396001 536788 424351
rect 538692 422294 538720 445182
rect 541714 445088 541770 445097
rect 541714 445023 541770 445032
rect 544198 445088 544254 445097
rect 544198 445023 544254 445032
rect 538692 422266 538904 422294
rect 538876 409170 538904 422266
rect 547340 412634 547368 445182
rect 547064 412606 547368 412634
rect 547064 409714 547092 412606
rect 546710 409686 547368 409714
rect 541714 409320 541770 409329
rect 544290 409320 544346 409329
rect 544226 409278 544290 409306
rect 541714 409255 541770 409264
rect 544290 409255 544346 409264
rect 538784 409142 539258 409170
rect 536746 395992 536802 396001
rect 536746 395927 536802 395936
rect 538784 393314 538812 409142
rect 547340 404977 547368 409686
rect 547326 404968 547382 404977
rect 547326 404903 547382 404912
rect 538692 393286 538812 393314
rect 536746 388376 536802 388385
rect 536746 388311 536802 388320
rect 536562 364712 536618 364721
rect 536562 364647 536618 364656
rect 536470 363352 536526 363361
rect 536470 363287 536526 363296
rect 536380 339448 536432 339454
rect 536380 339390 536432 339396
rect 536378 324592 536434 324601
rect 536378 324527 536434 324536
rect 536288 318776 536340 318782
rect 536288 318718 536340 318724
rect 536196 263560 536248 263566
rect 536196 263502 536248 263508
rect 536392 263498 536420 324527
rect 536484 303618 536512 363287
rect 536576 318714 536604 364647
rect 536760 359281 536788 388311
rect 538692 383654 538720 393286
rect 538692 383626 538812 383654
rect 538784 373266 538812 383626
rect 547340 373994 547368 404903
rect 547064 373966 547368 373994
rect 544474 373416 544530 373425
rect 544226 373374 544474 373402
rect 544474 373351 544530 373360
rect 547064 373266 547092 373966
rect 538784 373238 539258 373266
rect 546710 373238 547092 373266
rect 536746 359272 536802 359281
rect 536746 359207 536802 359216
rect 538784 354674 538812 373238
rect 541714 373144 541770 373153
rect 541714 373079 541770 373088
rect 547064 364334 547092 373238
rect 547064 364306 547368 364334
rect 538692 354646 538812 354674
rect 536746 352472 536802 352481
rect 536746 352407 536802 352416
rect 536654 327312 536710 327321
rect 536654 327247 536710 327256
rect 536564 318708 536616 318714
rect 536564 318650 536616 318656
rect 536472 303612 536524 303618
rect 536472 303554 536524 303560
rect 536668 303550 536696 327247
rect 536760 323241 536788 352407
rect 538692 345014 538720 354646
rect 547340 345014 547368 364306
rect 538692 344986 538904 345014
rect 538876 337770 538904 344986
rect 547064 344986 547368 345014
rect 541714 339552 541770 339561
rect 541714 339487 541770 339496
rect 544198 339552 544254 339561
rect 544198 339487 544254 339496
rect 538784 337742 539258 337770
rect 541728 337756 541756 339487
rect 544212 337756 544240 339487
rect 547064 337770 547092 344986
rect 546710 337742 547092 337770
rect 536746 323232 536802 323241
rect 536746 323167 536802 323176
rect 536746 316432 536802 316441
rect 536746 316367 536802 316376
rect 536656 303544 536708 303550
rect 536656 303486 536708 303492
rect 536760 287201 536788 316367
rect 538784 316034 538812 337742
rect 547064 335354 547092 337742
rect 547064 335326 547460 335354
rect 538784 316006 538904 316034
rect 538876 301730 538904 316006
rect 547432 306374 547460 335326
rect 547064 306346 547460 306374
rect 544198 303784 544254 303793
rect 544198 303719 544254 303728
rect 541714 303648 541770 303657
rect 541714 303583 541770 303592
rect 538692 301702 539258 301730
rect 541728 301716 541756 303583
rect 544212 301716 544240 303719
rect 547064 301730 547092 306346
rect 547326 303648 547382 303657
rect 547326 303583 547382 303592
rect 546710 301702 547092 301730
rect 536746 287192 536802 287201
rect 536746 287127 536802 287136
rect 536380 263492 536432 263498
rect 536380 263434 536432 263440
rect 538692 245585 538720 301702
rect 547340 300121 547368 303583
rect 547326 300112 547382 300121
rect 547326 300047 547382 300056
rect 580170 300112 580226 300121
rect 580170 300047 580226 300056
rect 580184 298761 580212 300047
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 538678 245576 538734 245585
rect 538678 245511 538734 245520
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 536104 69896 536156 69902
rect 536104 69838 536156 69844
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 470276 451183 470812 451479
rect 469036 450097 469572 450393
rect 470276 449012 470812 449308
rect 470276 432784 470812 433080
rect 477843 450200 477899 450256
rect 481160 450200 481216 450256
rect 484477 450200 484533 450256
rect 487793 450200 487849 450256
rect 474094 449656 474150 449712
rect 469036 431697 469572 431993
rect 470276 430612 470812 430908
rect 470276 411784 470812 412080
rect 483570 432248 483626 432304
rect 481270 432112 481326 432168
rect 474278 431840 474334 431896
rect 488078 431840 488134 431896
rect 478102 431568 478158 431624
rect 478970 427896 479026 427952
rect 485778 427896 485834 427952
rect 469036 410698 469572 410994
rect 470276 409612 470812 409908
rect 470276 390785 470812 391081
rect 473726 410896 473782 410952
rect 478418 410080 478474 410136
rect 484122 410352 484178 410408
rect 481362 410080 481418 410136
rect 487802 410080 487858 410136
rect 481822 407088 481878 407144
rect 485134 407088 485190 407144
rect 488538 390088 488594 390144
rect 469036 389702 469572 389998
rect 470276 388612 470812 388908
rect 470276 358185 470812 358481
rect 474922 389272 474978 389328
rect 478634 389272 478690 389328
rect 482098 389408 482154 389464
rect 486882 386416 486938 386472
rect 478878 357992 478934 358048
rect 481822 357992 481878 358048
rect 484950 357992 485006 358048
rect 488354 357992 488410 358048
rect 469036 357099 469572 357395
rect 470276 356012 470812 356308
rect 475014 357448 475070 357504
rect 470276 342184 470812 342480
rect 469036 341097 469572 341393
rect 470276 340012 470812 340308
rect 470276 322184 470812 322480
rect 477915 340992 477971 341048
rect 481232 340992 481288 341048
rect 484398 340992 484454 341048
rect 487894 340992 487950 341048
rect 474554 340448 474610 340504
rect 469036 321097 469572 321393
rect 470276 320012 470812 320308
rect 470276 306784 470812 307080
rect 474278 321272 474334 321328
rect 484582 321272 484638 321328
rect 488170 321000 488226 321056
rect 478142 320864 478198 320920
rect 481546 320864 481602 320920
rect 469036 305699 469572 305995
rect 470276 304612 470812 304908
rect 470276 287185 470812 287481
rect 487534 306176 487590 306232
rect 481004 306040 481060 306096
rect 473726 305904 473782 305960
rect 477739 305632 477795 305688
rect 484122 305496 484178 305552
rect 478633 286864 478689 286920
rect 474921 286592 474977 286648
rect 488630 286628 488632 286648
rect 488632 286628 488684 286648
rect 488684 286628 488686 286648
rect 488630 286592 488686 286628
rect 469036 286100 469572 286396
rect 470276 285012 470812 285308
rect 482345 285776 482401 285832
rect 485870 285776 485926 285832
rect 470276 267185 470812 267481
rect 469036 266099 469572 266395
rect 470276 265012 470812 265308
rect 479062 265920 479118 265976
rect 476486 264968 476542 265024
rect 479522 264968 479578 265024
rect 482834 264968 482890 265024
rect 488722 265512 488778 265568
rect 485686 264968 485742 265024
rect 535458 444760 535514 444816
rect 535458 443400 535514 443456
rect 535458 442040 535514 442096
rect 535458 440680 535514 440736
rect 535458 439320 535514 439376
rect 535458 437960 535514 438016
rect 535458 436600 535514 436656
rect 535458 435240 535514 435296
rect 535458 433880 535514 433936
rect 535458 432520 535514 432576
rect 536746 424360 536802 424416
rect 535458 409264 535514 409320
rect 535458 406544 535514 406600
rect 535458 404504 535514 404560
rect 535458 403144 535514 403200
rect 536378 401648 536434 401704
rect 536286 400288 536342 400344
rect 535458 399064 535514 399120
rect 536102 397432 536158 397488
rect 535458 396344 535514 396400
rect 535458 372816 535514 372872
rect 535458 371456 535514 371512
rect 535458 368736 535514 368792
rect 535458 367376 535514 367432
rect 535458 366016 535514 366072
rect 535458 361936 535514 361992
rect 535458 336776 535514 336832
rect 535458 331336 535514 331392
rect 535458 329976 535514 330032
rect 536010 328616 536066 328672
rect 535458 325896 535514 325952
rect 535458 300772 535460 300792
rect 535460 300772 535512 300792
rect 535512 300772 535514 300792
rect 535458 300736 535514 300772
rect 535458 299412 535460 299432
rect 535460 299412 535512 299432
rect 535512 299412 535514 299432
rect 535458 299376 535514 299412
rect 535458 298052 535460 298072
rect 535460 298052 535512 298072
rect 535512 298052 535514 298072
rect 535458 298016 535514 298052
rect 535458 296656 535514 296712
rect 535550 295296 535606 295352
rect 535458 293936 535514 293992
rect 535550 292576 535606 292632
rect 535458 291216 535514 291272
rect 535458 289876 535514 289912
rect 535458 289856 535460 289876
rect 535460 289856 535512 289876
rect 535512 289856 535514 289876
rect 535458 288496 535514 288552
rect 536194 360576 536250 360632
rect 536102 280336 536158 280392
rect 541714 445032 541770 445088
rect 544198 445032 544254 445088
rect 541714 409264 541770 409320
rect 544290 409264 544346 409320
rect 536746 395936 536802 395992
rect 547326 404912 547382 404968
rect 536746 388320 536802 388376
rect 536562 364656 536618 364712
rect 536470 363296 536526 363352
rect 536378 324536 536434 324592
rect 544474 373360 544530 373416
rect 536746 359216 536802 359272
rect 541714 373088 541770 373144
rect 536746 352416 536802 352472
rect 536654 327256 536710 327312
rect 541714 339496 541770 339552
rect 544198 339496 544254 339552
rect 536746 323176 536802 323232
rect 536746 316376 536802 316432
rect 544198 303728 544254 303784
rect 541714 303592 541770 303648
rect 547326 303592 547382 303648
rect 536746 287136 536802 287192
rect 547326 300056 547382 300112
rect 580170 300056 580226 300112
rect 580170 298696 580226 298752
rect 538678 245520 538734 245576
rect 580170 205672 580226 205728
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 470266 451483 470822 451484
rect 470266 451179 470272 451483
rect 470816 451179 470822 451483
rect 470266 451178 470822 451179
rect 469026 450397 469582 450398
rect 469026 450093 469032 450397
rect 469576 450093 469582 450397
rect 477838 450258 477904 450261
rect 481155 450260 481221 450261
rect 478454 450258 478460 450260
rect 477838 450256 478460 450258
rect 477838 450200 477843 450256
rect 477899 450200 478460 450256
rect 477838 450198 478460 450200
rect 477838 450195 477904 450198
rect 478454 450196 478460 450198
rect 478524 450196 478530 450260
rect 481155 450256 481220 450260
rect 481155 450200 481160 450256
rect 481216 450200 481220 450256
rect 481155 450196 481220 450200
rect 481284 450258 481290 450260
rect 481284 450198 481312 450258
rect 481284 450196 481290 450198
rect 484158 450196 484164 450260
rect 484228 450258 484234 450260
rect 484472 450258 484538 450261
rect 484228 450256 484538 450258
rect 484228 450200 484477 450256
rect 484533 450200 484538 450256
rect 484228 450198 484538 450200
rect 484228 450196 484234 450198
rect 481155 450195 481221 450196
rect 484472 450195 484538 450198
rect 487788 450260 487854 450261
rect 487788 450256 487844 450260
rect 487908 450258 487914 450260
rect 487788 450200 487793 450256
rect 487788 450196 487844 450200
rect 487908 450198 487945 450258
rect 487908 450196 487914 450198
rect 487788 450195 487854 450196
rect 469026 450092 469582 450093
rect -960 449428 480 449668
rect 473670 449652 473676 449716
rect 473740 449714 473746 449716
rect 474089 449714 474155 449717
rect 473740 449712 474155 449714
rect 473740 449656 474094 449712
rect 474150 449656 474155 449712
rect 473740 449654 474155 449656
rect 473740 449652 473746 449654
rect 474089 449651 474155 449654
rect 470266 449312 470822 449313
rect 470266 449008 470272 449312
rect 470816 449008 470822 449312
rect 470266 449007 470822 449008
rect 541566 445028 541572 445092
rect 541636 445090 541642 445092
rect 541709 445090 541775 445093
rect 541636 445088 541775 445090
rect 541636 445032 541714 445088
rect 541770 445032 541775 445088
rect 541636 445030 541775 445032
rect 541636 445028 541642 445030
rect 541709 445027 541775 445030
rect 544193 445090 544259 445093
rect 544326 445090 544332 445092
rect 544193 445088 544332 445090
rect 544193 445032 544198 445088
rect 544254 445032 544332 445088
rect 544193 445030 544332 445032
rect 544193 445027 544259 445030
rect 544326 445028 544332 445030
rect 544396 445028 544402 445092
rect 535453 444818 535519 444821
rect 535453 444816 538108 444818
rect 535453 444760 535458 444816
rect 535514 444760 538108 444816
rect 535453 444758 538108 444760
rect 535453 444755 535519 444758
rect 583520 444668 584960 444908
rect 535453 443458 535519 443461
rect 535453 443456 538108 443458
rect 535453 443400 535458 443456
rect 535514 443400 538108 443456
rect 535453 443398 538108 443400
rect 535453 443395 535519 443398
rect 535453 442098 535519 442101
rect 535453 442096 538108 442098
rect 535453 442040 535458 442096
rect 535514 442040 538108 442096
rect 535453 442038 538108 442040
rect 535453 442035 535519 442038
rect 535453 440738 535519 440741
rect 535453 440736 538108 440738
rect 535453 440680 535458 440736
rect 535514 440680 538108 440736
rect 535453 440678 538108 440680
rect 535453 440675 535519 440678
rect 535453 439378 535519 439381
rect 535453 439376 538108 439378
rect 535453 439320 535458 439376
rect 535514 439320 538108 439376
rect 535453 439318 538108 439320
rect 535453 439315 535519 439318
rect 535453 438018 535519 438021
rect 535453 438016 538108 438018
rect 535453 437960 535458 438016
rect 535514 437960 538108 438016
rect 535453 437958 538108 437960
rect 535453 437955 535519 437958
rect -960 436508 480 436748
rect 535453 436658 535519 436661
rect 535453 436656 538108 436658
rect 535453 436600 535458 436656
rect 535514 436600 538108 436656
rect 535453 436598 538108 436600
rect 535453 436595 535519 436598
rect 535453 435298 535519 435301
rect 535453 435296 538108 435298
rect 535453 435240 535458 435296
rect 535514 435240 538108 435296
rect 535453 435238 538108 435240
rect 535453 435235 535519 435238
rect 549294 434754 549300 434756
rect 547860 434694 549300 434754
rect 549294 434692 549300 434694
rect 549364 434692 549370 434756
rect 535453 433938 535519 433941
rect 535453 433936 538108 433938
rect 535453 433880 535458 433936
rect 535514 433880 538108 433936
rect 535453 433878 538108 433880
rect 535453 433875 535519 433878
rect 470266 433084 470822 433085
rect 470266 432780 470272 433084
rect 470816 432780 470822 433084
rect 470266 432779 470822 432780
rect 535453 432578 535519 432581
rect 535453 432576 538108 432578
rect 535453 432520 535458 432576
rect 535514 432520 538108 432576
rect 535453 432518 538108 432520
rect 535453 432515 535519 432518
rect 483565 432308 483631 432309
rect 483565 432306 483612 432308
rect 483520 432304 483612 432306
rect 483520 432248 483570 432304
rect 483520 432246 483612 432248
rect 483565 432244 483612 432246
rect 483676 432244 483682 432308
rect 483565 432243 483631 432244
rect 481265 432172 481331 432173
rect 481214 432108 481220 432172
rect 481284 432170 481331 432172
rect 481284 432168 481376 432170
rect 481326 432112 481376 432168
rect 481284 432110 481376 432112
rect 481284 432108 481331 432110
rect 481265 432107 481331 432108
rect 469026 431997 469582 431998
rect 469026 431693 469032 431997
rect 469576 431693 469582 431997
rect 473670 431836 473676 431900
rect 473740 431898 473746 431900
rect 474273 431898 474339 431901
rect 473740 431896 474339 431898
rect 473740 431840 474278 431896
rect 474334 431840 474339 431896
rect 473740 431838 474339 431840
rect 473740 431836 473746 431838
rect 474273 431835 474339 431838
rect 487654 431836 487660 431900
rect 487724 431898 487730 431900
rect 488073 431898 488139 431901
rect 487724 431896 488139 431898
rect 487724 431840 488078 431896
rect 488134 431840 488139 431896
rect 487724 431838 488139 431840
rect 487724 431836 487730 431838
rect 488073 431835 488139 431838
rect 469026 431692 469582 431693
rect 478097 431626 478163 431629
rect 478454 431626 478460 431628
rect 478097 431624 478460 431626
rect 478097 431568 478102 431624
rect 478158 431568 478460 431624
rect 478097 431566 478460 431568
rect 478097 431563 478163 431566
rect 478454 431564 478460 431566
rect 478524 431564 478530 431628
rect 583520 431476 584960 431716
rect 470266 430912 470822 430913
rect 470266 430608 470272 430912
rect 470816 430608 470822 430912
rect 470266 430607 470822 430608
rect 478965 427954 479031 427957
rect 480110 427954 480116 427956
rect 478965 427952 480116 427954
rect 478965 427896 478970 427952
rect 479026 427896 480116 427952
rect 478965 427894 480116 427896
rect 478965 427891 479031 427894
rect 480110 427892 480116 427894
rect 480180 427892 480186 427956
rect 485773 427954 485839 427957
rect 486550 427954 486556 427956
rect 485773 427952 486556 427954
rect 485773 427896 485778 427952
rect 485834 427896 486556 427952
rect 485773 427894 486556 427896
rect 485773 427891 485839 427894
rect 486550 427892 486556 427894
rect 486620 427892 486626 427956
rect 536741 424418 536807 424421
rect 538078 424418 538138 431188
rect 536741 424416 538138 424418
rect 536741 424360 536746 424416
rect 536802 424388 538138 424416
rect 536802 424360 538108 424388
rect 536741 424358 538108 424360
rect 536741 424355 536807 424358
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 470266 412084 470822 412085
rect 470266 411780 470272 412084
rect 470816 411780 470822 412084
rect 470266 411779 470822 411780
rect 469026 410998 469582 410999
rect 469026 410694 469032 410998
rect 469576 410694 469582 410998
rect 473721 410956 473787 410957
rect 473670 410892 473676 410956
rect 473740 410954 473787 410956
rect 473740 410952 473832 410954
rect 473782 410896 473832 410952
rect 473740 410894 473832 410896
rect 473740 410892 473787 410894
rect 473721 410891 473787 410892
rect 469026 410693 469582 410694
rect -960 410396 480 410636
rect 484117 410412 484183 410413
rect 484117 410410 484164 410412
rect 484072 410408 484164 410410
rect 484072 410352 484122 410408
rect 484072 410350 484164 410352
rect 484117 410348 484164 410350
rect 484228 410348 484234 410412
rect 484117 410347 484183 410348
rect 478413 410140 478479 410141
rect 481357 410140 481423 410141
rect 487797 410140 487863 410141
rect 478413 410138 478460 410140
rect 478368 410136 478460 410138
rect 478368 410080 478418 410136
rect 478368 410078 478460 410080
rect 478413 410076 478460 410078
rect 478524 410076 478530 410140
rect 481357 410138 481404 410140
rect 481312 410136 481404 410138
rect 481312 410080 481362 410136
rect 481312 410078 481404 410080
rect 481357 410076 481404 410078
rect 481468 410076 481474 410140
rect 487797 410138 487844 410140
rect 487756 410136 487844 410138
rect 487908 410138 487914 410140
rect 488390 410138 488396 410140
rect 487756 410080 487802 410136
rect 487756 410078 487844 410080
rect 487797 410076 487844 410078
rect 487908 410078 488396 410138
rect 487908 410076 487914 410078
rect 488390 410076 488396 410078
rect 488460 410076 488466 410140
rect 478413 410075 478479 410076
rect 481357 410075 481423 410076
rect 487797 410075 487863 410076
rect 470266 409912 470822 409913
rect 470266 409608 470272 409912
rect 470816 409608 470822 409912
rect 470266 409607 470822 409608
rect 535453 409322 535519 409325
rect 535453 409320 538138 409322
rect 535453 409264 535458 409320
rect 535514 409264 538138 409320
rect 535453 409262 538138 409264
rect 535453 409259 535519 409262
rect 538078 408816 538138 409262
rect 541566 409260 541572 409324
rect 541636 409322 541642 409324
rect 541709 409322 541775 409325
rect 544285 409324 544351 409325
rect 544285 409322 544332 409324
rect 541636 409320 541775 409322
rect 541636 409264 541714 409320
rect 541770 409264 541775 409320
rect 541636 409262 541775 409264
rect 544240 409320 544332 409322
rect 544240 409264 544290 409320
rect 544240 409262 544332 409264
rect 541636 409260 541642 409262
rect 541709 409259 541775 409262
rect 544285 409260 544332 409262
rect 544396 409260 544402 409324
rect 544285 409259 544351 409260
rect 480110 407492 480116 407556
rect 480180 407554 480186 407556
rect 480180 407494 538138 407554
rect 480180 407492 480186 407494
rect 538078 407456 538138 407494
rect 481817 407146 481883 407149
rect 482870 407146 482876 407148
rect 481817 407144 482876 407146
rect 481817 407088 481822 407144
rect 481878 407088 482876 407144
rect 481817 407086 482876 407088
rect 481817 407083 481883 407086
rect 482870 407084 482876 407086
rect 482940 407084 482946 407148
rect 485129 407146 485195 407149
rect 485630 407146 485636 407148
rect 485129 407144 485636 407146
rect 485129 407088 485134 407144
rect 485190 407088 485636 407144
rect 485129 407086 485636 407088
rect 485129 407083 485195 407086
rect 485630 407084 485636 407086
rect 485700 407084 485706 407148
rect 535453 406602 535519 406605
rect 535453 406600 538138 406602
rect 535453 406544 535458 406600
rect 535514 406544 538138 406600
rect 535453 406542 538138 406544
rect 535453 406539 535519 406542
rect 538078 406096 538138 406542
rect 547321 404970 547387 404973
rect 583520 404970 584960 405060
rect 547321 404968 584960 404970
rect 547321 404912 547326 404968
rect 547382 404912 584960 404968
rect 547321 404910 584960 404912
rect 547321 404907 547387 404910
rect 583520 404820 584960 404910
rect 535453 404562 535519 404565
rect 538078 404562 538138 404736
rect 535453 404560 538138 404562
rect 535453 404504 535458 404560
rect 535514 404504 538138 404560
rect 535453 404502 538138 404504
rect 535453 404499 535519 404502
rect 535453 403202 535519 403205
rect 538078 403202 538138 403376
rect 535453 403200 538138 403202
rect 535453 403144 535458 403200
rect 535514 403144 538138 403200
rect 535453 403142 538138 403144
rect 535453 403139 535519 403142
rect 536373 401706 536439 401709
rect 538078 401706 538138 402016
rect 536373 401704 538138 401706
rect 536373 401648 536378 401704
rect 536434 401648 538138 401704
rect 536373 401646 538138 401648
rect 536373 401643 536439 401646
rect 536281 400346 536347 400349
rect 538078 400346 538138 400656
rect 536281 400344 538138 400346
rect 536281 400288 536286 400344
rect 536342 400288 538138 400344
rect 536281 400286 538138 400288
rect 536281 400283 536347 400286
rect 535453 399122 535519 399125
rect 538078 399122 538138 399296
rect 535453 399120 538138 399122
rect 535453 399064 535458 399120
rect 535514 399064 538138 399120
rect 535453 399062 538138 399064
rect 535453 399059 535519 399062
rect 547830 398306 547890 398752
rect 549294 398306 549300 398308
rect 547830 398246 549300 398306
rect 549294 398244 549300 398246
rect 549364 398244 549370 398308
rect -960 397340 480 397580
rect 536097 397490 536163 397493
rect 538078 397490 538138 397936
rect 536097 397488 538138 397490
rect 536097 397432 536102 397488
rect 536158 397432 538138 397488
rect 536097 397430 538138 397432
rect 536097 397427 536163 397430
rect 535453 396402 535519 396405
rect 538078 396402 538138 396576
rect 535453 396400 538138 396402
rect 535453 396344 535458 396400
rect 535514 396344 538138 396400
rect 535453 396342 538138 396344
rect 535453 396339 535519 396342
rect 536741 395994 536807 395997
rect 536741 395992 538138 395994
rect 536741 395936 536746 395992
rect 536802 395936 538138 395992
rect 536741 395934 538138 395936
rect 536741 395931 536807 395934
rect 473670 391988 473676 392052
rect 473740 392050 473746 392052
rect 474958 392050 474964 392052
rect 473740 391990 474964 392050
rect 473740 391988 473746 391990
rect 474958 391988 474964 391990
rect 475028 391988 475034 392052
rect 470266 391085 470822 391086
rect 470266 390781 470272 391085
rect 470816 390781 470822 391085
rect 470266 390780 470822 390781
rect 484900 390297 484964 390303
rect 484900 390227 484964 390233
rect 488390 390084 488396 390148
rect 488460 390146 488466 390148
rect 488533 390146 488599 390149
rect 488460 390144 488599 390146
rect 488460 390088 488538 390144
rect 488594 390088 488599 390144
rect 488460 390086 488599 390088
rect 488460 390084 488466 390086
rect 488533 390083 488599 390086
rect 469026 390002 469582 390003
rect 469026 389698 469032 390002
rect 469576 389698 469582 390002
rect 469026 389697 469582 389698
rect 481766 389404 481772 389468
rect 481836 389466 481842 389468
rect 482093 389466 482159 389469
rect 481836 389464 482159 389466
rect 481836 389408 482098 389464
rect 482154 389408 482159 389464
rect 481836 389406 482159 389408
rect 481836 389404 481842 389406
rect 482093 389403 482159 389406
rect 474917 389332 474983 389333
rect 478629 389332 478695 389333
rect 474917 389330 474964 389332
rect 474872 389328 474964 389330
rect 474872 389272 474922 389328
rect 474872 389270 474964 389272
rect 474917 389268 474964 389270
rect 475028 389268 475034 389332
rect 478629 389330 478644 389332
rect 478552 389328 478644 389330
rect 478552 389272 478634 389328
rect 478552 389270 478644 389272
rect 478629 389268 478644 389270
rect 478708 389268 478714 389332
rect 474917 389267 474983 389268
rect 478629 389267 478695 389268
rect 470266 388912 470822 388913
rect 470266 388608 470272 388912
rect 470816 388608 470822 388912
rect 470266 388607 470822 388608
rect 536741 388378 536807 388381
rect 538078 388378 538138 395934
rect 583520 391628 584960 391868
rect 536741 388376 538138 388378
rect 536741 388320 536746 388376
rect 536802 388320 538138 388376
rect 536741 388318 538138 388320
rect 536741 388315 536807 388318
rect 486734 386412 486740 386476
rect 486804 386474 486810 386476
rect 486877 386474 486943 386477
rect 486804 386472 486943 386474
rect 486804 386416 486882 386472
rect 486938 386416 486943 386472
rect 486804 386414 486943 386416
rect 486804 386412 486810 386414
rect 486877 386411 486943 386414
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect 544469 373420 544535 373421
rect 544469 373418 544516 373420
rect 544424 373416 544516 373418
rect 544424 373360 544474 373416
rect 544424 373358 544516 373360
rect 544469 373356 544516 373358
rect 544580 373356 544586 373420
rect 544469 373355 544535 373356
rect 541566 373084 541572 373148
rect 541636 373146 541642 373148
rect 541709 373146 541775 373149
rect 541636 373144 541775 373146
rect 541636 373088 541714 373144
rect 541770 373088 541775 373144
rect 541636 373086 541775 373088
rect 541636 373084 541642 373086
rect 541709 373083 541775 373086
rect 535453 372874 535519 372877
rect 535453 372872 538108 372874
rect 535453 372816 535458 372872
rect 535514 372816 538108 372872
rect 535453 372814 538108 372816
rect 535453 372811 535519 372814
rect 535453 371514 535519 371517
rect 535453 371512 538108 371514
rect -960 371228 480 371468
rect 535453 371456 535458 371512
rect 535514 371456 538108 371512
rect 535453 371454 538108 371456
rect 535453 371451 535519 371454
rect 482870 370092 482876 370156
rect 482940 370154 482946 370156
rect 482940 370094 538108 370154
rect 482940 370092 482946 370094
rect 535453 368794 535519 368797
rect 535453 368792 538108 368794
rect 535453 368736 535458 368792
rect 535514 368736 538108 368792
rect 535453 368734 538108 368736
rect 535453 368731 535519 368734
rect 535453 367434 535519 367437
rect 535453 367432 538108 367434
rect 535453 367376 535458 367432
rect 535514 367376 538108 367432
rect 535453 367374 538108 367376
rect 535453 367371 535519 367374
rect 535453 366074 535519 366077
rect 535453 366072 538108 366074
rect 535453 366016 535458 366072
rect 535514 366016 538108 366072
rect 535453 366014 538108 366016
rect 535453 366011 535519 366014
rect 583520 364972 584960 365212
rect 536557 364714 536623 364717
rect 536557 364712 538108 364714
rect 536557 364656 536562 364712
rect 536618 364656 538108 364712
rect 536557 364654 538108 364656
rect 536557 364651 536623 364654
rect 536465 363354 536531 363357
rect 536465 363352 538108 363354
rect 536465 363296 536470 363352
rect 536526 363296 538108 363352
rect 536465 363294 538108 363296
rect 536465 363291 536531 363294
rect 549294 362810 549300 362812
rect 547860 362750 549300 362810
rect 549294 362748 549300 362750
rect 549364 362748 549370 362812
rect 535453 361994 535519 361997
rect 535453 361992 538108 361994
rect 535453 361936 535458 361992
rect 535514 361936 538108 361992
rect 535453 361934 538108 361936
rect 535453 361931 535519 361934
rect 536189 360634 536255 360637
rect 536189 360632 538108 360634
rect 536189 360576 536194 360632
rect 536250 360576 538108 360632
rect 536189 360574 538108 360576
rect 536189 360571 536255 360574
rect 536741 359274 536807 359277
rect 536741 359272 538108 359274
rect 536741 359216 536746 359272
rect 536802 359244 538108 359272
rect 536802 359216 538138 359244
rect 536741 359214 538138 359216
rect 536741 359211 536807 359214
rect -960 358308 480 358548
rect 470266 358485 470822 358486
rect 470266 358181 470272 358485
rect 470816 358181 470822 358485
rect 470266 358180 470822 358181
rect 478638 357988 478644 358052
rect 478708 358050 478714 358052
rect 478873 358050 478939 358053
rect 481817 358052 481883 358053
rect 484945 358052 485011 358053
rect 478708 358048 478939 358050
rect 478708 357992 478878 358048
rect 478934 357992 478939 358048
rect 478708 357990 478939 357992
rect 478708 357988 478714 357990
rect 478873 357987 478939 357990
rect 481766 357988 481772 358052
rect 481836 358050 481883 358052
rect 481836 358048 481928 358050
rect 481878 357992 481928 358048
rect 481836 357990 481928 357992
rect 481836 357988 481883 357990
rect 484894 357988 484900 358052
rect 484964 358050 485011 358052
rect 488349 358052 488415 358053
rect 488349 358050 488396 358052
rect 484964 358048 485056 358050
rect 485006 357992 485056 358048
rect 484964 357990 485056 357992
rect 488304 358048 488396 358050
rect 488304 357992 488354 358048
rect 488304 357990 488396 357992
rect 484964 357988 485011 357990
rect 481817 357987 481883 357988
rect 484945 357987 485011 357988
rect 488349 357988 488396 357990
rect 488460 357988 488466 358052
rect 488349 357987 488415 357988
rect 475009 357508 475075 357509
rect 474958 357444 474964 357508
rect 475028 357506 475075 357508
rect 475028 357504 475120 357506
rect 475070 357448 475120 357504
rect 475028 357446 475120 357448
rect 475028 357444 475075 357446
rect 475009 357443 475075 357444
rect 469026 357399 469582 357400
rect 469026 357095 469032 357399
rect 469576 357095 469582 357399
rect 469026 357094 469582 357095
rect 470266 356312 470822 356313
rect 470266 356008 470272 356312
rect 470816 356008 470822 356312
rect 470266 356007 470822 356008
rect 536741 352474 536807 352477
rect 538078 352474 538138 359214
rect 536741 352472 538138 352474
rect 536741 352416 536746 352472
rect 536802 352444 538138 352472
rect 536802 352416 538108 352444
rect 536741 352414 538108 352416
rect 536741 352411 536807 352414
rect 544326 351868 544332 351932
rect 544396 351930 544402 351932
rect 583520 351930 584960 352020
rect 544396 351870 584960 351930
rect 544396 351868 544402 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 473670 343708 473676 343772
rect 473740 343770 473746 343772
rect 474958 343770 474964 343772
rect 473740 343710 474964 343770
rect 473740 343708 473746 343710
rect 474958 343708 474964 343710
rect 475028 343708 475034 343772
rect 470266 342484 470822 342485
rect 470266 342180 470272 342484
rect 470816 342180 470822 342484
rect 470266 342179 470822 342180
rect 469026 341397 469582 341398
rect 469026 341093 469032 341397
rect 469576 341093 469582 341397
rect 469026 341092 469582 341093
rect 477910 341050 477976 341053
rect 478454 341050 478460 341052
rect 477910 341048 478460 341050
rect 477910 340992 477915 341048
rect 477971 340992 478460 341048
rect 477910 340990 478460 340992
rect 477910 340987 477976 340990
rect 478454 340988 478460 340990
rect 478524 340988 478530 341052
rect 481227 341050 481293 341053
rect 481398 341050 481404 341052
rect 481227 341048 481404 341050
rect 481227 340992 481232 341048
rect 481288 340992 481404 341048
rect 481227 340990 481404 340992
rect 481227 340987 481293 340990
rect 481398 340988 481404 340990
rect 481468 340988 481474 341052
rect 484158 340988 484164 341052
rect 484228 341050 484234 341052
rect 484393 341050 484459 341053
rect 484228 341048 484459 341050
rect 484228 340992 484398 341048
rect 484454 340992 484459 341048
rect 484228 340990 484459 340992
rect 484228 340988 484234 340990
rect 484393 340987 484459 340990
rect 487889 341050 487955 341053
rect 488022 341050 488028 341052
rect 487889 341048 488028 341050
rect 487889 340992 487894 341048
rect 487950 340992 488028 341048
rect 487889 340990 488028 340992
rect 487889 340987 487955 340990
rect 488022 340988 488028 340990
rect 488092 340988 488098 341052
rect 473670 340444 473676 340508
rect 473740 340506 473746 340508
rect 474549 340506 474615 340509
rect 473740 340504 474615 340506
rect 473740 340448 474554 340504
rect 474610 340448 474615 340504
rect 473740 340446 474615 340448
rect 473740 340444 473746 340446
rect 474549 340443 474615 340446
rect 470266 340312 470822 340313
rect 470266 340008 470272 340312
rect 470816 340008 470822 340312
rect 470266 340007 470822 340008
rect 541566 339492 541572 339556
rect 541636 339554 541642 339556
rect 541709 339554 541775 339557
rect 541636 339552 541775 339554
rect 541636 339496 541714 339552
rect 541770 339496 541775 339552
rect 541636 339494 541775 339496
rect 541636 339492 541642 339494
rect 541709 339491 541775 339494
rect 544193 339554 544259 339557
rect 544326 339554 544332 339556
rect 544193 339552 544332 339554
rect 544193 339496 544198 339552
rect 544254 339496 544332 339552
rect 544193 339494 544332 339496
rect 544193 339491 544259 339494
rect 544326 339492 544332 339494
rect 544396 339492 544402 339556
rect 583520 338452 584960 338692
rect 535453 336834 535519 336837
rect 535453 336832 538108 336834
rect 535453 336776 535458 336832
rect 535514 336776 538108 336832
rect 535453 336774 538108 336776
rect 535453 336771 535519 336774
rect 486550 335412 486556 335476
rect 486620 335474 486626 335476
rect 486620 335414 538108 335474
rect 486620 335412 486626 335414
rect 485630 334052 485636 334116
rect 485700 334114 485706 334116
rect 485700 334054 538108 334114
rect 485700 334052 485706 334054
rect 486734 332692 486740 332756
rect 486804 332754 486810 332756
rect 486804 332694 538108 332754
rect 486804 332692 486810 332694
rect -960 332196 480 332436
rect 535453 331394 535519 331397
rect 535453 331392 538108 331394
rect 535453 331336 535458 331392
rect 535514 331336 538108 331392
rect 535453 331334 538108 331336
rect 535453 331331 535519 331334
rect 535453 330034 535519 330037
rect 535453 330032 538108 330034
rect 535453 329976 535458 330032
rect 535514 329976 538108 330032
rect 535453 329974 538108 329976
rect 535453 329971 535519 329974
rect 536005 328674 536071 328677
rect 536005 328672 538108 328674
rect 536005 328616 536010 328672
rect 536066 328616 538108 328672
rect 536005 328614 538108 328616
rect 536005 328611 536071 328614
rect 536649 327314 536715 327317
rect 536649 327312 538108 327314
rect 536649 327256 536654 327312
rect 536710 327256 538108 327312
rect 536649 327254 538108 327256
rect 536649 327251 536715 327254
rect 549294 326770 549300 326772
rect 547860 326710 549300 326770
rect 549294 326708 549300 326710
rect 549364 326708 549370 326772
rect 535453 325954 535519 325957
rect 535453 325952 538108 325954
rect 535453 325896 535458 325952
rect 535514 325896 538108 325952
rect 535453 325894 538108 325896
rect 535453 325891 535519 325894
rect 583520 325124 584960 325364
rect 536373 324594 536439 324597
rect 536373 324592 538108 324594
rect 536373 324536 536378 324592
rect 536434 324536 538108 324592
rect 536373 324534 538108 324536
rect 536373 324531 536439 324534
rect 536741 323234 536807 323237
rect 536741 323232 538108 323234
rect 536741 323176 536746 323232
rect 536802 323204 538108 323232
rect 536802 323176 538138 323204
rect 536741 323174 538138 323176
rect 536741 323171 536807 323174
rect 470266 322484 470822 322485
rect 470266 322180 470272 322484
rect 470816 322180 470822 322484
rect 470266 322179 470822 322180
rect 469026 321397 469582 321398
rect 469026 321093 469032 321397
rect 469576 321093 469582 321397
rect 473670 321268 473676 321332
rect 473740 321330 473746 321332
rect 474273 321330 474339 321333
rect 473740 321328 474339 321330
rect 473740 321272 474278 321328
rect 474334 321272 474339 321328
rect 473740 321270 474339 321272
rect 473740 321268 473746 321270
rect 474273 321267 474339 321270
rect 484158 321268 484164 321332
rect 484228 321330 484234 321332
rect 484577 321330 484643 321333
rect 484228 321328 484643 321330
rect 484228 321272 484582 321328
rect 484638 321272 484643 321328
rect 484228 321270 484643 321272
rect 484228 321268 484234 321270
rect 484577 321267 484643 321270
rect 469026 321092 469582 321093
rect 488022 320996 488028 321060
rect 488092 321058 488098 321060
rect 488165 321058 488231 321061
rect 488092 321056 488231 321058
rect 488092 321000 488170 321056
rect 488226 321000 488231 321056
rect 488092 320998 488231 321000
rect 488092 320996 488098 320998
rect 488165 320995 488231 320998
rect 478137 320922 478203 320925
rect 481541 320924 481607 320925
rect 478638 320922 478644 320924
rect 478137 320920 478644 320922
rect 478137 320864 478142 320920
rect 478198 320864 478644 320920
rect 478137 320862 478644 320864
rect 478137 320859 478203 320862
rect 478638 320860 478644 320862
rect 478708 320860 478714 320924
rect 481541 320922 481588 320924
rect 481496 320920 481588 320922
rect 481496 320864 481546 320920
rect 481496 320862 481588 320864
rect 481541 320860 481588 320862
rect 481652 320860 481658 320924
rect 481541 320859 481607 320860
rect 470266 320312 470822 320313
rect 470266 320008 470272 320312
rect 470816 320008 470822 320312
rect 470266 320007 470822 320008
rect -960 319140 480 319380
rect 536741 316434 536807 316437
rect 538078 316434 538138 323174
rect 536741 316432 538138 316434
rect 536741 316376 536746 316432
rect 536802 316404 538138 316432
rect 536802 316376 538108 316404
rect 536741 316374 538108 316376
rect 536741 316371 536807 316374
rect 583520 311932 584960 312172
rect 470266 307084 470822 307085
rect 470266 306780 470272 307084
rect 470816 306780 470822 307084
rect 470266 306779 470822 306780
rect -960 306084 480 306324
rect 487654 306308 487660 306372
rect 487724 306308 487730 306372
rect 487529 306234 487595 306237
rect 487662 306234 487722 306308
rect 487529 306232 487722 306234
rect 487529 306176 487534 306232
rect 487590 306176 487722 306232
rect 487529 306174 487722 306176
rect 487529 306171 487595 306174
rect 480999 306098 481065 306101
rect 481582 306098 481588 306100
rect 480999 306096 481588 306098
rect 480999 306040 481004 306096
rect 481060 306040 481588 306096
rect 480999 306038 481588 306040
rect 480999 306035 481065 306038
rect 481582 306036 481588 306038
rect 481652 306036 481658 306100
rect 469026 305999 469582 306000
rect 469026 305695 469032 305999
rect 469576 305695 469582 305999
rect 473721 305964 473787 305965
rect 473670 305900 473676 305964
rect 473740 305962 473787 305964
rect 473740 305960 473832 305962
rect 473782 305904 473832 305960
rect 473740 305902 473832 305904
rect 473740 305900 473787 305902
rect 473721 305899 473787 305900
rect 469026 305694 469582 305695
rect 477734 305690 477800 305693
rect 478822 305690 478828 305692
rect 477734 305688 478828 305690
rect 477734 305632 477739 305688
rect 477795 305632 478828 305688
rect 477734 305630 478828 305632
rect 477734 305627 477800 305630
rect 478822 305628 478828 305630
rect 478892 305628 478898 305692
rect 484117 305556 484183 305557
rect 484117 305554 484164 305556
rect 484072 305552 484164 305554
rect 484072 305496 484122 305552
rect 484072 305494 484164 305496
rect 484117 305492 484164 305494
rect 484228 305492 484234 305556
rect 484117 305491 484183 305492
rect 470266 304912 470822 304913
rect 470266 304608 470272 304912
rect 470816 304608 470822 304912
rect 470266 304607 470822 304608
rect 544193 303786 544259 303789
rect 544326 303786 544332 303788
rect 544193 303784 544332 303786
rect 544193 303728 544198 303784
rect 544254 303728 544332 303784
rect 544193 303726 544332 303728
rect 544193 303723 544259 303726
rect 544326 303724 544332 303726
rect 544396 303724 544402 303788
rect 541566 303588 541572 303652
rect 541636 303650 541642 303652
rect 541709 303650 541775 303653
rect 547321 303650 547387 303653
rect 541636 303648 547387 303650
rect 541636 303592 541714 303648
rect 541770 303592 547326 303648
rect 547382 303592 547387 303648
rect 541636 303590 547387 303592
rect 541636 303588 541642 303590
rect 541709 303587 541775 303590
rect 547321 303587 547387 303590
rect 535453 300794 535519 300797
rect 535453 300792 538108 300794
rect 535453 300736 535458 300792
rect 535514 300736 538108 300792
rect 535453 300734 538108 300736
rect 535453 300731 535519 300734
rect 547321 300114 547387 300117
rect 580165 300114 580231 300117
rect 547321 300112 580231 300114
rect 547321 300056 547326 300112
rect 547382 300056 580170 300112
rect 580226 300056 580231 300112
rect 547321 300054 580231 300056
rect 547321 300051 547387 300054
rect 580165 300051 580231 300054
rect 535453 299434 535519 299437
rect 535453 299432 538108 299434
rect 535453 299376 535458 299432
rect 535514 299376 538108 299432
rect 535453 299374 538108 299376
rect 535453 299371 535519 299374
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 535453 298074 535519 298077
rect 535453 298072 538108 298074
rect 535453 298016 535458 298072
rect 535514 298016 538108 298072
rect 535453 298014 538108 298016
rect 535453 298011 535519 298014
rect 535453 296714 535519 296717
rect 535453 296712 538108 296714
rect 535453 296656 535458 296712
rect 535514 296656 538108 296712
rect 535453 296654 538108 296656
rect 535453 296651 535519 296654
rect 535545 295354 535611 295357
rect 535545 295352 538108 295354
rect 535545 295296 535550 295352
rect 535606 295296 538108 295352
rect 535545 295294 538108 295296
rect 535545 295291 535611 295294
rect 535453 293994 535519 293997
rect 535453 293992 538108 293994
rect 535453 293936 535458 293992
rect 535514 293936 538108 293992
rect 535453 293934 538108 293936
rect 535453 293931 535519 293934
rect -960 293028 480 293268
rect 535545 292634 535611 292637
rect 535545 292632 538108 292634
rect 535545 292576 535550 292632
rect 535606 292576 538108 292632
rect 535545 292574 538108 292576
rect 535545 292571 535611 292574
rect 535453 291274 535519 291277
rect 535453 291272 538108 291274
rect 535453 291216 535458 291272
rect 535514 291216 538108 291272
rect 535453 291214 538108 291216
rect 535453 291211 535519 291214
rect 549294 290730 549300 290732
rect 547860 290670 549300 290730
rect 549294 290668 549300 290670
rect 549364 290668 549370 290732
rect 535453 289914 535519 289917
rect 535453 289912 538108 289914
rect 535453 289856 535458 289912
rect 535514 289856 538108 289912
rect 535453 289854 538108 289856
rect 535453 289851 535519 289854
rect 473670 289716 473676 289780
rect 473740 289778 473746 289780
rect 476062 289778 476068 289780
rect 473740 289718 476068 289778
rect 473740 289716 473746 289718
rect 476062 289716 476068 289718
rect 476132 289716 476138 289780
rect 484158 289716 484164 289780
rect 484228 289778 484234 289780
rect 485814 289778 485820 289780
rect 484228 289718 485820 289778
rect 484228 289716 484234 289718
rect 485814 289716 485820 289718
rect 485884 289716 485890 289780
rect 535453 288554 535519 288557
rect 535453 288552 538108 288554
rect 535453 288496 535458 288552
rect 535514 288496 538108 288552
rect 535453 288494 538108 288496
rect 535453 288491 535519 288494
rect 470266 287485 470822 287486
rect 470266 287181 470272 287485
rect 470816 287181 470822 287485
rect 470266 287180 470822 287181
rect 536741 287194 536807 287197
rect 536741 287192 538108 287194
rect 536741 287136 536746 287192
rect 536802 287164 538108 287192
rect 536802 287136 538138 287164
rect 536741 287134 538138 287136
rect 536741 287131 536807 287134
rect 478628 286922 478694 286925
rect 478822 286922 478828 286924
rect 478628 286920 478828 286922
rect 478628 286864 478633 286920
rect 478689 286864 478828 286920
rect 478628 286862 478828 286864
rect 478628 286859 478694 286862
rect 478822 286860 478828 286862
rect 478892 286860 478898 286924
rect 488574 286724 488580 286788
rect 488644 286724 488650 286788
rect 488582 286653 488642 286724
rect 474916 286650 474982 286653
rect 476062 286650 476068 286652
rect 474916 286648 476068 286650
rect 474916 286592 474921 286648
rect 474977 286592 476068 286648
rect 474916 286590 476068 286592
rect 474916 286587 474982 286590
rect 476062 286588 476068 286590
rect 476132 286588 476138 286652
rect 488582 286648 488691 286653
rect 488582 286592 488630 286648
rect 488686 286592 488691 286648
rect 488582 286590 488691 286592
rect 488625 286587 488691 286590
rect 469026 286400 469582 286401
rect 469026 286096 469032 286400
rect 469576 286096 469582 286400
rect 469026 286095 469582 286096
rect 482340 285836 482406 285837
rect 485865 285836 485931 285837
rect 482318 285834 482324 285836
rect 482213 285774 482324 285834
rect 482388 285834 482406 285836
rect 482870 285834 482876 285836
rect 482388 285832 482876 285834
rect 482401 285776 482876 285832
rect 482318 285772 482324 285774
rect 482388 285774 482876 285776
rect 482388 285772 482406 285774
rect 482870 285772 482876 285774
rect 482940 285772 482946 285836
rect 485814 285772 485820 285836
rect 485884 285834 485931 285836
rect 485884 285832 485976 285834
rect 485926 285776 485976 285832
rect 485884 285774 485976 285776
rect 485884 285772 485931 285774
rect 482340 285771 482406 285772
rect 485865 285771 485931 285772
rect 470266 285312 470822 285313
rect 470266 285008 470272 285312
rect 470816 285008 470822 285312
rect 470266 285007 470822 285008
rect 536097 280394 536163 280397
rect 538078 280394 538138 287134
rect 583520 285276 584960 285516
rect 536097 280392 538138 280394
rect 536097 280336 536102 280392
rect 536158 280364 538138 280392
rect 536158 280336 538108 280364
rect 536097 280334 538108 280336
rect 536097 280331 536163 280334
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect 470266 267485 470822 267486
rect -960 267052 480 267292
rect 470266 267181 470272 267485
rect 470816 267181 470822 267485
rect 470266 267180 470822 267181
rect 469026 266399 469582 266400
rect 469026 266095 469032 266399
rect 469576 266095 469582 266399
rect 469026 266094 469582 266095
rect 479057 265980 479123 265981
rect 479006 265978 479012 265980
rect 478966 265918 479012 265978
rect 479076 265976 479123 265980
rect 479118 265920 479123 265976
rect 479006 265916 479012 265918
rect 479076 265916 479123 265920
rect 479057 265915 479123 265916
rect 488717 265570 488783 265573
rect 489126 265570 489132 265572
rect 488717 265568 489132 265570
rect 488717 265512 488722 265568
rect 488778 265512 489132 265568
rect 488717 265510 489132 265512
rect 488717 265507 488783 265510
rect 489126 265508 489132 265510
rect 489196 265508 489202 265572
rect 470266 265312 470822 265313
rect 470266 265008 470272 265312
rect 470816 265008 470822 265312
rect 476481 265028 476547 265029
rect 476430 265026 476436 265028
rect 470266 265007 470822 265008
rect 476354 264966 476436 265026
rect 476500 265026 476547 265028
rect 477350 265026 477356 265028
rect 476500 265024 477356 265026
rect 476542 264968 477356 265024
rect 476430 264964 476436 264966
rect 476500 264966 477356 264968
rect 476500 264964 476547 264966
rect 477350 264964 477356 264966
rect 477420 264964 477426 265028
rect 479517 265026 479583 265029
rect 482829 265028 482895 265029
rect 480110 265026 480116 265028
rect 479517 265024 480116 265026
rect 479517 264968 479522 265024
rect 479578 264968 480116 265024
rect 479517 264966 480116 264968
rect 476481 264963 476547 264964
rect 479517 264963 479583 264966
rect 480110 264964 480116 264966
rect 480180 264964 480186 265028
rect 482829 265026 482876 265028
rect 482784 265024 482876 265026
rect 482784 264968 482834 265024
rect 482784 264966 482876 264968
rect 482829 264964 482876 264966
rect 482940 264964 482946 265028
rect 485681 265026 485747 265029
rect 485814 265026 485820 265028
rect 485681 265024 485820 265026
rect 485681 264968 485686 265024
rect 485742 264968 485820 265024
rect 485681 264966 485820 264968
rect 482829 264963 482895 264964
rect 485681 264963 485747 264966
rect 485814 264964 485820 264966
rect 485884 265026 485890 265028
rect 486366 265026 486372 265028
rect 485884 264966 486372 265026
rect 485884 264964 485890 264966
rect 486366 264964 486372 264966
rect 486436 264964 486442 265028
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 538673 245578 538739 245581
rect 583520 245578 584960 245668
rect 538673 245576 584960 245578
rect 538673 245520 538678 245576
rect 538734 245520 584960 245576
rect 538673 245518 584960 245520
rect 538673 245515 538739 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 489126 165820 489132 165884
rect 489196 165882 489202 165884
rect 583520 165882 584960 165972
rect 489196 165822 584960 165882
rect 489196 165820 489202 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 486366 125972 486372 126036
rect 486436 126034 486442 126036
rect 583520 126034 584960 126124
rect 486436 125974 584960 126034
rect 486436 125972 486442 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 482870 86124 482876 86188
rect 482940 86186 482946 86188
rect 583520 86186 584960 86276
rect 482940 86126 584960 86186
rect 482940 86124 482946 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 480110 46276 480116 46340
rect 480180 46338 480186 46340
rect 583520 46338 584960 46428
rect 480180 46278 584960 46338
rect 480180 46276 480186 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 549294 19756 549300 19820
rect 549364 19818 549370 19820
rect 583520 19818 584960 19908
rect 549364 19758 584960 19818
rect 549364 19756 549370 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 477350 6564 477356 6628
rect 477420 6626 477426 6628
rect 583520 6626 584960 6716
rect 477420 6566 584960 6626
rect 477420 6564 477426 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 470272 451479 470816 451483
rect 470272 451183 470276 451479
rect 470276 451183 470812 451479
rect 470812 451183 470816 451479
rect 470272 451179 470816 451183
rect 469032 450393 469576 450397
rect 469032 450097 469036 450393
rect 469036 450097 469572 450393
rect 469572 450097 469576 450393
rect 469032 450093 469576 450097
rect 478460 450196 478524 450260
rect 481220 450196 481284 450260
rect 484164 450196 484228 450260
rect 487844 450256 487908 450260
rect 487844 450200 487849 450256
rect 487849 450200 487908 450256
rect 487844 450196 487908 450200
rect 473676 449652 473740 449716
rect 470272 449308 470816 449312
rect 470272 449012 470276 449308
rect 470276 449012 470812 449308
rect 470812 449012 470816 449308
rect 470272 449008 470816 449012
rect 541572 445028 541636 445092
rect 544332 445028 544396 445092
rect 549300 434692 549364 434756
rect 470272 433080 470816 433084
rect 470272 432784 470276 433080
rect 470276 432784 470812 433080
rect 470812 432784 470816 433080
rect 470272 432780 470816 432784
rect 483612 432304 483676 432308
rect 483612 432248 483626 432304
rect 483626 432248 483676 432304
rect 483612 432244 483676 432248
rect 481220 432168 481284 432172
rect 481220 432112 481270 432168
rect 481270 432112 481284 432168
rect 481220 432108 481284 432112
rect 469032 431993 469576 431997
rect 469032 431697 469036 431993
rect 469036 431697 469572 431993
rect 469572 431697 469576 431993
rect 469032 431693 469576 431697
rect 473676 431836 473740 431900
rect 487660 431836 487724 431900
rect 478460 431564 478524 431628
rect 470272 430908 470816 430912
rect 470272 430612 470276 430908
rect 470276 430612 470812 430908
rect 470812 430612 470816 430908
rect 470272 430608 470816 430612
rect 480116 427892 480180 427956
rect 486556 427892 486620 427956
rect 470272 412080 470816 412084
rect 470272 411784 470276 412080
rect 470276 411784 470812 412080
rect 470812 411784 470816 412080
rect 470272 411780 470816 411784
rect 469032 410994 469576 410998
rect 469032 410698 469036 410994
rect 469036 410698 469572 410994
rect 469572 410698 469576 410994
rect 469032 410694 469576 410698
rect 473676 410952 473740 410956
rect 473676 410896 473726 410952
rect 473726 410896 473740 410952
rect 473676 410892 473740 410896
rect 484164 410408 484228 410412
rect 484164 410352 484178 410408
rect 484178 410352 484228 410408
rect 484164 410348 484228 410352
rect 478460 410136 478524 410140
rect 478460 410080 478474 410136
rect 478474 410080 478524 410136
rect 478460 410076 478524 410080
rect 481404 410136 481468 410140
rect 481404 410080 481418 410136
rect 481418 410080 481468 410136
rect 481404 410076 481468 410080
rect 487844 410136 487908 410140
rect 487844 410080 487858 410136
rect 487858 410080 487908 410136
rect 487844 410076 487908 410080
rect 488396 410076 488460 410140
rect 470272 409908 470816 409912
rect 470272 409612 470276 409908
rect 470276 409612 470812 409908
rect 470812 409612 470816 409908
rect 470272 409608 470816 409612
rect 541572 409260 541636 409324
rect 544332 409320 544396 409324
rect 544332 409264 544346 409320
rect 544346 409264 544396 409320
rect 544332 409260 544396 409264
rect 480116 407492 480180 407556
rect 482876 407084 482940 407148
rect 485636 407084 485700 407148
rect 549300 398244 549364 398308
rect 473676 391988 473740 392052
rect 474964 391988 475028 392052
rect 470272 391081 470816 391085
rect 470272 390785 470276 391081
rect 470276 390785 470812 391081
rect 470812 390785 470816 391081
rect 470272 390781 470816 390785
rect 484900 390233 484964 390297
rect 488396 390084 488460 390148
rect 469032 389998 469576 390002
rect 469032 389702 469036 389998
rect 469036 389702 469572 389998
rect 469572 389702 469576 389998
rect 469032 389698 469576 389702
rect 481772 389404 481836 389468
rect 474964 389328 475028 389332
rect 474964 389272 474978 389328
rect 474978 389272 475028 389328
rect 474964 389268 475028 389272
rect 478644 389328 478708 389332
rect 478644 389272 478690 389328
rect 478690 389272 478708 389328
rect 478644 389268 478708 389272
rect 470272 388908 470816 388912
rect 470272 388612 470276 388908
rect 470276 388612 470812 388908
rect 470812 388612 470816 388908
rect 470272 388608 470816 388612
rect 486740 386412 486804 386476
rect 544516 373416 544580 373420
rect 544516 373360 544530 373416
rect 544530 373360 544580 373416
rect 544516 373356 544580 373360
rect 541572 373084 541636 373148
rect 482876 370092 482940 370156
rect 549300 362748 549364 362812
rect 470272 358481 470816 358485
rect 470272 358185 470276 358481
rect 470276 358185 470812 358481
rect 470812 358185 470816 358481
rect 470272 358181 470816 358185
rect 478644 357988 478708 358052
rect 481772 358048 481836 358052
rect 481772 357992 481822 358048
rect 481822 357992 481836 358048
rect 481772 357988 481836 357992
rect 484900 358048 484964 358052
rect 484900 357992 484950 358048
rect 484950 357992 484964 358048
rect 484900 357988 484964 357992
rect 488396 358048 488460 358052
rect 488396 357992 488410 358048
rect 488410 357992 488460 358048
rect 488396 357988 488460 357992
rect 474964 357504 475028 357508
rect 474964 357448 475014 357504
rect 475014 357448 475028 357504
rect 474964 357444 475028 357448
rect 469032 357395 469576 357399
rect 469032 357099 469036 357395
rect 469036 357099 469572 357395
rect 469572 357099 469576 357395
rect 469032 357095 469576 357099
rect 470272 356308 470816 356312
rect 470272 356012 470276 356308
rect 470276 356012 470812 356308
rect 470812 356012 470816 356308
rect 470272 356008 470816 356012
rect 544332 351868 544396 351932
rect 473676 343708 473740 343772
rect 474964 343708 475028 343772
rect 470272 342480 470816 342484
rect 470272 342184 470276 342480
rect 470276 342184 470812 342480
rect 470812 342184 470816 342480
rect 470272 342180 470816 342184
rect 469032 341393 469576 341397
rect 469032 341097 469036 341393
rect 469036 341097 469572 341393
rect 469572 341097 469576 341393
rect 469032 341093 469576 341097
rect 478460 340988 478524 341052
rect 481404 340988 481468 341052
rect 484164 340988 484228 341052
rect 488028 340988 488092 341052
rect 473676 340444 473740 340508
rect 470272 340308 470816 340312
rect 470272 340012 470276 340308
rect 470276 340012 470812 340308
rect 470812 340012 470816 340308
rect 470272 340008 470816 340012
rect 541572 339492 541636 339556
rect 544332 339492 544396 339556
rect 486556 335412 486620 335476
rect 485636 334052 485700 334116
rect 486740 332692 486804 332756
rect 549300 326708 549364 326772
rect 470272 322480 470816 322484
rect 470272 322184 470276 322480
rect 470276 322184 470812 322480
rect 470812 322184 470816 322480
rect 470272 322180 470816 322184
rect 469032 321393 469576 321397
rect 469032 321097 469036 321393
rect 469036 321097 469572 321393
rect 469572 321097 469576 321393
rect 469032 321093 469576 321097
rect 473676 321268 473740 321332
rect 484164 321268 484228 321332
rect 488028 320996 488092 321060
rect 478644 320860 478708 320924
rect 481588 320920 481652 320924
rect 481588 320864 481602 320920
rect 481602 320864 481652 320920
rect 481588 320860 481652 320864
rect 470272 320308 470816 320312
rect 470272 320012 470276 320308
rect 470276 320012 470812 320308
rect 470812 320012 470816 320308
rect 470272 320008 470816 320012
rect 470272 307080 470816 307084
rect 470272 306784 470276 307080
rect 470276 306784 470812 307080
rect 470812 306784 470816 307080
rect 470272 306780 470816 306784
rect 487660 306308 487724 306372
rect 481588 306036 481652 306100
rect 469032 305995 469576 305999
rect 469032 305699 469036 305995
rect 469036 305699 469572 305995
rect 469572 305699 469576 305995
rect 469032 305695 469576 305699
rect 473676 305960 473740 305964
rect 473676 305904 473726 305960
rect 473726 305904 473740 305960
rect 473676 305900 473740 305904
rect 478828 305628 478892 305692
rect 484164 305552 484228 305556
rect 484164 305496 484178 305552
rect 484178 305496 484228 305552
rect 484164 305492 484228 305496
rect 470272 304908 470816 304912
rect 470272 304612 470276 304908
rect 470276 304612 470812 304908
rect 470812 304612 470816 304908
rect 470272 304608 470816 304612
rect 544332 303724 544396 303788
rect 541572 303588 541636 303652
rect 549300 290668 549364 290732
rect 473676 289716 473740 289780
rect 476068 289716 476132 289780
rect 484164 289716 484228 289780
rect 485820 289716 485884 289780
rect 470272 287481 470816 287485
rect 470272 287185 470276 287481
rect 470276 287185 470812 287481
rect 470812 287185 470816 287481
rect 470272 287181 470816 287185
rect 478828 286860 478892 286924
rect 488580 286724 488644 286788
rect 476068 286588 476132 286652
rect 469032 286396 469576 286400
rect 469032 286100 469036 286396
rect 469036 286100 469572 286396
rect 469572 286100 469576 286396
rect 469032 286096 469576 286100
rect 482324 285832 482388 285836
rect 482324 285776 482345 285832
rect 482345 285776 482388 285832
rect 482324 285772 482388 285776
rect 482876 285772 482940 285836
rect 485820 285832 485884 285836
rect 485820 285776 485870 285832
rect 485870 285776 485884 285832
rect 485820 285772 485884 285776
rect 470272 285308 470816 285312
rect 470272 285012 470276 285308
rect 470276 285012 470812 285308
rect 470812 285012 470816 285308
rect 470272 285008 470816 285012
rect 470272 267481 470816 267485
rect 470272 267185 470276 267481
rect 470276 267185 470812 267481
rect 470812 267185 470816 267481
rect 470272 267181 470816 267185
rect 469032 266395 469576 266399
rect 469032 266099 469036 266395
rect 469036 266099 469572 266395
rect 469572 266099 469576 266395
rect 469032 266095 469576 266099
rect 479012 265976 479076 265980
rect 479012 265920 479062 265976
rect 479062 265920 479076 265976
rect 479012 265916 479076 265920
rect 489132 265508 489196 265572
rect 470272 265308 470816 265312
rect 470272 265012 470276 265308
rect 470276 265012 470812 265308
rect 470812 265012 470816 265308
rect 470272 265008 470816 265012
rect 476436 265024 476500 265028
rect 476436 264968 476486 265024
rect 476486 264968 476500 265024
rect 476436 264964 476500 264968
rect 477356 264964 477420 265028
rect 480116 264964 480180 265028
rect 482876 265024 482940 265028
rect 482876 264968 482890 265024
rect 482890 264968 482940 265024
rect 482876 264964 482940 264968
rect 485820 264964 485884 265028
rect 486372 264964 486436 265028
rect 489132 165820 489196 165884
rect 486372 125972 486436 126036
rect 482876 86124 482940 86188
rect 480116 46276 480180 46340
rect 549300 19756 549364 19820
rect 477356 6564 477420 6628
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 695334 -8106 711002
rect -8726 694778 -8694 695334
rect -8138 694778 -8106 695334
rect -8726 659334 -8106 694778
rect -8726 658778 -8694 659334
rect -8138 658778 -8106 659334
rect -8726 623334 -8106 658778
rect -8726 622778 -8694 623334
rect -8138 622778 -8106 623334
rect -8726 587334 -8106 622778
rect -8726 586778 -8694 587334
rect -8138 586778 -8106 587334
rect -8726 551334 -8106 586778
rect -8726 550778 -8694 551334
rect -8138 550778 -8106 551334
rect -8726 515334 -8106 550778
rect -8726 514778 -8694 515334
rect -8138 514778 -8106 515334
rect -8726 479334 -8106 514778
rect -8726 478778 -8694 479334
rect -8138 478778 -8106 479334
rect -8726 443334 -8106 478778
rect -8726 442778 -8694 443334
rect -8138 442778 -8106 443334
rect -8726 407334 -8106 442778
rect -8726 406778 -8694 407334
rect -8138 406778 -8106 407334
rect -8726 371334 -8106 406778
rect -8726 370778 -8694 371334
rect -8138 370778 -8106 371334
rect -8726 335334 -8106 370778
rect -8726 334778 -8694 335334
rect -8138 334778 -8106 335334
rect -8726 299334 -8106 334778
rect -8726 298778 -8694 299334
rect -8138 298778 -8106 299334
rect -8726 263334 -8106 298778
rect -8726 262778 -8694 263334
rect -8138 262778 -8106 263334
rect -8726 227334 -8106 262778
rect -8726 226778 -8694 227334
rect -8138 226778 -8106 227334
rect -8726 191334 -8106 226778
rect -8726 190778 -8694 191334
rect -8138 190778 -8106 191334
rect -8726 155334 -8106 190778
rect -8726 154778 -8694 155334
rect -8138 154778 -8106 155334
rect -8726 119334 -8106 154778
rect -8726 118778 -8694 119334
rect -8138 118778 -8106 119334
rect -8726 83334 -8106 118778
rect -8726 82778 -8694 83334
rect -8138 82778 -8106 83334
rect -8726 47334 -8106 82778
rect -8726 46778 -8694 47334
rect -8138 46778 -8106 47334
rect -8726 11334 -8106 46778
rect -8726 10778 -8694 11334
rect -8138 10778 -8106 11334
rect -8726 -7066 -8106 10778
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 694094 -7146 710042
rect -7766 693538 -7734 694094
rect -7178 693538 -7146 694094
rect -7766 658094 -7146 693538
rect -7766 657538 -7734 658094
rect -7178 657538 -7146 658094
rect -7766 622094 -7146 657538
rect -7766 621538 -7734 622094
rect -7178 621538 -7146 622094
rect -7766 586094 -7146 621538
rect -7766 585538 -7734 586094
rect -7178 585538 -7146 586094
rect -7766 550094 -7146 585538
rect -7766 549538 -7734 550094
rect -7178 549538 -7146 550094
rect -7766 514094 -7146 549538
rect -7766 513538 -7734 514094
rect -7178 513538 -7146 514094
rect -7766 478094 -7146 513538
rect -7766 477538 -7734 478094
rect -7178 477538 -7146 478094
rect -7766 442094 -7146 477538
rect -7766 441538 -7734 442094
rect -7178 441538 -7146 442094
rect -7766 406094 -7146 441538
rect -7766 405538 -7734 406094
rect -7178 405538 -7146 406094
rect -7766 370094 -7146 405538
rect -7766 369538 -7734 370094
rect -7178 369538 -7146 370094
rect -7766 334094 -7146 369538
rect -7766 333538 -7734 334094
rect -7178 333538 -7146 334094
rect -7766 298094 -7146 333538
rect -7766 297538 -7734 298094
rect -7178 297538 -7146 298094
rect -7766 262094 -7146 297538
rect -7766 261538 -7734 262094
rect -7178 261538 -7146 262094
rect -7766 226094 -7146 261538
rect -7766 225538 -7734 226094
rect -7178 225538 -7146 226094
rect -7766 190094 -7146 225538
rect -7766 189538 -7734 190094
rect -7178 189538 -7146 190094
rect -7766 154094 -7146 189538
rect -7766 153538 -7734 154094
rect -7178 153538 -7146 154094
rect -7766 118094 -7146 153538
rect -7766 117538 -7734 118094
rect -7178 117538 -7146 118094
rect -7766 82094 -7146 117538
rect -7766 81538 -7734 82094
rect -7178 81538 -7146 82094
rect -7766 46094 -7146 81538
rect -7766 45538 -7734 46094
rect -7178 45538 -7146 46094
rect -7766 10094 -7146 45538
rect -7766 9538 -7734 10094
rect -7178 9538 -7146 10094
rect -7766 -6106 -7146 9538
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 692854 -6186 709082
rect -6806 692298 -6774 692854
rect -6218 692298 -6186 692854
rect -6806 656854 -6186 692298
rect -6806 656298 -6774 656854
rect -6218 656298 -6186 656854
rect -6806 620854 -6186 656298
rect -6806 620298 -6774 620854
rect -6218 620298 -6186 620854
rect -6806 584854 -6186 620298
rect -6806 584298 -6774 584854
rect -6218 584298 -6186 584854
rect -6806 548854 -6186 584298
rect -6806 548298 -6774 548854
rect -6218 548298 -6186 548854
rect -6806 512854 -6186 548298
rect -6806 512298 -6774 512854
rect -6218 512298 -6186 512854
rect -6806 476854 -6186 512298
rect -6806 476298 -6774 476854
rect -6218 476298 -6186 476854
rect -6806 440854 -6186 476298
rect -6806 440298 -6774 440854
rect -6218 440298 -6186 440854
rect -6806 404854 -6186 440298
rect -6806 404298 -6774 404854
rect -6218 404298 -6186 404854
rect -6806 368854 -6186 404298
rect -6806 368298 -6774 368854
rect -6218 368298 -6186 368854
rect -6806 332854 -6186 368298
rect -6806 332298 -6774 332854
rect -6218 332298 -6186 332854
rect -6806 296854 -6186 332298
rect -6806 296298 -6774 296854
rect -6218 296298 -6186 296854
rect -6806 260854 -6186 296298
rect -6806 260298 -6774 260854
rect -6218 260298 -6186 260854
rect -6806 224854 -6186 260298
rect -6806 224298 -6774 224854
rect -6218 224298 -6186 224854
rect -6806 188854 -6186 224298
rect -6806 188298 -6774 188854
rect -6218 188298 -6186 188854
rect -6806 152854 -6186 188298
rect -6806 152298 -6774 152854
rect -6218 152298 -6186 152854
rect -6806 116854 -6186 152298
rect -6806 116298 -6774 116854
rect -6218 116298 -6186 116854
rect -6806 80854 -6186 116298
rect -6806 80298 -6774 80854
rect -6218 80298 -6186 80854
rect -6806 44854 -6186 80298
rect -6806 44298 -6774 44854
rect -6218 44298 -6186 44854
rect -6806 8854 -6186 44298
rect -6806 8298 -6774 8854
rect -6218 8298 -6186 8854
rect -6806 -5146 -6186 8298
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 691614 -5226 708122
rect -5846 691058 -5814 691614
rect -5258 691058 -5226 691614
rect -5846 655614 -5226 691058
rect -5846 655058 -5814 655614
rect -5258 655058 -5226 655614
rect -5846 619614 -5226 655058
rect -5846 619058 -5814 619614
rect -5258 619058 -5226 619614
rect -5846 583614 -5226 619058
rect -5846 583058 -5814 583614
rect -5258 583058 -5226 583614
rect -5846 547614 -5226 583058
rect -5846 547058 -5814 547614
rect -5258 547058 -5226 547614
rect -5846 511614 -5226 547058
rect -5846 511058 -5814 511614
rect -5258 511058 -5226 511614
rect -5846 475614 -5226 511058
rect -5846 475058 -5814 475614
rect -5258 475058 -5226 475614
rect -5846 439614 -5226 475058
rect -5846 439058 -5814 439614
rect -5258 439058 -5226 439614
rect -5846 403614 -5226 439058
rect -5846 403058 -5814 403614
rect -5258 403058 -5226 403614
rect -5846 367614 -5226 403058
rect -5846 367058 -5814 367614
rect -5258 367058 -5226 367614
rect -5846 331614 -5226 367058
rect -5846 331058 -5814 331614
rect -5258 331058 -5226 331614
rect -5846 295614 -5226 331058
rect -5846 295058 -5814 295614
rect -5258 295058 -5226 295614
rect -5846 259614 -5226 295058
rect -5846 259058 -5814 259614
rect -5258 259058 -5226 259614
rect -5846 223614 -5226 259058
rect -5846 223058 -5814 223614
rect -5258 223058 -5226 223614
rect -5846 187614 -5226 223058
rect -5846 187058 -5814 187614
rect -5258 187058 -5226 187614
rect -5846 151614 -5226 187058
rect -5846 151058 -5814 151614
rect -5258 151058 -5226 151614
rect -5846 115614 -5226 151058
rect -5846 115058 -5814 115614
rect -5258 115058 -5226 115614
rect -5846 79614 -5226 115058
rect -5846 79058 -5814 79614
rect -5258 79058 -5226 79614
rect -5846 43614 -5226 79058
rect -5846 43058 -5814 43614
rect -5258 43058 -5226 43614
rect -5846 7614 -5226 43058
rect -5846 7058 -5814 7614
rect -5258 7058 -5226 7614
rect -5846 -4186 -5226 7058
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 690374 -4266 707162
rect -4886 689818 -4854 690374
rect -4298 689818 -4266 690374
rect -4886 654374 -4266 689818
rect -4886 653818 -4854 654374
rect -4298 653818 -4266 654374
rect -4886 618374 -4266 653818
rect -4886 617818 -4854 618374
rect -4298 617818 -4266 618374
rect -4886 582374 -4266 617818
rect -4886 581818 -4854 582374
rect -4298 581818 -4266 582374
rect -4886 546374 -4266 581818
rect -4886 545818 -4854 546374
rect -4298 545818 -4266 546374
rect -4886 510374 -4266 545818
rect -4886 509818 -4854 510374
rect -4298 509818 -4266 510374
rect -4886 474374 -4266 509818
rect -4886 473818 -4854 474374
rect -4298 473818 -4266 474374
rect -4886 438374 -4266 473818
rect -4886 437818 -4854 438374
rect -4298 437818 -4266 438374
rect -4886 402374 -4266 437818
rect -4886 401818 -4854 402374
rect -4298 401818 -4266 402374
rect -4886 366374 -4266 401818
rect -4886 365818 -4854 366374
rect -4298 365818 -4266 366374
rect -4886 330374 -4266 365818
rect -4886 329818 -4854 330374
rect -4298 329818 -4266 330374
rect -4886 294374 -4266 329818
rect -4886 293818 -4854 294374
rect -4298 293818 -4266 294374
rect -4886 258374 -4266 293818
rect -4886 257818 -4854 258374
rect -4298 257818 -4266 258374
rect -4886 222374 -4266 257818
rect -4886 221818 -4854 222374
rect -4298 221818 -4266 222374
rect -4886 186374 -4266 221818
rect -4886 185818 -4854 186374
rect -4298 185818 -4266 186374
rect -4886 150374 -4266 185818
rect -4886 149818 -4854 150374
rect -4298 149818 -4266 150374
rect -4886 114374 -4266 149818
rect -4886 113818 -4854 114374
rect -4298 113818 -4266 114374
rect -4886 78374 -4266 113818
rect -4886 77818 -4854 78374
rect -4298 77818 -4266 78374
rect -4886 42374 -4266 77818
rect -4886 41818 -4854 42374
rect -4298 41818 -4266 42374
rect -4886 6374 -4266 41818
rect -4886 5818 -4854 6374
rect -4298 5818 -4266 6374
rect -4886 -3226 -4266 5818
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 689134 -3306 706202
rect -3926 688578 -3894 689134
rect -3338 688578 -3306 689134
rect -3926 653134 -3306 688578
rect -3926 652578 -3894 653134
rect -3338 652578 -3306 653134
rect -3926 617134 -3306 652578
rect -3926 616578 -3894 617134
rect -3338 616578 -3306 617134
rect -3926 581134 -3306 616578
rect -3926 580578 -3894 581134
rect -3338 580578 -3306 581134
rect -3926 545134 -3306 580578
rect -3926 544578 -3894 545134
rect -3338 544578 -3306 545134
rect -3926 509134 -3306 544578
rect -3926 508578 -3894 509134
rect -3338 508578 -3306 509134
rect -3926 473134 -3306 508578
rect -3926 472578 -3894 473134
rect -3338 472578 -3306 473134
rect -3926 437134 -3306 472578
rect -3926 436578 -3894 437134
rect -3338 436578 -3306 437134
rect -3926 401134 -3306 436578
rect -3926 400578 -3894 401134
rect -3338 400578 -3306 401134
rect -3926 365134 -3306 400578
rect -3926 364578 -3894 365134
rect -3338 364578 -3306 365134
rect -3926 329134 -3306 364578
rect -3926 328578 -3894 329134
rect -3338 328578 -3306 329134
rect -3926 293134 -3306 328578
rect -3926 292578 -3894 293134
rect -3338 292578 -3306 293134
rect -3926 257134 -3306 292578
rect -3926 256578 -3894 257134
rect -3338 256578 -3306 257134
rect -3926 221134 -3306 256578
rect -3926 220578 -3894 221134
rect -3338 220578 -3306 221134
rect -3926 185134 -3306 220578
rect -3926 184578 -3894 185134
rect -3338 184578 -3306 185134
rect -3926 149134 -3306 184578
rect -3926 148578 -3894 149134
rect -3338 148578 -3306 149134
rect -3926 113134 -3306 148578
rect -3926 112578 -3894 113134
rect -3338 112578 -3306 113134
rect -3926 77134 -3306 112578
rect -3926 76578 -3894 77134
rect -3338 76578 -3306 77134
rect -3926 41134 -3306 76578
rect -3926 40578 -3894 41134
rect -3338 40578 -3306 41134
rect -3926 5134 -3306 40578
rect -3926 4578 -3894 5134
rect -3338 4578 -3306 5134
rect -3926 -2266 -3306 4578
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 687894 -2346 705242
rect -2966 687338 -2934 687894
rect -2378 687338 -2346 687894
rect -2966 651894 -2346 687338
rect -2966 651338 -2934 651894
rect -2378 651338 -2346 651894
rect -2966 615894 -2346 651338
rect -2966 615338 -2934 615894
rect -2378 615338 -2346 615894
rect -2966 579894 -2346 615338
rect -2966 579338 -2934 579894
rect -2378 579338 -2346 579894
rect -2966 543894 -2346 579338
rect -2966 543338 -2934 543894
rect -2378 543338 -2346 543894
rect -2966 507894 -2346 543338
rect -2966 507338 -2934 507894
rect -2378 507338 -2346 507894
rect -2966 471894 -2346 507338
rect -2966 471338 -2934 471894
rect -2378 471338 -2346 471894
rect -2966 435894 -2346 471338
rect -2966 435338 -2934 435894
rect -2378 435338 -2346 435894
rect -2966 399894 -2346 435338
rect -2966 399338 -2934 399894
rect -2378 399338 -2346 399894
rect -2966 363894 -2346 399338
rect -2966 363338 -2934 363894
rect -2378 363338 -2346 363894
rect -2966 327894 -2346 363338
rect -2966 327338 -2934 327894
rect -2378 327338 -2346 327894
rect -2966 291894 -2346 327338
rect -2966 291338 -2934 291894
rect -2378 291338 -2346 291894
rect -2966 255894 -2346 291338
rect -2966 255338 -2934 255894
rect -2378 255338 -2346 255894
rect -2966 219894 -2346 255338
rect -2966 219338 -2934 219894
rect -2378 219338 -2346 219894
rect -2966 183894 -2346 219338
rect -2966 183338 -2934 183894
rect -2378 183338 -2346 183894
rect -2966 147894 -2346 183338
rect -2966 147338 -2934 147894
rect -2378 147338 -2346 147894
rect -2966 111894 -2346 147338
rect -2966 111338 -2934 111894
rect -2378 111338 -2346 111894
rect -2966 75894 -2346 111338
rect -2966 75338 -2934 75894
rect -2378 75338 -2346 75894
rect -2966 39894 -2346 75338
rect -2966 39338 -2934 39894
rect -2378 39338 -2346 39894
rect -2966 3894 -2346 39338
rect -2966 3338 -2934 3894
rect -2378 3338 -2346 3894
rect -2966 -1306 -2346 3338
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 686654 -1386 704282
rect -2006 686098 -1974 686654
rect -1418 686098 -1386 686654
rect -2006 650654 -1386 686098
rect -2006 650098 -1974 650654
rect -1418 650098 -1386 650654
rect -2006 614654 -1386 650098
rect -2006 614098 -1974 614654
rect -1418 614098 -1386 614654
rect -2006 578654 -1386 614098
rect -2006 578098 -1974 578654
rect -1418 578098 -1386 578654
rect -2006 542654 -1386 578098
rect -2006 542098 -1974 542654
rect -1418 542098 -1386 542654
rect -2006 506654 -1386 542098
rect -2006 506098 -1974 506654
rect -1418 506098 -1386 506654
rect -2006 470654 -1386 506098
rect -2006 470098 -1974 470654
rect -1418 470098 -1386 470654
rect -2006 434654 -1386 470098
rect -2006 434098 -1974 434654
rect -1418 434098 -1386 434654
rect -2006 398654 -1386 434098
rect -2006 398098 -1974 398654
rect -1418 398098 -1386 398654
rect -2006 362654 -1386 398098
rect -2006 362098 -1974 362654
rect -1418 362098 -1386 362654
rect -2006 326654 -1386 362098
rect -2006 326098 -1974 326654
rect -1418 326098 -1386 326654
rect -2006 290654 -1386 326098
rect -2006 290098 -1974 290654
rect -1418 290098 -1386 290654
rect -2006 254654 -1386 290098
rect -2006 254098 -1974 254654
rect -1418 254098 -1386 254654
rect -2006 218654 -1386 254098
rect -2006 218098 -1974 218654
rect -1418 218098 -1386 218654
rect -2006 182654 -1386 218098
rect -2006 182098 -1974 182654
rect -1418 182098 -1386 182654
rect -2006 146654 -1386 182098
rect -2006 146098 -1974 146654
rect -1418 146098 -1386 146654
rect -2006 110654 -1386 146098
rect -2006 110098 -1974 110654
rect -1418 110098 -1386 110654
rect -2006 74654 -1386 110098
rect -2006 74098 -1974 74654
rect -1418 74098 -1386 74654
rect -2006 38654 -1386 74098
rect -2006 38098 -1974 38654
rect -1418 38098 -1386 38654
rect -2006 2654 -1386 38098
rect -2006 2098 -1974 2654
rect -1418 2098 -1386 2654
rect -2006 -346 -1386 2098
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 994 704838 1614 711590
rect 994 704282 1026 704838
rect 1582 704282 1614 704838
rect 994 686654 1614 704282
rect 994 686098 1026 686654
rect 1582 686098 1614 686654
rect 994 650654 1614 686098
rect 994 650098 1026 650654
rect 1582 650098 1614 650654
rect 994 614654 1614 650098
rect 994 614098 1026 614654
rect 1582 614098 1614 614654
rect 994 578654 1614 614098
rect 994 578098 1026 578654
rect 1582 578098 1614 578654
rect 994 542654 1614 578098
rect 994 542098 1026 542654
rect 1582 542098 1614 542654
rect 994 506654 1614 542098
rect 994 506098 1026 506654
rect 1582 506098 1614 506654
rect 994 470654 1614 506098
rect 994 470098 1026 470654
rect 1582 470098 1614 470654
rect 994 434654 1614 470098
rect 994 434098 1026 434654
rect 1582 434098 1614 434654
rect 994 398654 1614 434098
rect 994 398098 1026 398654
rect 1582 398098 1614 398654
rect 994 362654 1614 398098
rect 994 362098 1026 362654
rect 1582 362098 1614 362654
rect 994 326654 1614 362098
rect 994 326098 1026 326654
rect 1582 326098 1614 326654
rect 994 290654 1614 326098
rect 994 290098 1026 290654
rect 1582 290098 1614 290654
rect 994 254654 1614 290098
rect 994 254098 1026 254654
rect 1582 254098 1614 254654
rect 994 218654 1614 254098
rect 994 218098 1026 218654
rect 1582 218098 1614 218654
rect 994 182654 1614 218098
rect 994 182098 1026 182654
rect 1582 182098 1614 182654
rect 994 146654 1614 182098
rect 994 146098 1026 146654
rect 1582 146098 1614 146654
rect 994 110654 1614 146098
rect 994 110098 1026 110654
rect 1582 110098 1614 110654
rect 994 74654 1614 110098
rect 994 74098 1026 74654
rect 1582 74098 1614 74654
rect 994 38654 1614 74098
rect 994 38098 1026 38654
rect 1582 38098 1614 38654
rect 994 2654 1614 38098
rect 994 2098 1026 2654
rect 1582 2098 1614 2654
rect 994 -346 1614 2098
rect 994 -902 1026 -346
rect 1582 -902 1614 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 994 -7654 1614 -902
rect 2234 705798 2854 711590
rect 2234 705242 2266 705798
rect 2822 705242 2854 705798
rect 2234 687894 2854 705242
rect 2234 687338 2266 687894
rect 2822 687338 2854 687894
rect 2234 651894 2854 687338
rect 2234 651338 2266 651894
rect 2822 651338 2854 651894
rect 2234 615894 2854 651338
rect 2234 615338 2266 615894
rect 2822 615338 2854 615894
rect 2234 579894 2854 615338
rect 2234 579338 2266 579894
rect 2822 579338 2854 579894
rect 2234 543894 2854 579338
rect 2234 543338 2266 543894
rect 2822 543338 2854 543894
rect 2234 507894 2854 543338
rect 2234 507338 2266 507894
rect 2822 507338 2854 507894
rect 2234 471894 2854 507338
rect 2234 471338 2266 471894
rect 2822 471338 2854 471894
rect 2234 435894 2854 471338
rect 2234 435338 2266 435894
rect 2822 435338 2854 435894
rect 2234 399894 2854 435338
rect 2234 399338 2266 399894
rect 2822 399338 2854 399894
rect 2234 363894 2854 399338
rect 2234 363338 2266 363894
rect 2822 363338 2854 363894
rect 2234 327894 2854 363338
rect 2234 327338 2266 327894
rect 2822 327338 2854 327894
rect 2234 291894 2854 327338
rect 2234 291338 2266 291894
rect 2822 291338 2854 291894
rect 2234 255894 2854 291338
rect 2234 255338 2266 255894
rect 2822 255338 2854 255894
rect 2234 219894 2854 255338
rect 2234 219338 2266 219894
rect 2822 219338 2854 219894
rect 2234 183894 2854 219338
rect 2234 183338 2266 183894
rect 2822 183338 2854 183894
rect 2234 147894 2854 183338
rect 2234 147338 2266 147894
rect 2822 147338 2854 147894
rect 2234 111894 2854 147338
rect 2234 111338 2266 111894
rect 2822 111338 2854 111894
rect 2234 75894 2854 111338
rect 2234 75338 2266 75894
rect 2822 75338 2854 75894
rect 2234 39894 2854 75338
rect 2234 39338 2266 39894
rect 2822 39338 2854 39894
rect 2234 3894 2854 39338
rect 2234 3338 2266 3894
rect 2822 3338 2854 3894
rect 2234 -1306 2854 3338
rect 2234 -1862 2266 -1306
rect 2822 -1862 2854 -1306
rect 2234 -7654 2854 -1862
rect 3474 706758 4094 711590
rect 3474 706202 3506 706758
rect 4062 706202 4094 706758
rect 3474 689134 4094 706202
rect 3474 688578 3506 689134
rect 4062 688578 4094 689134
rect 3474 653134 4094 688578
rect 3474 652578 3506 653134
rect 4062 652578 4094 653134
rect 3474 617134 4094 652578
rect 3474 616578 3506 617134
rect 4062 616578 4094 617134
rect 3474 581134 4094 616578
rect 3474 580578 3506 581134
rect 4062 580578 4094 581134
rect 3474 545134 4094 580578
rect 3474 544578 3506 545134
rect 4062 544578 4094 545134
rect 3474 509134 4094 544578
rect 3474 508578 3506 509134
rect 4062 508578 4094 509134
rect 3474 473134 4094 508578
rect 3474 472578 3506 473134
rect 4062 472578 4094 473134
rect 3474 437134 4094 472578
rect 3474 436578 3506 437134
rect 4062 436578 4094 437134
rect 3474 401134 4094 436578
rect 3474 400578 3506 401134
rect 4062 400578 4094 401134
rect 3474 365134 4094 400578
rect 3474 364578 3506 365134
rect 4062 364578 4094 365134
rect 3474 329134 4094 364578
rect 3474 328578 3506 329134
rect 4062 328578 4094 329134
rect 3474 293134 4094 328578
rect 3474 292578 3506 293134
rect 4062 292578 4094 293134
rect 3474 257134 4094 292578
rect 3474 256578 3506 257134
rect 4062 256578 4094 257134
rect 3474 221134 4094 256578
rect 3474 220578 3506 221134
rect 4062 220578 4094 221134
rect 3474 185134 4094 220578
rect 3474 184578 3506 185134
rect 4062 184578 4094 185134
rect 3474 149134 4094 184578
rect 3474 148578 3506 149134
rect 4062 148578 4094 149134
rect 3474 113134 4094 148578
rect 3474 112578 3506 113134
rect 4062 112578 4094 113134
rect 3474 77134 4094 112578
rect 3474 76578 3506 77134
rect 4062 76578 4094 77134
rect 3474 41134 4094 76578
rect 3474 40578 3506 41134
rect 4062 40578 4094 41134
rect 3474 5134 4094 40578
rect 3474 4578 3506 5134
rect 4062 4578 4094 5134
rect 3474 -2266 4094 4578
rect 3474 -2822 3506 -2266
rect 4062 -2822 4094 -2266
rect 3474 -7654 4094 -2822
rect 4714 707718 5334 711590
rect 4714 707162 4746 707718
rect 5302 707162 5334 707718
rect 4714 690374 5334 707162
rect 4714 689818 4746 690374
rect 5302 689818 5334 690374
rect 4714 654374 5334 689818
rect 4714 653818 4746 654374
rect 5302 653818 5334 654374
rect 4714 618374 5334 653818
rect 4714 617818 4746 618374
rect 5302 617818 5334 618374
rect 4714 582374 5334 617818
rect 4714 581818 4746 582374
rect 5302 581818 5334 582374
rect 4714 546374 5334 581818
rect 4714 545818 4746 546374
rect 5302 545818 5334 546374
rect 4714 510374 5334 545818
rect 4714 509818 4746 510374
rect 5302 509818 5334 510374
rect 4714 474374 5334 509818
rect 4714 473818 4746 474374
rect 5302 473818 5334 474374
rect 4714 438374 5334 473818
rect 4714 437818 4746 438374
rect 5302 437818 5334 438374
rect 4714 402374 5334 437818
rect 4714 401818 4746 402374
rect 5302 401818 5334 402374
rect 4714 366374 5334 401818
rect 4714 365818 4746 366374
rect 5302 365818 5334 366374
rect 4714 330374 5334 365818
rect 4714 329818 4746 330374
rect 5302 329818 5334 330374
rect 4714 294374 5334 329818
rect 4714 293818 4746 294374
rect 5302 293818 5334 294374
rect 4714 258374 5334 293818
rect 4714 257818 4746 258374
rect 5302 257818 5334 258374
rect 4714 222374 5334 257818
rect 4714 221818 4746 222374
rect 5302 221818 5334 222374
rect 4714 186374 5334 221818
rect 4714 185818 4746 186374
rect 5302 185818 5334 186374
rect 4714 150374 5334 185818
rect 4714 149818 4746 150374
rect 5302 149818 5334 150374
rect 4714 114374 5334 149818
rect 4714 113818 4746 114374
rect 5302 113818 5334 114374
rect 4714 78374 5334 113818
rect 4714 77818 4746 78374
rect 5302 77818 5334 78374
rect 4714 42374 5334 77818
rect 4714 41818 4746 42374
rect 5302 41818 5334 42374
rect 4714 6374 5334 41818
rect 4714 5818 4746 6374
rect 5302 5818 5334 6374
rect 4714 -3226 5334 5818
rect 4714 -3782 4746 -3226
rect 5302 -3782 5334 -3226
rect 4714 -7654 5334 -3782
rect 5954 708678 6574 711590
rect 5954 708122 5986 708678
rect 6542 708122 6574 708678
rect 5954 691614 6574 708122
rect 5954 691058 5986 691614
rect 6542 691058 6574 691614
rect 5954 655614 6574 691058
rect 5954 655058 5986 655614
rect 6542 655058 6574 655614
rect 5954 619614 6574 655058
rect 5954 619058 5986 619614
rect 6542 619058 6574 619614
rect 5954 583614 6574 619058
rect 5954 583058 5986 583614
rect 6542 583058 6574 583614
rect 5954 547614 6574 583058
rect 5954 547058 5986 547614
rect 6542 547058 6574 547614
rect 5954 511614 6574 547058
rect 5954 511058 5986 511614
rect 6542 511058 6574 511614
rect 5954 475614 6574 511058
rect 5954 475058 5986 475614
rect 6542 475058 6574 475614
rect 5954 439614 6574 475058
rect 5954 439058 5986 439614
rect 6542 439058 6574 439614
rect 5954 403614 6574 439058
rect 5954 403058 5986 403614
rect 6542 403058 6574 403614
rect 5954 367614 6574 403058
rect 5954 367058 5986 367614
rect 6542 367058 6574 367614
rect 5954 331614 6574 367058
rect 5954 331058 5986 331614
rect 6542 331058 6574 331614
rect 5954 295614 6574 331058
rect 5954 295058 5986 295614
rect 6542 295058 6574 295614
rect 5954 259614 6574 295058
rect 5954 259058 5986 259614
rect 6542 259058 6574 259614
rect 5954 223614 6574 259058
rect 5954 223058 5986 223614
rect 6542 223058 6574 223614
rect 5954 187614 6574 223058
rect 5954 187058 5986 187614
rect 6542 187058 6574 187614
rect 5954 151614 6574 187058
rect 5954 151058 5986 151614
rect 6542 151058 6574 151614
rect 5954 115614 6574 151058
rect 5954 115058 5986 115614
rect 6542 115058 6574 115614
rect 5954 79614 6574 115058
rect 5954 79058 5986 79614
rect 6542 79058 6574 79614
rect 5954 43614 6574 79058
rect 5954 43058 5986 43614
rect 6542 43058 6574 43614
rect 5954 7614 6574 43058
rect 5954 7058 5986 7614
rect 6542 7058 6574 7614
rect 5954 -4186 6574 7058
rect 5954 -4742 5986 -4186
rect 6542 -4742 6574 -4186
rect 5954 -7654 6574 -4742
rect 7194 709638 7814 711590
rect 7194 709082 7226 709638
rect 7782 709082 7814 709638
rect 7194 692854 7814 709082
rect 7194 692298 7226 692854
rect 7782 692298 7814 692854
rect 7194 656854 7814 692298
rect 7194 656298 7226 656854
rect 7782 656298 7814 656854
rect 7194 620854 7814 656298
rect 7194 620298 7226 620854
rect 7782 620298 7814 620854
rect 7194 584854 7814 620298
rect 7194 584298 7226 584854
rect 7782 584298 7814 584854
rect 7194 548854 7814 584298
rect 7194 548298 7226 548854
rect 7782 548298 7814 548854
rect 7194 512854 7814 548298
rect 7194 512298 7226 512854
rect 7782 512298 7814 512854
rect 7194 476854 7814 512298
rect 7194 476298 7226 476854
rect 7782 476298 7814 476854
rect 7194 440854 7814 476298
rect 7194 440298 7226 440854
rect 7782 440298 7814 440854
rect 7194 404854 7814 440298
rect 7194 404298 7226 404854
rect 7782 404298 7814 404854
rect 7194 368854 7814 404298
rect 7194 368298 7226 368854
rect 7782 368298 7814 368854
rect 7194 332854 7814 368298
rect 7194 332298 7226 332854
rect 7782 332298 7814 332854
rect 7194 296854 7814 332298
rect 7194 296298 7226 296854
rect 7782 296298 7814 296854
rect 7194 260854 7814 296298
rect 7194 260298 7226 260854
rect 7782 260298 7814 260854
rect 7194 224854 7814 260298
rect 7194 224298 7226 224854
rect 7782 224298 7814 224854
rect 7194 188854 7814 224298
rect 7194 188298 7226 188854
rect 7782 188298 7814 188854
rect 7194 152854 7814 188298
rect 7194 152298 7226 152854
rect 7782 152298 7814 152854
rect 7194 116854 7814 152298
rect 7194 116298 7226 116854
rect 7782 116298 7814 116854
rect 7194 80854 7814 116298
rect 7194 80298 7226 80854
rect 7782 80298 7814 80854
rect 7194 44854 7814 80298
rect 7194 44298 7226 44854
rect 7782 44298 7814 44854
rect 7194 8854 7814 44298
rect 7194 8298 7226 8854
rect 7782 8298 7814 8854
rect 7194 -5146 7814 8298
rect 7194 -5702 7226 -5146
rect 7782 -5702 7814 -5146
rect 7194 -7654 7814 -5702
rect 8434 710598 9054 711590
rect 8434 710042 8466 710598
rect 9022 710042 9054 710598
rect 8434 694094 9054 710042
rect 8434 693538 8466 694094
rect 9022 693538 9054 694094
rect 8434 658094 9054 693538
rect 8434 657538 8466 658094
rect 9022 657538 9054 658094
rect 8434 622094 9054 657538
rect 8434 621538 8466 622094
rect 9022 621538 9054 622094
rect 8434 586094 9054 621538
rect 8434 585538 8466 586094
rect 9022 585538 9054 586094
rect 8434 550094 9054 585538
rect 8434 549538 8466 550094
rect 9022 549538 9054 550094
rect 8434 514094 9054 549538
rect 8434 513538 8466 514094
rect 9022 513538 9054 514094
rect 8434 478094 9054 513538
rect 8434 477538 8466 478094
rect 9022 477538 9054 478094
rect 8434 442094 9054 477538
rect 8434 441538 8466 442094
rect 9022 441538 9054 442094
rect 8434 406094 9054 441538
rect 8434 405538 8466 406094
rect 9022 405538 9054 406094
rect 8434 370094 9054 405538
rect 8434 369538 8466 370094
rect 9022 369538 9054 370094
rect 8434 334094 9054 369538
rect 8434 333538 8466 334094
rect 9022 333538 9054 334094
rect 8434 298094 9054 333538
rect 8434 297538 8466 298094
rect 9022 297538 9054 298094
rect 8434 262094 9054 297538
rect 8434 261538 8466 262094
rect 9022 261538 9054 262094
rect 8434 226094 9054 261538
rect 8434 225538 8466 226094
rect 9022 225538 9054 226094
rect 8434 190094 9054 225538
rect 8434 189538 8466 190094
rect 9022 189538 9054 190094
rect 8434 154094 9054 189538
rect 8434 153538 8466 154094
rect 9022 153538 9054 154094
rect 8434 118094 9054 153538
rect 8434 117538 8466 118094
rect 9022 117538 9054 118094
rect 8434 82094 9054 117538
rect 8434 81538 8466 82094
rect 9022 81538 9054 82094
rect 8434 46094 9054 81538
rect 8434 45538 8466 46094
rect 9022 45538 9054 46094
rect 8434 10094 9054 45538
rect 8434 9538 8466 10094
rect 9022 9538 9054 10094
rect 8434 -6106 9054 9538
rect 8434 -6662 8466 -6106
rect 9022 -6662 9054 -6106
rect 8434 -7654 9054 -6662
rect 9674 711558 10294 711590
rect 9674 711002 9706 711558
rect 10262 711002 10294 711558
rect 9674 695334 10294 711002
rect 9674 694778 9706 695334
rect 10262 694778 10294 695334
rect 9674 659334 10294 694778
rect 9674 658778 9706 659334
rect 10262 658778 10294 659334
rect 9674 623334 10294 658778
rect 9674 622778 9706 623334
rect 10262 622778 10294 623334
rect 9674 587334 10294 622778
rect 9674 586778 9706 587334
rect 10262 586778 10294 587334
rect 9674 551334 10294 586778
rect 9674 550778 9706 551334
rect 10262 550778 10294 551334
rect 9674 515334 10294 550778
rect 9674 514778 9706 515334
rect 10262 514778 10294 515334
rect 9674 479334 10294 514778
rect 9674 478778 9706 479334
rect 10262 478778 10294 479334
rect 9674 443334 10294 478778
rect 9674 442778 9706 443334
rect 10262 442778 10294 443334
rect 9674 407334 10294 442778
rect 9674 406778 9706 407334
rect 10262 406778 10294 407334
rect 9674 371334 10294 406778
rect 9674 370778 9706 371334
rect 10262 370778 10294 371334
rect 9674 335334 10294 370778
rect 9674 334778 9706 335334
rect 10262 334778 10294 335334
rect 9674 299334 10294 334778
rect 9674 298778 9706 299334
rect 10262 298778 10294 299334
rect 9674 263334 10294 298778
rect 9674 262778 9706 263334
rect 10262 262778 10294 263334
rect 9674 227334 10294 262778
rect 9674 226778 9706 227334
rect 10262 226778 10294 227334
rect 9674 191334 10294 226778
rect 9674 190778 9706 191334
rect 10262 190778 10294 191334
rect 9674 155334 10294 190778
rect 9674 154778 9706 155334
rect 10262 154778 10294 155334
rect 9674 119334 10294 154778
rect 9674 118778 9706 119334
rect 10262 118778 10294 119334
rect 9674 83334 10294 118778
rect 9674 82778 9706 83334
rect 10262 82778 10294 83334
rect 9674 47334 10294 82778
rect 9674 46778 9706 47334
rect 10262 46778 10294 47334
rect 9674 11334 10294 46778
rect 9674 10778 9706 11334
rect 10262 10778 10294 11334
rect 9674 -7066 10294 10778
rect 9674 -7622 9706 -7066
rect 10262 -7622 10294 -7066
rect 9674 -7654 10294 -7622
rect 36994 704838 37614 711590
rect 36994 704282 37026 704838
rect 37582 704282 37614 704838
rect 36994 686654 37614 704282
rect 36994 686098 37026 686654
rect 37582 686098 37614 686654
rect 36994 650654 37614 686098
rect 36994 650098 37026 650654
rect 37582 650098 37614 650654
rect 36994 614654 37614 650098
rect 36994 614098 37026 614654
rect 37582 614098 37614 614654
rect 36994 578654 37614 614098
rect 36994 578098 37026 578654
rect 37582 578098 37614 578654
rect 36994 542654 37614 578098
rect 36994 542098 37026 542654
rect 37582 542098 37614 542654
rect 36994 506654 37614 542098
rect 36994 506098 37026 506654
rect 37582 506098 37614 506654
rect 36994 470654 37614 506098
rect 36994 470098 37026 470654
rect 37582 470098 37614 470654
rect 36994 434654 37614 470098
rect 36994 434098 37026 434654
rect 37582 434098 37614 434654
rect 36994 398654 37614 434098
rect 36994 398098 37026 398654
rect 37582 398098 37614 398654
rect 36994 362654 37614 398098
rect 36994 362098 37026 362654
rect 37582 362098 37614 362654
rect 36994 326654 37614 362098
rect 36994 326098 37026 326654
rect 37582 326098 37614 326654
rect 36994 290654 37614 326098
rect 36994 290098 37026 290654
rect 37582 290098 37614 290654
rect 36994 254654 37614 290098
rect 36994 254098 37026 254654
rect 37582 254098 37614 254654
rect 36994 218654 37614 254098
rect 36994 218098 37026 218654
rect 37582 218098 37614 218654
rect 36994 182654 37614 218098
rect 36994 182098 37026 182654
rect 37582 182098 37614 182654
rect 36994 146654 37614 182098
rect 36994 146098 37026 146654
rect 37582 146098 37614 146654
rect 36994 110654 37614 146098
rect 36994 110098 37026 110654
rect 37582 110098 37614 110654
rect 36994 74654 37614 110098
rect 36994 74098 37026 74654
rect 37582 74098 37614 74654
rect 36994 38654 37614 74098
rect 36994 38098 37026 38654
rect 37582 38098 37614 38654
rect 36994 2654 37614 38098
rect 36994 2098 37026 2654
rect 37582 2098 37614 2654
rect 36994 -346 37614 2098
rect 36994 -902 37026 -346
rect 37582 -902 37614 -346
rect 36994 -7654 37614 -902
rect 38234 705798 38854 711590
rect 38234 705242 38266 705798
rect 38822 705242 38854 705798
rect 38234 687894 38854 705242
rect 38234 687338 38266 687894
rect 38822 687338 38854 687894
rect 38234 651894 38854 687338
rect 38234 651338 38266 651894
rect 38822 651338 38854 651894
rect 38234 615894 38854 651338
rect 38234 615338 38266 615894
rect 38822 615338 38854 615894
rect 38234 579894 38854 615338
rect 38234 579338 38266 579894
rect 38822 579338 38854 579894
rect 38234 543894 38854 579338
rect 38234 543338 38266 543894
rect 38822 543338 38854 543894
rect 38234 507894 38854 543338
rect 38234 507338 38266 507894
rect 38822 507338 38854 507894
rect 38234 471894 38854 507338
rect 38234 471338 38266 471894
rect 38822 471338 38854 471894
rect 38234 435894 38854 471338
rect 38234 435338 38266 435894
rect 38822 435338 38854 435894
rect 38234 399894 38854 435338
rect 38234 399338 38266 399894
rect 38822 399338 38854 399894
rect 38234 363894 38854 399338
rect 38234 363338 38266 363894
rect 38822 363338 38854 363894
rect 38234 327894 38854 363338
rect 38234 327338 38266 327894
rect 38822 327338 38854 327894
rect 38234 291894 38854 327338
rect 38234 291338 38266 291894
rect 38822 291338 38854 291894
rect 38234 255894 38854 291338
rect 38234 255338 38266 255894
rect 38822 255338 38854 255894
rect 38234 219894 38854 255338
rect 38234 219338 38266 219894
rect 38822 219338 38854 219894
rect 38234 183894 38854 219338
rect 38234 183338 38266 183894
rect 38822 183338 38854 183894
rect 38234 147894 38854 183338
rect 38234 147338 38266 147894
rect 38822 147338 38854 147894
rect 38234 111894 38854 147338
rect 38234 111338 38266 111894
rect 38822 111338 38854 111894
rect 38234 75894 38854 111338
rect 38234 75338 38266 75894
rect 38822 75338 38854 75894
rect 38234 39894 38854 75338
rect 38234 39338 38266 39894
rect 38822 39338 38854 39894
rect 38234 3894 38854 39338
rect 38234 3338 38266 3894
rect 38822 3338 38854 3894
rect 38234 -1306 38854 3338
rect 38234 -1862 38266 -1306
rect 38822 -1862 38854 -1306
rect 38234 -7654 38854 -1862
rect 39474 706758 40094 711590
rect 39474 706202 39506 706758
rect 40062 706202 40094 706758
rect 39474 689134 40094 706202
rect 39474 688578 39506 689134
rect 40062 688578 40094 689134
rect 39474 653134 40094 688578
rect 39474 652578 39506 653134
rect 40062 652578 40094 653134
rect 39474 617134 40094 652578
rect 39474 616578 39506 617134
rect 40062 616578 40094 617134
rect 39474 581134 40094 616578
rect 39474 580578 39506 581134
rect 40062 580578 40094 581134
rect 39474 545134 40094 580578
rect 39474 544578 39506 545134
rect 40062 544578 40094 545134
rect 39474 509134 40094 544578
rect 39474 508578 39506 509134
rect 40062 508578 40094 509134
rect 39474 473134 40094 508578
rect 39474 472578 39506 473134
rect 40062 472578 40094 473134
rect 39474 437134 40094 472578
rect 39474 436578 39506 437134
rect 40062 436578 40094 437134
rect 39474 401134 40094 436578
rect 39474 400578 39506 401134
rect 40062 400578 40094 401134
rect 39474 365134 40094 400578
rect 39474 364578 39506 365134
rect 40062 364578 40094 365134
rect 39474 329134 40094 364578
rect 39474 328578 39506 329134
rect 40062 328578 40094 329134
rect 39474 293134 40094 328578
rect 39474 292578 39506 293134
rect 40062 292578 40094 293134
rect 39474 257134 40094 292578
rect 39474 256578 39506 257134
rect 40062 256578 40094 257134
rect 39474 221134 40094 256578
rect 39474 220578 39506 221134
rect 40062 220578 40094 221134
rect 39474 185134 40094 220578
rect 39474 184578 39506 185134
rect 40062 184578 40094 185134
rect 39474 149134 40094 184578
rect 39474 148578 39506 149134
rect 40062 148578 40094 149134
rect 39474 113134 40094 148578
rect 39474 112578 39506 113134
rect 40062 112578 40094 113134
rect 39474 77134 40094 112578
rect 39474 76578 39506 77134
rect 40062 76578 40094 77134
rect 39474 41134 40094 76578
rect 39474 40578 39506 41134
rect 40062 40578 40094 41134
rect 39474 5134 40094 40578
rect 39474 4578 39506 5134
rect 40062 4578 40094 5134
rect 39474 -2266 40094 4578
rect 39474 -2822 39506 -2266
rect 40062 -2822 40094 -2266
rect 39474 -7654 40094 -2822
rect 40714 707718 41334 711590
rect 40714 707162 40746 707718
rect 41302 707162 41334 707718
rect 40714 690374 41334 707162
rect 40714 689818 40746 690374
rect 41302 689818 41334 690374
rect 40714 654374 41334 689818
rect 40714 653818 40746 654374
rect 41302 653818 41334 654374
rect 40714 618374 41334 653818
rect 40714 617818 40746 618374
rect 41302 617818 41334 618374
rect 40714 582374 41334 617818
rect 40714 581818 40746 582374
rect 41302 581818 41334 582374
rect 40714 546374 41334 581818
rect 40714 545818 40746 546374
rect 41302 545818 41334 546374
rect 40714 510374 41334 545818
rect 40714 509818 40746 510374
rect 41302 509818 41334 510374
rect 40714 474374 41334 509818
rect 40714 473818 40746 474374
rect 41302 473818 41334 474374
rect 40714 438374 41334 473818
rect 40714 437818 40746 438374
rect 41302 437818 41334 438374
rect 40714 402374 41334 437818
rect 40714 401818 40746 402374
rect 41302 401818 41334 402374
rect 40714 366374 41334 401818
rect 40714 365818 40746 366374
rect 41302 365818 41334 366374
rect 40714 330374 41334 365818
rect 40714 329818 40746 330374
rect 41302 329818 41334 330374
rect 40714 294374 41334 329818
rect 40714 293818 40746 294374
rect 41302 293818 41334 294374
rect 40714 258374 41334 293818
rect 40714 257818 40746 258374
rect 41302 257818 41334 258374
rect 40714 222374 41334 257818
rect 40714 221818 40746 222374
rect 41302 221818 41334 222374
rect 40714 186374 41334 221818
rect 40714 185818 40746 186374
rect 41302 185818 41334 186374
rect 40714 150374 41334 185818
rect 40714 149818 40746 150374
rect 41302 149818 41334 150374
rect 40714 114374 41334 149818
rect 40714 113818 40746 114374
rect 41302 113818 41334 114374
rect 40714 78374 41334 113818
rect 40714 77818 40746 78374
rect 41302 77818 41334 78374
rect 40714 42374 41334 77818
rect 40714 41818 40746 42374
rect 41302 41818 41334 42374
rect 40714 6374 41334 41818
rect 40714 5818 40746 6374
rect 41302 5818 41334 6374
rect 40714 -3226 41334 5818
rect 40714 -3782 40746 -3226
rect 41302 -3782 41334 -3226
rect 40714 -7654 41334 -3782
rect 41954 708678 42574 711590
rect 41954 708122 41986 708678
rect 42542 708122 42574 708678
rect 41954 691614 42574 708122
rect 41954 691058 41986 691614
rect 42542 691058 42574 691614
rect 41954 655614 42574 691058
rect 41954 655058 41986 655614
rect 42542 655058 42574 655614
rect 41954 619614 42574 655058
rect 41954 619058 41986 619614
rect 42542 619058 42574 619614
rect 41954 583614 42574 619058
rect 41954 583058 41986 583614
rect 42542 583058 42574 583614
rect 41954 547614 42574 583058
rect 41954 547058 41986 547614
rect 42542 547058 42574 547614
rect 41954 511614 42574 547058
rect 41954 511058 41986 511614
rect 42542 511058 42574 511614
rect 41954 475614 42574 511058
rect 41954 475058 41986 475614
rect 42542 475058 42574 475614
rect 41954 439614 42574 475058
rect 41954 439058 41986 439614
rect 42542 439058 42574 439614
rect 41954 403614 42574 439058
rect 41954 403058 41986 403614
rect 42542 403058 42574 403614
rect 41954 367614 42574 403058
rect 41954 367058 41986 367614
rect 42542 367058 42574 367614
rect 41954 331614 42574 367058
rect 41954 331058 41986 331614
rect 42542 331058 42574 331614
rect 41954 295614 42574 331058
rect 41954 295058 41986 295614
rect 42542 295058 42574 295614
rect 41954 259614 42574 295058
rect 41954 259058 41986 259614
rect 42542 259058 42574 259614
rect 41954 223614 42574 259058
rect 41954 223058 41986 223614
rect 42542 223058 42574 223614
rect 41954 187614 42574 223058
rect 41954 187058 41986 187614
rect 42542 187058 42574 187614
rect 41954 151614 42574 187058
rect 41954 151058 41986 151614
rect 42542 151058 42574 151614
rect 41954 115614 42574 151058
rect 41954 115058 41986 115614
rect 42542 115058 42574 115614
rect 41954 79614 42574 115058
rect 41954 79058 41986 79614
rect 42542 79058 42574 79614
rect 41954 43614 42574 79058
rect 41954 43058 41986 43614
rect 42542 43058 42574 43614
rect 41954 7614 42574 43058
rect 41954 7058 41986 7614
rect 42542 7058 42574 7614
rect 41954 -4186 42574 7058
rect 41954 -4742 41986 -4186
rect 42542 -4742 42574 -4186
rect 41954 -7654 42574 -4742
rect 43194 709638 43814 711590
rect 43194 709082 43226 709638
rect 43782 709082 43814 709638
rect 43194 692854 43814 709082
rect 43194 692298 43226 692854
rect 43782 692298 43814 692854
rect 43194 656854 43814 692298
rect 43194 656298 43226 656854
rect 43782 656298 43814 656854
rect 43194 620854 43814 656298
rect 43194 620298 43226 620854
rect 43782 620298 43814 620854
rect 43194 584854 43814 620298
rect 43194 584298 43226 584854
rect 43782 584298 43814 584854
rect 43194 548854 43814 584298
rect 43194 548298 43226 548854
rect 43782 548298 43814 548854
rect 43194 512854 43814 548298
rect 43194 512298 43226 512854
rect 43782 512298 43814 512854
rect 43194 476854 43814 512298
rect 43194 476298 43226 476854
rect 43782 476298 43814 476854
rect 43194 440854 43814 476298
rect 43194 440298 43226 440854
rect 43782 440298 43814 440854
rect 43194 404854 43814 440298
rect 43194 404298 43226 404854
rect 43782 404298 43814 404854
rect 43194 368854 43814 404298
rect 43194 368298 43226 368854
rect 43782 368298 43814 368854
rect 43194 332854 43814 368298
rect 43194 332298 43226 332854
rect 43782 332298 43814 332854
rect 43194 296854 43814 332298
rect 43194 296298 43226 296854
rect 43782 296298 43814 296854
rect 43194 260854 43814 296298
rect 43194 260298 43226 260854
rect 43782 260298 43814 260854
rect 43194 224854 43814 260298
rect 43194 224298 43226 224854
rect 43782 224298 43814 224854
rect 43194 188854 43814 224298
rect 43194 188298 43226 188854
rect 43782 188298 43814 188854
rect 43194 152854 43814 188298
rect 43194 152298 43226 152854
rect 43782 152298 43814 152854
rect 43194 116854 43814 152298
rect 43194 116298 43226 116854
rect 43782 116298 43814 116854
rect 43194 80854 43814 116298
rect 43194 80298 43226 80854
rect 43782 80298 43814 80854
rect 43194 44854 43814 80298
rect 43194 44298 43226 44854
rect 43782 44298 43814 44854
rect 43194 8854 43814 44298
rect 43194 8298 43226 8854
rect 43782 8298 43814 8854
rect 43194 -5146 43814 8298
rect 43194 -5702 43226 -5146
rect 43782 -5702 43814 -5146
rect 43194 -7654 43814 -5702
rect 44434 710598 45054 711590
rect 44434 710042 44466 710598
rect 45022 710042 45054 710598
rect 44434 694094 45054 710042
rect 44434 693538 44466 694094
rect 45022 693538 45054 694094
rect 44434 658094 45054 693538
rect 44434 657538 44466 658094
rect 45022 657538 45054 658094
rect 44434 622094 45054 657538
rect 44434 621538 44466 622094
rect 45022 621538 45054 622094
rect 44434 586094 45054 621538
rect 44434 585538 44466 586094
rect 45022 585538 45054 586094
rect 44434 550094 45054 585538
rect 44434 549538 44466 550094
rect 45022 549538 45054 550094
rect 44434 514094 45054 549538
rect 44434 513538 44466 514094
rect 45022 513538 45054 514094
rect 44434 478094 45054 513538
rect 44434 477538 44466 478094
rect 45022 477538 45054 478094
rect 44434 442094 45054 477538
rect 44434 441538 44466 442094
rect 45022 441538 45054 442094
rect 44434 406094 45054 441538
rect 44434 405538 44466 406094
rect 45022 405538 45054 406094
rect 44434 370094 45054 405538
rect 44434 369538 44466 370094
rect 45022 369538 45054 370094
rect 44434 334094 45054 369538
rect 44434 333538 44466 334094
rect 45022 333538 45054 334094
rect 44434 298094 45054 333538
rect 44434 297538 44466 298094
rect 45022 297538 45054 298094
rect 44434 262094 45054 297538
rect 44434 261538 44466 262094
rect 45022 261538 45054 262094
rect 44434 226094 45054 261538
rect 44434 225538 44466 226094
rect 45022 225538 45054 226094
rect 44434 190094 45054 225538
rect 44434 189538 44466 190094
rect 45022 189538 45054 190094
rect 44434 154094 45054 189538
rect 44434 153538 44466 154094
rect 45022 153538 45054 154094
rect 44434 118094 45054 153538
rect 44434 117538 44466 118094
rect 45022 117538 45054 118094
rect 44434 82094 45054 117538
rect 44434 81538 44466 82094
rect 45022 81538 45054 82094
rect 44434 46094 45054 81538
rect 44434 45538 44466 46094
rect 45022 45538 45054 46094
rect 44434 10094 45054 45538
rect 44434 9538 44466 10094
rect 45022 9538 45054 10094
rect 44434 -6106 45054 9538
rect 44434 -6662 44466 -6106
rect 45022 -6662 45054 -6106
rect 44434 -7654 45054 -6662
rect 45674 711558 46294 711590
rect 45674 711002 45706 711558
rect 46262 711002 46294 711558
rect 45674 695334 46294 711002
rect 45674 694778 45706 695334
rect 46262 694778 46294 695334
rect 45674 659334 46294 694778
rect 45674 658778 45706 659334
rect 46262 658778 46294 659334
rect 45674 623334 46294 658778
rect 45674 622778 45706 623334
rect 46262 622778 46294 623334
rect 45674 587334 46294 622778
rect 45674 586778 45706 587334
rect 46262 586778 46294 587334
rect 45674 551334 46294 586778
rect 45674 550778 45706 551334
rect 46262 550778 46294 551334
rect 45674 515334 46294 550778
rect 45674 514778 45706 515334
rect 46262 514778 46294 515334
rect 45674 479334 46294 514778
rect 45674 478778 45706 479334
rect 46262 478778 46294 479334
rect 45674 443334 46294 478778
rect 45674 442778 45706 443334
rect 46262 442778 46294 443334
rect 45674 407334 46294 442778
rect 45674 406778 45706 407334
rect 46262 406778 46294 407334
rect 45674 371334 46294 406778
rect 45674 370778 45706 371334
rect 46262 370778 46294 371334
rect 45674 335334 46294 370778
rect 45674 334778 45706 335334
rect 46262 334778 46294 335334
rect 45674 299334 46294 334778
rect 45674 298778 45706 299334
rect 46262 298778 46294 299334
rect 45674 263334 46294 298778
rect 45674 262778 45706 263334
rect 46262 262778 46294 263334
rect 45674 227334 46294 262778
rect 45674 226778 45706 227334
rect 46262 226778 46294 227334
rect 45674 191334 46294 226778
rect 45674 190778 45706 191334
rect 46262 190778 46294 191334
rect 45674 155334 46294 190778
rect 45674 154778 45706 155334
rect 46262 154778 46294 155334
rect 45674 119334 46294 154778
rect 45674 118778 45706 119334
rect 46262 118778 46294 119334
rect 45674 83334 46294 118778
rect 45674 82778 45706 83334
rect 46262 82778 46294 83334
rect 45674 47334 46294 82778
rect 45674 46778 45706 47334
rect 46262 46778 46294 47334
rect 45674 11334 46294 46778
rect 45674 10778 45706 11334
rect 46262 10778 46294 11334
rect 45674 -7066 46294 10778
rect 45674 -7622 45706 -7066
rect 46262 -7622 46294 -7066
rect 45674 -7654 46294 -7622
rect 72994 704838 73614 711590
rect 72994 704282 73026 704838
rect 73582 704282 73614 704838
rect 72994 686654 73614 704282
rect 72994 686098 73026 686654
rect 73582 686098 73614 686654
rect 72994 650654 73614 686098
rect 72994 650098 73026 650654
rect 73582 650098 73614 650654
rect 72994 614654 73614 650098
rect 72994 614098 73026 614654
rect 73582 614098 73614 614654
rect 72994 578654 73614 614098
rect 72994 578098 73026 578654
rect 73582 578098 73614 578654
rect 72994 542654 73614 578098
rect 72994 542098 73026 542654
rect 73582 542098 73614 542654
rect 72994 506654 73614 542098
rect 72994 506098 73026 506654
rect 73582 506098 73614 506654
rect 72994 470654 73614 506098
rect 72994 470098 73026 470654
rect 73582 470098 73614 470654
rect 72994 434654 73614 470098
rect 72994 434098 73026 434654
rect 73582 434098 73614 434654
rect 72994 398654 73614 434098
rect 72994 398098 73026 398654
rect 73582 398098 73614 398654
rect 72994 362654 73614 398098
rect 72994 362098 73026 362654
rect 73582 362098 73614 362654
rect 72994 326654 73614 362098
rect 72994 326098 73026 326654
rect 73582 326098 73614 326654
rect 72994 290654 73614 326098
rect 72994 290098 73026 290654
rect 73582 290098 73614 290654
rect 72994 254654 73614 290098
rect 72994 254098 73026 254654
rect 73582 254098 73614 254654
rect 72994 218654 73614 254098
rect 72994 218098 73026 218654
rect 73582 218098 73614 218654
rect 72994 182654 73614 218098
rect 72994 182098 73026 182654
rect 73582 182098 73614 182654
rect 72994 146654 73614 182098
rect 72994 146098 73026 146654
rect 73582 146098 73614 146654
rect 72994 110654 73614 146098
rect 72994 110098 73026 110654
rect 73582 110098 73614 110654
rect 72994 74654 73614 110098
rect 72994 74098 73026 74654
rect 73582 74098 73614 74654
rect 72994 38654 73614 74098
rect 72994 38098 73026 38654
rect 73582 38098 73614 38654
rect 72994 2654 73614 38098
rect 72994 2098 73026 2654
rect 73582 2098 73614 2654
rect 72994 -346 73614 2098
rect 72994 -902 73026 -346
rect 73582 -902 73614 -346
rect 72994 -7654 73614 -902
rect 74234 705798 74854 711590
rect 74234 705242 74266 705798
rect 74822 705242 74854 705798
rect 74234 687894 74854 705242
rect 74234 687338 74266 687894
rect 74822 687338 74854 687894
rect 74234 651894 74854 687338
rect 74234 651338 74266 651894
rect 74822 651338 74854 651894
rect 74234 615894 74854 651338
rect 74234 615338 74266 615894
rect 74822 615338 74854 615894
rect 74234 579894 74854 615338
rect 74234 579338 74266 579894
rect 74822 579338 74854 579894
rect 74234 543894 74854 579338
rect 74234 543338 74266 543894
rect 74822 543338 74854 543894
rect 74234 507894 74854 543338
rect 74234 507338 74266 507894
rect 74822 507338 74854 507894
rect 74234 471894 74854 507338
rect 74234 471338 74266 471894
rect 74822 471338 74854 471894
rect 74234 435894 74854 471338
rect 74234 435338 74266 435894
rect 74822 435338 74854 435894
rect 74234 399894 74854 435338
rect 74234 399338 74266 399894
rect 74822 399338 74854 399894
rect 74234 363894 74854 399338
rect 74234 363338 74266 363894
rect 74822 363338 74854 363894
rect 74234 327894 74854 363338
rect 74234 327338 74266 327894
rect 74822 327338 74854 327894
rect 74234 291894 74854 327338
rect 74234 291338 74266 291894
rect 74822 291338 74854 291894
rect 74234 255894 74854 291338
rect 74234 255338 74266 255894
rect 74822 255338 74854 255894
rect 74234 219894 74854 255338
rect 74234 219338 74266 219894
rect 74822 219338 74854 219894
rect 74234 183894 74854 219338
rect 74234 183338 74266 183894
rect 74822 183338 74854 183894
rect 74234 147894 74854 183338
rect 74234 147338 74266 147894
rect 74822 147338 74854 147894
rect 74234 111894 74854 147338
rect 74234 111338 74266 111894
rect 74822 111338 74854 111894
rect 74234 75894 74854 111338
rect 74234 75338 74266 75894
rect 74822 75338 74854 75894
rect 74234 39894 74854 75338
rect 74234 39338 74266 39894
rect 74822 39338 74854 39894
rect 74234 3894 74854 39338
rect 74234 3338 74266 3894
rect 74822 3338 74854 3894
rect 74234 -1306 74854 3338
rect 74234 -1862 74266 -1306
rect 74822 -1862 74854 -1306
rect 74234 -7654 74854 -1862
rect 75474 706758 76094 711590
rect 75474 706202 75506 706758
rect 76062 706202 76094 706758
rect 75474 689134 76094 706202
rect 75474 688578 75506 689134
rect 76062 688578 76094 689134
rect 75474 653134 76094 688578
rect 75474 652578 75506 653134
rect 76062 652578 76094 653134
rect 75474 617134 76094 652578
rect 75474 616578 75506 617134
rect 76062 616578 76094 617134
rect 75474 581134 76094 616578
rect 75474 580578 75506 581134
rect 76062 580578 76094 581134
rect 75474 545134 76094 580578
rect 75474 544578 75506 545134
rect 76062 544578 76094 545134
rect 75474 509134 76094 544578
rect 75474 508578 75506 509134
rect 76062 508578 76094 509134
rect 75474 473134 76094 508578
rect 75474 472578 75506 473134
rect 76062 472578 76094 473134
rect 75474 437134 76094 472578
rect 75474 436578 75506 437134
rect 76062 436578 76094 437134
rect 75474 401134 76094 436578
rect 75474 400578 75506 401134
rect 76062 400578 76094 401134
rect 75474 365134 76094 400578
rect 75474 364578 75506 365134
rect 76062 364578 76094 365134
rect 75474 329134 76094 364578
rect 75474 328578 75506 329134
rect 76062 328578 76094 329134
rect 75474 293134 76094 328578
rect 75474 292578 75506 293134
rect 76062 292578 76094 293134
rect 75474 257134 76094 292578
rect 75474 256578 75506 257134
rect 76062 256578 76094 257134
rect 75474 221134 76094 256578
rect 75474 220578 75506 221134
rect 76062 220578 76094 221134
rect 75474 185134 76094 220578
rect 75474 184578 75506 185134
rect 76062 184578 76094 185134
rect 75474 149134 76094 184578
rect 75474 148578 75506 149134
rect 76062 148578 76094 149134
rect 75474 113134 76094 148578
rect 75474 112578 75506 113134
rect 76062 112578 76094 113134
rect 75474 77134 76094 112578
rect 75474 76578 75506 77134
rect 76062 76578 76094 77134
rect 75474 41134 76094 76578
rect 75474 40578 75506 41134
rect 76062 40578 76094 41134
rect 75474 5134 76094 40578
rect 75474 4578 75506 5134
rect 76062 4578 76094 5134
rect 75474 -2266 76094 4578
rect 75474 -2822 75506 -2266
rect 76062 -2822 76094 -2266
rect 75474 -7654 76094 -2822
rect 76714 707718 77334 711590
rect 76714 707162 76746 707718
rect 77302 707162 77334 707718
rect 76714 690374 77334 707162
rect 76714 689818 76746 690374
rect 77302 689818 77334 690374
rect 76714 654374 77334 689818
rect 76714 653818 76746 654374
rect 77302 653818 77334 654374
rect 76714 618374 77334 653818
rect 76714 617818 76746 618374
rect 77302 617818 77334 618374
rect 76714 582374 77334 617818
rect 76714 581818 76746 582374
rect 77302 581818 77334 582374
rect 76714 546374 77334 581818
rect 76714 545818 76746 546374
rect 77302 545818 77334 546374
rect 76714 510374 77334 545818
rect 76714 509818 76746 510374
rect 77302 509818 77334 510374
rect 76714 474374 77334 509818
rect 76714 473818 76746 474374
rect 77302 473818 77334 474374
rect 76714 438374 77334 473818
rect 76714 437818 76746 438374
rect 77302 437818 77334 438374
rect 76714 402374 77334 437818
rect 76714 401818 76746 402374
rect 77302 401818 77334 402374
rect 76714 366374 77334 401818
rect 76714 365818 76746 366374
rect 77302 365818 77334 366374
rect 76714 330374 77334 365818
rect 76714 329818 76746 330374
rect 77302 329818 77334 330374
rect 76714 294374 77334 329818
rect 76714 293818 76746 294374
rect 77302 293818 77334 294374
rect 76714 258374 77334 293818
rect 76714 257818 76746 258374
rect 77302 257818 77334 258374
rect 76714 222374 77334 257818
rect 76714 221818 76746 222374
rect 77302 221818 77334 222374
rect 76714 186374 77334 221818
rect 76714 185818 76746 186374
rect 77302 185818 77334 186374
rect 76714 150374 77334 185818
rect 76714 149818 76746 150374
rect 77302 149818 77334 150374
rect 76714 114374 77334 149818
rect 76714 113818 76746 114374
rect 77302 113818 77334 114374
rect 76714 78374 77334 113818
rect 76714 77818 76746 78374
rect 77302 77818 77334 78374
rect 76714 42374 77334 77818
rect 76714 41818 76746 42374
rect 77302 41818 77334 42374
rect 76714 6374 77334 41818
rect 76714 5818 76746 6374
rect 77302 5818 77334 6374
rect 76714 -3226 77334 5818
rect 76714 -3782 76746 -3226
rect 77302 -3782 77334 -3226
rect 76714 -7654 77334 -3782
rect 77954 708678 78574 711590
rect 77954 708122 77986 708678
rect 78542 708122 78574 708678
rect 77954 691614 78574 708122
rect 77954 691058 77986 691614
rect 78542 691058 78574 691614
rect 77954 655614 78574 691058
rect 77954 655058 77986 655614
rect 78542 655058 78574 655614
rect 77954 619614 78574 655058
rect 77954 619058 77986 619614
rect 78542 619058 78574 619614
rect 77954 583614 78574 619058
rect 77954 583058 77986 583614
rect 78542 583058 78574 583614
rect 77954 547614 78574 583058
rect 77954 547058 77986 547614
rect 78542 547058 78574 547614
rect 77954 511614 78574 547058
rect 77954 511058 77986 511614
rect 78542 511058 78574 511614
rect 77954 475614 78574 511058
rect 77954 475058 77986 475614
rect 78542 475058 78574 475614
rect 77954 439614 78574 475058
rect 77954 439058 77986 439614
rect 78542 439058 78574 439614
rect 77954 403614 78574 439058
rect 77954 403058 77986 403614
rect 78542 403058 78574 403614
rect 77954 367614 78574 403058
rect 77954 367058 77986 367614
rect 78542 367058 78574 367614
rect 77954 331614 78574 367058
rect 77954 331058 77986 331614
rect 78542 331058 78574 331614
rect 77954 295614 78574 331058
rect 77954 295058 77986 295614
rect 78542 295058 78574 295614
rect 77954 259614 78574 295058
rect 77954 259058 77986 259614
rect 78542 259058 78574 259614
rect 77954 223614 78574 259058
rect 77954 223058 77986 223614
rect 78542 223058 78574 223614
rect 77954 187614 78574 223058
rect 77954 187058 77986 187614
rect 78542 187058 78574 187614
rect 77954 151614 78574 187058
rect 77954 151058 77986 151614
rect 78542 151058 78574 151614
rect 77954 115614 78574 151058
rect 77954 115058 77986 115614
rect 78542 115058 78574 115614
rect 77954 79614 78574 115058
rect 77954 79058 77986 79614
rect 78542 79058 78574 79614
rect 77954 43614 78574 79058
rect 77954 43058 77986 43614
rect 78542 43058 78574 43614
rect 77954 7614 78574 43058
rect 77954 7058 77986 7614
rect 78542 7058 78574 7614
rect 77954 -4186 78574 7058
rect 77954 -4742 77986 -4186
rect 78542 -4742 78574 -4186
rect 77954 -7654 78574 -4742
rect 79194 709638 79814 711590
rect 79194 709082 79226 709638
rect 79782 709082 79814 709638
rect 79194 692854 79814 709082
rect 79194 692298 79226 692854
rect 79782 692298 79814 692854
rect 79194 656854 79814 692298
rect 79194 656298 79226 656854
rect 79782 656298 79814 656854
rect 79194 620854 79814 656298
rect 79194 620298 79226 620854
rect 79782 620298 79814 620854
rect 79194 584854 79814 620298
rect 79194 584298 79226 584854
rect 79782 584298 79814 584854
rect 79194 548854 79814 584298
rect 79194 548298 79226 548854
rect 79782 548298 79814 548854
rect 79194 512854 79814 548298
rect 79194 512298 79226 512854
rect 79782 512298 79814 512854
rect 79194 476854 79814 512298
rect 79194 476298 79226 476854
rect 79782 476298 79814 476854
rect 79194 440854 79814 476298
rect 79194 440298 79226 440854
rect 79782 440298 79814 440854
rect 79194 404854 79814 440298
rect 79194 404298 79226 404854
rect 79782 404298 79814 404854
rect 79194 368854 79814 404298
rect 79194 368298 79226 368854
rect 79782 368298 79814 368854
rect 79194 332854 79814 368298
rect 79194 332298 79226 332854
rect 79782 332298 79814 332854
rect 79194 296854 79814 332298
rect 79194 296298 79226 296854
rect 79782 296298 79814 296854
rect 79194 260854 79814 296298
rect 79194 260298 79226 260854
rect 79782 260298 79814 260854
rect 79194 224854 79814 260298
rect 79194 224298 79226 224854
rect 79782 224298 79814 224854
rect 79194 188854 79814 224298
rect 79194 188298 79226 188854
rect 79782 188298 79814 188854
rect 79194 152854 79814 188298
rect 79194 152298 79226 152854
rect 79782 152298 79814 152854
rect 79194 116854 79814 152298
rect 79194 116298 79226 116854
rect 79782 116298 79814 116854
rect 79194 80854 79814 116298
rect 79194 80298 79226 80854
rect 79782 80298 79814 80854
rect 79194 44854 79814 80298
rect 79194 44298 79226 44854
rect 79782 44298 79814 44854
rect 79194 8854 79814 44298
rect 79194 8298 79226 8854
rect 79782 8298 79814 8854
rect 79194 -5146 79814 8298
rect 79194 -5702 79226 -5146
rect 79782 -5702 79814 -5146
rect 79194 -7654 79814 -5702
rect 80434 710598 81054 711590
rect 80434 710042 80466 710598
rect 81022 710042 81054 710598
rect 80434 694094 81054 710042
rect 80434 693538 80466 694094
rect 81022 693538 81054 694094
rect 80434 658094 81054 693538
rect 80434 657538 80466 658094
rect 81022 657538 81054 658094
rect 80434 622094 81054 657538
rect 80434 621538 80466 622094
rect 81022 621538 81054 622094
rect 80434 586094 81054 621538
rect 80434 585538 80466 586094
rect 81022 585538 81054 586094
rect 80434 550094 81054 585538
rect 80434 549538 80466 550094
rect 81022 549538 81054 550094
rect 80434 514094 81054 549538
rect 80434 513538 80466 514094
rect 81022 513538 81054 514094
rect 80434 478094 81054 513538
rect 80434 477538 80466 478094
rect 81022 477538 81054 478094
rect 80434 442094 81054 477538
rect 80434 441538 80466 442094
rect 81022 441538 81054 442094
rect 80434 406094 81054 441538
rect 80434 405538 80466 406094
rect 81022 405538 81054 406094
rect 80434 370094 81054 405538
rect 80434 369538 80466 370094
rect 81022 369538 81054 370094
rect 80434 334094 81054 369538
rect 80434 333538 80466 334094
rect 81022 333538 81054 334094
rect 80434 298094 81054 333538
rect 80434 297538 80466 298094
rect 81022 297538 81054 298094
rect 80434 262094 81054 297538
rect 80434 261538 80466 262094
rect 81022 261538 81054 262094
rect 80434 226094 81054 261538
rect 80434 225538 80466 226094
rect 81022 225538 81054 226094
rect 80434 190094 81054 225538
rect 80434 189538 80466 190094
rect 81022 189538 81054 190094
rect 80434 154094 81054 189538
rect 80434 153538 80466 154094
rect 81022 153538 81054 154094
rect 80434 118094 81054 153538
rect 80434 117538 80466 118094
rect 81022 117538 81054 118094
rect 80434 82094 81054 117538
rect 80434 81538 80466 82094
rect 81022 81538 81054 82094
rect 80434 46094 81054 81538
rect 80434 45538 80466 46094
rect 81022 45538 81054 46094
rect 80434 10094 81054 45538
rect 80434 9538 80466 10094
rect 81022 9538 81054 10094
rect 80434 -6106 81054 9538
rect 80434 -6662 80466 -6106
rect 81022 -6662 81054 -6106
rect 80434 -7654 81054 -6662
rect 81674 711558 82294 711590
rect 81674 711002 81706 711558
rect 82262 711002 82294 711558
rect 81674 695334 82294 711002
rect 81674 694778 81706 695334
rect 82262 694778 82294 695334
rect 81674 659334 82294 694778
rect 81674 658778 81706 659334
rect 82262 658778 82294 659334
rect 81674 623334 82294 658778
rect 81674 622778 81706 623334
rect 82262 622778 82294 623334
rect 81674 587334 82294 622778
rect 81674 586778 81706 587334
rect 82262 586778 82294 587334
rect 81674 551334 82294 586778
rect 81674 550778 81706 551334
rect 82262 550778 82294 551334
rect 81674 515334 82294 550778
rect 81674 514778 81706 515334
rect 82262 514778 82294 515334
rect 81674 479334 82294 514778
rect 81674 478778 81706 479334
rect 82262 478778 82294 479334
rect 81674 443334 82294 478778
rect 81674 442778 81706 443334
rect 82262 442778 82294 443334
rect 81674 407334 82294 442778
rect 81674 406778 81706 407334
rect 82262 406778 82294 407334
rect 81674 371334 82294 406778
rect 81674 370778 81706 371334
rect 82262 370778 82294 371334
rect 81674 335334 82294 370778
rect 81674 334778 81706 335334
rect 82262 334778 82294 335334
rect 81674 299334 82294 334778
rect 81674 298778 81706 299334
rect 82262 298778 82294 299334
rect 81674 263334 82294 298778
rect 81674 262778 81706 263334
rect 82262 262778 82294 263334
rect 81674 227334 82294 262778
rect 81674 226778 81706 227334
rect 82262 226778 82294 227334
rect 81674 191334 82294 226778
rect 81674 190778 81706 191334
rect 82262 190778 82294 191334
rect 81674 155334 82294 190778
rect 81674 154778 81706 155334
rect 82262 154778 82294 155334
rect 81674 119334 82294 154778
rect 81674 118778 81706 119334
rect 82262 118778 82294 119334
rect 81674 83334 82294 118778
rect 81674 82778 81706 83334
rect 82262 82778 82294 83334
rect 81674 47334 82294 82778
rect 81674 46778 81706 47334
rect 82262 46778 82294 47334
rect 81674 11334 82294 46778
rect 81674 10778 81706 11334
rect 82262 10778 82294 11334
rect 81674 -7066 82294 10778
rect 81674 -7622 81706 -7066
rect 82262 -7622 82294 -7066
rect 81674 -7654 82294 -7622
rect 108994 704838 109614 711590
rect 108994 704282 109026 704838
rect 109582 704282 109614 704838
rect 108994 686654 109614 704282
rect 108994 686098 109026 686654
rect 109582 686098 109614 686654
rect 108994 650654 109614 686098
rect 108994 650098 109026 650654
rect 109582 650098 109614 650654
rect 108994 614654 109614 650098
rect 108994 614098 109026 614654
rect 109582 614098 109614 614654
rect 108994 578654 109614 614098
rect 108994 578098 109026 578654
rect 109582 578098 109614 578654
rect 108994 542654 109614 578098
rect 108994 542098 109026 542654
rect 109582 542098 109614 542654
rect 108994 506654 109614 542098
rect 108994 506098 109026 506654
rect 109582 506098 109614 506654
rect 108994 470654 109614 506098
rect 108994 470098 109026 470654
rect 109582 470098 109614 470654
rect 108994 434654 109614 470098
rect 108994 434098 109026 434654
rect 109582 434098 109614 434654
rect 108994 398654 109614 434098
rect 108994 398098 109026 398654
rect 109582 398098 109614 398654
rect 108994 362654 109614 398098
rect 108994 362098 109026 362654
rect 109582 362098 109614 362654
rect 108994 326654 109614 362098
rect 108994 326098 109026 326654
rect 109582 326098 109614 326654
rect 108994 290654 109614 326098
rect 108994 290098 109026 290654
rect 109582 290098 109614 290654
rect 108994 254654 109614 290098
rect 108994 254098 109026 254654
rect 109582 254098 109614 254654
rect 108994 218654 109614 254098
rect 108994 218098 109026 218654
rect 109582 218098 109614 218654
rect 108994 182654 109614 218098
rect 108994 182098 109026 182654
rect 109582 182098 109614 182654
rect 108994 146654 109614 182098
rect 108994 146098 109026 146654
rect 109582 146098 109614 146654
rect 108994 110654 109614 146098
rect 108994 110098 109026 110654
rect 109582 110098 109614 110654
rect 108994 74654 109614 110098
rect 108994 74098 109026 74654
rect 109582 74098 109614 74654
rect 108994 38654 109614 74098
rect 108994 38098 109026 38654
rect 109582 38098 109614 38654
rect 108994 2654 109614 38098
rect 108994 2098 109026 2654
rect 109582 2098 109614 2654
rect 108994 -346 109614 2098
rect 108994 -902 109026 -346
rect 109582 -902 109614 -346
rect 108994 -7654 109614 -902
rect 110234 705798 110854 711590
rect 110234 705242 110266 705798
rect 110822 705242 110854 705798
rect 110234 687894 110854 705242
rect 110234 687338 110266 687894
rect 110822 687338 110854 687894
rect 110234 651894 110854 687338
rect 110234 651338 110266 651894
rect 110822 651338 110854 651894
rect 110234 615894 110854 651338
rect 110234 615338 110266 615894
rect 110822 615338 110854 615894
rect 110234 579894 110854 615338
rect 110234 579338 110266 579894
rect 110822 579338 110854 579894
rect 110234 543894 110854 579338
rect 110234 543338 110266 543894
rect 110822 543338 110854 543894
rect 110234 507894 110854 543338
rect 110234 507338 110266 507894
rect 110822 507338 110854 507894
rect 110234 471894 110854 507338
rect 110234 471338 110266 471894
rect 110822 471338 110854 471894
rect 110234 435894 110854 471338
rect 110234 435338 110266 435894
rect 110822 435338 110854 435894
rect 110234 399894 110854 435338
rect 110234 399338 110266 399894
rect 110822 399338 110854 399894
rect 110234 363894 110854 399338
rect 110234 363338 110266 363894
rect 110822 363338 110854 363894
rect 110234 327894 110854 363338
rect 110234 327338 110266 327894
rect 110822 327338 110854 327894
rect 110234 291894 110854 327338
rect 110234 291338 110266 291894
rect 110822 291338 110854 291894
rect 110234 255894 110854 291338
rect 110234 255338 110266 255894
rect 110822 255338 110854 255894
rect 110234 219894 110854 255338
rect 110234 219338 110266 219894
rect 110822 219338 110854 219894
rect 110234 183894 110854 219338
rect 110234 183338 110266 183894
rect 110822 183338 110854 183894
rect 110234 147894 110854 183338
rect 110234 147338 110266 147894
rect 110822 147338 110854 147894
rect 110234 111894 110854 147338
rect 110234 111338 110266 111894
rect 110822 111338 110854 111894
rect 110234 75894 110854 111338
rect 110234 75338 110266 75894
rect 110822 75338 110854 75894
rect 110234 39894 110854 75338
rect 110234 39338 110266 39894
rect 110822 39338 110854 39894
rect 110234 3894 110854 39338
rect 110234 3338 110266 3894
rect 110822 3338 110854 3894
rect 110234 -1306 110854 3338
rect 110234 -1862 110266 -1306
rect 110822 -1862 110854 -1306
rect 110234 -7654 110854 -1862
rect 111474 706758 112094 711590
rect 111474 706202 111506 706758
rect 112062 706202 112094 706758
rect 111474 689134 112094 706202
rect 111474 688578 111506 689134
rect 112062 688578 112094 689134
rect 111474 653134 112094 688578
rect 111474 652578 111506 653134
rect 112062 652578 112094 653134
rect 111474 617134 112094 652578
rect 111474 616578 111506 617134
rect 112062 616578 112094 617134
rect 111474 581134 112094 616578
rect 111474 580578 111506 581134
rect 112062 580578 112094 581134
rect 111474 545134 112094 580578
rect 111474 544578 111506 545134
rect 112062 544578 112094 545134
rect 111474 509134 112094 544578
rect 111474 508578 111506 509134
rect 112062 508578 112094 509134
rect 111474 473134 112094 508578
rect 111474 472578 111506 473134
rect 112062 472578 112094 473134
rect 111474 437134 112094 472578
rect 111474 436578 111506 437134
rect 112062 436578 112094 437134
rect 111474 401134 112094 436578
rect 111474 400578 111506 401134
rect 112062 400578 112094 401134
rect 111474 365134 112094 400578
rect 111474 364578 111506 365134
rect 112062 364578 112094 365134
rect 111474 329134 112094 364578
rect 111474 328578 111506 329134
rect 112062 328578 112094 329134
rect 111474 293134 112094 328578
rect 111474 292578 111506 293134
rect 112062 292578 112094 293134
rect 111474 257134 112094 292578
rect 111474 256578 111506 257134
rect 112062 256578 112094 257134
rect 111474 221134 112094 256578
rect 111474 220578 111506 221134
rect 112062 220578 112094 221134
rect 111474 185134 112094 220578
rect 111474 184578 111506 185134
rect 112062 184578 112094 185134
rect 111474 149134 112094 184578
rect 111474 148578 111506 149134
rect 112062 148578 112094 149134
rect 111474 113134 112094 148578
rect 111474 112578 111506 113134
rect 112062 112578 112094 113134
rect 111474 77134 112094 112578
rect 111474 76578 111506 77134
rect 112062 76578 112094 77134
rect 111474 41134 112094 76578
rect 111474 40578 111506 41134
rect 112062 40578 112094 41134
rect 111474 5134 112094 40578
rect 111474 4578 111506 5134
rect 112062 4578 112094 5134
rect 111474 -2266 112094 4578
rect 111474 -2822 111506 -2266
rect 112062 -2822 112094 -2266
rect 111474 -7654 112094 -2822
rect 112714 707718 113334 711590
rect 112714 707162 112746 707718
rect 113302 707162 113334 707718
rect 112714 690374 113334 707162
rect 112714 689818 112746 690374
rect 113302 689818 113334 690374
rect 112714 654374 113334 689818
rect 112714 653818 112746 654374
rect 113302 653818 113334 654374
rect 112714 618374 113334 653818
rect 112714 617818 112746 618374
rect 113302 617818 113334 618374
rect 112714 582374 113334 617818
rect 112714 581818 112746 582374
rect 113302 581818 113334 582374
rect 112714 546374 113334 581818
rect 112714 545818 112746 546374
rect 113302 545818 113334 546374
rect 112714 510374 113334 545818
rect 112714 509818 112746 510374
rect 113302 509818 113334 510374
rect 112714 474374 113334 509818
rect 112714 473818 112746 474374
rect 113302 473818 113334 474374
rect 112714 438374 113334 473818
rect 112714 437818 112746 438374
rect 113302 437818 113334 438374
rect 112714 402374 113334 437818
rect 112714 401818 112746 402374
rect 113302 401818 113334 402374
rect 112714 366374 113334 401818
rect 112714 365818 112746 366374
rect 113302 365818 113334 366374
rect 112714 330374 113334 365818
rect 112714 329818 112746 330374
rect 113302 329818 113334 330374
rect 112714 294374 113334 329818
rect 112714 293818 112746 294374
rect 113302 293818 113334 294374
rect 112714 258374 113334 293818
rect 112714 257818 112746 258374
rect 113302 257818 113334 258374
rect 112714 222374 113334 257818
rect 112714 221818 112746 222374
rect 113302 221818 113334 222374
rect 112714 186374 113334 221818
rect 112714 185818 112746 186374
rect 113302 185818 113334 186374
rect 112714 150374 113334 185818
rect 112714 149818 112746 150374
rect 113302 149818 113334 150374
rect 112714 114374 113334 149818
rect 112714 113818 112746 114374
rect 113302 113818 113334 114374
rect 112714 78374 113334 113818
rect 112714 77818 112746 78374
rect 113302 77818 113334 78374
rect 112714 42374 113334 77818
rect 112714 41818 112746 42374
rect 113302 41818 113334 42374
rect 112714 6374 113334 41818
rect 112714 5818 112746 6374
rect 113302 5818 113334 6374
rect 112714 -3226 113334 5818
rect 112714 -3782 112746 -3226
rect 113302 -3782 113334 -3226
rect 112714 -7654 113334 -3782
rect 113954 708678 114574 711590
rect 113954 708122 113986 708678
rect 114542 708122 114574 708678
rect 113954 691614 114574 708122
rect 113954 691058 113986 691614
rect 114542 691058 114574 691614
rect 113954 655614 114574 691058
rect 113954 655058 113986 655614
rect 114542 655058 114574 655614
rect 113954 619614 114574 655058
rect 113954 619058 113986 619614
rect 114542 619058 114574 619614
rect 113954 583614 114574 619058
rect 113954 583058 113986 583614
rect 114542 583058 114574 583614
rect 113954 547614 114574 583058
rect 113954 547058 113986 547614
rect 114542 547058 114574 547614
rect 113954 511614 114574 547058
rect 113954 511058 113986 511614
rect 114542 511058 114574 511614
rect 113954 475614 114574 511058
rect 113954 475058 113986 475614
rect 114542 475058 114574 475614
rect 113954 439614 114574 475058
rect 113954 439058 113986 439614
rect 114542 439058 114574 439614
rect 113954 403614 114574 439058
rect 113954 403058 113986 403614
rect 114542 403058 114574 403614
rect 113954 367614 114574 403058
rect 113954 367058 113986 367614
rect 114542 367058 114574 367614
rect 113954 331614 114574 367058
rect 113954 331058 113986 331614
rect 114542 331058 114574 331614
rect 113954 295614 114574 331058
rect 113954 295058 113986 295614
rect 114542 295058 114574 295614
rect 113954 259614 114574 295058
rect 113954 259058 113986 259614
rect 114542 259058 114574 259614
rect 113954 223614 114574 259058
rect 113954 223058 113986 223614
rect 114542 223058 114574 223614
rect 113954 187614 114574 223058
rect 113954 187058 113986 187614
rect 114542 187058 114574 187614
rect 113954 151614 114574 187058
rect 113954 151058 113986 151614
rect 114542 151058 114574 151614
rect 113954 115614 114574 151058
rect 113954 115058 113986 115614
rect 114542 115058 114574 115614
rect 113954 79614 114574 115058
rect 113954 79058 113986 79614
rect 114542 79058 114574 79614
rect 113954 43614 114574 79058
rect 113954 43058 113986 43614
rect 114542 43058 114574 43614
rect 113954 7614 114574 43058
rect 113954 7058 113986 7614
rect 114542 7058 114574 7614
rect 113954 -4186 114574 7058
rect 113954 -4742 113986 -4186
rect 114542 -4742 114574 -4186
rect 113954 -7654 114574 -4742
rect 115194 709638 115814 711590
rect 115194 709082 115226 709638
rect 115782 709082 115814 709638
rect 115194 692854 115814 709082
rect 115194 692298 115226 692854
rect 115782 692298 115814 692854
rect 115194 656854 115814 692298
rect 115194 656298 115226 656854
rect 115782 656298 115814 656854
rect 115194 620854 115814 656298
rect 115194 620298 115226 620854
rect 115782 620298 115814 620854
rect 115194 584854 115814 620298
rect 115194 584298 115226 584854
rect 115782 584298 115814 584854
rect 115194 548854 115814 584298
rect 115194 548298 115226 548854
rect 115782 548298 115814 548854
rect 115194 512854 115814 548298
rect 115194 512298 115226 512854
rect 115782 512298 115814 512854
rect 115194 476854 115814 512298
rect 115194 476298 115226 476854
rect 115782 476298 115814 476854
rect 115194 440854 115814 476298
rect 115194 440298 115226 440854
rect 115782 440298 115814 440854
rect 115194 404854 115814 440298
rect 115194 404298 115226 404854
rect 115782 404298 115814 404854
rect 115194 368854 115814 404298
rect 115194 368298 115226 368854
rect 115782 368298 115814 368854
rect 115194 332854 115814 368298
rect 115194 332298 115226 332854
rect 115782 332298 115814 332854
rect 115194 296854 115814 332298
rect 115194 296298 115226 296854
rect 115782 296298 115814 296854
rect 115194 260854 115814 296298
rect 115194 260298 115226 260854
rect 115782 260298 115814 260854
rect 115194 224854 115814 260298
rect 115194 224298 115226 224854
rect 115782 224298 115814 224854
rect 115194 188854 115814 224298
rect 115194 188298 115226 188854
rect 115782 188298 115814 188854
rect 115194 152854 115814 188298
rect 115194 152298 115226 152854
rect 115782 152298 115814 152854
rect 115194 116854 115814 152298
rect 115194 116298 115226 116854
rect 115782 116298 115814 116854
rect 115194 80854 115814 116298
rect 115194 80298 115226 80854
rect 115782 80298 115814 80854
rect 115194 44854 115814 80298
rect 115194 44298 115226 44854
rect 115782 44298 115814 44854
rect 115194 8854 115814 44298
rect 115194 8298 115226 8854
rect 115782 8298 115814 8854
rect 115194 -5146 115814 8298
rect 115194 -5702 115226 -5146
rect 115782 -5702 115814 -5146
rect 115194 -7654 115814 -5702
rect 116434 710598 117054 711590
rect 116434 710042 116466 710598
rect 117022 710042 117054 710598
rect 116434 694094 117054 710042
rect 116434 693538 116466 694094
rect 117022 693538 117054 694094
rect 116434 658094 117054 693538
rect 116434 657538 116466 658094
rect 117022 657538 117054 658094
rect 116434 622094 117054 657538
rect 116434 621538 116466 622094
rect 117022 621538 117054 622094
rect 116434 586094 117054 621538
rect 116434 585538 116466 586094
rect 117022 585538 117054 586094
rect 116434 550094 117054 585538
rect 116434 549538 116466 550094
rect 117022 549538 117054 550094
rect 116434 514094 117054 549538
rect 116434 513538 116466 514094
rect 117022 513538 117054 514094
rect 116434 478094 117054 513538
rect 116434 477538 116466 478094
rect 117022 477538 117054 478094
rect 116434 442094 117054 477538
rect 116434 441538 116466 442094
rect 117022 441538 117054 442094
rect 116434 406094 117054 441538
rect 116434 405538 116466 406094
rect 117022 405538 117054 406094
rect 116434 370094 117054 405538
rect 116434 369538 116466 370094
rect 117022 369538 117054 370094
rect 116434 334094 117054 369538
rect 116434 333538 116466 334094
rect 117022 333538 117054 334094
rect 116434 298094 117054 333538
rect 116434 297538 116466 298094
rect 117022 297538 117054 298094
rect 116434 262094 117054 297538
rect 116434 261538 116466 262094
rect 117022 261538 117054 262094
rect 116434 226094 117054 261538
rect 116434 225538 116466 226094
rect 117022 225538 117054 226094
rect 116434 190094 117054 225538
rect 116434 189538 116466 190094
rect 117022 189538 117054 190094
rect 116434 154094 117054 189538
rect 116434 153538 116466 154094
rect 117022 153538 117054 154094
rect 116434 118094 117054 153538
rect 116434 117538 116466 118094
rect 117022 117538 117054 118094
rect 116434 82094 117054 117538
rect 116434 81538 116466 82094
rect 117022 81538 117054 82094
rect 116434 46094 117054 81538
rect 116434 45538 116466 46094
rect 117022 45538 117054 46094
rect 116434 10094 117054 45538
rect 116434 9538 116466 10094
rect 117022 9538 117054 10094
rect 116434 -6106 117054 9538
rect 116434 -6662 116466 -6106
rect 117022 -6662 117054 -6106
rect 116434 -7654 117054 -6662
rect 117674 711558 118294 711590
rect 117674 711002 117706 711558
rect 118262 711002 118294 711558
rect 117674 695334 118294 711002
rect 117674 694778 117706 695334
rect 118262 694778 118294 695334
rect 117674 659334 118294 694778
rect 117674 658778 117706 659334
rect 118262 658778 118294 659334
rect 117674 623334 118294 658778
rect 117674 622778 117706 623334
rect 118262 622778 118294 623334
rect 117674 587334 118294 622778
rect 117674 586778 117706 587334
rect 118262 586778 118294 587334
rect 117674 551334 118294 586778
rect 117674 550778 117706 551334
rect 118262 550778 118294 551334
rect 117674 515334 118294 550778
rect 117674 514778 117706 515334
rect 118262 514778 118294 515334
rect 117674 479334 118294 514778
rect 117674 478778 117706 479334
rect 118262 478778 118294 479334
rect 117674 443334 118294 478778
rect 117674 442778 117706 443334
rect 118262 442778 118294 443334
rect 117674 407334 118294 442778
rect 117674 406778 117706 407334
rect 118262 406778 118294 407334
rect 117674 371334 118294 406778
rect 117674 370778 117706 371334
rect 118262 370778 118294 371334
rect 117674 335334 118294 370778
rect 117674 334778 117706 335334
rect 118262 334778 118294 335334
rect 117674 299334 118294 334778
rect 117674 298778 117706 299334
rect 118262 298778 118294 299334
rect 117674 263334 118294 298778
rect 117674 262778 117706 263334
rect 118262 262778 118294 263334
rect 117674 227334 118294 262778
rect 117674 226778 117706 227334
rect 118262 226778 118294 227334
rect 117674 191334 118294 226778
rect 117674 190778 117706 191334
rect 118262 190778 118294 191334
rect 117674 155334 118294 190778
rect 117674 154778 117706 155334
rect 118262 154778 118294 155334
rect 117674 119334 118294 154778
rect 117674 118778 117706 119334
rect 118262 118778 118294 119334
rect 117674 83334 118294 118778
rect 117674 82778 117706 83334
rect 118262 82778 118294 83334
rect 117674 47334 118294 82778
rect 117674 46778 117706 47334
rect 118262 46778 118294 47334
rect 117674 11334 118294 46778
rect 117674 10778 117706 11334
rect 118262 10778 118294 11334
rect 117674 -7066 118294 10778
rect 117674 -7622 117706 -7066
rect 118262 -7622 118294 -7066
rect 117674 -7654 118294 -7622
rect 144994 704838 145614 711590
rect 144994 704282 145026 704838
rect 145582 704282 145614 704838
rect 144994 686654 145614 704282
rect 144994 686098 145026 686654
rect 145582 686098 145614 686654
rect 144994 650654 145614 686098
rect 144994 650098 145026 650654
rect 145582 650098 145614 650654
rect 144994 614654 145614 650098
rect 144994 614098 145026 614654
rect 145582 614098 145614 614654
rect 144994 578654 145614 614098
rect 144994 578098 145026 578654
rect 145582 578098 145614 578654
rect 144994 542654 145614 578098
rect 144994 542098 145026 542654
rect 145582 542098 145614 542654
rect 144994 506654 145614 542098
rect 144994 506098 145026 506654
rect 145582 506098 145614 506654
rect 144994 470654 145614 506098
rect 144994 470098 145026 470654
rect 145582 470098 145614 470654
rect 144994 434654 145614 470098
rect 144994 434098 145026 434654
rect 145582 434098 145614 434654
rect 144994 398654 145614 434098
rect 144994 398098 145026 398654
rect 145582 398098 145614 398654
rect 144994 362654 145614 398098
rect 144994 362098 145026 362654
rect 145582 362098 145614 362654
rect 144994 326654 145614 362098
rect 144994 326098 145026 326654
rect 145582 326098 145614 326654
rect 144994 290654 145614 326098
rect 144994 290098 145026 290654
rect 145582 290098 145614 290654
rect 144994 254654 145614 290098
rect 144994 254098 145026 254654
rect 145582 254098 145614 254654
rect 144994 218654 145614 254098
rect 144994 218098 145026 218654
rect 145582 218098 145614 218654
rect 144994 182654 145614 218098
rect 144994 182098 145026 182654
rect 145582 182098 145614 182654
rect 144994 146654 145614 182098
rect 144994 146098 145026 146654
rect 145582 146098 145614 146654
rect 144994 110654 145614 146098
rect 144994 110098 145026 110654
rect 145582 110098 145614 110654
rect 144994 74654 145614 110098
rect 144994 74098 145026 74654
rect 145582 74098 145614 74654
rect 144994 38654 145614 74098
rect 144994 38098 145026 38654
rect 145582 38098 145614 38654
rect 144994 2654 145614 38098
rect 144994 2098 145026 2654
rect 145582 2098 145614 2654
rect 144994 -346 145614 2098
rect 144994 -902 145026 -346
rect 145582 -902 145614 -346
rect 144994 -7654 145614 -902
rect 146234 705798 146854 711590
rect 146234 705242 146266 705798
rect 146822 705242 146854 705798
rect 146234 687894 146854 705242
rect 146234 687338 146266 687894
rect 146822 687338 146854 687894
rect 146234 651894 146854 687338
rect 146234 651338 146266 651894
rect 146822 651338 146854 651894
rect 146234 615894 146854 651338
rect 146234 615338 146266 615894
rect 146822 615338 146854 615894
rect 146234 579894 146854 615338
rect 146234 579338 146266 579894
rect 146822 579338 146854 579894
rect 146234 543894 146854 579338
rect 146234 543338 146266 543894
rect 146822 543338 146854 543894
rect 146234 507894 146854 543338
rect 146234 507338 146266 507894
rect 146822 507338 146854 507894
rect 146234 471894 146854 507338
rect 146234 471338 146266 471894
rect 146822 471338 146854 471894
rect 146234 435894 146854 471338
rect 146234 435338 146266 435894
rect 146822 435338 146854 435894
rect 146234 399894 146854 435338
rect 146234 399338 146266 399894
rect 146822 399338 146854 399894
rect 146234 363894 146854 399338
rect 146234 363338 146266 363894
rect 146822 363338 146854 363894
rect 146234 327894 146854 363338
rect 146234 327338 146266 327894
rect 146822 327338 146854 327894
rect 146234 291894 146854 327338
rect 146234 291338 146266 291894
rect 146822 291338 146854 291894
rect 146234 255894 146854 291338
rect 146234 255338 146266 255894
rect 146822 255338 146854 255894
rect 146234 219894 146854 255338
rect 146234 219338 146266 219894
rect 146822 219338 146854 219894
rect 146234 183894 146854 219338
rect 146234 183338 146266 183894
rect 146822 183338 146854 183894
rect 146234 147894 146854 183338
rect 146234 147338 146266 147894
rect 146822 147338 146854 147894
rect 146234 111894 146854 147338
rect 146234 111338 146266 111894
rect 146822 111338 146854 111894
rect 146234 75894 146854 111338
rect 146234 75338 146266 75894
rect 146822 75338 146854 75894
rect 146234 39894 146854 75338
rect 146234 39338 146266 39894
rect 146822 39338 146854 39894
rect 146234 3894 146854 39338
rect 146234 3338 146266 3894
rect 146822 3338 146854 3894
rect 146234 -1306 146854 3338
rect 146234 -1862 146266 -1306
rect 146822 -1862 146854 -1306
rect 146234 -7654 146854 -1862
rect 147474 706758 148094 711590
rect 147474 706202 147506 706758
rect 148062 706202 148094 706758
rect 147474 689134 148094 706202
rect 147474 688578 147506 689134
rect 148062 688578 148094 689134
rect 147474 653134 148094 688578
rect 147474 652578 147506 653134
rect 148062 652578 148094 653134
rect 147474 617134 148094 652578
rect 147474 616578 147506 617134
rect 148062 616578 148094 617134
rect 147474 581134 148094 616578
rect 147474 580578 147506 581134
rect 148062 580578 148094 581134
rect 147474 545134 148094 580578
rect 147474 544578 147506 545134
rect 148062 544578 148094 545134
rect 147474 509134 148094 544578
rect 147474 508578 147506 509134
rect 148062 508578 148094 509134
rect 147474 473134 148094 508578
rect 147474 472578 147506 473134
rect 148062 472578 148094 473134
rect 147474 437134 148094 472578
rect 147474 436578 147506 437134
rect 148062 436578 148094 437134
rect 147474 401134 148094 436578
rect 147474 400578 147506 401134
rect 148062 400578 148094 401134
rect 147474 365134 148094 400578
rect 147474 364578 147506 365134
rect 148062 364578 148094 365134
rect 147474 329134 148094 364578
rect 147474 328578 147506 329134
rect 148062 328578 148094 329134
rect 147474 293134 148094 328578
rect 147474 292578 147506 293134
rect 148062 292578 148094 293134
rect 147474 257134 148094 292578
rect 147474 256578 147506 257134
rect 148062 256578 148094 257134
rect 147474 221134 148094 256578
rect 147474 220578 147506 221134
rect 148062 220578 148094 221134
rect 147474 185134 148094 220578
rect 147474 184578 147506 185134
rect 148062 184578 148094 185134
rect 147474 149134 148094 184578
rect 147474 148578 147506 149134
rect 148062 148578 148094 149134
rect 147474 113134 148094 148578
rect 147474 112578 147506 113134
rect 148062 112578 148094 113134
rect 147474 77134 148094 112578
rect 147474 76578 147506 77134
rect 148062 76578 148094 77134
rect 147474 41134 148094 76578
rect 147474 40578 147506 41134
rect 148062 40578 148094 41134
rect 147474 5134 148094 40578
rect 147474 4578 147506 5134
rect 148062 4578 148094 5134
rect 147474 -2266 148094 4578
rect 147474 -2822 147506 -2266
rect 148062 -2822 148094 -2266
rect 147474 -7654 148094 -2822
rect 148714 707718 149334 711590
rect 148714 707162 148746 707718
rect 149302 707162 149334 707718
rect 148714 690374 149334 707162
rect 148714 689818 148746 690374
rect 149302 689818 149334 690374
rect 148714 654374 149334 689818
rect 148714 653818 148746 654374
rect 149302 653818 149334 654374
rect 148714 618374 149334 653818
rect 148714 617818 148746 618374
rect 149302 617818 149334 618374
rect 148714 582374 149334 617818
rect 148714 581818 148746 582374
rect 149302 581818 149334 582374
rect 148714 546374 149334 581818
rect 148714 545818 148746 546374
rect 149302 545818 149334 546374
rect 148714 510374 149334 545818
rect 148714 509818 148746 510374
rect 149302 509818 149334 510374
rect 148714 474374 149334 509818
rect 148714 473818 148746 474374
rect 149302 473818 149334 474374
rect 148714 438374 149334 473818
rect 148714 437818 148746 438374
rect 149302 437818 149334 438374
rect 148714 402374 149334 437818
rect 148714 401818 148746 402374
rect 149302 401818 149334 402374
rect 148714 366374 149334 401818
rect 148714 365818 148746 366374
rect 149302 365818 149334 366374
rect 148714 330374 149334 365818
rect 148714 329818 148746 330374
rect 149302 329818 149334 330374
rect 148714 294374 149334 329818
rect 148714 293818 148746 294374
rect 149302 293818 149334 294374
rect 148714 258374 149334 293818
rect 148714 257818 148746 258374
rect 149302 257818 149334 258374
rect 148714 222374 149334 257818
rect 148714 221818 148746 222374
rect 149302 221818 149334 222374
rect 148714 186374 149334 221818
rect 148714 185818 148746 186374
rect 149302 185818 149334 186374
rect 148714 150374 149334 185818
rect 148714 149818 148746 150374
rect 149302 149818 149334 150374
rect 148714 114374 149334 149818
rect 148714 113818 148746 114374
rect 149302 113818 149334 114374
rect 148714 78374 149334 113818
rect 148714 77818 148746 78374
rect 149302 77818 149334 78374
rect 148714 42374 149334 77818
rect 148714 41818 148746 42374
rect 149302 41818 149334 42374
rect 148714 6374 149334 41818
rect 148714 5818 148746 6374
rect 149302 5818 149334 6374
rect 148714 -3226 149334 5818
rect 148714 -3782 148746 -3226
rect 149302 -3782 149334 -3226
rect 148714 -7654 149334 -3782
rect 149954 708678 150574 711590
rect 149954 708122 149986 708678
rect 150542 708122 150574 708678
rect 149954 691614 150574 708122
rect 149954 691058 149986 691614
rect 150542 691058 150574 691614
rect 149954 655614 150574 691058
rect 149954 655058 149986 655614
rect 150542 655058 150574 655614
rect 149954 619614 150574 655058
rect 149954 619058 149986 619614
rect 150542 619058 150574 619614
rect 149954 583614 150574 619058
rect 149954 583058 149986 583614
rect 150542 583058 150574 583614
rect 149954 547614 150574 583058
rect 149954 547058 149986 547614
rect 150542 547058 150574 547614
rect 149954 511614 150574 547058
rect 149954 511058 149986 511614
rect 150542 511058 150574 511614
rect 149954 475614 150574 511058
rect 149954 475058 149986 475614
rect 150542 475058 150574 475614
rect 149954 439614 150574 475058
rect 149954 439058 149986 439614
rect 150542 439058 150574 439614
rect 149954 403614 150574 439058
rect 149954 403058 149986 403614
rect 150542 403058 150574 403614
rect 149954 367614 150574 403058
rect 149954 367058 149986 367614
rect 150542 367058 150574 367614
rect 149954 331614 150574 367058
rect 149954 331058 149986 331614
rect 150542 331058 150574 331614
rect 149954 295614 150574 331058
rect 149954 295058 149986 295614
rect 150542 295058 150574 295614
rect 149954 259614 150574 295058
rect 149954 259058 149986 259614
rect 150542 259058 150574 259614
rect 149954 223614 150574 259058
rect 149954 223058 149986 223614
rect 150542 223058 150574 223614
rect 149954 187614 150574 223058
rect 149954 187058 149986 187614
rect 150542 187058 150574 187614
rect 149954 151614 150574 187058
rect 149954 151058 149986 151614
rect 150542 151058 150574 151614
rect 149954 115614 150574 151058
rect 149954 115058 149986 115614
rect 150542 115058 150574 115614
rect 149954 79614 150574 115058
rect 149954 79058 149986 79614
rect 150542 79058 150574 79614
rect 149954 43614 150574 79058
rect 149954 43058 149986 43614
rect 150542 43058 150574 43614
rect 149954 7614 150574 43058
rect 149954 7058 149986 7614
rect 150542 7058 150574 7614
rect 149954 -4186 150574 7058
rect 149954 -4742 149986 -4186
rect 150542 -4742 150574 -4186
rect 149954 -7654 150574 -4742
rect 151194 709638 151814 711590
rect 151194 709082 151226 709638
rect 151782 709082 151814 709638
rect 151194 692854 151814 709082
rect 151194 692298 151226 692854
rect 151782 692298 151814 692854
rect 151194 656854 151814 692298
rect 151194 656298 151226 656854
rect 151782 656298 151814 656854
rect 151194 620854 151814 656298
rect 151194 620298 151226 620854
rect 151782 620298 151814 620854
rect 151194 584854 151814 620298
rect 151194 584298 151226 584854
rect 151782 584298 151814 584854
rect 151194 548854 151814 584298
rect 151194 548298 151226 548854
rect 151782 548298 151814 548854
rect 151194 512854 151814 548298
rect 151194 512298 151226 512854
rect 151782 512298 151814 512854
rect 151194 476854 151814 512298
rect 151194 476298 151226 476854
rect 151782 476298 151814 476854
rect 151194 440854 151814 476298
rect 151194 440298 151226 440854
rect 151782 440298 151814 440854
rect 151194 404854 151814 440298
rect 151194 404298 151226 404854
rect 151782 404298 151814 404854
rect 151194 368854 151814 404298
rect 151194 368298 151226 368854
rect 151782 368298 151814 368854
rect 151194 332854 151814 368298
rect 151194 332298 151226 332854
rect 151782 332298 151814 332854
rect 151194 296854 151814 332298
rect 151194 296298 151226 296854
rect 151782 296298 151814 296854
rect 151194 260854 151814 296298
rect 151194 260298 151226 260854
rect 151782 260298 151814 260854
rect 151194 224854 151814 260298
rect 151194 224298 151226 224854
rect 151782 224298 151814 224854
rect 151194 188854 151814 224298
rect 151194 188298 151226 188854
rect 151782 188298 151814 188854
rect 151194 152854 151814 188298
rect 151194 152298 151226 152854
rect 151782 152298 151814 152854
rect 151194 116854 151814 152298
rect 151194 116298 151226 116854
rect 151782 116298 151814 116854
rect 151194 80854 151814 116298
rect 151194 80298 151226 80854
rect 151782 80298 151814 80854
rect 151194 44854 151814 80298
rect 151194 44298 151226 44854
rect 151782 44298 151814 44854
rect 151194 8854 151814 44298
rect 151194 8298 151226 8854
rect 151782 8298 151814 8854
rect 151194 -5146 151814 8298
rect 151194 -5702 151226 -5146
rect 151782 -5702 151814 -5146
rect 151194 -7654 151814 -5702
rect 152434 710598 153054 711590
rect 152434 710042 152466 710598
rect 153022 710042 153054 710598
rect 152434 694094 153054 710042
rect 152434 693538 152466 694094
rect 153022 693538 153054 694094
rect 152434 658094 153054 693538
rect 152434 657538 152466 658094
rect 153022 657538 153054 658094
rect 152434 622094 153054 657538
rect 152434 621538 152466 622094
rect 153022 621538 153054 622094
rect 152434 586094 153054 621538
rect 152434 585538 152466 586094
rect 153022 585538 153054 586094
rect 152434 550094 153054 585538
rect 152434 549538 152466 550094
rect 153022 549538 153054 550094
rect 152434 514094 153054 549538
rect 152434 513538 152466 514094
rect 153022 513538 153054 514094
rect 152434 478094 153054 513538
rect 152434 477538 152466 478094
rect 153022 477538 153054 478094
rect 152434 442094 153054 477538
rect 152434 441538 152466 442094
rect 153022 441538 153054 442094
rect 152434 406094 153054 441538
rect 152434 405538 152466 406094
rect 153022 405538 153054 406094
rect 152434 370094 153054 405538
rect 152434 369538 152466 370094
rect 153022 369538 153054 370094
rect 152434 334094 153054 369538
rect 152434 333538 152466 334094
rect 153022 333538 153054 334094
rect 152434 298094 153054 333538
rect 152434 297538 152466 298094
rect 153022 297538 153054 298094
rect 152434 262094 153054 297538
rect 152434 261538 152466 262094
rect 153022 261538 153054 262094
rect 152434 226094 153054 261538
rect 152434 225538 152466 226094
rect 153022 225538 153054 226094
rect 152434 190094 153054 225538
rect 152434 189538 152466 190094
rect 153022 189538 153054 190094
rect 152434 154094 153054 189538
rect 152434 153538 152466 154094
rect 153022 153538 153054 154094
rect 152434 118094 153054 153538
rect 152434 117538 152466 118094
rect 153022 117538 153054 118094
rect 152434 82094 153054 117538
rect 152434 81538 152466 82094
rect 153022 81538 153054 82094
rect 152434 46094 153054 81538
rect 152434 45538 152466 46094
rect 153022 45538 153054 46094
rect 152434 10094 153054 45538
rect 152434 9538 152466 10094
rect 153022 9538 153054 10094
rect 152434 -6106 153054 9538
rect 152434 -6662 152466 -6106
rect 153022 -6662 153054 -6106
rect 152434 -7654 153054 -6662
rect 153674 711558 154294 711590
rect 153674 711002 153706 711558
rect 154262 711002 154294 711558
rect 153674 695334 154294 711002
rect 153674 694778 153706 695334
rect 154262 694778 154294 695334
rect 153674 659334 154294 694778
rect 153674 658778 153706 659334
rect 154262 658778 154294 659334
rect 153674 623334 154294 658778
rect 153674 622778 153706 623334
rect 154262 622778 154294 623334
rect 153674 587334 154294 622778
rect 153674 586778 153706 587334
rect 154262 586778 154294 587334
rect 153674 551334 154294 586778
rect 153674 550778 153706 551334
rect 154262 550778 154294 551334
rect 153674 515334 154294 550778
rect 153674 514778 153706 515334
rect 154262 514778 154294 515334
rect 153674 479334 154294 514778
rect 153674 478778 153706 479334
rect 154262 478778 154294 479334
rect 153674 443334 154294 478778
rect 153674 442778 153706 443334
rect 154262 442778 154294 443334
rect 153674 407334 154294 442778
rect 153674 406778 153706 407334
rect 154262 406778 154294 407334
rect 153674 371334 154294 406778
rect 153674 370778 153706 371334
rect 154262 370778 154294 371334
rect 153674 335334 154294 370778
rect 153674 334778 153706 335334
rect 154262 334778 154294 335334
rect 153674 299334 154294 334778
rect 153674 298778 153706 299334
rect 154262 298778 154294 299334
rect 153674 263334 154294 298778
rect 153674 262778 153706 263334
rect 154262 262778 154294 263334
rect 153674 227334 154294 262778
rect 153674 226778 153706 227334
rect 154262 226778 154294 227334
rect 153674 191334 154294 226778
rect 153674 190778 153706 191334
rect 154262 190778 154294 191334
rect 153674 155334 154294 190778
rect 153674 154778 153706 155334
rect 154262 154778 154294 155334
rect 153674 119334 154294 154778
rect 153674 118778 153706 119334
rect 154262 118778 154294 119334
rect 153674 83334 154294 118778
rect 153674 82778 153706 83334
rect 154262 82778 154294 83334
rect 153674 47334 154294 82778
rect 153674 46778 153706 47334
rect 154262 46778 154294 47334
rect 153674 11334 154294 46778
rect 153674 10778 153706 11334
rect 154262 10778 154294 11334
rect 153674 -7066 154294 10778
rect 153674 -7622 153706 -7066
rect 154262 -7622 154294 -7066
rect 153674 -7654 154294 -7622
rect 180994 704838 181614 711590
rect 180994 704282 181026 704838
rect 181582 704282 181614 704838
rect 180994 686654 181614 704282
rect 180994 686098 181026 686654
rect 181582 686098 181614 686654
rect 180994 650654 181614 686098
rect 180994 650098 181026 650654
rect 181582 650098 181614 650654
rect 180994 614654 181614 650098
rect 180994 614098 181026 614654
rect 181582 614098 181614 614654
rect 180994 578654 181614 614098
rect 180994 578098 181026 578654
rect 181582 578098 181614 578654
rect 180994 542654 181614 578098
rect 180994 542098 181026 542654
rect 181582 542098 181614 542654
rect 180994 506654 181614 542098
rect 180994 506098 181026 506654
rect 181582 506098 181614 506654
rect 180994 470654 181614 506098
rect 180994 470098 181026 470654
rect 181582 470098 181614 470654
rect 180994 434654 181614 470098
rect 180994 434098 181026 434654
rect 181582 434098 181614 434654
rect 180994 398654 181614 434098
rect 180994 398098 181026 398654
rect 181582 398098 181614 398654
rect 180994 362654 181614 398098
rect 180994 362098 181026 362654
rect 181582 362098 181614 362654
rect 180994 326654 181614 362098
rect 180994 326098 181026 326654
rect 181582 326098 181614 326654
rect 180994 290654 181614 326098
rect 180994 290098 181026 290654
rect 181582 290098 181614 290654
rect 180994 254654 181614 290098
rect 180994 254098 181026 254654
rect 181582 254098 181614 254654
rect 180994 218654 181614 254098
rect 180994 218098 181026 218654
rect 181582 218098 181614 218654
rect 180994 182654 181614 218098
rect 180994 182098 181026 182654
rect 181582 182098 181614 182654
rect 180994 146654 181614 182098
rect 180994 146098 181026 146654
rect 181582 146098 181614 146654
rect 180994 110654 181614 146098
rect 180994 110098 181026 110654
rect 181582 110098 181614 110654
rect 180994 74654 181614 110098
rect 180994 74098 181026 74654
rect 181582 74098 181614 74654
rect 180994 38654 181614 74098
rect 180994 38098 181026 38654
rect 181582 38098 181614 38654
rect 180994 2654 181614 38098
rect 180994 2098 181026 2654
rect 181582 2098 181614 2654
rect 180994 -346 181614 2098
rect 180994 -902 181026 -346
rect 181582 -902 181614 -346
rect 180994 -7654 181614 -902
rect 182234 705798 182854 711590
rect 182234 705242 182266 705798
rect 182822 705242 182854 705798
rect 182234 687894 182854 705242
rect 182234 687338 182266 687894
rect 182822 687338 182854 687894
rect 182234 651894 182854 687338
rect 182234 651338 182266 651894
rect 182822 651338 182854 651894
rect 182234 615894 182854 651338
rect 182234 615338 182266 615894
rect 182822 615338 182854 615894
rect 182234 579894 182854 615338
rect 182234 579338 182266 579894
rect 182822 579338 182854 579894
rect 182234 543894 182854 579338
rect 182234 543338 182266 543894
rect 182822 543338 182854 543894
rect 182234 507894 182854 543338
rect 182234 507338 182266 507894
rect 182822 507338 182854 507894
rect 182234 471894 182854 507338
rect 182234 471338 182266 471894
rect 182822 471338 182854 471894
rect 182234 435894 182854 471338
rect 182234 435338 182266 435894
rect 182822 435338 182854 435894
rect 182234 399894 182854 435338
rect 182234 399338 182266 399894
rect 182822 399338 182854 399894
rect 182234 363894 182854 399338
rect 182234 363338 182266 363894
rect 182822 363338 182854 363894
rect 182234 327894 182854 363338
rect 182234 327338 182266 327894
rect 182822 327338 182854 327894
rect 182234 291894 182854 327338
rect 182234 291338 182266 291894
rect 182822 291338 182854 291894
rect 182234 255894 182854 291338
rect 182234 255338 182266 255894
rect 182822 255338 182854 255894
rect 182234 219894 182854 255338
rect 182234 219338 182266 219894
rect 182822 219338 182854 219894
rect 182234 183894 182854 219338
rect 182234 183338 182266 183894
rect 182822 183338 182854 183894
rect 182234 147894 182854 183338
rect 182234 147338 182266 147894
rect 182822 147338 182854 147894
rect 182234 111894 182854 147338
rect 182234 111338 182266 111894
rect 182822 111338 182854 111894
rect 182234 75894 182854 111338
rect 182234 75338 182266 75894
rect 182822 75338 182854 75894
rect 182234 39894 182854 75338
rect 182234 39338 182266 39894
rect 182822 39338 182854 39894
rect 182234 3894 182854 39338
rect 182234 3338 182266 3894
rect 182822 3338 182854 3894
rect 182234 -1306 182854 3338
rect 182234 -1862 182266 -1306
rect 182822 -1862 182854 -1306
rect 182234 -7654 182854 -1862
rect 183474 706758 184094 711590
rect 183474 706202 183506 706758
rect 184062 706202 184094 706758
rect 183474 689134 184094 706202
rect 183474 688578 183506 689134
rect 184062 688578 184094 689134
rect 183474 653134 184094 688578
rect 183474 652578 183506 653134
rect 184062 652578 184094 653134
rect 183474 617134 184094 652578
rect 183474 616578 183506 617134
rect 184062 616578 184094 617134
rect 183474 581134 184094 616578
rect 183474 580578 183506 581134
rect 184062 580578 184094 581134
rect 183474 545134 184094 580578
rect 183474 544578 183506 545134
rect 184062 544578 184094 545134
rect 183474 509134 184094 544578
rect 183474 508578 183506 509134
rect 184062 508578 184094 509134
rect 183474 473134 184094 508578
rect 183474 472578 183506 473134
rect 184062 472578 184094 473134
rect 183474 437134 184094 472578
rect 183474 436578 183506 437134
rect 184062 436578 184094 437134
rect 183474 401134 184094 436578
rect 183474 400578 183506 401134
rect 184062 400578 184094 401134
rect 183474 365134 184094 400578
rect 183474 364578 183506 365134
rect 184062 364578 184094 365134
rect 183474 329134 184094 364578
rect 183474 328578 183506 329134
rect 184062 328578 184094 329134
rect 183474 293134 184094 328578
rect 183474 292578 183506 293134
rect 184062 292578 184094 293134
rect 183474 257134 184094 292578
rect 183474 256578 183506 257134
rect 184062 256578 184094 257134
rect 183474 221134 184094 256578
rect 183474 220578 183506 221134
rect 184062 220578 184094 221134
rect 183474 185134 184094 220578
rect 183474 184578 183506 185134
rect 184062 184578 184094 185134
rect 183474 149134 184094 184578
rect 183474 148578 183506 149134
rect 184062 148578 184094 149134
rect 183474 113134 184094 148578
rect 183474 112578 183506 113134
rect 184062 112578 184094 113134
rect 183474 77134 184094 112578
rect 183474 76578 183506 77134
rect 184062 76578 184094 77134
rect 183474 41134 184094 76578
rect 183474 40578 183506 41134
rect 184062 40578 184094 41134
rect 183474 5134 184094 40578
rect 183474 4578 183506 5134
rect 184062 4578 184094 5134
rect 183474 -2266 184094 4578
rect 183474 -2822 183506 -2266
rect 184062 -2822 184094 -2266
rect 183474 -7654 184094 -2822
rect 184714 707718 185334 711590
rect 184714 707162 184746 707718
rect 185302 707162 185334 707718
rect 184714 690374 185334 707162
rect 184714 689818 184746 690374
rect 185302 689818 185334 690374
rect 184714 654374 185334 689818
rect 184714 653818 184746 654374
rect 185302 653818 185334 654374
rect 184714 618374 185334 653818
rect 184714 617818 184746 618374
rect 185302 617818 185334 618374
rect 184714 582374 185334 617818
rect 184714 581818 184746 582374
rect 185302 581818 185334 582374
rect 184714 546374 185334 581818
rect 184714 545818 184746 546374
rect 185302 545818 185334 546374
rect 184714 510374 185334 545818
rect 184714 509818 184746 510374
rect 185302 509818 185334 510374
rect 184714 474374 185334 509818
rect 184714 473818 184746 474374
rect 185302 473818 185334 474374
rect 184714 438374 185334 473818
rect 184714 437818 184746 438374
rect 185302 437818 185334 438374
rect 184714 402374 185334 437818
rect 184714 401818 184746 402374
rect 185302 401818 185334 402374
rect 184714 366374 185334 401818
rect 184714 365818 184746 366374
rect 185302 365818 185334 366374
rect 184714 330374 185334 365818
rect 184714 329818 184746 330374
rect 185302 329818 185334 330374
rect 184714 294374 185334 329818
rect 184714 293818 184746 294374
rect 185302 293818 185334 294374
rect 184714 258374 185334 293818
rect 184714 257818 184746 258374
rect 185302 257818 185334 258374
rect 184714 222374 185334 257818
rect 184714 221818 184746 222374
rect 185302 221818 185334 222374
rect 184714 186374 185334 221818
rect 184714 185818 184746 186374
rect 185302 185818 185334 186374
rect 184714 150374 185334 185818
rect 184714 149818 184746 150374
rect 185302 149818 185334 150374
rect 184714 114374 185334 149818
rect 184714 113818 184746 114374
rect 185302 113818 185334 114374
rect 184714 78374 185334 113818
rect 184714 77818 184746 78374
rect 185302 77818 185334 78374
rect 184714 42374 185334 77818
rect 184714 41818 184746 42374
rect 185302 41818 185334 42374
rect 184714 6374 185334 41818
rect 184714 5818 184746 6374
rect 185302 5818 185334 6374
rect 184714 -3226 185334 5818
rect 184714 -3782 184746 -3226
rect 185302 -3782 185334 -3226
rect 184714 -7654 185334 -3782
rect 185954 708678 186574 711590
rect 185954 708122 185986 708678
rect 186542 708122 186574 708678
rect 185954 691614 186574 708122
rect 185954 691058 185986 691614
rect 186542 691058 186574 691614
rect 185954 655614 186574 691058
rect 185954 655058 185986 655614
rect 186542 655058 186574 655614
rect 185954 619614 186574 655058
rect 185954 619058 185986 619614
rect 186542 619058 186574 619614
rect 185954 583614 186574 619058
rect 185954 583058 185986 583614
rect 186542 583058 186574 583614
rect 185954 547614 186574 583058
rect 185954 547058 185986 547614
rect 186542 547058 186574 547614
rect 185954 511614 186574 547058
rect 185954 511058 185986 511614
rect 186542 511058 186574 511614
rect 185954 475614 186574 511058
rect 185954 475058 185986 475614
rect 186542 475058 186574 475614
rect 185954 439614 186574 475058
rect 185954 439058 185986 439614
rect 186542 439058 186574 439614
rect 185954 403614 186574 439058
rect 185954 403058 185986 403614
rect 186542 403058 186574 403614
rect 185954 367614 186574 403058
rect 185954 367058 185986 367614
rect 186542 367058 186574 367614
rect 185954 331614 186574 367058
rect 185954 331058 185986 331614
rect 186542 331058 186574 331614
rect 185954 295614 186574 331058
rect 185954 295058 185986 295614
rect 186542 295058 186574 295614
rect 185954 259614 186574 295058
rect 185954 259058 185986 259614
rect 186542 259058 186574 259614
rect 185954 223614 186574 259058
rect 185954 223058 185986 223614
rect 186542 223058 186574 223614
rect 185954 187614 186574 223058
rect 185954 187058 185986 187614
rect 186542 187058 186574 187614
rect 185954 151614 186574 187058
rect 185954 151058 185986 151614
rect 186542 151058 186574 151614
rect 185954 115614 186574 151058
rect 185954 115058 185986 115614
rect 186542 115058 186574 115614
rect 185954 79614 186574 115058
rect 185954 79058 185986 79614
rect 186542 79058 186574 79614
rect 185954 43614 186574 79058
rect 185954 43058 185986 43614
rect 186542 43058 186574 43614
rect 185954 7614 186574 43058
rect 185954 7058 185986 7614
rect 186542 7058 186574 7614
rect 185954 -4186 186574 7058
rect 185954 -4742 185986 -4186
rect 186542 -4742 186574 -4186
rect 185954 -7654 186574 -4742
rect 187194 709638 187814 711590
rect 187194 709082 187226 709638
rect 187782 709082 187814 709638
rect 187194 692854 187814 709082
rect 187194 692298 187226 692854
rect 187782 692298 187814 692854
rect 187194 656854 187814 692298
rect 187194 656298 187226 656854
rect 187782 656298 187814 656854
rect 187194 620854 187814 656298
rect 187194 620298 187226 620854
rect 187782 620298 187814 620854
rect 187194 584854 187814 620298
rect 187194 584298 187226 584854
rect 187782 584298 187814 584854
rect 187194 548854 187814 584298
rect 187194 548298 187226 548854
rect 187782 548298 187814 548854
rect 187194 512854 187814 548298
rect 187194 512298 187226 512854
rect 187782 512298 187814 512854
rect 187194 476854 187814 512298
rect 187194 476298 187226 476854
rect 187782 476298 187814 476854
rect 187194 440854 187814 476298
rect 187194 440298 187226 440854
rect 187782 440298 187814 440854
rect 187194 404854 187814 440298
rect 187194 404298 187226 404854
rect 187782 404298 187814 404854
rect 187194 368854 187814 404298
rect 187194 368298 187226 368854
rect 187782 368298 187814 368854
rect 187194 332854 187814 368298
rect 187194 332298 187226 332854
rect 187782 332298 187814 332854
rect 187194 296854 187814 332298
rect 187194 296298 187226 296854
rect 187782 296298 187814 296854
rect 187194 260854 187814 296298
rect 187194 260298 187226 260854
rect 187782 260298 187814 260854
rect 187194 224854 187814 260298
rect 187194 224298 187226 224854
rect 187782 224298 187814 224854
rect 187194 188854 187814 224298
rect 187194 188298 187226 188854
rect 187782 188298 187814 188854
rect 187194 152854 187814 188298
rect 187194 152298 187226 152854
rect 187782 152298 187814 152854
rect 187194 116854 187814 152298
rect 187194 116298 187226 116854
rect 187782 116298 187814 116854
rect 187194 80854 187814 116298
rect 187194 80298 187226 80854
rect 187782 80298 187814 80854
rect 187194 44854 187814 80298
rect 187194 44298 187226 44854
rect 187782 44298 187814 44854
rect 187194 8854 187814 44298
rect 187194 8298 187226 8854
rect 187782 8298 187814 8854
rect 187194 -5146 187814 8298
rect 187194 -5702 187226 -5146
rect 187782 -5702 187814 -5146
rect 187194 -7654 187814 -5702
rect 188434 710598 189054 711590
rect 188434 710042 188466 710598
rect 189022 710042 189054 710598
rect 188434 694094 189054 710042
rect 188434 693538 188466 694094
rect 189022 693538 189054 694094
rect 188434 658094 189054 693538
rect 188434 657538 188466 658094
rect 189022 657538 189054 658094
rect 188434 622094 189054 657538
rect 188434 621538 188466 622094
rect 189022 621538 189054 622094
rect 188434 586094 189054 621538
rect 188434 585538 188466 586094
rect 189022 585538 189054 586094
rect 188434 550094 189054 585538
rect 188434 549538 188466 550094
rect 189022 549538 189054 550094
rect 188434 514094 189054 549538
rect 188434 513538 188466 514094
rect 189022 513538 189054 514094
rect 188434 478094 189054 513538
rect 188434 477538 188466 478094
rect 189022 477538 189054 478094
rect 188434 442094 189054 477538
rect 188434 441538 188466 442094
rect 189022 441538 189054 442094
rect 188434 406094 189054 441538
rect 188434 405538 188466 406094
rect 189022 405538 189054 406094
rect 188434 370094 189054 405538
rect 188434 369538 188466 370094
rect 189022 369538 189054 370094
rect 188434 334094 189054 369538
rect 188434 333538 188466 334094
rect 189022 333538 189054 334094
rect 188434 298094 189054 333538
rect 188434 297538 188466 298094
rect 189022 297538 189054 298094
rect 188434 262094 189054 297538
rect 188434 261538 188466 262094
rect 189022 261538 189054 262094
rect 188434 226094 189054 261538
rect 188434 225538 188466 226094
rect 189022 225538 189054 226094
rect 188434 190094 189054 225538
rect 188434 189538 188466 190094
rect 189022 189538 189054 190094
rect 188434 154094 189054 189538
rect 188434 153538 188466 154094
rect 189022 153538 189054 154094
rect 188434 118094 189054 153538
rect 188434 117538 188466 118094
rect 189022 117538 189054 118094
rect 188434 82094 189054 117538
rect 188434 81538 188466 82094
rect 189022 81538 189054 82094
rect 188434 46094 189054 81538
rect 188434 45538 188466 46094
rect 189022 45538 189054 46094
rect 188434 10094 189054 45538
rect 188434 9538 188466 10094
rect 189022 9538 189054 10094
rect 188434 -6106 189054 9538
rect 188434 -6662 188466 -6106
rect 189022 -6662 189054 -6106
rect 188434 -7654 189054 -6662
rect 189674 711558 190294 711590
rect 189674 711002 189706 711558
rect 190262 711002 190294 711558
rect 189674 695334 190294 711002
rect 189674 694778 189706 695334
rect 190262 694778 190294 695334
rect 189674 659334 190294 694778
rect 189674 658778 189706 659334
rect 190262 658778 190294 659334
rect 189674 623334 190294 658778
rect 189674 622778 189706 623334
rect 190262 622778 190294 623334
rect 189674 587334 190294 622778
rect 189674 586778 189706 587334
rect 190262 586778 190294 587334
rect 189674 551334 190294 586778
rect 189674 550778 189706 551334
rect 190262 550778 190294 551334
rect 189674 515334 190294 550778
rect 189674 514778 189706 515334
rect 190262 514778 190294 515334
rect 189674 479334 190294 514778
rect 189674 478778 189706 479334
rect 190262 478778 190294 479334
rect 189674 443334 190294 478778
rect 189674 442778 189706 443334
rect 190262 442778 190294 443334
rect 189674 407334 190294 442778
rect 189674 406778 189706 407334
rect 190262 406778 190294 407334
rect 189674 371334 190294 406778
rect 189674 370778 189706 371334
rect 190262 370778 190294 371334
rect 189674 335334 190294 370778
rect 189674 334778 189706 335334
rect 190262 334778 190294 335334
rect 189674 299334 190294 334778
rect 189674 298778 189706 299334
rect 190262 298778 190294 299334
rect 189674 263334 190294 298778
rect 189674 262778 189706 263334
rect 190262 262778 190294 263334
rect 189674 227334 190294 262778
rect 189674 226778 189706 227334
rect 190262 226778 190294 227334
rect 189674 191334 190294 226778
rect 189674 190778 189706 191334
rect 190262 190778 190294 191334
rect 189674 155334 190294 190778
rect 189674 154778 189706 155334
rect 190262 154778 190294 155334
rect 189674 119334 190294 154778
rect 189674 118778 189706 119334
rect 190262 118778 190294 119334
rect 189674 83334 190294 118778
rect 189674 82778 189706 83334
rect 190262 82778 190294 83334
rect 189674 47334 190294 82778
rect 189674 46778 189706 47334
rect 190262 46778 190294 47334
rect 189674 11334 190294 46778
rect 189674 10778 189706 11334
rect 190262 10778 190294 11334
rect 189674 -7066 190294 10778
rect 189674 -7622 189706 -7066
rect 190262 -7622 190294 -7066
rect 189674 -7654 190294 -7622
rect 216994 704838 217614 711590
rect 216994 704282 217026 704838
rect 217582 704282 217614 704838
rect 216994 686654 217614 704282
rect 216994 686098 217026 686654
rect 217582 686098 217614 686654
rect 216994 650654 217614 686098
rect 216994 650098 217026 650654
rect 217582 650098 217614 650654
rect 216994 614654 217614 650098
rect 216994 614098 217026 614654
rect 217582 614098 217614 614654
rect 216994 578654 217614 614098
rect 216994 578098 217026 578654
rect 217582 578098 217614 578654
rect 216994 542654 217614 578098
rect 216994 542098 217026 542654
rect 217582 542098 217614 542654
rect 216994 506654 217614 542098
rect 216994 506098 217026 506654
rect 217582 506098 217614 506654
rect 216994 470654 217614 506098
rect 216994 470098 217026 470654
rect 217582 470098 217614 470654
rect 216994 434654 217614 470098
rect 216994 434098 217026 434654
rect 217582 434098 217614 434654
rect 216994 398654 217614 434098
rect 216994 398098 217026 398654
rect 217582 398098 217614 398654
rect 216994 362654 217614 398098
rect 216994 362098 217026 362654
rect 217582 362098 217614 362654
rect 216994 326654 217614 362098
rect 216994 326098 217026 326654
rect 217582 326098 217614 326654
rect 216994 290654 217614 326098
rect 216994 290098 217026 290654
rect 217582 290098 217614 290654
rect 216994 254654 217614 290098
rect 216994 254098 217026 254654
rect 217582 254098 217614 254654
rect 216994 218654 217614 254098
rect 216994 218098 217026 218654
rect 217582 218098 217614 218654
rect 216994 182654 217614 218098
rect 216994 182098 217026 182654
rect 217582 182098 217614 182654
rect 216994 146654 217614 182098
rect 216994 146098 217026 146654
rect 217582 146098 217614 146654
rect 216994 110654 217614 146098
rect 216994 110098 217026 110654
rect 217582 110098 217614 110654
rect 216994 74654 217614 110098
rect 216994 74098 217026 74654
rect 217582 74098 217614 74654
rect 216994 38654 217614 74098
rect 216994 38098 217026 38654
rect 217582 38098 217614 38654
rect 216994 2654 217614 38098
rect 216994 2098 217026 2654
rect 217582 2098 217614 2654
rect 216994 -346 217614 2098
rect 216994 -902 217026 -346
rect 217582 -902 217614 -346
rect 216994 -7654 217614 -902
rect 218234 705798 218854 711590
rect 218234 705242 218266 705798
rect 218822 705242 218854 705798
rect 218234 687894 218854 705242
rect 218234 687338 218266 687894
rect 218822 687338 218854 687894
rect 218234 651894 218854 687338
rect 218234 651338 218266 651894
rect 218822 651338 218854 651894
rect 218234 615894 218854 651338
rect 218234 615338 218266 615894
rect 218822 615338 218854 615894
rect 218234 579894 218854 615338
rect 218234 579338 218266 579894
rect 218822 579338 218854 579894
rect 218234 543894 218854 579338
rect 218234 543338 218266 543894
rect 218822 543338 218854 543894
rect 218234 507894 218854 543338
rect 218234 507338 218266 507894
rect 218822 507338 218854 507894
rect 218234 471894 218854 507338
rect 218234 471338 218266 471894
rect 218822 471338 218854 471894
rect 218234 435894 218854 471338
rect 218234 435338 218266 435894
rect 218822 435338 218854 435894
rect 218234 399894 218854 435338
rect 218234 399338 218266 399894
rect 218822 399338 218854 399894
rect 218234 363894 218854 399338
rect 218234 363338 218266 363894
rect 218822 363338 218854 363894
rect 218234 327894 218854 363338
rect 218234 327338 218266 327894
rect 218822 327338 218854 327894
rect 218234 291894 218854 327338
rect 218234 291338 218266 291894
rect 218822 291338 218854 291894
rect 218234 255894 218854 291338
rect 218234 255338 218266 255894
rect 218822 255338 218854 255894
rect 218234 219894 218854 255338
rect 218234 219338 218266 219894
rect 218822 219338 218854 219894
rect 218234 183894 218854 219338
rect 218234 183338 218266 183894
rect 218822 183338 218854 183894
rect 218234 147894 218854 183338
rect 218234 147338 218266 147894
rect 218822 147338 218854 147894
rect 218234 111894 218854 147338
rect 218234 111338 218266 111894
rect 218822 111338 218854 111894
rect 218234 75894 218854 111338
rect 218234 75338 218266 75894
rect 218822 75338 218854 75894
rect 218234 39894 218854 75338
rect 218234 39338 218266 39894
rect 218822 39338 218854 39894
rect 218234 3894 218854 39338
rect 218234 3338 218266 3894
rect 218822 3338 218854 3894
rect 218234 -1306 218854 3338
rect 218234 -1862 218266 -1306
rect 218822 -1862 218854 -1306
rect 218234 -7654 218854 -1862
rect 219474 706758 220094 711590
rect 219474 706202 219506 706758
rect 220062 706202 220094 706758
rect 219474 689134 220094 706202
rect 219474 688578 219506 689134
rect 220062 688578 220094 689134
rect 219474 653134 220094 688578
rect 219474 652578 219506 653134
rect 220062 652578 220094 653134
rect 219474 617134 220094 652578
rect 219474 616578 219506 617134
rect 220062 616578 220094 617134
rect 219474 581134 220094 616578
rect 219474 580578 219506 581134
rect 220062 580578 220094 581134
rect 219474 545134 220094 580578
rect 219474 544578 219506 545134
rect 220062 544578 220094 545134
rect 219474 509134 220094 544578
rect 219474 508578 219506 509134
rect 220062 508578 220094 509134
rect 219474 473134 220094 508578
rect 219474 472578 219506 473134
rect 220062 472578 220094 473134
rect 219474 437134 220094 472578
rect 219474 436578 219506 437134
rect 220062 436578 220094 437134
rect 219474 401134 220094 436578
rect 219474 400578 219506 401134
rect 220062 400578 220094 401134
rect 219474 365134 220094 400578
rect 219474 364578 219506 365134
rect 220062 364578 220094 365134
rect 219474 329134 220094 364578
rect 219474 328578 219506 329134
rect 220062 328578 220094 329134
rect 219474 293134 220094 328578
rect 219474 292578 219506 293134
rect 220062 292578 220094 293134
rect 219474 257134 220094 292578
rect 219474 256578 219506 257134
rect 220062 256578 220094 257134
rect 219474 221134 220094 256578
rect 219474 220578 219506 221134
rect 220062 220578 220094 221134
rect 219474 185134 220094 220578
rect 219474 184578 219506 185134
rect 220062 184578 220094 185134
rect 219474 149134 220094 184578
rect 219474 148578 219506 149134
rect 220062 148578 220094 149134
rect 219474 113134 220094 148578
rect 219474 112578 219506 113134
rect 220062 112578 220094 113134
rect 219474 77134 220094 112578
rect 219474 76578 219506 77134
rect 220062 76578 220094 77134
rect 219474 41134 220094 76578
rect 219474 40578 219506 41134
rect 220062 40578 220094 41134
rect 219474 5134 220094 40578
rect 219474 4578 219506 5134
rect 220062 4578 220094 5134
rect 219474 -2266 220094 4578
rect 219474 -2822 219506 -2266
rect 220062 -2822 220094 -2266
rect 219474 -7654 220094 -2822
rect 220714 707718 221334 711590
rect 220714 707162 220746 707718
rect 221302 707162 221334 707718
rect 220714 690374 221334 707162
rect 220714 689818 220746 690374
rect 221302 689818 221334 690374
rect 220714 654374 221334 689818
rect 220714 653818 220746 654374
rect 221302 653818 221334 654374
rect 220714 618374 221334 653818
rect 220714 617818 220746 618374
rect 221302 617818 221334 618374
rect 220714 582374 221334 617818
rect 220714 581818 220746 582374
rect 221302 581818 221334 582374
rect 220714 546374 221334 581818
rect 220714 545818 220746 546374
rect 221302 545818 221334 546374
rect 220714 510374 221334 545818
rect 220714 509818 220746 510374
rect 221302 509818 221334 510374
rect 220714 474374 221334 509818
rect 220714 473818 220746 474374
rect 221302 473818 221334 474374
rect 220714 438374 221334 473818
rect 220714 437818 220746 438374
rect 221302 437818 221334 438374
rect 220714 402374 221334 437818
rect 220714 401818 220746 402374
rect 221302 401818 221334 402374
rect 220714 366374 221334 401818
rect 220714 365818 220746 366374
rect 221302 365818 221334 366374
rect 220714 330374 221334 365818
rect 220714 329818 220746 330374
rect 221302 329818 221334 330374
rect 220714 294374 221334 329818
rect 220714 293818 220746 294374
rect 221302 293818 221334 294374
rect 220714 258374 221334 293818
rect 220714 257818 220746 258374
rect 221302 257818 221334 258374
rect 220714 222374 221334 257818
rect 220714 221818 220746 222374
rect 221302 221818 221334 222374
rect 220714 186374 221334 221818
rect 220714 185818 220746 186374
rect 221302 185818 221334 186374
rect 220714 150374 221334 185818
rect 220714 149818 220746 150374
rect 221302 149818 221334 150374
rect 220714 114374 221334 149818
rect 220714 113818 220746 114374
rect 221302 113818 221334 114374
rect 220714 78374 221334 113818
rect 220714 77818 220746 78374
rect 221302 77818 221334 78374
rect 220714 42374 221334 77818
rect 220714 41818 220746 42374
rect 221302 41818 221334 42374
rect 220714 6374 221334 41818
rect 220714 5818 220746 6374
rect 221302 5818 221334 6374
rect 220714 -3226 221334 5818
rect 220714 -3782 220746 -3226
rect 221302 -3782 221334 -3226
rect 220714 -7654 221334 -3782
rect 221954 708678 222574 711590
rect 221954 708122 221986 708678
rect 222542 708122 222574 708678
rect 221954 691614 222574 708122
rect 221954 691058 221986 691614
rect 222542 691058 222574 691614
rect 221954 655614 222574 691058
rect 221954 655058 221986 655614
rect 222542 655058 222574 655614
rect 221954 619614 222574 655058
rect 221954 619058 221986 619614
rect 222542 619058 222574 619614
rect 221954 583614 222574 619058
rect 221954 583058 221986 583614
rect 222542 583058 222574 583614
rect 221954 547614 222574 583058
rect 221954 547058 221986 547614
rect 222542 547058 222574 547614
rect 221954 511614 222574 547058
rect 221954 511058 221986 511614
rect 222542 511058 222574 511614
rect 221954 475614 222574 511058
rect 221954 475058 221986 475614
rect 222542 475058 222574 475614
rect 221954 439614 222574 475058
rect 221954 439058 221986 439614
rect 222542 439058 222574 439614
rect 221954 403614 222574 439058
rect 221954 403058 221986 403614
rect 222542 403058 222574 403614
rect 221954 367614 222574 403058
rect 221954 367058 221986 367614
rect 222542 367058 222574 367614
rect 221954 331614 222574 367058
rect 221954 331058 221986 331614
rect 222542 331058 222574 331614
rect 221954 295614 222574 331058
rect 221954 295058 221986 295614
rect 222542 295058 222574 295614
rect 221954 259614 222574 295058
rect 221954 259058 221986 259614
rect 222542 259058 222574 259614
rect 221954 223614 222574 259058
rect 221954 223058 221986 223614
rect 222542 223058 222574 223614
rect 221954 187614 222574 223058
rect 221954 187058 221986 187614
rect 222542 187058 222574 187614
rect 221954 151614 222574 187058
rect 221954 151058 221986 151614
rect 222542 151058 222574 151614
rect 221954 115614 222574 151058
rect 221954 115058 221986 115614
rect 222542 115058 222574 115614
rect 221954 79614 222574 115058
rect 221954 79058 221986 79614
rect 222542 79058 222574 79614
rect 221954 43614 222574 79058
rect 221954 43058 221986 43614
rect 222542 43058 222574 43614
rect 221954 7614 222574 43058
rect 221954 7058 221986 7614
rect 222542 7058 222574 7614
rect 221954 -4186 222574 7058
rect 221954 -4742 221986 -4186
rect 222542 -4742 222574 -4186
rect 221954 -7654 222574 -4742
rect 223194 709638 223814 711590
rect 223194 709082 223226 709638
rect 223782 709082 223814 709638
rect 223194 692854 223814 709082
rect 223194 692298 223226 692854
rect 223782 692298 223814 692854
rect 223194 656854 223814 692298
rect 223194 656298 223226 656854
rect 223782 656298 223814 656854
rect 223194 620854 223814 656298
rect 223194 620298 223226 620854
rect 223782 620298 223814 620854
rect 223194 584854 223814 620298
rect 223194 584298 223226 584854
rect 223782 584298 223814 584854
rect 223194 548854 223814 584298
rect 223194 548298 223226 548854
rect 223782 548298 223814 548854
rect 223194 512854 223814 548298
rect 223194 512298 223226 512854
rect 223782 512298 223814 512854
rect 223194 476854 223814 512298
rect 223194 476298 223226 476854
rect 223782 476298 223814 476854
rect 223194 440854 223814 476298
rect 223194 440298 223226 440854
rect 223782 440298 223814 440854
rect 223194 404854 223814 440298
rect 223194 404298 223226 404854
rect 223782 404298 223814 404854
rect 223194 368854 223814 404298
rect 223194 368298 223226 368854
rect 223782 368298 223814 368854
rect 223194 332854 223814 368298
rect 223194 332298 223226 332854
rect 223782 332298 223814 332854
rect 223194 296854 223814 332298
rect 223194 296298 223226 296854
rect 223782 296298 223814 296854
rect 223194 260854 223814 296298
rect 223194 260298 223226 260854
rect 223782 260298 223814 260854
rect 223194 224854 223814 260298
rect 223194 224298 223226 224854
rect 223782 224298 223814 224854
rect 223194 188854 223814 224298
rect 223194 188298 223226 188854
rect 223782 188298 223814 188854
rect 223194 152854 223814 188298
rect 223194 152298 223226 152854
rect 223782 152298 223814 152854
rect 223194 116854 223814 152298
rect 223194 116298 223226 116854
rect 223782 116298 223814 116854
rect 223194 80854 223814 116298
rect 223194 80298 223226 80854
rect 223782 80298 223814 80854
rect 223194 44854 223814 80298
rect 223194 44298 223226 44854
rect 223782 44298 223814 44854
rect 223194 8854 223814 44298
rect 223194 8298 223226 8854
rect 223782 8298 223814 8854
rect 223194 -5146 223814 8298
rect 223194 -5702 223226 -5146
rect 223782 -5702 223814 -5146
rect 223194 -7654 223814 -5702
rect 224434 710598 225054 711590
rect 224434 710042 224466 710598
rect 225022 710042 225054 710598
rect 224434 694094 225054 710042
rect 224434 693538 224466 694094
rect 225022 693538 225054 694094
rect 224434 658094 225054 693538
rect 224434 657538 224466 658094
rect 225022 657538 225054 658094
rect 224434 622094 225054 657538
rect 224434 621538 224466 622094
rect 225022 621538 225054 622094
rect 224434 586094 225054 621538
rect 224434 585538 224466 586094
rect 225022 585538 225054 586094
rect 224434 550094 225054 585538
rect 224434 549538 224466 550094
rect 225022 549538 225054 550094
rect 224434 514094 225054 549538
rect 224434 513538 224466 514094
rect 225022 513538 225054 514094
rect 224434 478094 225054 513538
rect 224434 477538 224466 478094
rect 225022 477538 225054 478094
rect 224434 442094 225054 477538
rect 224434 441538 224466 442094
rect 225022 441538 225054 442094
rect 224434 406094 225054 441538
rect 224434 405538 224466 406094
rect 225022 405538 225054 406094
rect 224434 370094 225054 405538
rect 224434 369538 224466 370094
rect 225022 369538 225054 370094
rect 224434 334094 225054 369538
rect 224434 333538 224466 334094
rect 225022 333538 225054 334094
rect 224434 298094 225054 333538
rect 224434 297538 224466 298094
rect 225022 297538 225054 298094
rect 224434 262094 225054 297538
rect 224434 261538 224466 262094
rect 225022 261538 225054 262094
rect 224434 226094 225054 261538
rect 224434 225538 224466 226094
rect 225022 225538 225054 226094
rect 224434 190094 225054 225538
rect 224434 189538 224466 190094
rect 225022 189538 225054 190094
rect 224434 154094 225054 189538
rect 224434 153538 224466 154094
rect 225022 153538 225054 154094
rect 224434 118094 225054 153538
rect 224434 117538 224466 118094
rect 225022 117538 225054 118094
rect 224434 82094 225054 117538
rect 224434 81538 224466 82094
rect 225022 81538 225054 82094
rect 224434 46094 225054 81538
rect 224434 45538 224466 46094
rect 225022 45538 225054 46094
rect 224434 10094 225054 45538
rect 224434 9538 224466 10094
rect 225022 9538 225054 10094
rect 224434 -6106 225054 9538
rect 224434 -6662 224466 -6106
rect 225022 -6662 225054 -6106
rect 224434 -7654 225054 -6662
rect 225674 711558 226294 711590
rect 225674 711002 225706 711558
rect 226262 711002 226294 711558
rect 225674 695334 226294 711002
rect 225674 694778 225706 695334
rect 226262 694778 226294 695334
rect 225674 659334 226294 694778
rect 225674 658778 225706 659334
rect 226262 658778 226294 659334
rect 225674 623334 226294 658778
rect 225674 622778 225706 623334
rect 226262 622778 226294 623334
rect 225674 587334 226294 622778
rect 225674 586778 225706 587334
rect 226262 586778 226294 587334
rect 225674 551334 226294 586778
rect 225674 550778 225706 551334
rect 226262 550778 226294 551334
rect 225674 515334 226294 550778
rect 225674 514778 225706 515334
rect 226262 514778 226294 515334
rect 225674 479334 226294 514778
rect 225674 478778 225706 479334
rect 226262 478778 226294 479334
rect 225674 443334 226294 478778
rect 225674 442778 225706 443334
rect 226262 442778 226294 443334
rect 225674 407334 226294 442778
rect 225674 406778 225706 407334
rect 226262 406778 226294 407334
rect 225674 371334 226294 406778
rect 225674 370778 225706 371334
rect 226262 370778 226294 371334
rect 225674 335334 226294 370778
rect 225674 334778 225706 335334
rect 226262 334778 226294 335334
rect 225674 299334 226294 334778
rect 225674 298778 225706 299334
rect 226262 298778 226294 299334
rect 225674 263334 226294 298778
rect 225674 262778 225706 263334
rect 226262 262778 226294 263334
rect 225674 227334 226294 262778
rect 225674 226778 225706 227334
rect 226262 226778 226294 227334
rect 225674 191334 226294 226778
rect 225674 190778 225706 191334
rect 226262 190778 226294 191334
rect 225674 155334 226294 190778
rect 225674 154778 225706 155334
rect 226262 154778 226294 155334
rect 225674 119334 226294 154778
rect 225674 118778 225706 119334
rect 226262 118778 226294 119334
rect 225674 83334 226294 118778
rect 225674 82778 225706 83334
rect 226262 82778 226294 83334
rect 225674 47334 226294 82778
rect 225674 46778 225706 47334
rect 226262 46778 226294 47334
rect 225674 11334 226294 46778
rect 225674 10778 225706 11334
rect 226262 10778 226294 11334
rect 225674 -7066 226294 10778
rect 225674 -7622 225706 -7066
rect 226262 -7622 226294 -7066
rect 225674 -7654 226294 -7622
rect 252994 704838 253614 711590
rect 252994 704282 253026 704838
rect 253582 704282 253614 704838
rect 252994 686654 253614 704282
rect 252994 686098 253026 686654
rect 253582 686098 253614 686654
rect 252994 650654 253614 686098
rect 252994 650098 253026 650654
rect 253582 650098 253614 650654
rect 252994 614654 253614 650098
rect 252994 614098 253026 614654
rect 253582 614098 253614 614654
rect 252994 578654 253614 614098
rect 252994 578098 253026 578654
rect 253582 578098 253614 578654
rect 252994 542654 253614 578098
rect 252994 542098 253026 542654
rect 253582 542098 253614 542654
rect 252994 506654 253614 542098
rect 252994 506098 253026 506654
rect 253582 506098 253614 506654
rect 252994 470654 253614 506098
rect 252994 470098 253026 470654
rect 253582 470098 253614 470654
rect 252994 434654 253614 470098
rect 252994 434098 253026 434654
rect 253582 434098 253614 434654
rect 252994 398654 253614 434098
rect 252994 398098 253026 398654
rect 253582 398098 253614 398654
rect 252994 362654 253614 398098
rect 252994 362098 253026 362654
rect 253582 362098 253614 362654
rect 252994 326654 253614 362098
rect 252994 326098 253026 326654
rect 253582 326098 253614 326654
rect 252994 290654 253614 326098
rect 252994 290098 253026 290654
rect 253582 290098 253614 290654
rect 252994 254654 253614 290098
rect 252994 254098 253026 254654
rect 253582 254098 253614 254654
rect 252994 218654 253614 254098
rect 252994 218098 253026 218654
rect 253582 218098 253614 218654
rect 252994 182654 253614 218098
rect 252994 182098 253026 182654
rect 253582 182098 253614 182654
rect 252994 146654 253614 182098
rect 252994 146098 253026 146654
rect 253582 146098 253614 146654
rect 252994 110654 253614 146098
rect 252994 110098 253026 110654
rect 253582 110098 253614 110654
rect 252994 74654 253614 110098
rect 252994 74098 253026 74654
rect 253582 74098 253614 74654
rect 252994 38654 253614 74098
rect 252994 38098 253026 38654
rect 253582 38098 253614 38654
rect 252994 2654 253614 38098
rect 252994 2098 253026 2654
rect 253582 2098 253614 2654
rect 252994 -346 253614 2098
rect 252994 -902 253026 -346
rect 253582 -902 253614 -346
rect 252994 -7654 253614 -902
rect 254234 705798 254854 711590
rect 254234 705242 254266 705798
rect 254822 705242 254854 705798
rect 254234 687894 254854 705242
rect 254234 687338 254266 687894
rect 254822 687338 254854 687894
rect 254234 651894 254854 687338
rect 254234 651338 254266 651894
rect 254822 651338 254854 651894
rect 254234 615894 254854 651338
rect 254234 615338 254266 615894
rect 254822 615338 254854 615894
rect 254234 579894 254854 615338
rect 254234 579338 254266 579894
rect 254822 579338 254854 579894
rect 254234 543894 254854 579338
rect 254234 543338 254266 543894
rect 254822 543338 254854 543894
rect 254234 507894 254854 543338
rect 254234 507338 254266 507894
rect 254822 507338 254854 507894
rect 254234 471894 254854 507338
rect 254234 471338 254266 471894
rect 254822 471338 254854 471894
rect 254234 435894 254854 471338
rect 254234 435338 254266 435894
rect 254822 435338 254854 435894
rect 254234 399894 254854 435338
rect 254234 399338 254266 399894
rect 254822 399338 254854 399894
rect 254234 363894 254854 399338
rect 254234 363338 254266 363894
rect 254822 363338 254854 363894
rect 254234 327894 254854 363338
rect 254234 327338 254266 327894
rect 254822 327338 254854 327894
rect 254234 291894 254854 327338
rect 254234 291338 254266 291894
rect 254822 291338 254854 291894
rect 254234 255894 254854 291338
rect 254234 255338 254266 255894
rect 254822 255338 254854 255894
rect 254234 219894 254854 255338
rect 254234 219338 254266 219894
rect 254822 219338 254854 219894
rect 254234 183894 254854 219338
rect 254234 183338 254266 183894
rect 254822 183338 254854 183894
rect 254234 147894 254854 183338
rect 254234 147338 254266 147894
rect 254822 147338 254854 147894
rect 254234 111894 254854 147338
rect 254234 111338 254266 111894
rect 254822 111338 254854 111894
rect 254234 75894 254854 111338
rect 254234 75338 254266 75894
rect 254822 75338 254854 75894
rect 254234 39894 254854 75338
rect 254234 39338 254266 39894
rect 254822 39338 254854 39894
rect 254234 3894 254854 39338
rect 254234 3338 254266 3894
rect 254822 3338 254854 3894
rect 254234 -1306 254854 3338
rect 254234 -1862 254266 -1306
rect 254822 -1862 254854 -1306
rect 254234 -7654 254854 -1862
rect 255474 706758 256094 711590
rect 255474 706202 255506 706758
rect 256062 706202 256094 706758
rect 255474 689134 256094 706202
rect 255474 688578 255506 689134
rect 256062 688578 256094 689134
rect 255474 653134 256094 688578
rect 255474 652578 255506 653134
rect 256062 652578 256094 653134
rect 255474 617134 256094 652578
rect 255474 616578 255506 617134
rect 256062 616578 256094 617134
rect 255474 581134 256094 616578
rect 255474 580578 255506 581134
rect 256062 580578 256094 581134
rect 255474 545134 256094 580578
rect 255474 544578 255506 545134
rect 256062 544578 256094 545134
rect 255474 509134 256094 544578
rect 255474 508578 255506 509134
rect 256062 508578 256094 509134
rect 255474 473134 256094 508578
rect 255474 472578 255506 473134
rect 256062 472578 256094 473134
rect 255474 437134 256094 472578
rect 255474 436578 255506 437134
rect 256062 436578 256094 437134
rect 255474 401134 256094 436578
rect 255474 400578 255506 401134
rect 256062 400578 256094 401134
rect 255474 365134 256094 400578
rect 255474 364578 255506 365134
rect 256062 364578 256094 365134
rect 255474 329134 256094 364578
rect 255474 328578 255506 329134
rect 256062 328578 256094 329134
rect 255474 293134 256094 328578
rect 255474 292578 255506 293134
rect 256062 292578 256094 293134
rect 255474 257134 256094 292578
rect 255474 256578 255506 257134
rect 256062 256578 256094 257134
rect 255474 221134 256094 256578
rect 255474 220578 255506 221134
rect 256062 220578 256094 221134
rect 255474 185134 256094 220578
rect 255474 184578 255506 185134
rect 256062 184578 256094 185134
rect 255474 149134 256094 184578
rect 255474 148578 255506 149134
rect 256062 148578 256094 149134
rect 255474 113134 256094 148578
rect 255474 112578 255506 113134
rect 256062 112578 256094 113134
rect 255474 77134 256094 112578
rect 255474 76578 255506 77134
rect 256062 76578 256094 77134
rect 255474 41134 256094 76578
rect 255474 40578 255506 41134
rect 256062 40578 256094 41134
rect 255474 5134 256094 40578
rect 255474 4578 255506 5134
rect 256062 4578 256094 5134
rect 255474 -2266 256094 4578
rect 255474 -2822 255506 -2266
rect 256062 -2822 256094 -2266
rect 255474 -7654 256094 -2822
rect 256714 707718 257334 711590
rect 256714 707162 256746 707718
rect 257302 707162 257334 707718
rect 256714 690374 257334 707162
rect 256714 689818 256746 690374
rect 257302 689818 257334 690374
rect 256714 654374 257334 689818
rect 256714 653818 256746 654374
rect 257302 653818 257334 654374
rect 256714 618374 257334 653818
rect 256714 617818 256746 618374
rect 257302 617818 257334 618374
rect 256714 582374 257334 617818
rect 256714 581818 256746 582374
rect 257302 581818 257334 582374
rect 256714 546374 257334 581818
rect 256714 545818 256746 546374
rect 257302 545818 257334 546374
rect 256714 510374 257334 545818
rect 256714 509818 256746 510374
rect 257302 509818 257334 510374
rect 256714 474374 257334 509818
rect 256714 473818 256746 474374
rect 257302 473818 257334 474374
rect 256714 438374 257334 473818
rect 256714 437818 256746 438374
rect 257302 437818 257334 438374
rect 256714 402374 257334 437818
rect 256714 401818 256746 402374
rect 257302 401818 257334 402374
rect 256714 366374 257334 401818
rect 256714 365818 256746 366374
rect 257302 365818 257334 366374
rect 256714 330374 257334 365818
rect 256714 329818 256746 330374
rect 257302 329818 257334 330374
rect 256714 294374 257334 329818
rect 256714 293818 256746 294374
rect 257302 293818 257334 294374
rect 256714 258374 257334 293818
rect 256714 257818 256746 258374
rect 257302 257818 257334 258374
rect 256714 222374 257334 257818
rect 256714 221818 256746 222374
rect 257302 221818 257334 222374
rect 256714 186374 257334 221818
rect 256714 185818 256746 186374
rect 257302 185818 257334 186374
rect 256714 150374 257334 185818
rect 256714 149818 256746 150374
rect 257302 149818 257334 150374
rect 256714 114374 257334 149818
rect 256714 113818 256746 114374
rect 257302 113818 257334 114374
rect 256714 78374 257334 113818
rect 256714 77818 256746 78374
rect 257302 77818 257334 78374
rect 256714 42374 257334 77818
rect 256714 41818 256746 42374
rect 257302 41818 257334 42374
rect 256714 6374 257334 41818
rect 256714 5818 256746 6374
rect 257302 5818 257334 6374
rect 256714 -3226 257334 5818
rect 256714 -3782 256746 -3226
rect 257302 -3782 257334 -3226
rect 256714 -7654 257334 -3782
rect 257954 708678 258574 711590
rect 257954 708122 257986 708678
rect 258542 708122 258574 708678
rect 257954 691614 258574 708122
rect 257954 691058 257986 691614
rect 258542 691058 258574 691614
rect 257954 655614 258574 691058
rect 257954 655058 257986 655614
rect 258542 655058 258574 655614
rect 257954 619614 258574 655058
rect 257954 619058 257986 619614
rect 258542 619058 258574 619614
rect 257954 583614 258574 619058
rect 257954 583058 257986 583614
rect 258542 583058 258574 583614
rect 257954 547614 258574 583058
rect 257954 547058 257986 547614
rect 258542 547058 258574 547614
rect 257954 511614 258574 547058
rect 257954 511058 257986 511614
rect 258542 511058 258574 511614
rect 257954 475614 258574 511058
rect 257954 475058 257986 475614
rect 258542 475058 258574 475614
rect 257954 439614 258574 475058
rect 257954 439058 257986 439614
rect 258542 439058 258574 439614
rect 257954 403614 258574 439058
rect 257954 403058 257986 403614
rect 258542 403058 258574 403614
rect 257954 367614 258574 403058
rect 257954 367058 257986 367614
rect 258542 367058 258574 367614
rect 257954 331614 258574 367058
rect 257954 331058 257986 331614
rect 258542 331058 258574 331614
rect 257954 295614 258574 331058
rect 257954 295058 257986 295614
rect 258542 295058 258574 295614
rect 257954 259614 258574 295058
rect 257954 259058 257986 259614
rect 258542 259058 258574 259614
rect 257954 223614 258574 259058
rect 257954 223058 257986 223614
rect 258542 223058 258574 223614
rect 257954 187614 258574 223058
rect 257954 187058 257986 187614
rect 258542 187058 258574 187614
rect 257954 151614 258574 187058
rect 257954 151058 257986 151614
rect 258542 151058 258574 151614
rect 257954 115614 258574 151058
rect 257954 115058 257986 115614
rect 258542 115058 258574 115614
rect 257954 79614 258574 115058
rect 257954 79058 257986 79614
rect 258542 79058 258574 79614
rect 257954 43614 258574 79058
rect 257954 43058 257986 43614
rect 258542 43058 258574 43614
rect 257954 7614 258574 43058
rect 257954 7058 257986 7614
rect 258542 7058 258574 7614
rect 257954 -4186 258574 7058
rect 257954 -4742 257986 -4186
rect 258542 -4742 258574 -4186
rect 257954 -7654 258574 -4742
rect 259194 709638 259814 711590
rect 259194 709082 259226 709638
rect 259782 709082 259814 709638
rect 259194 692854 259814 709082
rect 259194 692298 259226 692854
rect 259782 692298 259814 692854
rect 259194 656854 259814 692298
rect 259194 656298 259226 656854
rect 259782 656298 259814 656854
rect 259194 620854 259814 656298
rect 259194 620298 259226 620854
rect 259782 620298 259814 620854
rect 259194 584854 259814 620298
rect 259194 584298 259226 584854
rect 259782 584298 259814 584854
rect 259194 548854 259814 584298
rect 259194 548298 259226 548854
rect 259782 548298 259814 548854
rect 259194 512854 259814 548298
rect 259194 512298 259226 512854
rect 259782 512298 259814 512854
rect 259194 476854 259814 512298
rect 259194 476298 259226 476854
rect 259782 476298 259814 476854
rect 259194 440854 259814 476298
rect 259194 440298 259226 440854
rect 259782 440298 259814 440854
rect 259194 404854 259814 440298
rect 259194 404298 259226 404854
rect 259782 404298 259814 404854
rect 259194 368854 259814 404298
rect 259194 368298 259226 368854
rect 259782 368298 259814 368854
rect 259194 332854 259814 368298
rect 259194 332298 259226 332854
rect 259782 332298 259814 332854
rect 259194 296854 259814 332298
rect 259194 296298 259226 296854
rect 259782 296298 259814 296854
rect 259194 260854 259814 296298
rect 259194 260298 259226 260854
rect 259782 260298 259814 260854
rect 259194 224854 259814 260298
rect 259194 224298 259226 224854
rect 259782 224298 259814 224854
rect 259194 188854 259814 224298
rect 259194 188298 259226 188854
rect 259782 188298 259814 188854
rect 259194 152854 259814 188298
rect 259194 152298 259226 152854
rect 259782 152298 259814 152854
rect 259194 116854 259814 152298
rect 259194 116298 259226 116854
rect 259782 116298 259814 116854
rect 259194 80854 259814 116298
rect 259194 80298 259226 80854
rect 259782 80298 259814 80854
rect 259194 44854 259814 80298
rect 259194 44298 259226 44854
rect 259782 44298 259814 44854
rect 259194 8854 259814 44298
rect 259194 8298 259226 8854
rect 259782 8298 259814 8854
rect 259194 -5146 259814 8298
rect 259194 -5702 259226 -5146
rect 259782 -5702 259814 -5146
rect 259194 -7654 259814 -5702
rect 260434 710598 261054 711590
rect 260434 710042 260466 710598
rect 261022 710042 261054 710598
rect 260434 694094 261054 710042
rect 260434 693538 260466 694094
rect 261022 693538 261054 694094
rect 260434 658094 261054 693538
rect 260434 657538 260466 658094
rect 261022 657538 261054 658094
rect 260434 622094 261054 657538
rect 260434 621538 260466 622094
rect 261022 621538 261054 622094
rect 260434 586094 261054 621538
rect 260434 585538 260466 586094
rect 261022 585538 261054 586094
rect 260434 550094 261054 585538
rect 260434 549538 260466 550094
rect 261022 549538 261054 550094
rect 260434 514094 261054 549538
rect 260434 513538 260466 514094
rect 261022 513538 261054 514094
rect 260434 478094 261054 513538
rect 260434 477538 260466 478094
rect 261022 477538 261054 478094
rect 260434 442094 261054 477538
rect 260434 441538 260466 442094
rect 261022 441538 261054 442094
rect 260434 406094 261054 441538
rect 260434 405538 260466 406094
rect 261022 405538 261054 406094
rect 260434 370094 261054 405538
rect 260434 369538 260466 370094
rect 261022 369538 261054 370094
rect 260434 334094 261054 369538
rect 260434 333538 260466 334094
rect 261022 333538 261054 334094
rect 260434 298094 261054 333538
rect 260434 297538 260466 298094
rect 261022 297538 261054 298094
rect 260434 262094 261054 297538
rect 260434 261538 260466 262094
rect 261022 261538 261054 262094
rect 260434 226094 261054 261538
rect 260434 225538 260466 226094
rect 261022 225538 261054 226094
rect 260434 190094 261054 225538
rect 260434 189538 260466 190094
rect 261022 189538 261054 190094
rect 260434 154094 261054 189538
rect 260434 153538 260466 154094
rect 261022 153538 261054 154094
rect 260434 118094 261054 153538
rect 260434 117538 260466 118094
rect 261022 117538 261054 118094
rect 260434 82094 261054 117538
rect 260434 81538 260466 82094
rect 261022 81538 261054 82094
rect 260434 46094 261054 81538
rect 260434 45538 260466 46094
rect 261022 45538 261054 46094
rect 260434 10094 261054 45538
rect 260434 9538 260466 10094
rect 261022 9538 261054 10094
rect 260434 -6106 261054 9538
rect 260434 -6662 260466 -6106
rect 261022 -6662 261054 -6106
rect 260434 -7654 261054 -6662
rect 261674 711558 262294 711590
rect 261674 711002 261706 711558
rect 262262 711002 262294 711558
rect 261674 695334 262294 711002
rect 261674 694778 261706 695334
rect 262262 694778 262294 695334
rect 261674 659334 262294 694778
rect 261674 658778 261706 659334
rect 262262 658778 262294 659334
rect 261674 623334 262294 658778
rect 261674 622778 261706 623334
rect 262262 622778 262294 623334
rect 261674 587334 262294 622778
rect 261674 586778 261706 587334
rect 262262 586778 262294 587334
rect 261674 551334 262294 586778
rect 261674 550778 261706 551334
rect 262262 550778 262294 551334
rect 261674 515334 262294 550778
rect 261674 514778 261706 515334
rect 262262 514778 262294 515334
rect 261674 479334 262294 514778
rect 261674 478778 261706 479334
rect 262262 478778 262294 479334
rect 261674 443334 262294 478778
rect 261674 442778 261706 443334
rect 262262 442778 262294 443334
rect 261674 407334 262294 442778
rect 261674 406778 261706 407334
rect 262262 406778 262294 407334
rect 261674 371334 262294 406778
rect 261674 370778 261706 371334
rect 262262 370778 262294 371334
rect 261674 335334 262294 370778
rect 261674 334778 261706 335334
rect 262262 334778 262294 335334
rect 261674 299334 262294 334778
rect 261674 298778 261706 299334
rect 262262 298778 262294 299334
rect 261674 263334 262294 298778
rect 261674 262778 261706 263334
rect 262262 262778 262294 263334
rect 261674 227334 262294 262778
rect 261674 226778 261706 227334
rect 262262 226778 262294 227334
rect 261674 191334 262294 226778
rect 261674 190778 261706 191334
rect 262262 190778 262294 191334
rect 261674 155334 262294 190778
rect 261674 154778 261706 155334
rect 262262 154778 262294 155334
rect 261674 119334 262294 154778
rect 261674 118778 261706 119334
rect 262262 118778 262294 119334
rect 261674 83334 262294 118778
rect 261674 82778 261706 83334
rect 262262 82778 262294 83334
rect 261674 47334 262294 82778
rect 261674 46778 261706 47334
rect 262262 46778 262294 47334
rect 261674 11334 262294 46778
rect 261674 10778 261706 11334
rect 262262 10778 262294 11334
rect 261674 -7066 262294 10778
rect 261674 -7622 261706 -7066
rect 262262 -7622 262294 -7066
rect 261674 -7654 262294 -7622
rect 288994 704838 289614 711590
rect 288994 704282 289026 704838
rect 289582 704282 289614 704838
rect 288994 686654 289614 704282
rect 288994 686098 289026 686654
rect 289582 686098 289614 686654
rect 288994 650654 289614 686098
rect 288994 650098 289026 650654
rect 289582 650098 289614 650654
rect 288994 614654 289614 650098
rect 288994 614098 289026 614654
rect 289582 614098 289614 614654
rect 288994 578654 289614 614098
rect 288994 578098 289026 578654
rect 289582 578098 289614 578654
rect 288994 542654 289614 578098
rect 288994 542098 289026 542654
rect 289582 542098 289614 542654
rect 288994 506654 289614 542098
rect 288994 506098 289026 506654
rect 289582 506098 289614 506654
rect 288994 470654 289614 506098
rect 288994 470098 289026 470654
rect 289582 470098 289614 470654
rect 288994 434654 289614 470098
rect 288994 434098 289026 434654
rect 289582 434098 289614 434654
rect 288994 398654 289614 434098
rect 288994 398098 289026 398654
rect 289582 398098 289614 398654
rect 288994 362654 289614 398098
rect 288994 362098 289026 362654
rect 289582 362098 289614 362654
rect 288994 326654 289614 362098
rect 288994 326098 289026 326654
rect 289582 326098 289614 326654
rect 288994 290654 289614 326098
rect 288994 290098 289026 290654
rect 289582 290098 289614 290654
rect 288994 254654 289614 290098
rect 288994 254098 289026 254654
rect 289582 254098 289614 254654
rect 288994 218654 289614 254098
rect 288994 218098 289026 218654
rect 289582 218098 289614 218654
rect 288994 182654 289614 218098
rect 288994 182098 289026 182654
rect 289582 182098 289614 182654
rect 288994 146654 289614 182098
rect 288994 146098 289026 146654
rect 289582 146098 289614 146654
rect 288994 110654 289614 146098
rect 288994 110098 289026 110654
rect 289582 110098 289614 110654
rect 288994 74654 289614 110098
rect 288994 74098 289026 74654
rect 289582 74098 289614 74654
rect 288994 38654 289614 74098
rect 288994 38098 289026 38654
rect 289582 38098 289614 38654
rect 288994 2654 289614 38098
rect 288994 2098 289026 2654
rect 289582 2098 289614 2654
rect 288994 -346 289614 2098
rect 288994 -902 289026 -346
rect 289582 -902 289614 -346
rect 288994 -7654 289614 -902
rect 290234 705798 290854 711590
rect 290234 705242 290266 705798
rect 290822 705242 290854 705798
rect 290234 687894 290854 705242
rect 290234 687338 290266 687894
rect 290822 687338 290854 687894
rect 290234 651894 290854 687338
rect 290234 651338 290266 651894
rect 290822 651338 290854 651894
rect 290234 615894 290854 651338
rect 290234 615338 290266 615894
rect 290822 615338 290854 615894
rect 290234 579894 290854 615338
rect 290234 579338 290266 579894
rect 290822 579338 290854 579894
rect 290234 543894 290854 579338
rect 290234 543338 290266 543894
rect 290822 543338 290854 543894
rect 290234 507894 290854 543338
rect 290234 507338 290266 507894
rect 290822 507338 290854 507894
rect 290234 471894 290854 507338
rect 290234 471338 290266 471894
rect 290822 471338 290854 471894
rect 290234 435894 290854 471338
rect 290234 435338 290266 435894
rect 290822 435338 290854 435894
rect 290234 399894 290854 435338
rect 290234 399338 290266 399894
rect 290822 399338 290854 399894
rect 290234 363894 290854 399338
rect 290234 363338 290266 363894
rect 290822 363338 290854 363894
rect 290234 327894 290854 363338
rect 290234 327338 290266 327894
rect 290822 327338 290854 327894
rect 290234 291894 290854 327338
rect 290234 291338 290266 291894
rect 290822 291338 290854 291894
rect 290234 255894 290854 291338
rect 290234 255338 290266 255894
rect 290822 255338 290854 255894
rect 290234 219894 290854 255338
rect 290234 219338 290266 219894
rect 290822 219338 290854 219894
rect 290234 183894 290854 219338
rect 290234 183338 290266 183894
rect 290822 183338 290854 183894
rect 290234 147894 290854 183338
rect 290234 147338 290266 147894
rect 290822 147338 290854 147894
rect 290234 111894 290854 147338
rect 290234 111338 290266 111894
rect 290822 111338 290854 111894
rect 290234 75894 290854 111338
rect 290234 75338 290266 75894
rect 290822 75338 290854 75894
rect 290234 39894 290854 75338
rect 290234 39338 290266 39894
rect 290822 39338 290854 39894
rect 290234 3894 290854 39338
rect 290234 3338 290266 3894
rect 290822 3338 290854 3894
rect 290234 -1306 290854 3338
rect 290234 -1862 290266 -1306
rect 290822 -1862 290854 -1306
rect 290234 -7654 290854 -1862
rect 291474 706758 292094 711590
rect 291474 706202 291506 706758
rect 292062 706202 292094 706758
rect 291474 689134 292094 706202
rect 291474 688578 291506 689134
rect 292062 688578 292094 689134
rect 291474 653134 292094 688578
rect 291474 652578 291506 653134
rect 292062 652578 292094 653134
rect 291474 617134 292094 652578
rect 291474 616578 291506 617134
rect 292062 616578 292094 617134
rect 291474 581134 292094 616578
rect 291474 580578 291506 581134
rect 292062 580578 292094 581134
rect 291474 545134 292094 580578
rect 291474 544578 291506 545134
rect 292062 544578 292094 545134
rect 291474 509134 292094 544578
rect 291474 508578 291506 509134
rect 292062 508578 292094 509134
rect 291474 473134 292094 508578
rect 291474 472578 291506 473134
rect 292062 472578 292094 473134
rect 291474 437134 292094 472578
rect 291474 436578 291506 437134
rect 292062 436578 292094 437134
rect 291474 401134 292094 436578
rect 291474 400578 291506 401134
rect 292062 400578 292094 401134
rect 291474 365134 292094 400578
rect 291474 364578 291506 365134
rect 292062 364578 292094 365134
rect 291474 329134 292094 364578
rect 291474 328578 291506 329134
rect 292062 328578 292094 329134
rect 291474 293134 292094 328578
rect 291474 292578 291506 293134
rect 292062 292578 292094 293134
rect 291474 257134 292094 292578
rect 291474 256578 291506 257134
rect 292062 256578 292094 257134
rect 291474 221134 292094 256578
rect 291474 220578 291506 221134
rect 292062 220578 292094 221134
rect 291474 185134 292094 220578
rect 291474 184578 291506 185134
rect 292062 184578 292094 185134
rect 291474 149134 292094 184578
rect 291474 148578 291506 149134
rect 292062 148578 292094 149134
rect 291474 113134 292094 148578
rect 291474 112578 291506 113134
rect 292062 112578 292094 113134
rect 291474 77134 292094 112578
rect 291474 76578 291506 77134
rect 292062 76578 292094 77134
rect 291474 41134 292094 76578
rect 291474 40578 291506 41134
rect 292062 40578 292094 41134
rect 291474 5134 292094 40578
rect 291474 4578 291506 5134
rect 292062 4578 292094 5134
rect 291474 -2266 292094 4578
rect 291474 -2822 291506 -2266
rect 292062 -2822 292094 -2266
rect 291474 -7654 292094 -2822
rect 292714 707718 293334 711590
rect 292714 707162 292746 707718
rect 293302 707162 293334 707718
rect 292714 690374 293334 707162
rect 292714 689818 292746 690374
rect 293302 689818 293334 690374
rect 292714 654374 293334 689818
rect 292714 653818 292746 654374
rect 293302 653818 293334 654374
rect 292714 618374 293334 653818
rect 292714 617818 292746 618374
rect 293302 617818 293334 618374
rect 292714 582374 293334 617818
rect 292714 581818 292746 582374
rect 293302 581818 293334 582374
rect 292714 546374 293334 581818
rect 292714 545818 292746 546374
rect 293302 545818 293334 546374
rect 292714 510374 293334 545818
rect 292714 509818 292746 510374
rect 293302 509818 293334 510374
rect 292714 474374 293334 509818
rect 292714 473818 292746 474374
rect 293302 473818 293334 474374
rect 292714 438374 293334 473818
rect 292714 437818 292746 438374
rect 293302 437818 293334 438374
rect 292714 402374 293334 437818
rect 292714 401818 292746 402374
rect 293302 401818 293334 402374
rect 292714 366374 293334 401818
rect 292714 365818 292746 366374
rect 293302 365818 293334 366374
rect 292714 330374 293334 365818
rect 292714 329818 292746 330374
rect 293302 329818 293334 330374
rect 292714 294374 293334 329818
rect 292714 293818 292746 294374
rect 293302 293818 293334 294374
rect 292714 258374 293334 293818
rect 292714 257818 292746 258374
rect 293302 257818 293334 258374
rect 292714 222374 293334 257818
rect 292714 221818 292746 222374
rect 293302 221818 293334 222374
rect 292714 186374 293334 221818
rect 292714 185818 292746 186374
rect 293302 185818 293334 186374
rect 292714 150374 293334 185818
rect 292714 149818 292746 150374
rect 293302 149818 293334 150374
rect 292714 114374 293334 149818
rect 292714 113818 292746 114374
rect 293302 113818 293334 114374
rect 292714 78374 293334 113818
rect 292714 77818 292746 78374
rect 293302 77818 293334 78374
rect 292714 42374 293334 77818
rect 292714 41818 292746 42374
rect 293302 41818 293334 42374
rect 292714 6374 293334 41818
rect 292714 5818 292746 6374
rect 293302 5818 293334 6374
rect 292714 -3226 293334 5818
rect 292714 -3782 292746 -3226
rect 293302 -3782 293334 -3226
rect 292714 -7654 293334 -3782
rect 293954 708678 294574 711590
rect 293954 708122 293986 708678
rect 294542 708122 294574 708678
rect 293954 691614 294574 708122
rect 293954 691058 293986 691614
rect 294542 691058 294574 691614
rect 293954 655614 294574 691058
rect 293954 655058 293986 655614
rect 294542 655058 294574 655614
rect 293954 619614 294574 655058
rect 293954 619058 293986 619614
rect 294542 619058 294574 619614
rect 293954 583614 294574 619058
rect 293954 583058 293986 583614
rect 294542 583058 294574 583614
rect 293954 547614 294574 583058
rect 293954 547058 293986 547614
rect 294542 547058 294574 547614
rect 293954 511614 294574 547058
rect 293954 511058 293986 511614
rect 294542 511058 294574 511614
rect 293954 475614 294574 511058
rect 293954 475058 293986 475614
rect 294542 475058 294574 475614
rect 293954 439614 294574 475058
rect 293954 439058 293986 439614
rect 294542 439058 294574 439614
rect 293954 403614 294574 439058
rect 293954 403058 293986 403614
rect 294542 403058 294574 403614
rect 293954 367614 294574 403058
rect 293954 367058 293986 367614
rect 294542 367058 294574 367614
rect 293954 331614 294574 367058
rect 293954 331058 293986 331614
rect 294542 331058 294574 331614
rect 293954 295614 294574 331058
rect 293954 295058 293986 295614
rect 294542 295058 294574 295614
rect 293954 259614 294574 295058
rect 293954 259058 293986 259614
rect 294542 259058 294574 259614
rect 293954 223614 294574 259058
rect 293954 223058 293986 223614
rect 294542 223058 294574 223614
rect 293954 187614 294574 223058
rect 293954 187058 293986 187614
rect 294542 187058 294574 187614
rect 293954 151614 294574 187058
rect 293954 151058 293986 151614
rect 294542 151058 294574 151614
rect 293954 115614 294574 151058
rect 293954 115058 293986 115614
rect 294542 115058 294574 115614
rect 293954 79614 294574 115058
rect 293954 79058 293986 79614
rect 294542 79058 294574 79614
rect 293954 43614 294574 79058
rect 293954 43058 293986 43614
rect 294542 43058 294574 43614
rect 293954 7614 294574 43058
rect 293954 7058 293986 7614
rect 294542 7058 294574 7614
rect 293954 -4186 294574 7058
rect 293954 -4742 293986 -4186
rect 294542 -4742 294574 -4186
rect 293954 -7654 294574 -4742
rect 295194 709638 295814 711590
rect 295194 709082 295226 709638
rect 295782 709082 295814 709638
rect 295194 692854 295814 709082
rect 295194 692298 295226 692854
rect 295782 692298 295814 692854
rect 295194 656854 295814 692298
rect 295194 656298 295226 656854
rect 295782 656298 295814 656854
rect 295194 620854 295814 656298
rect 295194 620298 295226 620854
rect 295782 620298 295814 620854
rect 295194 584854 295814 620298
rect 295194 584298 295226 584854
rect 295782 584298 295814 584854
rect 295194 548854 295814 584298
rect 295194 548298 295226 548854
rect 295782 548298 295814 548854
rect 295194 512854 295814 548298
rect 295194 512298 295226 512854
rect 295782 512298 295814 512854
rect 295194 476854 295814 512298
rect 295194 476298 295226 476854
rect 295782 476298 295814 476854
rect 295194 440854 295814 476298
rect 295194 440298 295226 440854
rect 295782 440298 295814 440854
rect 295194 404854 295814 440298
rect 295194 404298 295226 404854
rect 295782 404298 295814 404854
rect 295194 368854 295814 404298
rect 295194 368298 295226 368854
rect 295782 368298 295814 368854
rect 295194 332854 295814 368298
rect 295194 332298 295226 332854
rect 295782 332298 295814 332854
rect 295194 296854 295814 332298
rect 295194 296298 295226 296854
rect 295782 296298 295814 296854
rect 295194 260854 295814 296298
rect 295194 260298 295226 260854
rect 295782 260298 295814 260854
rect 295194 224854 295814 260298
rect 295194 224298 295226 224854
rect 295782 224298 295814 224854
rect 295194 188854 295814 224298
rect 295194 188298 295226 188854
rect 295782 188298 295814 188854
rect 295194 152854 295814 188298
rect 295194 152298 295226 152854
rect 295782 152298 295814 152854
rect 295194 116854 295814 152298
rect 295194 116298 295226 116854
rect 295782 116298 295814 116854
rect 295194 80854 295814 116298
rect 295194 80298 295226 80854
rect 295782 80298 295814 80854
rect 295194 44854 295814 80298
rect 295194 44298 295226 44854
rect 295782 44298 295814 44854
rect 295194 8854 295814 44298
rect 295194 8298 295226 8854
rect 295782 8298 295814 8854
rect 295194 -5146 295814 8298
rect 295194 -5702 295226 -5146
rect 295782 -5702 295814 -5146
rect 295194 -7654 295814 -5702
rect 296434 710598 297054 711590
rect 296434 710042 296466 710598
rect 297022 710042 297054 710598
rect 296434 694094 297054 710042
rect 296434 693538 296466 694094
rect 297022 693538 297054 694094
rect 296434 658094 297054 693538
rect 296434 657538 296466 658094
rect 297022 657538 297054 658094
rect 296434 622094 297054 657538
rect 296434 621538 296466 622094
rect 297022 621538 297054 622094
rect 296434 586094 297054 621538
rect 296434 585538 296466 586094
rect 297022 585538 297054 586094
rect 296434 550094 297054 585538
rect 296434 549538 296466 550094
rect 297022 549538 297054 550094
rect 296434 514094 297054 549538
rect 296434 513538 296466 514094
rect 297022 513538 297054 514094
rect 296434 478094 297054 513538
rect 296434 477538 296466 478094
rect 297022 477538 297054 478094
rect 296434 442094 297054 477538
rect 296434 441538 296466 442094
rect 297022 441538 297054 442094
rect 296434 406094 297054 441538
rect 296434 405538 296466 406094
rect 297022 405538 297054 406094
rect 296434 370094 297054 405538
rect 296434 369538 296466 370094
rect 297022 369538 297054 370094
rect 296434 334094 297054 369538
rect 296434 333538 296466 334094
rect 297022 333538 297054 334094
rect 296434 298094 297054 333538
rect 296434 297538 296466 298094
rect 297022 297538 297054 298094
rect 296434 262094 297054 297538
rect 296434 261538 296466 262094
rect 297022 261538 297054 262094
rect 296434 226094 297054 261538
rect 296434 225538 296466 226094
rect 297022 225538 297054 226094
rect 296434 190094 297054 225538
rect 296434 189538 296466 190094
rect 297022 189538 297054 190094
rect 296434 154094 297054 189538
rect 296434 153538 296466 154094
rect 297022 153538 297054 154094
rect 296434 118094 297054 153538
rect 296434 117538 296466 118094
rect 297022 117538 297054 118094
rect 296434 82094 297054 117538
rect 296434 81538 296466 82094
rect 297022 81538 297054 82094
rect 296434 46094 297054 81538
rect 296434 45538 296466 46094
rect 297022 45538 297054 46094
rect 296434 10094 297054 45538
rect 296434 9538 296466 10094
rect 297022 9538 297054 10094
rect 296434 -6106 297054 9538
rect 296434 -6662 296466 -6106
rect 297022 -6662 297054 -6106
rect 296434 -7654 297054 -6662
rect 297674 711558 298294 711590
rect 297674 711002 297706 711558
rect 298262 711002 298294 711558
rect 297674 695334 298294 711002
rect 297674 694778 297706 695334
rect 298262 694778 298294 695334
rect 297674 659334 298294 694778
rect 297674 658778 297706 659334
rect 298262 658778 298294 659334
rect 297674 623334 298294 658778
rect 297674 622778 297706 623334
rect 298262 622778 298294 623334
rect 297674 587334 298294 622778
rect 297674 586778 297706 587334
rect 298262 586778 298294 587334
rect 297674 551334 298294 586778
rect 297674 550778 297706 551334
rect 298262 550778 298294 551334
rect 297674 515334 298294 550778
rect 297674 514778 297706 515334
rect 298262 514778 298294 515334
rect 297674 479334 298294 514778
rect 297674 478778 297706 479334
rect 298262 478778 298294 479334
rect 297674 443334 298294 478778
rect 297674 442778 297706 443334
rect 298262 442778 298294 443334
rect 297674 407334 298294 442778
rect 297674 406778 297706 407334
rect 298262 406778 298294 407334
rect 297674 371334 298294 406778
rect 297674 370778 297706 371334
rect 298262 370778 298294 371334
rect 297674 335334 298294 370778
rect 297674 334778 297706 335334
rect 298262 334778 298294 335334
rect 297674 299334 298294 334778
rect 297674 298778 297706 299334
rect 298262 298778 298294 299334
rect 297674 263334 298294 298778
rect 297674 262778 297706 263334
rect 298262 262778 298294 263334
rect 297674 227334 298294 262778
rect 297674 226778 297706 227334
rect 298262 226778 298294 227334
rect 297674 191334 298294 226778
rect 297674 190778 297706 191334
rect 298262 190778 298294 191334
rect 297674 155334 298294 190778
rect 297674 154778 297706 155334
rect 298262 154778 298294 155334
rect 297674 119334 298294 154778
rect 297674 118778 297706 119334
rect 298262 118778 298294 119334
rect 297674 83334 298294 118778
rect 297674 82778 297706 83334
rect 298262 82778 298294 83334
rect 297674 47334 298294 82778
rect 297674 46778 297706 47334
rect 298262 46778 298294 47334
rect 297674 11334 298294 46778
rect 297674 10778 297706 11334
rect 298262 10778 298294 11334
rect 297674 -7066 298294 10778
rect 297674 -7622 297706 -7066
rect 298262 -7622 298294 -7066
rect 297674 -7654 298294 -7622
rect 324994 704838 325614 711590
rect 324994 704282 325026 704838
rect 325582 704282 325614 704838
rect 324994 686654 325614 704282
rect 324994 686098 325026 686654
rect 325582 686098 325614 686654
rect 324994 650654 325614 686098
rect 324994 650098 325026 650654
rect 325582 650098 325614 650654
rect 324994 614654 325614 650098
rect 324994 614098 325026 614654
rect 325582 614098 325614 614654
rect 324994 578654 325614 614098
rect 324994 578098 325026 578654
rect 325582 578098 325614 578654
rect 324994 542654 325614 578098
rect 324994 542098 325026 542654
rect 325582 542098 325614 542654
rect 324994 506654 325614 542098
rect 324994 506098 325026 506654
rect 325582 506098 325614 506654
rect 324994 470654 325614 506098
rect 324994 470098 325026 470654
rect 325582 470098 325614 470654
rect 324994 434654 325614 470098
rect 324994 434098 325026 434654
rect 325582 434098 325614 434654
rect 324994 398654 325614 434098
rect 324994 398098 325026 398654
rect 325582 398098 325614 398654
rect 324994 362654 325614 398098
rect 324994 362098 325026 362654
rect 325582 362098 325614 362654
rect 324994 326654 325614 362098
rect 324994 326098 325026 326654
rect 325582 326098 325614 326654
rect 324994 290654 325614 326098
rect 324994 290098 325026 290654
rect 325582 290098 325614 290654
rect 324994 254654 325614 290098
rect 324994 254098 325026 254654
rect 325582 254098 325614 254654
rect 324994 218654 325614 254098
rect 324994 218098 325026 218654
rect 325582 218098 325614 218654
rect 324994 182654 325614 218098
rect 324994 182098 325026 182654
rect 325582 182098 325614 182654
rect 324994 146654 325614 182098
rect 324994 146098 325026 146654
rect 325582 146098 325614 146654
rect 324994 110654 325614 146098
rect 324994 110098 325026 110654
rect 325582 110098 325614 110654
rect 324994 74654 325614 110098
rect 324994 74098 325026 74654
rect 325582 74098 325614 74654
rect 324994 38654 325614 74098
rect 324994 38098 325026 38654
rect 325582 38098 325614 38654
rect 324994 2654 325614 38098
rect 324994 2098 325026 2654
rect 325582 2098 325614 2654
rect 324994 -346 325614 2098
rect 324994 -902 325026 -346
rect 325582 -902 325614 -346
rect 324994 -7654 325614 -902
rect 326234 705798 326854 711590
rect 326234 705242 326266 705798
rect 326822 705242 326854 705798
rect 326234 687894 326854 705242
rect 326234 687338 326266 687894
rect 326822 687338 326854 687894
rect 326234 651894 326854 687338
rect 326234 651338 326266 651894
rect 326822 651338 326854 651894
rect 326234 615894 326854 651338
rect 326234 615338 326266 615894
rect 326822 615338 326854 615894
rect 326234 579894 326854 615338
rect 326234 579338 326266 579894
rect 326822 579338 326854 579894
rect 326234 543894 326854 579338
rect 326234 543338 326266 543894
rect 326822 543338 326854 543894
rect 326234 507894 326854 543338
rect 326234 507338 326266 507894
rect 326822 507338 326854 507894
rect 326234 471894 326854 507338
rect 326234 471338 326266 471894
rect 326822 471338 326854 471894
rect 326234 435894 326854 471338
rect 326234 435338 326266 435894
rect 326822 435338 326854 435894
rect 326234 399894 326854 435338
rect 326234 399338 326266 399894
rect 326822 399338 326854 399894
rect 326234 363894 326854 399338
rect 326234 363338 326266 363894
rect 326822 363338 326854 363894
rect 326234 327894 326854 363338
rect 326234 327338 326266 327894
rect 326822 327338 326854 327894
rect 326234 291894 326854 327338
rect 326234 291338 326266 291894
rect 326822 291338 326854 291894
rect 326234 255894 326854 291338
rect 326234 255338 326266 255894
rect 326822 255338 326854 255894
rect 326234 219894 326854 255338
rect 326234 219338 326266 219894
rect 326822 219338 326854 219894
rect 326234 183894 326854 219338
rect 326234 183338 326266 183894
rect 326822 183338 326854 183894
rect 326234 147894 326854 183338
rect 326234 147338 326266 147894
rect 326822 147338 326854 147894
rect 326234 111894 326854 147338
rect 326234 111338 326266 111894
rect 326822 111338 326854 111894
rect 326234 75894 326854 111338
rect 326234 75338 326266 75894
rect 326822 75338 326854 75894
rect 326234 39894 326854 75338
rect 326234 39338 326266 39894
rect 326822 39338 326854 39894
rect 326234 3894 326854 39338
rect 326234 3338 326266 3894
rect 326822 3338 326854 3894
rect 326234 -1306 326854 3338
rect 326234 -1862 326266 -1306
rect 326822 -1862 326854 -1306
rect 326234 -7654 326854 -1862
rect 327474 706758 328094 711590
rect 327474 706202 327506 706758
rect 328062 706202 328094 706758
rect 327474 689134 328094 706202
rect 327474 688578 327506 689134
rect 328062 688578 328094 689134
rect 327474 653134 328094 688578
rect 327474 652578 327506 653134
rect 328062 652578 328094 653134
rect 327474 617134 328094 652578
rect 327474 616578 327506 617134
rect 328062 616578 328094 617134
rect 327474 581134 328094 616578
rect 327474 580578 327506 581134
rect 328062 580578 328094 581134
rect 327474 545134 328094 580578
rect 327474 544578 327506 545134
rect 328062 544578 328094 545134
rect 327474 509134 328094 544578
rect 327474 508578 327506 509134
rect 328062 508578 328094 509134
rect 327474 473134 328094 508578
rect 327474 472578 327506 473134
rect 328062 472578 328094 473134
rect 327474 437134 328094 472578
rect 327474 436578 327506 437134
rect 328062 436578 328094 437134
rect 327474 401134 328094 436578
rect 327474 400578 327506 401134
rect 328062 400578 328094 401134
rect 327474 365134 328094 400578
rect 327474 364578 327506 365134
rect 328062 364578 328094 365134
rect 327474 329134 328094 364578
rect 327474 328578 327506 329134
rect 328062 328578 328094 329134
rect 327474 293134 328094 328578
rect 327474 292578 327506 293134
rect 328062 292578 328094 293134
rect 327474 257134 328094 292578
rect 327474 256578 327506 257134
rect 328062 256578 328094 257134
rect 327474 221134 328094 256578
rect 327474 220578 327506 221134
rect 328062 220578 328094 221134
rect 327474 185134 328094 220578
rect 327474 184578 327506 185134
rect 328062 184578 328094 185134
rect 327474 149134 328094 184578
rect 327474 148578 327506 149134
rect 328062 148578 328094 149134
rect 327474 113134 328094 148578
rect 327474 112578 327506 113134
rect 328062 112578 328094 113134
rect 327474 77134 328094 112578
rect 327474 76578 327506 77134
rect 328062 76578 328094 77134
rect 327474 41134 328094 76578
rect 327474 40578 327506 41134
rect 328062 40578 328094 41134
rect 327474 5134 328094 40578
rect 327474 4578 327506 5134
rect 328062 4578 328094 5134
rect 327474 -2266 328094 4578
rect 327474 -2822 327506 -2266
rect 328062 -2822 328094 -2266
rect 327474 -7654 328094 -2822
rect 328714 707718 329334 711590
rect 328714 707162 328746 707718
rect 329302 707162 329334 707718
rect 328714 690374 329334 707162
rect 328714 689818 328746 690374
rect 329302 689818 329334 690374
rect 328714 654374 329334 689818
rect 328714 653818 328746 654374
rect 329302 653818 329334 654374
rect 328714 618374 329334 653818
rect 328714 617818 328746 618374
rect 329302 617818 329334 618374
rect 328714 582374 329334 617818
rect 328714 581818 328746 582374
rect 329302 581818 329334 582374
rect 328714 546374 329334 581818
rect 328714 545818 328746 546374
rect 329302 545818 329334 546374
rect 328714 510374 329334 545818
rect 328714 509818 328746 510374
rect 329302 509818 329334 510374
rect 328714 474374 329334 509818
rect 328714 473818 328746 474374
rect 329302 473818 329334 474374
rect 328714 438374 329334 473818
rect 328714 437818 328746 438374
rect 329302 437818 329334 438374
rect 328714 402374 329334 437818
rect 328714 401818 328746 402374
rect 329302 401818 329334 402374
rect 328714 366374 329334 401818
rect 328714 365818 328746 366374
rect 329302 365818 329334 366374
rect 328714 330374 329334 365818
rect 328714 329818 328746 330374
rect 329302 329818 329334 330374
rect 328714 294374 329334 329818
rect 328714 293818 328746 294374
rect 329302 293818 329334 294374
rect 328714 258374 329334 293818
rect 328714 257818 328746 258374
rect 329302 257818 329334 258374
rect 328714 222374 329334 257818
rect 328714 221818 328746 222374
rect 329302 221818 329334 222374
rect 328714 186374 329334 221818
rect 328714 185818 328746 186374
rect 329302 185818 329334 186374
rect 328714 150374 329334 185818
rect 328714 149818 328746 150374
rect 329302 149818 329334 150374
rect 328714 114374 329334 149818
rect 328714 113818 328746 114374
rect 329302 113818 329334 114374
rect 328714 78374 329334 113818
rect 328714 77818 328746 78374
rect 329302 77818 329334 78374
rect 328714 42374 329334 77818
rect 328714 41818 328746 42374
rect 329302 41818 329334 42374
rect 328714 6374 329334 41818
rect 328714 5818 328746 6374
rect 329302 5818 329334 6374
rect 328714 -3226 329334 5818
rect 328714 -3782 328746 -3226
rect 329302 -3782 329334 -3226
rect 328714 -7654 329334 -3782
rect 329954 708678 330574 711590
rect 329954 708122 329986 708678
rect 330542 708122 330574 708678
rect 329954 691614 330574 708122
rect 329954 691058 329986 691614
rect 330542 691058 330574 691614
rect 329954 655614 330574 691058
rect 329954 655058 329986 655614
rect 330542 655058 330574 655614
rect 329954 619614 330574 655058
rect 329954 619058 329986 619614
rect 330542 619058 330574 619614
rect 329954 583614 330574 619058
rect 329954 583058 329986 583614
rect 330542 583058 330574 583614
rect 329954 547614 330574 583058
rect 329954 547058 329986 547614
rect 330542 547058 330574 547614
rect 329954 511614 330574 547058
rect 329954 511058 329986 511614
rect 330542 511058 330574 511614
rect 329954 475614 330574 511058
rect 329954 475058 329986 475614
rect 330542 475058 330574 475614
rect 329954 439614 330574 475058
rect 329954 439058 329986 439614
rect 330542 439058 330574 439614
rect 329954 403614 330574 439058
rect 329954 403058 329986 403614
rect 330542 403058 330574 403614
rect 329954 367614 330574 403058
rect 329954 367058 329986 367614
rect 330542 367058 330574 367614
rect 329954 331614 330574 367058
rect 329954 331058 329986 331614
rect 330542 331058 330574 331614
rect 329954 295614 330574 331058
rect 329954 295058 329986 295614
rect 330542 295058 330574 295614
rect 329954 259614 330574 295058
rect 329954 259058 329986 259614
rect 330542 259058 330574 259614
rect 329954 223614 330574 259058
rect 329954 223058 329986 223614
rect 330542 223058 330574 223614
rect 329954 187614 330574 223058
rect 329954 187058 329986 187614
rect 330542 187058 330574 187614
rect 329954 151614 330574 187058
rect 329954 151058 329986 151614
rect 330542 151058 330574 151614
rect 329954 115614 330574 151058
rect 329954 115058 329986 115614
rect 330542 115058 330574 115614
rect 329954 79614 330574 115058
rect 329954 79058 329986 79614
rect 330542 79058 330574 79614
rect 329954 43614 330574 79058
rect 329954 43058 329986 43614
rect 330542 43058 330574 43614
rect 329954 7614 330574 43058
rect 329954 7058 329986 7614
rect 330542 7058 330574 7614
rect 329954 -4186 330574 7058
rect 329954 -4742 329986 -4186
rect 330542 -4742 330574 -4186
rect 329954 -7654 330574 -4742
rect 331194 709638 331814 711590
rect 331194 709082 331226 709638
rect 331782 709082 331814 709638
rect 331194 692854 331814 709082
rect 331194 692298 331226 692854
rect 331782 692298 331814 692854
rect 331194 656854 331814 692298
rect 331194 656298 331226 656854
rect 331782 656298 331814 656854
rect 331194 620854 331814 656298
rect 331194 620298 331226 620854
rect 331782 620298 331814 620854
rect 331194 584854 331814 620298
rect 331194 584298 331226 584854
rect 331782 584298 331814 584854
rect 331194 548854 331814 584298
rect 331194 548298 331226 548854
rect 331782 548298 331814 548854
rect 331194 512854 331814 548298
rect 331194 512298 331226 512854
rect 331782 512298 331814 512854
rect 331194 476854 331814 512298
rect 331194 476298 331226 476854
rect 331782 476298 331814 476854
rect 331194 440854 331814 476298
rect 331194 440298 331226 440854
rect 331782 440298 331814 440854
rect 331194 404854 331814 440298
rect 331194 404298 331226 404854
rect 331782 404298 331814 404854
rect 331194 368854 331814 404298
rect 331194 368298 331226 368854
rect 331782 368298 331814 368854
rect 331194 332854 331814 368298
rect 331194 332298 331226 332854
rect 331782 332298 331814 332854
rect 331194 296854 331814 332298
rect 331194 296298 331226 296854
rect 331782 296298 331814 296854
rect 331194 260854 331814 296298
rect 331194 260298 331226 260854
rect 331782 260298 331814 260854
rect 331194 224854 331814 260298
rect 331194 224298 331226 224854
rect 331782 224298 331814 224854
rect 331194 188854 331814 224298
rect 331194 188298 331226 188854
rect 331782 188298 331814 188854
rect 331194 152854 331814 188298
rect 331194 152298 331226 152854
rect 331782 152298 331814 152854
rect 331194 116854 331814 152298
rect 331194 116298 331226 116854
rect 331782 116298 331814 116854
rect 331194 80854 331814 116298
rect 331194 80298 331226 80854
rect 331782 80298 331814 80854
rect 331194 44854 331814 80298
rect 331194 44298 331226 44854
rect 331782 44298 331814 44854
rect 331194 8854 331814 44298
rect 331194 8298 331226 8854
rect 331782 8298 331814 8854
rect 331194 -5146 331814 8298
rect 331194 -5702 331226 -5146
rect 331782 -5702 331814 -5146
rect 331194 -7654 331814 -5702
rect 332434 710598 333054 711590
rect 332434 710042 332466 710598
rect 333022 710042 333054 710598
rect 332434 694094 333054 710042
rect 332434 693538 332466 694094
rect 333022 693538 333054 694094
rect 332434 658094 333054 693538
rect 332434 657538 332466 658094
rect 333022 657538 333054 658094
rect 332434 622094 333054 657538
rect 332434 621538 332466 622094
rect 333022 621538 333054 622094
rect 332434 586094 333054 621538
rect 332434 585538 332466 586094
rect 333022 585538 333054 586094
rect 332434 550094 333054 585538
rect 332434 549538 332466 550094
rect 333022 549538 333054 550094
rect 332434 514094 333054 549538
rect 332434 513538 332466 514094
rect 333022 513538 333054 514094
rect 332434 478094 333054 513538
rect 332434 477538 332466 478094
rect 333022 477538 333054 478094
rect 332434 442094 333054 477538
rect 332434 441538 332466 442094
rect 333022 441538 333054 442094
rect 332434 406094 333054 441538
rect 332434 405538 332466 406094
rect 333022 405538 333054 406094
rect 332434 370094 333054 405538
rect 332434 369538 332466 370094
rect 333022 369538 333054 370094
rect 332434 334094 333054 369538
rect 332434 333538 332466 334094
rect 333022 333538 333054 334094
rect 332434 298094 333054 333538
rect 332434 297538 332466 298094
rect 333022 297538 333054 298094
rect 332434 262094 333054 297538
rect 332434 261538 332466 262094
rect 333022 261538 333054 262094
rect 332434 226094 333054 261538
rect 332434 225538 332466 226094
rect 333022 225538 333054 226094
rect 332434 190094 333054 225538
rect 332434 189538 332466 190094
rect 333022 189538 333054 190094
rect 332434 154094 333054 189538
rect 332434 153538 332466 154094
rect 333022 153538 333054 154094
rect 332434 118094 333054 153538
rect 332434 117538 332466 118094
rect 333022 117538 333054 118094
rect 332434 82094 333054 117538
rect 332434 81538 332466 82094
rect 333022 81538 333054 82094
rect 332434 46094 333054 81538
rect 332434 45538 332466 46094
rect 333022 45538 333054 46094
rect 332434 10094 333054 45538
rect 332434 9538 332466 10094
rect 333022 9538 333054 10094
rect 332434 -6106 333054 9538
rect 332434 -6662 332466 -6106
rect 333022 -6662 333054 -6106
rect 332434 -7654 333054 -6662
rect 333674 711558 334294 711590
rect 333674 711002 333706 711558
rect 334262 711002 334294 711558
rect 333674 695334 334294 711002
rect 333674 694778 333706 695334
rect 334262 694778 334294 695334
rect 333674 659334 334294 694778
rect 333674 658778 333706 659334
rect 334262 658778 334294 659334
rect 333674 623334 334294 658778
rect 333674 622778 333706 623334
rect 334262 622778 334294 623334
rect 333674 587334 334294 622778
rect 333674 586778 333706 587334
rect 334262 586778 334294 587334
rect 333674 551334 334294 586778
rect 333674 550778 333706 551334
rect 334262 550778 334294 551334
rect 333674 515334 334294 550778
rect 333674 514778 333706 515334
rect 334262 514778 334294 515334
rect 333674 479334 334294 514778
rect 333674 478778 333706 479334
rect 334262 478778 334294 479334
rect 333674 443334 334294 478778
rect 333674 442778 333706 443334
rect 334262 442778 334294 443334
rect 333674 407334 334294 442778
rect 333674 406778 333706 407334
rect 334262 406778 334294 407334
rect 333674 371334 334294 406778
rect 333674 370778 333706 371334
rect 334262 370778 334294 371334
rect 333674 335334 334294 370778
rect 333674 334778 333706 335334
rect 334262 334778 334294 335334
rect 333674 299334 334294 334778
rect 333674 298778 333706 299334
rect 334262 298778 334294 299334
rect 333674 263334 334294 298778
rect 333674 262778 333706 263334
rect 334262 262778 334294 263334
rect 333674 227334 334294 262778
rect 333674 226778 333706 227334
rect 334262 226778 334294 227334
rect 333674 191334 334294 226778
rect 333674 190778 333706 191334
rect 334262 190778 334294 191334
rect 333674 155334 334294 190778
rect 333674 154778 333706 155334
rect 334262 154778 334294 155334
rect 333674 119334 334294 154778
rect 333674 118778 333706 119334
rect 334262 118778 334294 119334
rect 333674 83334 334294 118778
rect 333674 82778 333706 83334
rect 334262 82778 334294 83334
rect 333674 47334 334294 82778
rect 333674 46778 333706 47334
rect 334262 46778 334294 47334
rect 333674 11334 334294 46778
rect 333674 10778 333706 11334
rect 334262 10778 334294 11334
rect 333674 -7066 334294 10778
rect 333674 -7622 333706 -7066
rect 334262 -7622 334294 -7066
rect 333674 -7654 334294 -7622
rect 360994 704838 361614 711590
rect 360994 704282 361026 704838
rect 361582 704282 361614 704838
rect 360994 686654 361614 704282
rect 360994 686098 361026 686654
rect 361582 686098 361614 686654
rect 360994 650654 361614 686098
rect 360994 650098 361026 650654
rect 361582 650098 361614 650654
rect 360994 614654 361614 650098
rect 360994 614098 361026 614654
rect 361582 614098 361614 614654
rect 360994 578654 361614 614098
rect 360994 578098 361026 578654
rect 361582 578098 361614 578654
rect 360994 542654 361614 578098
rect 360994 542098 361026 542654
rect 361582 542098 361614 542654
rect 360994 506654 361614 542098
rect 360994 506098 361026 506654
rect 361582 506098 361614 506654
rect 360994 470654 361614 506098
rect 360994 470098 361026 470654
rect 361582 470098 361614 470654
rect 360994 434654 361614 470098
rect 360994 434098 361026 434654
rect 361582 434098 361614 434654
rect 360994 398654 361614 434098
rect 360994 398098 361026 398654
rect 361582 398098 361614 398654
rect 360994 362654 361614 398098
rect 360994 362098 361026 362654
rect 361582 362098 361614 362654
rect 360994 326654 361614 362098
rect 360994 326098 361026 326654
rect 361582 326098 361614 326654
rect 360994 290654 361614 326098
rect 360994 290098 361026 290654
rect 361582 290098 361614 290654
rect 360994 254654 361614 290098
rect 360994 254098 361026 254654
rect 361582 254098 361614 254654
rect 360994 218654 361614 254098
rect 360994 218098 361026 218654
rect 361582 218098 361614 218654
rect 360994 182654 361614 218098
rect 360994 182098 361026 182654
rect 361582 182098 361614 182654
rect 360994 146654 361614 182098
rect 360994 146098 361026 146654
rect 361582 146098 361614 146654
rect 360994 110654 361614 146098
rect 360994 110098 361026 110654
rect 361582 110098 361614 110654
rect 360994 74654 361614 110098
rect 360994 74098 361026 74654
rect 361582 74098 361614 74654
rect 360994 38654 361614 74098
rect 360994 38098 361026 38654
rect 361582 38098 361614 38654
rect 360994 2654 361614 38098
rect 360994 2098 361026 2654
rect 361582 2098 361614 2654
rect 360994 -346 361614 2098
rect 360994 -902 361026 -346
rect 361582 -902 361614 -346
rect 360994 -7654 361614 -902
rect 362234 705798 362854 711590
rect 362234 705242 362266 705798
rect 362822 705242 362854 705798
rect 362234 687894 362854 705242
rect 362234 687338 362266 687894
rect 362822 687338 362854 687894
rect 362234 651894 362854 687338
rect 362234 651338 362266 651894
rect 362822 651338 362854 651894
rect 362234 615894 362854 651338
rect 362234 615338 362266 615894
rect 362822 615338 362854 615894
rect 362234 579894 362854 615338
rect 362234 579338 362266 579894
rect 362822 579338 362854 579894
rect 362234 543894 362854 579338
rect 362234 543338 362266 543894
rect 362822 543338 362854 543894
rect 362234 507894 362854 543338
rect 362234 507338 362266 507894
rect 362822 507338 362854 507894
rect 362234 471894 362854 507338
rect 362234 471338 362266 471894
rect 362822 471338 362854 471894
rect 362234 435894 362854 471338
rect 362234 435338 362266 435894
rect 362822 435338 362854 435894
rect 362234 399894 362854 435338
rect 362234 399338 362266 399894
rect 362822 399338 362854 399894
rect 362234 363894 362854 399338
rect 362234 363338 362266 363894
rect 362822 363338 362854 363894
rect 362234 327894 362854 363338
rect 362234 327338 362266 327894
rect 362822 327338 362854 327894
rect 362234 291894 362854 327338
rect 362234 291338 362266 291894
rect 362822 291338 362854 291894
rect 362234 255894 362854 291338
rect 362234 255338 362266 255894
rect 362822 255338 362854 255894
rect 362234 219894 362854 255338
rect 362234 219338 362266 219894
rect 362822 219338 362854 219894
rect 362234 183894 362854 219338
rect 362234 183338 362266 183894
rect 362822 183338 362854 183894
rect 362234 147894 362854 183338
rect 362234 147338 362266 147894
rect 362822 147338 362854 147894
rect 362234 111894 362854 147338
rect 362234 111338 362266 111894
rect 362822 111338 362854 111894
rect 362234 75894 362854 111338
rect 362234 75338 362266 75894
rect 362822 75338 362854 75894
rect 362234 39894 362854 75338
rect 362234 39338 362266 39894
rect 362822 39338 362854 39894
rect 362234 3894 362854 39338
rect 362234 3338 362266 3894
rect 362822 3338 362854 3894
rect 362234 -1306 362854 3338
rect 362234 -1862 362266 -1306
rect 362822 -1862 362854 -1306
rect 362234 -7654 362854 -1862
rect 363474 706758 364094 711590
rect 363474 706202 363506 706758
rect 364062 706202 364094 706758
rect 363474 689134 364094 706202
rect 363474 688578 363506 689134
rect 364062 688578 364094 689134
rect 363474 653134 364094 688578
rect 363474 652578 363506 653134
rect 364062 652578 364094 653134
rect 363474 617134 364094 652578
rect 363474 616578 363506 617134
rect 364062 616578 364094 617134
rect 363474 581134 364094 616578
rect 363474 580578 363506 581134
rect 364062 580578 364094 581134
rect 363474 545134 364094 580578
rect 363474 544578 363506 545134
rect 364062 544578 364094 545134
rect 363474 509134 364094 544578
rect 363474 508578 363506 509134
rect 364062 508578 364094 509134
rect 363474 473134 364094 508578
rect 363474 472578 363506 473134
rect 364062 472578 364094 473134
rect 363474 437134 364094 472578
rect 363474 436578 363506 437134
rect 364062 436578 364094 437134
rect 363474 401134 364094 436578
rect 363474 400578 363506 401134
rect 364062 400578 364094 401134
rect 363474 365134 364094 400578
rect 363474 364578 363506 365134
rect 364062 364578 364094 365134
rect 363474 329134 364094 364578
rect 363474 328578 363506 329134
rect 364062 328578 364094 329134
rect 363474 293134 364094 328578
rect 363474 292578 363506 293134
rect 364062 292578 364094 293134
rect 363474 257134 364094 292578
rect 363474 256578 363506 257134
rect 364062 256578 364094 257134
rect 363474 221134 364094 256578
rect 363474 220578 363506 221134
rect 364062 220578 364094 221134
rect 363474 185134 364094 220578
rect 363474 184578 363506 185134
rect 364062 184578 364094 185134
rect 363474 149134 364094 184578
rect 363474 148578 363506 149134
rect 364062 148578 364094 149134
rect 363474 113134 364094 148578
rect 363474 112578 363506 113134
rect 364062 112578 364094 113134
rect 363474 77134 364094 112578
rect 363474 76578 363506 77134
rect 364062 76578 364094 77134
rect 363474 41134 364094 76578
rect 363474 40578 363506 41134
rect 364062 40578 364094 41134
rect 363474 5134 364094 40578
rect 363474 4578 363506 5134
rect 364062 4578 364094 5134
rect 363474 -2266 364094 4578
rect 363474 -2822 363506 -2266
rect 364062 -2822 364094 -2266
rect 363474 -7654 364094 -2822
rect 364714 707718 365334 711590
rect 364714 707162 364746 707718
rect 365302 707162 365334 707718
rect 364714 690374 365334 707162
rect 364714 689818 364746 690374
rect 365302 689818 365334 690374
rect 364714 654374 365334 689818
rect 364714 653818 364746 654374
rect 365302 653818 365334 654374
rect 364714 618374 365334 653818
rect 364714 617818 364746 618374
rect 365302 617818 365334 618374
rect 364714 582374 365334 617818
rect 364714 581818 364746 582374
rect 365302 581818 365334 582374
rect 364714 546374 365334 581818
rect 364714 545818 364746 546374
rect 365302 545818 365334 546374
rect 364714 510374 365334 545818
rect 364714 509818 364746 510374
rect 365302 509818 365334 510374
rect 364714 474374 365334 509818
rect 364714 473818 364746 474374
rect 365302 473818 365334 474374
rect 364714 438374 365334 473818
rect 364714 437818 364746 438374
rect 365302 437818 365334 438374
rect 364714 402374 365334 437818
rect 364714 401818 364746 402374
rect 365302 401818 365334 402374
rect 364714 366374 365334 401818
rect 364714 365818 364746 366374
rect 365302 365818 365334 366374
rect 364714 330374 365334 365818
rect 364714 329818 364746 330374
rect 365302 329818 365334 330374
rect 364714 294374 365334 329818
rect 364714 293818 364746 294374
rect 365302 293818 365334 294374
rect 364714 258374 365334 293818
rect 364714 257818 364746 258374
rect 365302 257818 365334 258374
rect 364714 222374 365334 257818
rect 364714 221818 364746 222374
rect 365302 221818 365334 222374
rect 364714 186374 365334 221818
rect 364714 185818 364746 186374
rect 365302 185818 365334 186374
rect 364714 150374 365334 185818
rect 364714 149818 364746 150374
rect 365302 149818 365334 150374
rect 364714 114374 365334 149818
rect 364714 113818 364746 114374
rect 365302 113818 365334 114374
rect 364714 78374 365334 113818
rect 364714 77818 364746 78374
rect 365302 77818 365334 78374
rect 364714 42374 365334 77818
rect 364714 41818 364746 42374
rect 365302 41818 365334 42374
rect 364714 6374 365334 41818
rect 364714 5818 364746 6374
rect 365302 5818 365334 6374
rect 364714 -3226 365334 5818
rect 364714 -3782 364746 -3226
rect 365302 -3782 365334 -3226
rect 364714 -7654 365334 -3782
rect 365954 708678 366574 711590
rect 365954 708122 365986 708678
rect 366542 708122 366574 708678
rect 365954 691614 366574 708122
rect 365954 691058 365986 691614
rect 366542 691058 366574 691614
rect 365954 655614 366574 691058
rect 365954 655058 365986 655614
rect 366542 655058 366574 655614
rect 365954 619614 366574 655058
rect 365954 619058 365986 619614
rect 366542 619058 366574 619614
rect 365954 583614 366574 619058
rect 365954 583058 365986 583614
rect 366542 583058 366574 583614
rect 365954 547614 366574 583058
rect 365954 547058 365986 547614
rect 366542 547058 366574 547614
rect 365954 511614 366574 547058
rect 365954 511058 365986 511614
rect 366542 511058 366574 511614
rect 365954 475614 366574 511058
rect 365954 475058 365986 475614
rect 366542 475058 366574 475614
rect 365954 439614 366574 475058
rect 365954 439058 365986 439614
rect 366542 439058 366574 439614
rect 365954 403614 366574 439058
rect 365954 403058 365986 403614
rect 366542 403058 366574 403614
rect 365954 367614 366574 403058
rect 365954 367058 365986 367614
rect 366542 367058 366574 367614
rect 365954 331614 366574 367058
rect 365954 331058 365986 331614
rect 366542 331058 366574 331614
rect 365954 295614 366574 331058
rect 365954 295058 365986 295614
rect 366542 295058 366574 295614
rect 365954 259614 366574 295058
rect 365954 259058 365986 259614
rect 366542 259058 366574 259614
rect 365954 223614 366574 259058
rect 365954 223058 365986 223614
rect 366542 223058 366574 223614
rect 365954 187614 366574 223058
rect 365954 187058 365986 187614
rect 366542 187058 366574 187614
rect 365954 151614 366574 187058
rect 365954 151058 365986 151614
rect 366542 151058 366574 151614
rect 365954 115614 366574 151058
rect 365954 115058 365986 115614
rect 366542 115058 366574 115614
rect 365954 79614 366574 115058
rect 365954 79058 365986 79614
rect 366542 79058 366574 79614
rect 365954 43614 366574 79058
rect 365954 43058 365986 43614
rect 366542 43058 366574 43614
rect 365954 7614 366574 43058
rect 365954 7058 365986 7614
rect 366542 7058 366574 7614
rect 365954 -4186 366574 7058
rect 365954 -4742 365986 -4186
rect 366542 -4742 366574 -4186
rect 365954 -7654 366574 -4742
rect 367194 709638 367814 711590
rect 367194 709082 367226 709638
rect 367782 709082 367814 709638
rect 367194 692854 367814 709082
rect 367194 692298 367226 692854
rect 367782 692298 367814 692854
rect 367194 656854 367814 692298
rect 367194 656298 367226 656854
rect 367782 656298 367814 656854
rect 367194 620854 367814 656298
rect 367194 620298 367226 620854
rect 367782 620298 367814 620854
rect 367194 584854 367814 620298
rect 367194 584298 367226 584854
rect 367782 584298 367814 584854
rect 367194 548854 367814 584298
rect 367194 548298 367226 548854
rect 367782 548298 367814 548854
rect 367194 512854 367814 548298
rect 367194 512298 367226 512854
rect 367782 512298 367814 512854
rect 367194 476854 367814 512298
rect 367194 476298 367226 476854
rect 367782 476298 367814 476854
rect 367194 440854 367814 476298
rect 367194 440298 367226 440854
rect 367782 440298 367814 440854
rect 367194 404854 367814 440298
rect 367194 404298 367226 404854
rect 367782 404298 367814 404854
rect 367194 368854 367814 404298
rect 367194 368298 367226 368854
rect 367782 368298 367814 368854
rect 367194 332854 367814 368298
rect 367194 332298 367226 332854
rect 367782 332298 367814 332854
rect 367194 296854 367814 332298
rect 367194 296298 367226 296854
rect 367782 296298 367814 296854
rect 367194 260854 367814 296298
rect 367194 260298 367226 260854
rect 367782 260298 367814 260854
rect 367194 224854 367814 260298
rect 367194 224298 367226 224854
rect 367782 224298 367814 224854
rect 367194 188854 367814 224298
rect 367194 188298 367226 188854
rect 367782 188298 367814 188854
rect 367194 152854 367814 188298
rect 367194 152298 367226 152854
rect 367782 152298 367814 152854
rect 367194 116854 367814 152298
rect 367194 116298 367226 116854
rect 367782 116298 367814 116854
rect 367194 80854 367814 116298
rect 367194 80298 367226 80854
rect 367782 80298 367814 80854
rect 367194 44854 367814 80298
rect 367194 44298 367226 44854
rect 367782 44298 367814 44854
rect 367194 8854 367814 44298
rect 367194 8298 367226 8854
rect 367782 8298 367814 8854
rect 367194 -5146 367814 8298
rect 367194 -5702 367226 -5146
rect 367782 -5702 367814 -5146
rect 367194 -7654 367814 -5702
rect 368434 710598 369054 711590
rect 368434 710042 368466 710598
rect 369022 710042 369054 710598
rect 368434 694094 369054 710042
rect 368434 693538 368466 694094
rect 369022 693538 369054 694094
rect 368434 658094 369054 693538
rect 368434 657538 368466 658094
rect 369022 657538 369054 658094
rect 368434 622094 369054 657538
rect 368434 621538 368466 622094
rect 369022 621538 369054 622094
rect 368434 586094 369054 621538
rect 368434 585538 368466 586094
rect 369022 585538 369054 586094
rect 368434 550094 369054 585538
rect 368434 549538 368466 550094
rect 369022 549538 369054 550094
rect 368434 514094 369054 549538
rect 368434 513538 368466 514094
rect 369022 513538 369054 514094
rect 368434 478094 369054 513538
rect 368434 477538 368466 478094
rect 369022 477538 369054 478094
rect 368434 442094 369054 477538
rect 368434 441538 368466 442094
rect 369022 441538 369054 442094
rect 368434 406094 369054 441538
rect 368434 405538 368466 406094
rect 369022 405538 369054 406094
rect 368434 370094 369054 405538
rect 368434 369538 368466 370094
rect 369022 369538 369054 370094
rect 368434 334094 369054 369538
rect 368434 333538 368466 334094
rect 369022 333538 369054 334094
rect 368434 298094 369054 333538
rect 368434 297538 368466 298094
rect 369022 297538 369054 298094
rect 368434 262094 369054 297538
rect 368434 261538 368466 262094
rect 369022 261538 369054 262094
rect 368434 226094 369054 261538
rect 368434 225538 368466 226094
rect 369022 225538 369054 226094
rect 368434 190094 369054 225538
rect 368434 189538 368466 190094
rect 369022 189538 369054 190094
rect 368434 154094 369054 189538
rect 368434 153538 368466 154094
rect 369022 153538 369054 154094
rect 368434 118094 369054 153538
rect 368434 117538 368466 118094
rect 369022 117538 369054 118094
rect 368434 82094 369054 117538
rect 368434 81538 368466 82094
rect 369022 81538 369054 82094
rect 368434 46094 369054 81538
rect 368434 45538 368466 46094
rect 369022 45538 369054 46094
rect 368434 10094 369054 45538
rect 368434 9538 368466 10094
rect 369022 9538 369054 10094
rect 368434 -6106 369054 9538
rect 368434 -6662 368466 -6106
rect 369022 -6662 369054 -6106
rect 368434 -7654 369054 -6662
rect 369674 711558 370294 711590
rect 369674 711002 369706 711558
rect 370262 711002 370294 711558
rect 369674 695334 370294 711002
rect 369674 694778 369706 695334
rect 370262 694778 370294 695334
rect 369674 659334 370294 694778
rect 369674 658778 369706 659334
rect 370262 658778 370294 659334
rect 369674 623334 370294 658778
rect 369674 622778 369706 623334
rect 370262 622778 370294 623334
rect 369674 587334 370294 622778
rect 369674 586778 369706 587334
rect 370262 586778 370294 587334
rect 369674 551334 370294 586778
rect 369674 550778 369706 551334
rect 370262 550778 370294 551334
rect 369674 515334 370294 550778
rect 369674 514778 369706 515334
rect 370262 514778 370294 515334
rect 369674 479334 370294 514778
rect 369674 478778 369706 479334
rect 370262 478778 370294 479334
rect 369674 443334 370294 478778
rect 369674 442778 369706 443334
rect 370262 442778 370294 443334
rect 369674 407334 370294 442778
rect 369674 406778 369706 407334
rect 370262 406778 370294 407334
rect 369674 371334 370294 406778
rect 369674 370778 369706 371334
rect 370262 370778 370294 371334
rect 369674 335334 370294 370778
rect 369674 334778 369706 335334
rect 370262 334778 370294 335334
rect 369674 299334 370294 334778
rect 369674 298778 369706 299334
rect 370262 298778 370294 299334
rect 369674 263334 370294 298778
rect 369674 262778 369706 263334
rect 370262 262778 370294 263334
rect 369674 227334 370294 262778
rect 369674 226778 369706 227334
rect 370262 226778 370294 227334
rect 369674 191334 370294 226778
rect 369674 190778 369706 191334
rect 370262 190778 370294 191334
rect 369674 155334 370294 190778
rect 369674 154778 369706 155334
rect 370262 154778 370294 155334
rect 369674 119334 370294 154778
rect 369674 118778 369706 119334
rect 370262 118778 370294 119334
rect 369674 83334 370294 118778
rect 369674 82778 369706 83334
rect 370262 82778 370294 83334
rect 369674 47334 370294 82778
rect 369674 46778 369706 47334
rect 370262 46778 370294 47334
rect 369674 11334 370294 46778
rect 369674 10778 369706 11334
rect 370262 10778 370294 11334
rect 369674 -7066 370294 10778
rect 369674 -7622 369706 -7066
rect 370262 -7622 370294 -7066
rect 369674 -7654 370294 -7622
rect 396994 704838 397614 711590
rect 396994 704282 397026 704838
rect 397582 704282 397614 704838
rect 396994 686654 397614 704282
rect 396994 686098 397026 686654
rect 397582 686098 397614 686654
rect 396994 650654 397614 686098
rect 396994 650098 397026 650654
rect 397582 650098 397614 650654
rect 396994 614654 397614 650098
rect 396994 614098 397026 614654
rect 397582 614098 397614 614654
rect 396994 578654 397614 614098
rect 396994 578098 397026 578654
rect 397582 578098 397614 578654
rect 396994 542654 397614 578098
rect 396994 542098 397026 542654
rect 397582 542098 397614 542654
rect 396994 506654 397614 542098
rect 396994 506098 397026 506654
rect 397582 506098 397614 506654
rect 396994 470654 397614 506098
rect 396994 470098 397026 470654
rect 397582 470098 397614 470654
rect 396994 434654 397614 470098
rect 396994 434098 397026 434654
rect 397582 434098 397614 434654
rect 396994 398654 397614 434098
rect 396994 398098 397026 398654
rect 397582 398098 397614 398654
rect 396994 362654 397614 398098
rect 396994 362098 397026 362654
rect 397582 362098 397614 362654
rect 396994 326654 397614 362098
rect 396994 326098 397026 326654
rect 397582 326098 397614 326654
rect 396994 290654 397614 326098
rect 396994 290098 397026 290654
rect 397582 290098 397614 290654
rect 396994 254654 397614 290098
rect 396994 254098 397026 254654
rect 397582 254098 397614 254654
rect 396994 218654 397614 254098
rect 396994 218098 397026 218654
rect 397582 218098 397614 218654
rect 396994 182654 397614 218098
rect 396994 182098 397026 182654
rect 397582 182098 397614 182654
rect 396994 146654 397614 182098
rect 396994 146098 397026 146654
rect 397582 146098 397614 146654
rect 396994 110654 397614 146098
rect 396994 110098 397026 110654
rect 397582 110098 397614 110654
rect 396994 74654 397614 110098
rect 396994 74098 397026 74654
rect 397582 74098 397614 74654
rect 396994 38654 397614 74098
rect 396994 38098 397026 38654
rect 397582 38098 397614 38654
rect 396994 2654 397614 38098
rect 396994 2098 397026 2654
rect 397582 2098 397614 2654
rect 396994 -346 397614 2098
rect 396994 -902 397026 -346
rect 397582 -902 397614 -346
rect 396994 -7654 397614 -902
rect 398234 705798 398854 711590
rect 398234 705242 398266 705798
rect 398822 705242 398854 705798
rect 398234 687894 398854 705242
rect 398234 687338 398266 687894
rect 398822 687338 398854 687894
rect 398234 651894 398854 687338
rect 398234 651338 398266 651894
rect 398822 651338 398854 651894
rect 398234 615894 398854 651338
rect 398234 615338 398266 615894
rect 398822 615338 398854 615894
rect 398234 579894 398854 615338
rect 398234 579338 398266 579894
rect 398822 579338 398854 579894
rect 398234 543894 398854 579338
rect 398234 543338 398266 543894
rect 398822 543338 398854 543894
rect 398234 507894 398854 543338
rect 398234 507338 398266 507894
rect 398822 507338 398854 507894
rect 398234 471894 398854 507338
rect 398234 471338 398266 471894
rect 398822 471338 398854 471894
rect 398234 435894 398854 471338
rect 398234 435338 398266 435894
rect 398822 435338 398854 435894
rect 398234 399894 398854 435338
rect 398234 399338 398266 399894
rect 398822 399338 398854 399894
rect 398234 363894 398854 399338
rect 398234 363338 398266 363894
rect 398822 363338 398854 363894
rect 398234 327894 398854 363338
rect 398234 327338 398266 327894
rect 398822 327338 398854 327894
rect 398234 291894 398854 327338
rect 398234 291338 398266 291894
rect 398822 291338 398854 291894
rect 398234 255894 398854 291338
rect 398234 255338 398266 255894
rect 398822 255338 398854 255894
rect 398234 219894 398854 255338
rect 398234 219338 398266 219894
rect 398822 219338 398854 219894
rect 398234 183894 398854 219338
rect 398234 183338 398266 183894
rect 398822 183338 398854 183894
rect 398234 147894 398854 183338
rect 398234 147338 398266 147894
rect 398822 147338 398854 147894
rect 398234 111894 398854 147338
rect 398234 111338 398266 111894
rect 398822 111338 398854 111894
rect 398234 75894 398854 111338
rect 398234 75338 398266 75894
rect 398822 75338 398854 75894
rect 398234 39894 398854 75338
rect 398234 39338 398266 39894
rect 398822 39338 398854 39894
rect 398234 3894 398854 39338
rect 398234 3338 398266 3894
rect 398822 3338 398854 3894
rect 398234 -1306 398854 3338
rect 398234 -1862 398266 -1306
rect 398822 -1862 398854 -1306
rect 398234 -7654 398854 -1862
rect 399474 706758 400094 711590
rect 399474 706202 399506 706758
rect 400062 706202 400094 706758
rect 399474 689134 400094 706202
rect 399474 688578 399506 689134
rect 400062 688578 400094 689134
rect 399474 653134 400094 688578
rect 399474 652578 399506 653134
rect 400062 652578 400094 653134
rect 399474 617134 400094 652578
rect 399474 616578 399506 617134
rect 400062 616578 400094 617134
rect 399474 581134 400094 616578
rect 399474 580578 399506 581134
rect 400062 580578 400094 581134
rect 399474 545134 400094 580578
rect 399474 544578 399506 545134
rect 400062 544578 400094 545134
rect 399474 509134 400094 544578
rect 399474 508578 399506 509134
rect 400062 508578 400094 509134
rect 399474 473134 400094 508578
rect 399474 472578 399506 473134
rect 400062 472578 400094 473134
rect 399474 437134 400094 472578
rect 399474 436578 399506 437134
rect 400062 436578 400094 437134
rect 399474 401134 400094 436578
rect 399474 400578 399506 401134
rect 400062 400578 400094 401134
rect 399474 365134 400094 400578
rect 399474 364578 399506 365134
rect 400062 364578 400094 365134
rect 399474 329134 400094 364578
rect 399474 328578 399506 329134
rect 400062 328578 400094 329134
rect 399474 293134 400094 328578
rect 399474 292578 399506 293134
rect 400062 292578 400094 293134
rect 399474 257134 400094 292578
rect 399474 256578 399506 257134
rect 400062 256578 400094 257134
rect 399474 221134 400094 256578
rect 399474 220578 399506 221134
rect 400062 220578 400094 221134
rect 399474 185134 400094 220578
rect 399474 184578 399506 185134
rect 400062 184578 400094 185134
rect 399474 149134 400094 184578
rect 399474 148578 399506 149134
rect 400062 148578 400094 149134
rect 399474 113134 400094 148578
rect 399474 112578 399506 113134
rect 400062 112578 400094 113134
rect 399474 77134 400094 112578
rect 399474 76578 399506 77134
rect 400062 76578 400094 77134
rect 399474 41134 400094 76578
rect 399474 40578 399506 41134
rect 400062 40578 400094 41134
rect 399474 5134 400094 40578
rect 399474 4578 399506 5134
rect 400062 4578 400094 5134
rect 399474 -2266 400094 4578
rect 399474 -2822 399506 -2266
rect 400062 -2822 400094 -2266
rect 399474 -7654 400094 -2822
rect 400714 707718 401334 711590
rect 400714 707162 400746 707718
rect 401302 707162 401334 707718
rect 400714 690374 401334 707162
rect 400714 689818 400746 690374
rect 401302 689818 401334 690374
rect 400714 654374 401334 689818
rect 400714 653818 400746 654374
rect 401302 653818 401334 654374
rect 400714 618374 401334 653818
rect 400714 617818 400746 618374
rect 401302 617818 401334 618374
rect 400714 582374 401334 617818
rect 400714 581818 400746 582374
rect 401302 581818 401334 582374
rect 400714 546374 401334 581818
rect 400714 545818 400746 546374
rect 401302 545818 401334 546374
rect 400714 510374 401334 545818
rect 400714 509818 400746 510374
rect 401302 509818 401334 510374
rect 400714 474374 401334 509818
rect 400714 473818 400746 474374
rect 401302 473818 401334 474374
rect 400714 438374 401334 473818
rect 400714 437818 400746 438374
rect 401302 437818 401334 438374
rect 400714 402374 401334 437818
rect 400714 401818 400746 402374
rect 401302 401818 401334 402374
rect 400714 366374 401334 401818
rect 400714 365818 400746 366374
rect 401302 365818 401334 366374
rect 400714 330374 401334 365818
rect 400714 329818 400746 330374
rect 401302 329818 401334 330374
rect 400714 294374 401334 329818
rect 400714 293818 400746 294374
rect 401302 293818 401334 294374
rect 400714 258374 401334 293818
rect 400714 257818 400746 258374
rect 401302 257818 401334 258374
rect 400714 222374 401334 257818
rect 400714 221818 400746 222374
rect 401302 221818 401334 222374
rect 400714 186374 401334 221818
rect 400714 185818 400746 186374
rect 401302 185818 401334 186374
rect 400714 150374 401334 185818
rect 400714 149818 400746 150374
rect 401302 149818 401334 150374
rect 400714 114374 401334 149818
rect 400714 113818 400746 114374
rect 401302 113818 401334 114374
rect 400714 78374 401334 113818
rect 400714 77818 400746 78374
rect 401302 77818 401334 78374
rect 400714 42374 401334 77818
rect 400714 41818 400746 42374
rect 401302 41818 401334 42374
rect 400714 6374 401334 41818
rect 400714 5818 400746 6374
rect 401302 5818 401334 6374
rect 400714 -3226 401334 5818
rect 400714 -3782 400746 -3226
rect 401302 -3782 401334 -3226
rect 400714 -7654 401334 -3782
rect 401954 708678 402574 711590
rect 401954 708122 401986 708678
rect 402542 708122 402574 708678
rect 401954 691614 402574 708122
rect 401954 691058 401986 691614
rect 402542 691058 402574 691614
rect 401954 655614 402574 691058
rect 401954 655058 401986 655614
rect 402542 655058 402574 655614
rect 401954 619614 402574 655058
rect 401954 619058 401986 619614
rect 402542 619058 402574 619614
rect 401954 583614 402574 619058
rect 401954 583058 401986 583614
rect 402542 583058 402574 583614
rect 401954 547614 402574 583058
rect 401954 547058 401986 547614
rect 402542 547058 402574 547614
rect 401954 511614 402574 547058
rect 401954 511058 401986 511614
rect 402542 511058 402574 511614
rect 401954 475614 402574 511058
rect 401954 475058 401986 475614
rect 402542 475058 402574 475614
rect 401954 439614 402574 475058
rect 401954 439058 401986 439614
rect 402542 439058 402574 439614
rect 401954 403614 402574 439058
rect 401954 403058 401986 403614
rect 402542 403058 402574 403614
rect 401954 367614 402574 403058
rect 401954 367058 401986 367614
rect 402542 367058 402574 367614
rect 401954 331614 402574 367058
rect 401954 331058 401986 331614
rect 402542 331058 402574 331614
rect 401954 295614 402574 331058
rect 401954 295058 401986 295614
rect 402542 295058 402574 295614
rect 401954 259614 402574 295058
rect 401954 259058 401986 259614
rect 402542 259058 402574 259614
rect 401954 223614 402574 259058
rect 401954 223058 401986 223614
rect 402542 223058 402574 223614
rect 401954 187614 402574 223058
rect 401954 187058 401986 187614
rect 402542 187058 402574 187614
rect 401954 151614 402574 187058
rect 401954 151058 401986 151614
rect 402542 151058 402574 151614
rect 401954 115614 402574 151058
rect 401954 115058 401986 115614
rect 402542 115058 402574 115614
rect 401954 79614 402574 115058
rect 401954 79058 401986 79614
rect 402542 79058 402574 79614
rect 401954 43614 402574 79058
rect 401954 43058 401986 43614
rect 402542 43058 402574 43614
rect 401954 7614 402574 43058
rect 401954 7058 401986 7614
rect 402542 7058 402574 7614
rect 401954 -4186 402574 7058
rect 401954 -4742 401986 -4186
rect 402542 -4742 402574 -4186
rect 401954 -7654 402574 -4742
rect 403194 709638 403814 711590
rect 403194 709082 403226 709638
rect 403782 709082 403814 709638
rect 403194 692854 403814 709082
rect 403194 692298 403226 692854
rect 403782 692298 403814 692854
rect 403194 656854 403814 692298
rect 403194 656298 403226 656854
rect 403782 656298 403814 656854
rect 403194 620854 403814 656298
rect 403194 620298 403226 620854
rect 403782 620298 403814 620854
rect 403194 584854 403814 620298
rect 403194 584298 403226 584854
rect 403782 584298 403814 584854
rect 403194 548854 403814 584298
rect 403194 548298 403226 548854
rect 403782 548298 403814 548854
rect 403194 512854 403814 548298
rect 403194 512298 403226 512854
rect 403782 512298 403814 512854
rect 403194 476854 403814 512298
rect 403194 476298 403226 476854
rect 403782 476298 403814 476854
rect 403194 440854 403814 476298
rect 403194 440298 403226 440854
rect 403782 440298 403814 440854
rect 403194 404854 403814 440298
rect 403194 404298 403226 404854
rect 403782 404298 403814 404854
rect 403194 368854 403814 404298
rect 403194 368298 403226 368854
rect 403782 368298 403814 368854
rect 403194 332854 403814 368298
rect 403194 332298 403226 332854
rect 403782 332298 403814 332854
rect 403194 296854 403814 332298
rect 403194 296298 403226 296854
rect 403782 296298 403814 296854
rect 403194 260854 403814 296298
rect 403194 260298 403226 260854
rect 403782 260298 403814 260854
rect 403194 224854 403814 260298
rect 403194 224298 403226 224854
rect 403782 224298 403814 224854
rect 403194 188854 403814 224298
rect 403194 188298 403226 188854
rect 403782 188298 403814 188854
rect 403194 152854 403814 188298
rect 403194 152298 403226 152854
rect 403782 152298 403814 152854
rect 403194 116854 403814 152298
rect 403194 116298 403226 116854
rect 403782 116298 403814 116854
rect 403194 80854 403814 116298
rect 403194 80298 403226 80854
rect 403782 80298 403814 80854
rect 403194 44854 403814 80298
rect 403194 44298 403226 44854
rect 403782 44298 403814 44854
rect 403194 8854 403814 44298
rect 403194 8298 403226 8854
rect 403782 8298 403814 8854
rect 403194 -5146 403814 8298
rect 403194 -5702 403226 -5146
rect 403782 -5702 403814 -5146
rect 403194 -7654 403814 -5702
rect 404434 710598 405054 711590
rect 404434 710042 404466 710598
rect 405022 710042 405054 710598
rect 404434 694094 405054 710042
rect 404434 693538 404466 694094
rect 405022 693538 405054 694094
rect 404434 658094 405054 693538
rect 404434 657538 404466 658094
rect 405022 657538 405054 658094
rect 404434 622094 405054 657538
rect 404434 621538 404466 622094
rect 405022 621538 405054 622094
rect 404434 586094 405054 621538
rect 404434 585538 404466 586094
rect 405022 585538 405054 586094
rect 404434 550094 405054 585538
rect 404434 549538 404466 550094
rect 405022 549538 405054 550094
rect 404434 514094 405054 549538
rect 404434 513538 404466 514094
rect 405022 513538 405054 514094
rect 404434 478094 405054 513538
rect 404434 477538 404466 478094
rect 405022 477538 405054 478094
rect 404434 442094 405054 477538
rect 404434 441538 404466 442094
rect 405022 441538 405054 442094
rect 404434 406094 405054 441538
rect 404434 405538 404466 406094
rect 405022 405538 405054 406094
rect 404434 370094 405054 405538
rect 404434 369538 404466 370094
rect 405022 369538 405054 370094
rect 404434 334094 405054 369538
rect 404434 333538 404466 334094
rect 405022 333538 405054 334094
rect 404434 298094 405054 333538
rect 404434 297538 404466 298094
rect 405022 297538 405054 298094
rect 404434 262094 405054 297538
rect 404434 261538 404466 262094
rect 405022 261538 405054 262094
rect 404434 226094 405054 261538
rect 404434 225538 404466 226094
rect 405022 225538 405054 226094
rect 404434 190094 405054 225538
rect 404434 189538 404466 190094
rect 405022 189538 405054 190094
rect 404434 154094 405054 189538
rect 404434 153538 404466 154094
rect 405022 153538 405054 154094
rect 404434 118094 405054 153538
rect 404434 117538 404466 118094
rect 405022 117538 405054 118094
rect 404434 82094 405054 117538
rect 404434 81538 404466 82094
rect 405022 81538 405054 82094
rect 404434 46094 405054 81538
rect 404434 45538 404466 46094
rect 405022 45538 405054 46094
rect 404434 10094 405054 45538
rect 404434 9538 404466 10094
rect 405022 9538 405054 10094
rect 404434 -6106 405054 9538
rect 404434 -6662 404466 -6106
rect 405022 -6662 405054 -6106
rect 404434 -7654 405054 -6662
rect 405674 711558 406294 711590
rect 405674 711002 405706 711558
rect 406262 711002 406294 711558
rect 405674 695334 406294 711002
rect 405674 694778 405706 695334
rect 406262 694778 406294 695334
rect 405674 659334 406294 694778
rect 405674 658778 405706 659334
rect 406262 658778 406294 659334
rect 405674 623334 406294 658778
rect 405674 622778 405706 623334
rect 406262 622778 406294 623334
rect 405674 587334 406294 622778
rect 405674 586778 405706 587334
rect 406262 586778 406294 587334
rect 405674 551334 406294 586778
rect 405674 550778 405706 551334
rect 406262 550778 406294 551334
rect 405674 515334 406294 550778
rect 405674 514778 405706 515334
rect 406262 514778 406294 515334
rect 405674 479334 406294 514778
rect 405674 478778 405706 479334
rect 406262 478778 406294 479334
rect 405674 443334 406294 478778
rect 405674 442778 405706 443334
rect 406262 442778 406294 443334
rect 405674 407334 406294 442778
rect 405674 406778 405706 407334
rect 406262 406778 406294 407334
rect 405674 371334 406294 406778
rect 405674 370778 405706 371334
rect 406262 370778 406294 371334
rect 405674 335334 406294 370778
rect 405674 334778 405706 335334
rect 406262 334778 406294 335334
rect 405674 299334 406294 334778
rect 405674 298778 405706 299334
rect 406262 298778 406294 299334
rect 405674 263334 406294 298778
rect 405674 262778 405706 263334
rect 406262 262778 406294 263334
rect 405674 227334 406294 262778
rect 405674 226778 405706 227334
rect 406262 226778 406294 227334
rect 405674 191334 406294 226778
rect 405674 190778 405706 191334
rect 406262 190778 406294 191334
rect 405674 155334 406294 190778
rect 405674 154778 405706 155334
rect 406262 154778 406294 155334
rect 405674 119334 406294 154778
rect 405674 118778 405706 119334
rect 406262 118778 406294 119334
rect 405674 83334 406294 118778
rect 405674 82778 405706 83334
rect 406262 82778 406294 83334
rect 405674 47334 406294 82778
rect 405674 46778 405706 47334
rect 406262 46778 406294 47334
rect 405674 11334 406294 46778
rect 405674 10778 405706 11334
rect 406262 10778 406294 11334
rect 405674 -7066 406294 10778
rect 405674 -7622 405706 -7066
rect 406262 -7622 406294 -7066
rect 405674 -7654 406294 -7622
rect 432994 704838 433614 711590
rect 432994 704282 433026 704838
rect 433582 704282 433614 704838
rect 432994 686654 433614 704282
rect 432994 686098 433026 686654
rect 433582 686098 433614 686654
rect 432994 650654 433614 686098
rect 432994 650098 433026 650654
rect 433582 650098 433614 650654
rect 432994 614654 433614 650098
rect 432994 614098 433026 614654
rect 433582 614098 433614 614654
rect 432994 578654 433614 614098
rect 432994 578098 433026 578654
rect 433582 578098 433614 578654
rect 432994 542654 433614 578098
rect 432994 542098 433026 542654
rect 433582 542098 433614 542654
rect 432994 506654 433614 542098
rect 432994 506098 433026 506654
rect 433582 506098 433614 506654
rect 432994 470654 433614 506098
rect 432994 470098 433026 470654
rect 433582 470098 433614 470654
rect 432994 434654 433614 470098
rect 432994 434098 433026 434654
rect 433582 434098 433614 434654
rect 432994 398654 433614 434098
rect 432994 398098 433026 398654
rect 433582 398098 433614 398654
rect 432994 362654 433614 398098
rect 432994 362098 433026 362654
rect 433582 362098 433614 362654
rect 432994 326654 433614 362098
rect 432994 326098 433026 326654
rect 433582 326098 433614 326654
rect 432994 290654 433614 326098
rect 432994 290098 433026 290654
rect 433582 290098 433614 290654
rect 432994 254654 433614 290098
rect 432994 254098 433026 254654
rect 433582 254098 433614 254654
rect 432994 218654 433614 254098
rect 432994 218098 433026 218654
rect 433582 218098 433614 218654
rect 432994 182654 433614 218098
rect 432994 182098 433026 182654
rect 433582 182098 433614 182654
rect 432994 146654 433614 182098
rect 432994 146098 433026 146654
rect 433582 146098 433614 146654
rect 432994 110654 433614 146098
rect 432994 110098 433026 110654
rect 433582 110098 433614 110654
rect 432994 74654 433614 110098
rect 432994 74098 433026 74654
rect 433582 74098 433614 74654
rect 432994 38654 433614 74098
rect 432994 38098 433026 38654
rect 433582 38098 433614 38654
rect 432994 2654 433614 38098
rect 432994 2098 433026 2654
rect 433582 2098 433614 2654
rect 432994 -346 433614 2098
rect 432994 -902 433026 -346
rect 433582 -902 433614 -346
rect 432994 -7654 433614 -902
rect 434234 705798 434854 711590
rect 434234 705242 434266 705798
rect 434822 705242 434854 705798
rect 434234 687894 434854 705242
rect 434234 687338 434266 687894
rect 434822 687338 434854 687894
rect 434234 651894 434854 687338
rect 434234 651338 434266 651894
rect 434822 651338 434854 651894
rect 434234 615894 434854 651338
rect 434234 615338 434266 615894
rect 434822 615338 434854 615894
rect 434234 579894 434854 615338
rect 434234 579338 434266 579894
rect 434822 579338 434854 579894
rect 434234 543894 434854 579338
rect 434234 543338 434266 543894
rect 434822 543338 434854 543894
rect 434234 507894 434854 543338
rect 434234 507338 434266 507894
rect 434822 507338 434854 507894
rect 434234 471894 434854 507338
rect 434234 471338 434266 471894
rect 434822 471338 434854 471894
rect 434234 435894 434854 471338
rect 434234 435338 434266 435894
rect 434822 435338 434854 435894
rect 434234 399894 434854 435338
rect 434234 399338 434266 399894
rect 434822 399338 434854 399894
rect 434234 363894 434854 399338
rect 434234 363338 434266 363894
rect 434822 363338 434854 363894
rect 434234 327894 434854 363338
rect 434234 327338 434266 327894
rect 434822 327338 434854 327894
rect 434234 291894 434854 327338
rect 434234 291338 434266 291894
rect 434822 291338 434854 291894
rect 434234 255894 434854 291338
rect 434234 255338 434266 255894
rect 434822 255338 434854 255894
rect 434234 219894 434854 255338
rect 434234 219338 434266 219894
rect 434822 219338 434854 219894
rect 434234 183894 434854 219338
rect 434234 183338 434266 183894
rect 434822 183338 434854 183894
rect 434234 147894 434854 183338
rect 434234 147338 434266 147894
rect 434822 147338 434854 147894
rect 434234 111894 434854 147338
rect 434234 111338 434266 111894
rect 434822 111338 434854 111894
rect 434234 75894 434854 111338
rect 434234 75338 434266 75894
rect 434822 75338 434854 75894
rect 434234 39894 434854 75338
rect 434234 39338 434266 39894
rect 434822 39338 434854 39894
rect 434234 3894 434854 39338
rect 434234 3338 434266 3894
rect 434822 3338 434854 3894
rect 434234 -1306 434854 3338
rect 434234 -1862 434266 -1306
rect 434822 -1862 434854 -1306
rect 434234 -7654 434854 -1862
rect 435474 706758 436094 711590
rect 435474 706202 435506 706758
rect 436062 706202 436094 706758
rect 435474 689134 436094 706202
rect 435474 688578 435506 689134
rect 436062 688578 436094 689134
rect 435474 653134 436094 688578
rect 435474 652578 435506 653134
rect 436062 652578 436094 653134
rect 435474 617134 436094 652578
rect 435474 616578 435506 617134
rect 436062 616578 436094 617134
rect 435474 581134 436094 616578
rect 435474 580578 435506 581134
rect 436062 580578 436094 581134
rect 435474 545134 436094 580578
rect 435474 544578 435506 545134
rect 436062 544578 436094 545134
rect 435474 509134 436094 544578
rect 435474 508578 435506 509134
rect 436062 508578 436094 509134
rect 435474 473134 436094 508578
rect 435474 472578 435506 473134
rect 436062 472578 436094 473134
rect 435474 437134 436094 472578
rect 435474 436578 435506 437134
rect 436062 436578 436094 437134
rect 435474 401134 436094 436578
rect 435474 400578 435506 401134
rect 436062 400578 436094 401134
rect 435474 365134 436094 400578
rect 435474 364578 435506 365134
rect 436062 364578 436094 365134
rect 435474 329134 436094 364578
rect 435474 328578 435506 329134
rect 436062 328578 436094 329134
rect 435474 293134 436094 328578
rect 435474 292578 435506 293134
rect 436062 292578 436094 293134
rect 435474 257134 436094 292578
rect 435474 256578 435506 257134
rect 436062 256578 436094 257134
rect 435474 221134 436094 256578
rect 435474 220578 435506 221134
rect 436062 220578 436094 221134
rect 435474 185134 436094 220578
rect 435474 184578 435506 185134
rect 436062 184578 436094 185134
rect 435474 149134 436094 184578
rect 435474 148578 435506 149134
rect 436062 148578 436094 149134
rect 435474 113134 436094 148578
rect 435474 112578 435506 113134
rect 436062 112578 436094 113134
rect 435474 77134 436094 112578
rect 435474 76578 435506 77134
rect 436062 76578 436094 77134
rect 435474 41134 436094 76578
rect 435474 40578 435506 41134
rect 436062 40578 436094 41134
rect 435474 5134 436094 40578
rect 435474 4578 435506 5134
rect 436062 4578 436094 5134
rect 435474 -2266 436094 4578
rect 435474 -2822 435506 -2266
rect 436062 -2822 436094 -2266
rect 435474 -7654 436094 -2822
rect 436714 707718 437334 711590
rect 436714 707162 436746 707718
rect 437302 707162 437334 707718
rect 436714 690374 437334 707162
rect 436714 689818 436746 690374
rect 437302 689818 437334 690374
rect 436714 654374 437334 689818
rect 436714 653818 436746 654374
rect 437302 653818 437334 654374
rect 436714 618374 437334 653818
rect 436714 617818 436746 618374
rect 437302 617818 437334 618374
rect 436714 582374 437334 617818
rect 436714 581818 436746 582374
rect 437302 581818 437334 582374
rect 436714 546374 437334 581818
rect 436714 545818 436746 546374
rect 437302 545818 437334 546374
rect 436714 510374 437334 545818
rect 436714 509818 436746 510374
rect 437302 509818 437334 510374
rect 436714 474374 437334 509818
rect 436714 473818 436746 474374
rect 437302 473818 437334 474374
rect 436714 438374 437334 473818
rect 436714 437818 436746 438374
rect 437302 437818 437334 438374
rect 436714 402374 437334 437818
rect 436714 401818 436746 402374
rect 437302 401818 437334 402374
rect 436714 366374 437334 401818
rect 436714 365818 436746 366374
rect 437302 365818 437334 366374
rect 436714 330374 437334 365818
rect 436714 329818 436746 330374
rect 437302 329818 437334 330374
rect 436714 294374 437334 329818
rect 436714 293818 436746 294374
rect 437302 293818 437334 294374
rect 436714 258374 437334 293818
rect 436714 257818 436746 258374
rect 437302 257818 437334 258374
rect 436714 222374 437334 257818
rect 436714 221818 436746 222374
rect 437302 221818 437334 222374
rect 436714 186374 437334 221818
rect 436714 185818 436746 186374
rect 437302 185818 437334 186374
rect 436714 150374 437334 185818
rect 436714 149818 436746 150374
rect 437302 149818 437334 150374
rect 436714 114374 437334 149818
rect 436714 113818 436746 114374
rect 437302 113818 437334 114374
rect 436714 78374 437334 113818
rect 436714 77818 436746 78374
rect 437302 77818 437334 78374
rect 436714 42374 437334 77818
rect 436714 41818 436746 42374
rect 437302 41818 437334 42374
rect 436714 6374 437334 41818
rect 436714 5818 436746 6374
rect 437302 5818 437334 6374
rect 436714 -3226 437334 5818
rect 436714 -3782 436746 -3226
rect 437302 -3782 437334 -3226
rect 436714 -7654 437334 -3782
rect 437954 708678 438574 711590
rect 437954 708122 437986 708678
rect 438542 708122 438574 708678
rect 437954 691614 438574 708122
rect 437954 691058 437986 691614
rect 438542 691058 438574 691614
rect 437954 655614 438574 691058
rect 437954 655058 437986 655614
rect 438542 655058 438574 655614
rect 437954 619614 438574 655058
rect 437954 619058 437986 619614
rect 438542 619058 438574 619614
rect 437954 583614 438574 619058
rect 437954 583058 437986 583614
rect 438542 583058 438574 583614
rect 437954 547614 438574 583058
rect 437954 547058 437986 547614
rect 438542 547058 438574 547614
rect 437954 511614 438574 547058
rect 437954 511058 437986 511614
rect 438542 511058 438574 511614
rect 437954 475614 438574 511058
rect 437954 475058 437986 475614
rect 438542 475058 438574 475614
rect 437954 439614 438574 475058
rect 437954 439058 437986 439614
rect 438542 439058 438574 439614
rect 437954 403614 438574 439058
rect 437954 403058 437986 403614
rect 438542 403058 438574 403614
rect 437954 367614 438574 403058
rect 437954 367058 437986 367614
rect 438542 367058 438574 367614
rect 437954 331614 438574 367058
rect 437954 331058 437986 331614
rect 438542 331058 438574 331614
rect 437954 295614 438574 331058
rect 437954 295058 437986 295614
rect 438542 295058 438574 295614
rect 437954 259614 438574 295058
rect 437954 259058 437986 259614
rect 438542 259058 438574 259614
rect 437954 223614 438574 259058
rect 437954 223058 437986 223614
rect 438542 223058 438574 223614
rect 437954 187614 438574 223058
rect 437954 187058 437986 187614
rect 438542 187058 438574 187614
rect 437954 151614 438574 187058
rect 437954 151058 437986 151614
rect 438542 151058 438574 151614
rect 437954 115614 438574 151058
rect 437954 115058 437986 115614
rect 438542 115058 438574 115614
rect 437954 79614 438574 115058
rect 437954 79058 437986 79614
rect 438542 79058 438574 79614
rect 437954 43614 438574 79058
rect 437954 43058 437986 43614
rect 438542 43058 438574 43614
rect 437954 7614 438574 43058
rect 437954 7058 437986 7614
rect 438542 7058 438574 7614
rect 437954 -4186 438574 7058
rect 437954 -4742 437986 -4186
rect 438542 -4742 438574 -4186
rect 437954 -7654 438574 -4742
rect 439194 709638 439814 711590
rect 439194 709082 439226 709638
rect 439782 709082 439814 709638
rect 439194 692854 439814 709082
rect 439194 692298 439226 692854
rect 439782 692298 439814 692854
rect 439194 656854 439814 692298
rect 439194 656298 439226 656854
rect 439782 656298 439814 656854
rect 439194 620854 439814 656298
rect 439194 620298 439226 620854
rect 439782 620298 439814 620854
rect 439194 584854 439814 620298
rect 439194 584298 439226 584854
rect 439782 584298 439814 584854
rect 439194 548854 439814 584298
rect 439194 548298 439226 548854
rect 439782 548298 439814 548854
rect 439194 512854 439814 548298
rect 439194 512298 439226 512854
rect 439782 512298 439814 512854
rect 439194 476854 439814 512298
rect 439194 476298 439226 476854
rect 439782 476298 439814 476854
rect 439194 440854 439814 476298
rect 439194 440298 439226 440854
rect 439782 440298 439814 440854
rect 439194 404854 439814 440298
rect 439194 404298 439226 404854
rect 439782 404298 439814 404854
rect 439194 368854 439814 404298
rect 439194 368298 439226 368854
rect 439782 368298 439814 368854
rect 439194 332854 439814 368298
rect 439194 332298 439226 332854
rect 439782 332298 439814 332854
rect 439194 296854 439814 332298
rect 439194 296298 439226 296854
rect 439782 296298 439814 296854
rect 439194 260854 439814 296298
rect 439194 260298 439226 260854
rect 439782 260298 439814 260854
rect 439194 224854 439814 260298
rect 439194 224298 439226 224854
rect 439782 224298 439814 224854
rect 439194 188854 439814 224298
rect 439194 188298 439226 188854
rect 439782 188298 439814 188854
rect 439194 152854 439814 188298
rect 439194 152298 439226 152854
rect 439782 152298 439814 152854
rect 439194 116854 439814 152298
rect 439194 116298 439226 116854
rect 439782 116298 439814 116854
rect 439194 80854 439814 116298
rect 439194 80298 439226 80854
rect 439782 80298 439814 80854
rect 439194 44854 439814 80298
rect 439194 44298 439226 44854
rect 439782 44298 439814 44854
rect 439194 8854 439814 44298
rect 439194 8298 439226 8854
rect 439782 8298 439814 8854
rect 439194 -5146 439814 8298
rect 439194 -5702 439226 -5146
rect 439782 -5702 439814 -5146
rect 439194 -7654 439814 -5702
rect 440434 710598 441054 711590
rect 440434 710042 440466 710598
rect 441022 710042 441054 710598
rect 440434 694094 441054 710042
rect 440434 693538 440466 694094
rect 441022 693538 441054 694094
rect 440434 658094 441054 693538
rect 440434 657538 440466 658094
rect 441022 657538 441054 658094
rect 440434 622094 441054 657538
rect 440434 621538 440466 622094
rect 441022 621538 441054 622094
rect 440434 586094 441054 621538
rect 440434 585538 440466 586094
rect 441022 585538 441054 586094
rect 440434 550094 441054 585538
rect 440434 549538 440466 550094
rect 441022 549538 441054 550094
rect 440434 514094 441054 549538
rect 440434 513538 440466 514094
rect 441022 513538 441054 514094
rect 440434 478094 441054 513538
rect 440434 477538 440466 478094
rect 441022 477538 441054 478094
rect 440434 442094 441054 477538
rect 440434 441538 440466 442094
rect 441022 441538 441054 442094
rect 440434 406094 441054 441538
rect 440434 405538 440466 406094
rect 441022 405538 441054 406094
rect 440434 370094 441054 405538
rect 440434 369538 440466 370094
rect 441022 369538 441054 370094
rect 440434 334094 441054 369538
rect 440434 333538 440466 334094
rect 441022 333538 441054 334094
rect 440434 298094 441054 333538
rect 440434 297538 440466 298094
rect 441022 297538 441054 298094
rect 440434 262094 441054 297538
rect 440434 261538 440466 262094
rect 441022 261538 441054 262094
rect 440434 226094 441054 261538
rect 440434 225538 440466 226094
rect 441022 225538 441054 226094
rect 440434 190094 441054 225538
rect 440434 189538 440466 190094
rect 441022 189538 441054 190094
rect 440434 154094 441054 189538
rect 440434 153538 440466 154094
rect 441022 153538 441054 154094
rect 440434 118094 441054 153538
rect 440434 117538 440466 118094
rect 441022 117538 441054 118094
rect 440434 82094 441054 117538
rect 440434 81538 440466 82094
rect 441022 81538 441054 82094
rect 440434 46094 441054 81538
rect 440434 45538 440466 46094
rect 441022 45538 441054 46094
rect 440434 10094 441054 45538
rect 440434 9538 440466 10094
rect 441022 9538 441054 10094
rect 440434 -6106 441054 9538
rect 440434 -6662 440466 -6106
rect 441022 -6662 441054 -6106
rect 440434 -7654 441054 -6662
rect 441674 711558 442294 711590
rect 441674 711002 441706 711558
rect 442262 711002 442294 711558
rect 441674 695334 442294 711002
rect 441674 694778 441706 695334
rect 442262 694778 442294 695334
rect 441674 659334 442294 694778
rect 441674 658778 441706 659334
rect 442262 658778 442294 659334
rect 441674 623334 442294 658778
rect 441674 622778 441706 623334
rect 442262 622778 442294 623334
rect 441674 587334 442294 622778
rect 441674 586778 441706 587334
rect 442262 586778 442294 587334
rect 441674 551334 442294 586778
rect 441674 550778 441706 551334
rect 442262 550778 442294 551334
rect 441674 515334 442294 550778
rect 441674 514778 441706 515334
rect 442262 514778 442294 515334
rect 441674 479334 442294 514778
rect 441674 478778 441706 479334
rect 442262 478778 442294 479334
rect 441674 443334 442294 478778
rect 441674 442778 441706 443334
rect 442262 442778 442294 443334
rect 441674 407334 442294 442778
rect 441674 406778 441706 407334
rect 442262 406778 442294 407334
rect 441674 371334 442294 406778
rect 441674 370778 441706 371334
rect 442262 370778 442294 371334
rect 441674 335334 442294 370778
rect 441674 334778 441706 335334
rect 442262 334778 442294 335334
rect 441674 299334 442294 334778
rect 441674 298778 441706 299334
rect 442262 298778 442294 299334
rect 441674 263334 442294 298778
rect 441674 262778 441706 263334
rect 442262 262778 442294 263334
rect 441674 227334 442294 262778
rect 441674 226778 441706 227334
rect 442262 226778 442294 227334
rect 441674 191334 442294 226778
rect 441674 190778 441706 191334
rect 442262 190778 442294 191334
rect 441674 155334 442294 190778
rect 441674 154778 441706 155334
rect 442262 154778 442294 155334
rect 441674 119334 442294 154778
rect 441674 118778 441706 119334
rect 442262 118778 442294 119334
rect 441674 83334 442294 118778
rect 441674 82778 441706 83334
rect 442262 82778 442294 83334
rect 441674 47334 442294 82778
rect 441674 46778 441706 47334
rect 442262 46778 442294 47334
rect 441674 11334 442294 46778
rect 441674 10778 441706 11334
rect 442262 10778 442294 11334
rect 441674 -7066 442294 10778
rect 441674 -7622 441706 -7066
rect 442262 -7622 442294 -7066
rect 441674 -7654 442294 -7622
rect 468994 704838 469614 711590
rect 468994 704282 469026 704838
rect 469582 704282 469614 704838
rect 468994 686654 469614 704282
rect 468994 686098 469026 686654
rect 469582 686098 469614 686654
rect 468994 650654 469614 686098
rect 468994 650098 469026 650654
rect 469582 650098 469614 650654
rect 468994 614654 469614 650098
rect 468994 614098 469026 614654
rect 469582 614098 469614 614654
rect 468994 578654 469614 614098
rect 468994 578098 469026 578654
rect 469582 578098 469614 578654
rect 468994 542654 469614 578098
rect 468994 542098 469026 542654
rect 469582 542098 469614 542654
rect 468994 506654 469614 542098
rect 468994 506098 469026 506654
rect 469582 506098 469614 506654
rect 468994 470654 469614 506098
rect 468994 470098 469026 470654
rect 469582 470098 469614 470654
rect 468994 450397 469614 470098
rect 468994 450093 469032 450397
rect 469576 450093 469614 450397
rect 468994 434654 469614 450093
rect 468994 434098 469026 434654
rect 469582 434098 469614 434654
rect 468994 431997 469614 434098
rect 468994 431693 469032 431997
rect 469576 431693 469614 431997
rect 468994 410998 469614 431693
rect 468994 410694 469032 410998
rect 469576 410694 469614 410998
rect 468994 398654 469614 410694
rect 468994 398098 469026 398654
rect 469582 398098 469614 398654
rect 468994 390002 469614 398098
rect 468994 389698 469032 390002
rect 469576 389698 469614 390002
rect 468994 362654 469614 389698
rect 468994 362098 469026 362654
rect 469582 362098 469614 362654
rect 468994 357399 469614 362098
rect 468994 357095 469032 357399
rect 469576 357095 469614 357399
rect 468994 341397 469614 357095
rect 468994 341093 469032 341397
rect 469576 341093 469614 341397
rect 468994 326654 469614 341093
rect 468994 326098 469026 326654
rect 469582 326098 469614 326654
rect 468994 321397 469614 326098
rect 468994 321093 469032 321397
rect 469576 321093 469614 321397
rect 468994 305999 469614 321093
rect 468994 305695 469032 305999
rect 469576 305695 469614 305999
rect 468994 290654 469614 305695
rect 468994 290098 469026 290654
rect 469582 290098 469614 290654
rect 468994 286400 469614 290098
rect 468994 286096 469032 286400
rect 469576 286096 469614 286400
rect 468994 266399 469614 286096
rect 468994 266095 469032 266399
rect 469576 266095 469614 266399
rect 468994 254654 469614 266095
rect 468994 254098 469026 254654
rect 469582 254098 469614 254654
rect 468994 218654 469614 254098
rect 468994 218098 469026 218654
rect 469582 218098 469614 218654
rect 468994 182654 469614 218098
rect 468994 182098 469026 182654
rect 469582 182098 469614 182654
rect 468994 146654 469614 182098
rect 468994 146098 469026 146654
rect 469582 146098 469614 146654
rect 468994 110654 469614 146098
rect 468994 110098 469026 110654
rect 469582 110098 469614 110654
rect 468994 74654 469614 110098
rect 468994 74098 469026 74654
rect 469582 74098 469614 74654
rect 468994 38654 469614 74098
rect 468994 38098 469026 38654
rect 469582 38098 469614 38654
rect 468994 2654 469614 38098
rect 468994 2098 469026 2654
rect 469582 2098 469614 2654
rect 468994 -346 469614 2098
rect 468994 -902 469026 -346
rect 469582 -902 469614 -346
rect 468994 -7654 469614 -902
rect 470234 705798 470854 711590
rect 470234 705242 470266 705798
rect 470822 705242 470854 705798
rect 470234 687894 470854 705242
rect 470234 687338 470266 687894
rect 470822 687338 470854 687894
rect 470234 651894 470854 687338
rect 470234 651338 470266 651894
rect 470822 651338 470854 651894
rect 470234 615894 470854 651338
rect 470234 615338 470266 615894
rect 470822 615338 470854 615894
rect 470234 579894 470854 615338
rect 470234 579338 470266 579894
rect 470822 579338 470854 579894
rect 470234 543894 470854 579338
rect 470234 543338 470266 543894
rect 470822 543338 470854 543894
rect 470234 507894 470854 543338
rect 470234 507338 470266 507894
rect 470822 507338 470854 507894
rect 470234 471894 470854 507338
rect 470234 471338 470266 471894
rect 470822 471338 470854 471894
rect 470234 451483 470854 471338
rect 470234 451179 470272 451483
rect 470816 451179 470854 451483
rect 470234 449312 470854 451179
rect 470234 449008 470272 449312
rect 470816 449008 470854 449312
rect 470234 435894 470854 449008
rect 470234 435338 470266 435894
rect 470822 435338 470854 435894
rect 470234 433084 470854 435338
rect 470234 432780 470272 433084
rect 470816 432780 470854 433084
rect 470234 430912 470854 432780
rect 470234 430608 470272 430912
rect 470816 430608 470854 430912
rect 470234 412084 470854 430608
rect 470234 411780 470272 412084
rect 470816 411780 470854 412084
rect 470234 409912 470854 411780
rect 470234 409608 470272 409912
rect 470816 409608 470854 409912
rect 470234 399894 470854 409608
rect 470234 399338 470266 399894
rect 470822 399338 470854 399894
rect 470234 391085 470854 399338
rect 470234 390781 470272 391085
rect 470816 390781 470854 391085
rect 470234 388912 470854 390781
rect 470234 388608 470272 388912
rect 470816 388608 470854 388912
rect 470234 363894 470854 388608
rect 470234 363338 470266 363894
rect 470822 363338 470854 363894
rect 470234 358485 470854 363338
rect 470234 358181 470272 358485
rect 470816 358181 470854 358485
rect 470234 356312 470854 358181
rect 470234 356008 470272 356312
rect 470816 356008 470854 356312
rect 470234 342484 470854 356008
rect 470234 342180 470272 342484
rect 470816 342180 470854 342484
rect 470234 340312 470854 342180
rect 470234 340008 470272 340312
rect 470816 340008 470854 340312
rect 470234 327894 470854 340008
rect 470234 327338 470266 327894
rect 470822 327338 470854 327894
rect 470234 322484 470854 327338
rect 470234 322180 470272 322484
rect 470816 322180 470854 322484
rect 470234 320312 470854 322180
rect 470234 320008 470272 320312
rect 470816 320008 470854 320312
rect 470234 307084 470854 320008
rect 470234 306780 470272 307084
rect 470816 306780 470854 307084
rect 470234 304912 470854 306780
rect 470234 304608 470272 304912
rect 470816 304608 470854 304912
rect 470234 291894 470854 304608
rect 470234 291338 470266 291894
rect 470822 291338 470854 291894
rect 470234 287485 470854 291338
rect 470234 287181 470272 287485
rect 470816 287181 470854 287485
rect 470234 285312 470854 287181
rect 470234 285008 470272 285312
rect 470816 285008 470854 285312
rect 470234 267485 470854 285008
rect 470234 267181 470272 267485
rect 470816 267181 470854 267485
rect 470234 265312 470854 267181
rect 470234 265008 470272 265312
rect 470816 265008 470854 265312
rect 470234 255894 470854 265008
rect 470234 255338 470266 255894
rect 470822 255338 470854 255894
rect 470234 219894 470854 255338
rect 470234 219338 470266 219894
rect 470822 219338 470854 219894
rect 470234 183894 470854 219338
rect 470234 183338 470266 183894
rect 470822 183338 470854 183894
rect 470234 147894 470854 183338
rect 470234 147338 470266 147894
rect 470822 147338 470854 147894
rect 470234 111894 470854 147338
rect 470234 111338 470266 111894
rect 470822 111338 470854 111894
rect 470234 75894 470854 111338
rect 470234 75338 470266 75894
rect 470822 75338 470854 75894
rect 470234 39894 470854 75338
rect 470234 39338 470266 39894
rect 470822 39338 470854 39894
rect 470234 3894 470854 39338
rect 470234 3338 470266 3894
rect 470822 3338 470854 3894
rect 470234 -1306 470854 3338
rect 470234 -1862 470266 -1306
rect 470822 -1862 470854 -1306
rect 470234 -7654 470854 -1862
rect 471474 706758 472094 711590
rect 471474 706202 471506 706758
rect 472062 706202 472094 706758
rect 471474 689134 472094 706202
rect 471474 688578 471506 689134
rect 472062 688578 472094 689134
rect 471474 653134 472094 688578
rect 471474 652578 471506 653134
rect 472062 652578 472094 653134
rect 471474 617134 472094 652578
rect 471474 616578 471506 617134
rect 472062 616578 472094 617134
rect 471474 581134 472094 616578
rect 471474 580578 471506 581134
rect 472062 580578 472094 581134
rect 471474 545134 472094 580578
rect 471474 544578 471506 545134
rect 472062 544578 472094 545134
rect 471474 509134 472094 544578
rect 471474 508578 471506 509134
rect 472062 508578 472094 509134
rect 471474 473134 472094 508578
rect 471474 472578 471506 473134
rect 472062 472578 472094 473134
rect 471474 437134 472094 472578
rect 471474 436578 471506 437134
rect 472062 436578 472094 437134
rect 471474 401134 472094 436578
rect 471474 400578 471506 401134
rect 472062 400578 472094 401134
rect 471474 365134 472094 400578
rect 471474 364578 471506 365134
rect 472062 364578 472094 365134
rect 471474 329134 472094 364578
rect 472714 707718 473334 711590
rect 472714 707162 472746 707718
rect 473302 707162 473334 707718
rect 472714 690374 473334 707162
rect 472714 689818 472746 690374
rect 473302 689818 473334 690374
rect 472714 654374 473334 689818
rect 472714 653818 472746 654374
rect 473302 653818 473334 654374
rect 472714 618374 473334 653818
rect 472714 617818 472746 618374
rect 473302 617818 473334 618374
rect 472714 582374 473334 617818
rect 472714 581818 472746 582374
rect 473302 581818 473334 582374
rect 472714 546374 473334 581818
rect 472714 545818 472746 546374
rect 473302 545818 473334 546374
rect 472714 510374 473334 545818
rect 472714 509818 472746 510374
rect 473302 509818 473334 510374
rect 472714 474374 473334 509818
rect 472714 473818 472746 474374
rect 473302 473818 473334 474374
rect 472714 438374 473334 473818
rect 473954 708678 474574 711590
rect 473954 708122 473986 708678
rect 474542 708122 474574 708678
rect 473954 691614 474574 708122
rect 473954 691058 473986 691614
rect 474542 691058 474574 691614
rect 473954 655614 474574 691058
rect 473954 655058 473986 655614
rect 474542 655058 474574 655614
rect 473954 619614 474574 655058
rect 473954 619058 473986 619614
rect 474542 619058 474574 619614
rect 473954 583614 474574 619058
rect 473954 583058 473986 583614
rect 474542 583058 474574 583614
rect 473954 547614 474574 583058
rect 473954 547058 473986 547614
rect 474542 547058 474574 547614
rect 473954 511614 474574 547058
rect 473954 511058 473986 511614
rect 474542 511058 474574 511614
rect 473954 475614 474574 511058
rect 473954 475058 473986 475614
rect 474542 475058 474574 475614
rect 473675 449716 473741 449717
rect 473675 449652 473676 449716
rect 473740 449652 473741 449716
rect 473675 449651 473741 449652
rect 472714 437818 472746 438374
rect 473302 437818 473334 438374
rect 472714 402374 473334 437818
rect 473678 431901 473738 449651
rect 473954 439614 474574 475058
rect 473954 439058 473986 439614
rect 474542 439058 474574 439614
rect 473675 431900 473741 431901
rect 473675 431836 473676 431900
rect 473740 431836 473741 431900
rect 473675 431835 473741 431836
rect 473678 410957 473738 431835
rect 473675 410956 473741 410957
rect 473675 410892 473676 410956
rect 473740 410892 473741 410956
rect 473675 410891 473741 410892
rect 472714 401818 472746 402374
rect 473302 401818 473334 402374
rect 472714 366374 473334 401818
rect 473678 392053 473738 410891
rect 473954 403614 474574 439058
rect 473954 403058 473986 403614
rect 474542 403058 474574 403614
rect 473675 392052 473741 392053
rect 473675 391988 473676 392052
rect 473740 391988 473741 392052
rect 473675 391987 473741 391988
rect 472714 365818 472746 366374
rect 473302 365818 473334 366374
rect 472714 359060 473334 365818
rect 473954 367614 474574 403058
rect 475194 709638 475814 711590
rect 475194 709082 475226 709638
rect 475782 709082 475814 709638
rect 475194 692854 475814 709082
rect 475194 692298 475226 692854
rect 475782 692298 475814 692854
rect 475194 656854 475814 692298
rect 475194 656298 475226 656854
rect 475782 656298 475814 656854
rect 475194 620854 475814 656298
rect 475194 620298 475226 620854
rect 475782 620298 475814 620854
rect 475194 584854 475814 620298
rect 475194 584298 475226 584854
rect 475782 584298 475814 584854
rect 475194 548854 475814 584298
rect 475194 548298 475226 548854
rect 475782 548298 475814 548854
rect 475194 512854 475814 548298
rect 475194 512298 475226 512854
rect 475782 512298 475814 512854
rect 475194 476854 475814 512298
rect 475194 476298 475226 476854
rect 475782 476298 475814 476854
rect 475194 440854 475814 476298
rect 475194 440298 475226 440854
rect 475782 440298 475814 440854
rect 475194 404854 475814 440298
rect 475194 404298 475226 404854
rect 475782 404298 475814 404854
rect 474963 392052 475029 392053
rect 474963 391988 474964 392052
rect 475028 391988 475029 392052
rect 474963 391987 475029 391988
rect 474966 389333 475026 391987
rect 474963 389332 475029 389333
rect 474963 389268 474964 389332
rect 475028 389268 475029 389332
rect 474963 389267 475029 389268
rect 473954 367058 473986 367614
rect 474542 367058 474574 367614
rect 473954 359060 474574 367058
rect 474966 357509 475026 389267
rect 475194 368854 475814 404298
rect 475194 368298 475226 368854
rect 475782 368298 475814 368854
rect 475194 359060 475814 368298
rect 476434 710598 477054 711590
rect 476434 710042 476466 710598
rect 477022 710042 477054 710598
rect 476434 694094 477054 710042
rect 476434 693538 476466 694094
rect 477022 693538 477054 694094
rect 476434 658094 477054 693538
rect 476434 657538 476466 658094
rect 477022 657538 477054 658094
rect 476434 622094 477054 657538
rect 476434 621538 476466 622094
rect 477022 621538 477054 622094
rect 476434 586094 477054 621538
rect 476434 585538 476466 586094
rect 477022 585538 477054 586094
rect 476434 550094 477054 585538
rect 476434 549538 476466 550094
rect 477022 549538 477054 550094
rect 476434 514094 477054 549538
rect 476434 513538 476466 514094
rect 477022 513538 477054 514094
rect 476434 478094 477054 513538
rect 476434 477538 476466 478094
rect 477022 477538 477054 478094
rect 476434 442094 477054 477538
rect 476434 441538 476466 442094
rect 477022 441538 477054 442094
rect 476434 406094 477054 441538
rect 476434 405538 476466 406094
rect 477022 405538 477054 406094
rect 476434 370094 477054 405538
rect 476434 369538 476466 370094
rect 477022 369538 477054 370094
rect 476434 359060 477054 369538
rect 477674 711558 478294 711590
rect 477674 711002 477706 711558
rect 478262 711002 478294 711558
rect 477674 695334 478294 711002
rect 477674 694778 477706 695334
rect 478262 694778 478294 695334
rect 477674 659334 478294 694778
rect 477674 658778 477706 659334
rect 478262 658778 478294 659334
rect 477674 623334 478294 658778
rect 477674 622778 477706 623334
rect 478262 622778 478294 623334
rect 477674 587334 478294 622778
rect 477674 586778 477706 587334
rect 478262 586778 478294 587334
rect 477674 551334 478294 586778
rect 477674 550778 477706 551334
rect 478262 550778 478294 551334
rect 477674 515334 478294 550778
rect 477674 514778 477706 515334
rect 478262 514778 478294 515334
rect 477674 479334 478294 514778
rect 477674 478778 477706 479334
rect 478262 478778 478294 479334
rect 477674 443334 478294 478778
rect 504994 704838 505614 711590
rect 504994 704282 505026 704838
rect 505582 704282 505614 704838
rect 504994 686654 505614 704282
rect 504994 686098 505026 686654
rect 505582 686098 505614 686654
rect 504994 650654 505614 686098
rect 504994 650098 505026 650654
rect 505582 650098 505614 650654
rect 504994 614654 505614 650098
rect 504994 614098 505026 614654
rect 505582 614098 505614 614654
rect 504994 578654 505614 614098
rect 504994 578098 505026 578654
rect 505582 578098 505614 578654
rect 504994 542654 505614 578098
rect 504994 542098 505026 542654
rect 505582 542098 505614 542654
rect 504994 506654 505614 542098
rect 504994 506098 505026 506654
rect 505582 506098 505614 506654
rect 504994 470654 505614 506098
rect 504994 470098 505026 470654
rect 505582 470098 505614 470654
rect 478459 450260 478525 450261
rect 478459 450196 478460 450260
rect 478524 450196 478525 450260
rect 478459 450195 478525 450196
rect 481219 450260 481285 450261
rect 481219 450196 481220 450260
rect 481284 450196 481285 450260
rect 481219 450195 481285 450196
rect 484163 450260 484229 450261
rect 484163 450196 484164 450260
rect 484228 450196 484229 450260
rect 484163 450195 484229 450196
rect 487843 450260 487909 450261
rect 487843 450196 487844 450260
rect 487908 450196 487909 450260
rect 487843 450195 487909 450196
rect 477674 442778 477706 443334
rect 478262 442778 478294 443334
rect 477674 407334 478294 442778
rect 478462 431629 478522 450195
rect 481222 432173 481282 450195
rect 483611 432308 483677 432309
rect 483611 432244 483612 432308
rect 483676 432244 483677 432308
rect 483611 432243 483677 432244
rect 481219 432172 481285 432173
rect 481219 432108 481220 432172
rect 481284 432108 481285 432172
rect 481219 432107 481285 432108
rect 481222 431970 481282 432107
rect 481038 431910 481282 431970
rect 483614 431970 483674 432243
rect 484166 431970 484226 450195
rect 487846 441630 487906 450195
rect 483614 431910 484226 431970
rect 487662 441570 487906 441630
rect 478459 431628 478525 431629
rect 478459 431564 478460 431628
rect 478524 431564 478525 431628
rect 478459 431563 478525 431564
rect 478462 410141 478522 431563
rect 480115 427956 480181 427957
rect 480115 427892 480116 427956
rect 480180 427892 480181 427956
rect 480115 427891 480181 427892
rect 478459 410140 478525 410141
rect 478459 410076 478460 410140
rect 478524 410076 478525 410140
rect 478459 410075 478525 410076
rect 477674 406778 477706 407334
rect 478262 406778 478294 407334
rect 477674 371334 478294 406778
rect 478462 402990 478522 410075
rect 480118 407557 480178 427891
rect 481038 422310 481098 431910
rect 483614 422310 483674 431910
rect 487662 431901 487722 441570
rect 504994 434654 505614 470098
rect 504994 434098 505026 434654
rect 505582 434098 505614 434654
rect 487659 431900 487725 431901
rect 487659 431836 487660 431900
rect 487724 431836 487725 431900
rect 487659 431835 487725 431836
rect 486555 427956 486621 427957
rect 486555 427892 486556 427956
rect 486620 427892 486621 427956
rect 486555 427891 486621 427892
rect 481038 422250 481466 422310
rect 483614 422250 484226 422310
rect 481406 410141 481466 422250
rect 484166 410413 484226 422250
rect 484163 410412 484229 410413
rect 484163 410348 484164 410412
rect 484228 410348 484229 410412
rect 484163 410347 484229 410348
rect 481403 410140 481469 410141
rect 481403 410076 481404 410140
rect 481468 410076 481469 410140
rect 481403 410075 481469 410076
rect 480115 407556 480181 407557
rect 480115 407492 480116 407556
rect 480180 407492 480181 407556
rect 480115 407491 480181 407492
rect 478462 402930 478706 402990
rect 478646 389333 478706 402930
rect 481406 393330 481466 410075
rect 482875 407148 482941 407149
rect 482875 407084 482876 407148
rect 482940 407084 482941 407148
rect 482875 407083 482941 407084
rect 481406 393270 481834 393330
rect 481774 389469 481834 393270
rect 481771 389468 481837 389469
rect 481771 389404 481772 389468
rect 481836 389404 481837 389468
rect 481771 389403 481837 389404
rect 478643 389332 478709 389333
rect 478643 389268 478644 389332
rect 478708 389268 478709 389332
rect 478643 389267 478709 389268
rect 477674 370778 477706 371334
rect 478262 370778 478294 371334
rect 477674 359060 478294 370778
rect 478646 358053 478706 389267
rect 481774 358053 481834 389403
rect 482878 370157 482938 407083
rect 484166 393330 484226 410347
rect 485635 407148 485701 407149
rect 485635 407084 485636 407148
rect 485700 407084 485701 407148
rect 485635 407083 485701 407084
rect 484166 393270 484962 393330
rect 484902 390298 484962 393270
rect 484899 390297 484965 390298
rect 484899 390233 484900 390297
rect 484964 390233 484965 390297
rect 484899 390232 484965 390233
rect 482875 370156 482941 370157
rect 482875 370092 482876 370156
rect 482940 370092 482941 370156
rect 482875 370091 482941 370092
rect 484902 358053 484962 390232
rect 478643 358052 478709 358053
rect 478643 357988 478644 358052
rect 478708 357988 478709 358052
rect 478643 357987 478709 357988
rect 481771 358052 481837 358053
rect 481771 357988 481772 358052
rect 481836 357988 481837 358052
rect 481771 357987 481837 357988
rect 484899 358052 484965 358053
rect 484899 357988 484900 358052
rect 484964 357988 484965 358052
rect 484899 357987 484965 357988
rect 474963 357508 475029 357509
rect 474963 357444 474964 357508
rect 475028 357444 475029 357508
rect 474963 357443 475029 357444
rect 474966 357370 475026 357443
rect 474966 357310 475394 357370
rect 475334 356690 475394 357310
rect 474966 356630 475394 356690
rect 471474 328578 471506 329134
rect 472062 328578 472094 329134
rect 471474 293134 472094 328578
rect 471474 292578 471506 293134
rect 472062 292578 472094 293134
rect 471474 257134 472094 292578
rect 472714 330374 473334 354615
rect 473675 343772 473741 343773
rect 473675 343708 473676 343772
rect 473740 343708 473741 343772
rect 473675 343707 473741 343708
rect 473678 340509 473738 343707
rect 473675 340508 473741 340509
rect 473675 340444 473676 340508
rect 473740 340444 473741 340508
rect 473675 340443 473741 340444
rect 472714 329818 472746 330374
rect 473302 329818 473334 330374
rect 472714 294374 473334 329818
rect 473678 321333 473738 340443
rect 473954 331614 474574 354615
rect 474966 343773 475026 356630
rect 474963 343772 475029 343773
rect 474963 343708 474964 343772
rect 475028 343708 475029 343772
rect 474963 343707 475029 343708
rect 473954 331058 473986 331614
rect 474542 331058 474574 331614
rect 473675 321332 473741 321333
rect 473675 321268 473676 321332
rect 473740 321268 473741 321332
rect 473675 321267 473741 321268
rect 473678 305965 473738 321267
rect 473675 305964 473741 305965
rect 473675 305900 473676 305964
rect 473740 305900 473741 305964
rect 473675 305899 473741 305900
rect 472714 293818 472746 294374
rect 473302 293818 473334 294374
rect 472714 268060 473334 293818
rect 473678 289781 473738 305899
rect 473954 295614 474574 331058
rect 473954 295058 473986 295614
rect 474542 295058 474574 295614
rect 473675 289780 473741 289781
rect 473675 289716 473676 289780
rect 473740 289716 473741 289780
rect 473675 289715 473741 289716
rect 473954 268060 474574 295058
rect 475194 332854 475814 354615
rect 475194 332298 475226 332854
rect 475782 332298 475814 332854
rect 475194 296854 475814 332298
rect 475194 296298 475226 296854
rect 475782 296298 475814 296854
rect 475194 268060 475814 296298
rect 476434 334094 477054 354615
rect 476434 333538 476466 334094
rect 477022 333538 477054 334094
rect 476434 298094 477054 333538
rect 476434 297538 476466 298094
rect 477022 297538 477054 298094
rect 476067 289780 476133 289781
rect 476067 289716 476068 289780
rect 476132 289716 476133 289780
rect 476067 289715 476133 289716
rect 476070 286653 476130 289715
rect 476067 286652 476133 286653
rect 476067 286588 476068 286652
rect 476132 286588 476133 286652
rect 476067 286587 476133 286588
rect 476070 267750 476130 286587
rect 476434 268060 477054 297538
rect 477674 335334 478294 354615
rect 478646 345030 478706 357987
rect 481774 354690 481834 357987
rect 484902 354690 484962 357987
rect 481590 354630 481834 354690
rect 484534 354630 484962 354690
rect 481590 345030 481650 354630
rect 484534 345030 484594 354630
rect 478462 344970 478706 345030
rect 481406 344970 481650 345030
rect 484166 344970 484594 345030
rect 478462 341053 478522 344970
rect 481406 341053 481466 344970
rect 484166 341053 484226 344970
rect 478459 341052 478525 341053
rect 478459 340988 478460 341052
rect 478524 340988 478525 341052
rect 478459 340987 478525 340988
rect 481403 341052 481469 341053
rect 481403 340988 481404 341052
rect 481468 340988 481469 341052
rect 481403 340987 481469 340988
rect 484163 341052 484229 341053
rect 484163 340988 484164 341052
rect 484228 340988 484229 341052
rect 484163 340987 484229 340988
rect 477674 334778 477706 335334
rect 478262 334778 478294 335334
rect 477674 299334 478294 334778
rect 478462 325710 478522 340987
rect 481406 325710 481466 340987
rect 478462 325650 478706 325710
rect 481406 325650 481650 325710
rect 478646 320925 478706 325650
rect 481590 320925 481650 325650
rect 484166 321333 484226 340987
rect 485638 334117 485698 407083
rect 486558 335477 486618 427891
rect 487662 422310 487722 431835
rect 487662 422250 487906 422310
rect 487846 410141 487906 422250
rect 487843 410140 487909 410141
rect 487843 410076 487844 410140
rect 487908 410076 487909 410140
rect 487843 410075 487909 410076
rect 488395 410140 488461 410141
rect 488395 410076 488396 410140
rect 488460 410076 488461 410140
rect 488395 410075 488461 410076
rect 488398 390149 488458 410075
rect 504994 398654 505614 434098
rect 504994 398098 505026 398654
rect 505582 398098 505614 398654
rect 488395 390148 488461 390149
rect 488395 390084 488396 390148
rect 488460 390084 488461 390148
rect 488395 390083 488461 390084
rect 486739 386476 486805 386477
rect 486739 386412 486740 386476
rect 486804 386412 486805 386476
rect 486739 386411 486805 386412
rect 486555 335476 486621 335477
rect 486555 335412 486556 335476
rect 486620 335412 486621 335476
rect 486555 335411 486621 335412
rect 485635 334116 485701 334117
rect 485635 334052 485636 334116
rect 485700 334052 485701 334116
rect 485635 334051 485701 334052
rect 486742 332757 486802 386411
rect 488398 358053 488458 390083
rect 504994 362654 505614 398098
rect 504994 362098 505026 362654
rect 505582 362098 505614 362654
rect 488395 358052 488461 358053
rect 488395 357988 488396 358052
rect 488460 357988 488461 358052
rect 488395 357987 488461 357988
rect 488398 354690 488458 357987
rect 487662 354630 488458 354690
rect 487662 345030 487722 354630
rect 487662 344970 488090 345030
rect 488030 341053 488090 344970
rect 488027 341052 488093 341053
rect 488027 340988 488028 341052
rect 488092 340988 488093 341052
rect 488027 340987 488093 340988
rect 486739 332756 486805 332757
rect 486739 332692 486740 332756
rect 486804 332692 486805 332756
rect 486739 332691 486805 332692
rect 484163 321332 484229 321333
rect 484163 321268 484164 321332
rect 484228 321268 484229 321332
rect 484163 321267 484229 321268
rect 478643 320924 478709 320925
rect 478643 320860 478644 320924
rect 478708 320860 478709 320924
rect 478643 320859 478709 320860
rect 481587 320924 481653 320925
rect 481587 320860 481588 320924
rect 481652 320860 481653 320924
rect 481587 320859 481653 320860
rect 478646 306390 478706 320859
rect 481590 306390 481650 320859
rect 478646 306330 478890 306390
rect 478830 305693 478890 306330
rect 481590 306330 482202 306390
rect 481590 306101 481650 306330
rect 481587 306100 481653 306101
rect 481587 306036 481588 306100
rect 481652 306036 481653 306100
rect 481587 306035 481653 306036
rect 478827 305692 478893 305693
rect 478827 305628 478828 305692
rect 478892 305628 478893 305692
rect 478827 305627 478893 305628
rect 477674 298778 477706 299334
rect 478262 298778 478294 299334
rect 477674 268060 478294 298778
rect 478830 287070 478890 305627
rect 482142 287070 482202 306330
rect 484166 305557 484226 321267
rect 488030 321061 488090 340987
rect 504994 326654 505614 362098
rect 504994 326098 505026 326654
rect 505582 326098 505614 326654
rect 488027 321060 488093 321061
rect 488027 320996 488028 321060
rect 488092 320996 488093 321060
rect 488027 320995 488093 320996
rect 488030 316050 488090 320995
rect 487662 315990 488090 316050
rect 487662 306390 487722 315990
rect 487662 306373 488458 306390
rect 487659 306372 488458 306373
rect 487659 306308 487660 306372
rect 487724 306330 488458 306372
rect 487724 306308 487725 306330
rect 487659 306307 487725 306308
rect 484163 305556 484229 305557
rect 484163 305492 484164 305556
rect 484228 305492 484229 305556
rect 484163 305491 484229 305492
rect 484166 289781 484226 305491
rect 484163 289780 484229 289781
rect 484163 289716 484164 289780
rect 484228 289716 484229 289780
rect 484163 289715 484229 289716
rect 485819 289780 485885 289781
rect 485819 289716 485820 289780
rect 485884 289716 485885 289780
rect 485819 289715 485885 289716
rect 478830 287010 479074 287070
rect 482142 287010 482386 287070
rect 478830 286925 478890 287010
rect 478827 286924 478893 286925
rect 478827 286860 478828 286924
rect 478892 286860 478893 286924
rect 478827 286859 478893 286860
rect 476070 267690 476498 267750
rect 476438 265029 476498 267690
rect 479014 265981 479074 287010
rect 482326 285837 482386 287010
rect 485822 285837 485882 289715
rect 488398 288690 488458 306330
rect 504994 290654 505614 326098
rect 504994 290098 505026 290654
rect 505582 290098 505614 290654
rect 488398 288630 488642 288690
rect 488582 286789 488642 288630
rect 488579 286788 488645 286789
rect 488579 286724 488580 286788
rect 488644 286724 488645 286788
rect 488579 286723 488645 286724
rect 482323 285836 482389 285837
rect 482323 285772 482324 285836
rect 482388 285772 482389 285836
rect 482323 285771 482389 285772
rect 482875 285836 482941 285837
rect 482875 285772 482876 285836
rect 482940 285772 482941 285836
rect 482875 285771 482941 285772
rect 485819 285836 485885 285837
rect 485819 285772 485820 285836
rect 485884 285772 485885 285836
rect 485819 285771 485885 285772
rect 479011 265980 479077 265981
rect 479011 265916 479012 265980
rect 479076 265916 479077 265980
rect 479011 265915 479077 265916
rect 482878 265029 482938 285771
rect 485822 265029 485882 285771
rect 488582 267750 488642 286723
rect 488582 267690 489194 267750
rect 489134 265573 489194 267690
rect 489131 265572 489197 265573
rect 489131 265508 489132 265572
rect 489196 265508 489197 265572
rect 489131 265507 489197 265508
rect 476435 265028 476501 265029
rect 476435 264964 476436 265028
rect 476500 264964 476501 265028
rect 476435 264963 476501 264964
rect 477355 265028 477421 265029
rect 477355 264964 477356 265028
rect 477420 264964 477421 265028
rect 477355 264963 477421 264964
rect 480115 265028 480181 265029
rect 480115 264964 480116 265028
rect 480180 264964 480181 265028
rect 480115 264963 480181 264964
rect 482875 265028 482941 265029
rect 482875 264964 482876 265028
rect 482940 264964 482941 265028
rect 482875 264963 482941 264964
rect 485819 265028 485885 265029
rect 485819 264964 485820 265028
rect 485884 264964 485885 265028
rect 485819 264963 485885 264964
rect 486371 265028 486437 265029
rect 486371 264964 486372 265028
rect 486436 264964 486437 265028
rect 486371 264963 486437 264964
rect 471474 256578 471506 257134
rect 472062 256578 472094 257134
rect 471474 221134 472094 256578
rect 471474 220578 471506 221134
rect 472062 220578 472094 221134
rect 471474 185134 472094 220578
rect 471474 184578 471506 185134
rect 472062 184578 472094 185134
rect 471474 149134 472094 184578
rect 471474 148578 471506 149134
rect 472062 148578 472094 149134
rect 471474 113134 472094 148578
rect 471474 112578 471506 113134
rect 472062 112578 472094 113134
rect 471474 77134 472094 112578
rect 471474 76578 471506 77134
rect 472062 76578 472094 77134
rect 471474 41134 472094 76578
rect 471474 40578 471506 41134
rect 472062 40578 472094 41134
rect 471474 5134 472094 40578
rect 471474 4578 471506 5134
rect 472062 4578 472094 5134
rect 471474 -2266 472094 4578
rect 471474 -2822 471506 -2266
rect 472062 -2822 472094 -2266
rect 471474 -7654 472094 -2822
rect 472714 258374 473334 263615
rect 472714 257818 472746 258374
rect 473302 257818 473334 258374
rect 472714 222374 473334 257818
rect 472714 221818 472746 222374
rect 473302 221818 473334 222374
rect 472714 186374 473334 221818
rect 472714 185818 472746 186374
rect 473302 185818 473334 186374
rect 472714 150374 473334 185818
rect 472714 149818 472746 150374
rect 473302 149818 473334 150374
rect 472714 114374 473334 149818
rect 472714 113818 472746 114374
rect 473302 113818 473334 114374
rect 472714 78374 473334 113818
rect 472714 77818 472746 78374
rect 473302 77818 473334 78374
rect 472714 42374 473334 77818
rect 472714 41818 472746 42374
rect 473302 41818 473334 42374
rect 472714 6374 473334 41818
rect 472714 5818 472746 6374
rect 473302 5818 473334 6374
rect 472714 -3226 473334 5818
rect 472714 -3782 472746 -3226
rect 473302 -3782 473334 -3226
rect 472714 -7654 473334 -3782
rect 473954 259614 474574 263615
rect 473954 259058 473986 259614
rect 474542 259058 474574 259614
rect 473954 223614 474574 259058
rect 473954 223058 473986 223614
rect 474542 223058 474574 223614
rect 473954 187614 474574 223058
rect 473954 187058 473986 187614
rect 474542 187058 474574 187614
rect 473954 151614 474574 187058
rect 473954 151058 473986 151614
rect 474542 151058 474574 151614
rect 473954 115614 474574 151058
rect 473954 115058 473986 115614
rect 474542 115058 474574 115614
rect 473954 79614 474574 115058
rect 473954 79058 473986 79614
rect 474542 79058 474574 79614
rect 473954 43614 474574 79058
rect 473954 43058 473986 43614
rect 474542 43058 474574 43614
rect 473954 7614 474574 43058
rect 473954 7058 473986 7614
rect 474542 7058 474574 7614
rect 473954 -4186 474574 7058
rect 473954 -4742 473986 -4186
rect 474542 -4742 474574 -4186
rect 473954 -7654 474574 -4742
rect 475194 260854 475814 263615
rect 475194 260298 475226 260854
rect 475782 260298 475814 260854
rect 475194 224854 475814 260298
rect 475194 224298 475226 224854
rect 475782 224298 475814 224854
rect 475194 188854 475814 224298
rect 475194 188298 475226 188854
rect 475782 188298 475814 188854
rect 475194 152854 475814 188298
rect 475194 152298 475226 152854
rect 475782 152298 475814 152854
rect 475194 116854 475814 152298
rect 475194 116298 475226 116854
rect 475782 116298 475814 116854
rect 475194 80854 475814 116298
rect 475194 80298 475226 80854
rect 475782 80298 475814 80854
rect 475194 44854 475814 80298
rect 475194 44298 475226 44854
rect 475782 44298 475814 44854
rect 475194 8854 475814 44298
rect 475194 8298 475226 8854
rect 475782 8298 475814 8854
rect 475194 -5146 475814 8298
rect 475194 -5702 475226 -5146
rect 475782 -5702 475814 -5146
rect 475194 -7654 475814 -5702
rect 476434 262094 477054 263615
rect 476434 261538 476466 262094
rect 477022 261538 477054 262094
rect 476434 226094 477054 261538
rect 476434 225538 476466 226094
rect 477022 225538 477054 226094
rect 476434 190094 477054 225538
rect 476434 189538 476466 190094
rect 477022 189538 477054 190094
rect 476434 154094 477054 189538
rect 476434 153538 476466 154094
rect 477022 153538 477054 154094
rect 476434 118094 477054 153538
rect 476434 117538 476466 118094
rect 477022 117538 477054 118094
rect 476434 82094 477054 117538
rect 476434 81538 476466 82094
rect 477022 81538 477054 82094
rect 476434 46094 477054 81538
rect 476434 45538 476466 46094
rect 477022 45538 477054 46094
rect 476434 10094 477054 45538
rect 476434 9538 476466 10094
rect 477022 9538 477054 10094
rect 476434 -6106 477054 9538
rect 477358 6629 477418 264963
rect 477674 263334 478294 263615
rect 477674 262778 477706 263334
rect 478262 262778 478294 263334
rect 477674 227334 478294 262778
rect 477674 226778 477706 227334
rect 478262 226778 478294 227334
rect 477674 191334 478294 226778
rect 477674 190778 477706 191334
rect 478262 190778 478294 191334
rect 477674 155334 478294 190778
rect 477674 154778 477706 155334
rect 478262 154778 478294 155334
rect 477674 119334 478294 154778
rect 477674 118778 477706 119334
rect 478262 118778 478294 119334
rect 477674 83334 478294 118778
rect 477674 82778 477706 83334
rect 478262 82778 478294 83334
rect 477674 47334 478294 82778
rect 477674 46778 477706 47334
rect 478262 46778 478294 47334
rect 477674 11334 478294 46778
rect 480118 46341 480178 264963
rect 482878 86189 482938 264963
rect 486374 126037 486434 264963
rect 489134 165885 489194 265507
rect 504994 254654 505614 290098
rect 504994 254098 505026 254654
rect 505582 254098 505614 254654
rect 504994 218654 505614 254098
rect 504994 218098 505026 218654
rect 505582 218098 505614 218654
rect 504994 182654 505614 218098
rect 504994 182098 505026 182654
rect 505582 182098 505614 182654
rect 489131 165884 489197 165885
rect 489131 165820 489132 165884
rect 489196 165820 489197 165884
rect 489131 165819 489197 165820
rect 504994 146654 505614 182098
rect 504994 146098 505026 146654
rect 505582 146098 505614 146654
rect 486371 126036 486437 126037
rect 486371 125972 486372 126036
rect 486436 125972 486437 126036
rect 486371 125971 486437 125972
rect 504994 110654 505614 146098
rect 504994 110098 505026 110654
rect 505582 110098 505614 110654
rect 482875 86188 482941 86189
rect 482875 86124 482876 86188
rect 482940 86124 482941 86188
rect 482875 86123 482941 86124
rect 504994 74654 505614 110098
rect 504994 74098 505026 74654
rect 505582 74098 505614 74654
rect 480115 46340 480181 46341
rect 480115 46276 480116 46340
rect 480180 46276 480181 46340
rect 480115 46275 480181 46276
rect 477674 10778 477706 11334
rect 478262 10778 478294 11334
rect 477355 6628 477421 6629
rect 477355 6564 477356 6628
rect 477420 6564 477421 6628
rect 477355 6563 477421 6564
rect 476434 -6662 476466 -6106
rect 477022 -6662 477054 -6106
rect 476434 -7654 477054 -6662
rect 477674 -7066 478294 10778
rect 477674 -7622 477706 -7066
rect 478262 -7622 478294 -7066
rect 477674 -7654 478294 -7622
rect 504994 38654 505614 74098
rect 504994 38098 505026 38654
rect 505582 38098 505614 38654
rect 504994 2654 505614 38098
rect 504994 2098 505026 2654
rect 505582 2098 505614 2654
rect 504994 -346 505614 2098
rect 504994 -902 505026 -346
rect 505582 -902 505614 -346
rect 504994 -7654 505614 -902
rect 506234 705798 506854 711590
rect 506234 705242 506266 705798
rect 506822 705242 506854 705798
rect 506234 687894 506854 705242
rect 506234 687338 506266 687894
rect 506822 687338 506854 687894
rect 506234 651894 506854 687338
rect 506234 651338 506266 651894
rect 506822 651338 506854 651894
rect 506234 615894 506854 651338
rect 506234 615338 506266 615894
rect 506822 615338 506854 615894
rect 506234 579894 506854 615338
rect 506234 579338 506266 579894
rect 506822 579338 506854 579894
rect 506234 543894 506854 579338
rect 506234 543338 506266 543894
rect 506822 543338 506854 543894
rect 506234 507894 506854 543338
rect 506234 507338 506266 507894
rect 506822 507338 506854 507894
rect 506234 471894 506854 507338
rect 506234 471338 506266 471894
rect 506822 471338 506854 471894
rect 506234 435894 506854 471338
rect 506234 435338 506266 435894
rect 506822 435338 506854 435894
rect 506234 399894 506854 435338
rect 506234 399338 506266 399894
rect 506822 399338 506854 399894
rect 506234 363894 506854 399338
rect 506234 363338 506266 363894
rect 506822 363338 506854 363894
rect 506234 327894 506854 363338
rect 506234 327338 506266 327894
rect 506822 327338 506854 327894
rect 506234 291894 506854 327338
rect 506234 291338 506266 291894
rect 506822 291338 506854 291894
rect 506234 255894 506854 291338
rect 506234 255338 506266 255894
rect 506822 255338 506854 255894
rect 506234 219894 506854 255338
rect 506234 219338 506266 219894
rect 506822 219338 506854 219894
rect 506234 183894 506854 219338
rect 506234 183338 506266 183894
rect 506822 183338 506854 183894
rect 506234 147894 506854 183338
rect 506234 147338 506266 147894
rect 506822 147338 506854 147894
rect 506234 111894 506854 147338
rect 506234 111338 506266 111894
rect 506822 111338 506854 111894
rect 506234 75894 506854 111338
rect 506234 75338 506266 75894
rect 506822 75338 506854 75894
rect 506234 39894 506854 75338
rect 506234 39338 506266 39894
rect 506822 39338 506854 39894
rect 506234 3894 506854 39338
rect 506234 3338 506266 3894
rect 506822 3338 506854 3894
rect 506234 -1306 506854 3338
rect 506234 -1862 506266 -1306
rect 506822 -1862 506854 -1306
rect 506234 -7654 506854 -1862
rect 507474 706758 508094 711590
rect 507474 706202 507506 706758
rect 508062 706202 508094 706758
rect 507474 689134 508094 706202
rect 507474 688578 507506 689134
rect 508062 688578 508094 689134
rect 507474 653134 508094 688578
rect 507474 652578 507506 653134
rect 508062 652578 508094 653134
rect 507474 617134 508094 652578
rect 507474 616578 507506 617134
rect 508062 616578 508094 617134
rect 507474 581134 508094 616578
rect 507474 580578 507506 581134
rect 508062 580578 508094 581134
rect 507474 545134 508094 580578
rect 507474 544578 507506 545134
rect 508062 544578 508094 545134
rect 507474 509134 508094 544578
rect 507474 508578 507506 509134
rect 508062 508578 508094 509134
rect 507474 473134 508094 508578
rect 507474 472578 507506 473134
rect 508062 472578 508094 473134
rect 507474 437134 508094 472578
rect 507474 436578 507506 437134
rect 508062 436578 508094 437134
rect 507474 401134 508094 436578
rect 507474 400578 507506 401134
rect 508062 400578 508094 401134
rect 507474 365134 508094 400578
rect 507474 364578 507506 365134
rect 508062 364578 508094 365134
rect 507474 329134 508094 364578
rect 507474 328578 507506 329134
rect 508062 328578 508094 329134
rect 507474 293134 508094 328578
rect 507474 292578 507506 293134
rect 508062 292578 508094 293134
rect 507474 257134 508094 292578
rect 507474 256578 507506 257134
rect 508062 256578 508094 257134
rect 507474 221134 508094 256578
rect 507474 220578 507506 221134
rect 508062 220578 508094 221134
rect 507474 185134 508094 220578
rect 507474 184578 507506 185134
rect 508062 184578 508094 185134
rect 507474 149134 508094 184578
rect 507474 148578 507506 149134
rect 508062 148578 508094 149134
rect 507474 113134 508094 148578
rect 507474 112578 507506 113134
rect 508062 112578 508094 113134
rect 507474 77134 508094 112578
rect 507474 76578 507506 77134
rect 508062 76578 508094 77134
rect 507474 41134 508094 76578
rect 507474 40578 507506 41134
rect 508062 40578 508094 41134
rect 507474 5134 508094 40578
rect 507474 4578 507506 5134
rect 508062 4578 508094 5134
rect 507474 -2266 508094 4578
rect 507474 -2822 507506 -2266
rect 508062 -2822 508094 -2266
rect 507474 -7654 508094 -2822
rect 508714 707718 509334 711590
rect 508714 707162 508746 707718
rect 509302 707162 509334 707718
rect 508714 690374 509334 707162
rect 508714 689818 508746 690374
rect 509302 689818 509334 690374
rect 508714 654374 509334 689818
rect 508714 653818 508746 654374
rect 509302 653818 509334 654374
rect 508714 618374 509334 653818
rect 508714 617818 508746 618374
rect 509302 617818 509334 618374
rect 508714 582374 509334 617818
rect 508714 581818 508746 582374
rect 509302 581818 509334 582374
rect 508714 546374 509334 581818
rect 508714 545818 508746 546374
rect 509302 545818 509334 546374
rect 508714 510374 509334 545818
rect 508714 509818 508746 510374
rect 509302 509818 509334 510374
rect 508714 474374 509334 509818
rect 508714 473818 508746 474374
rect 509302 473818 509334 474374
rect 508714 438374 509334 473818
rect 508714 437818 508746 438374
rect 509302 437818 509334 438374
rect 508714 402374 509334 437818
rect 508714 401818 508746 402374
rect 509302 401818 509334 402374
rect 508714 366374 509334 401818
rect 508714 365818 508746 366374
rect 509302 365818 509334 366374
rect 508714 330374 509334 365818
rect 508714 329818 508746 330374
rect 509302 329818 509334 330374
rect 508714 294374 509334 329818
rect 508714 293818 508746 294374
rect 509302 293818 509334 294374
rect 508714 258374 509334 293818
rect 508714 257818 508746 258374
rect 509302 257818 509334 258374
rect 508714 222374 509334 257818
rect 508714 221818 508746 222374
rect 509302 221818 509334 222374
rect 508714 186374 509334 221818
rect 508714 185818 508746 186374
rect 509302 185818 509334 186374
rect 508714 150374 509334 185818
rect 508714 149818 508746 150374
rect 509302 149818 509334 150374
rect 508714 114374 509334 149818
rect 508714 113818 508746 114374
rect 509302 113818 509334 114374
rect 508714 78374 509334 113818
rect 508714 77818 508746 78374
rect 509302 77818 509334 78374
rect 508714 42374 509334 77818
rect 508714 41818 508746 42374
rect 509302 41818 509334 42374
rect 508714 6374 509334 41818
rect 508714 5818 508746 6374
rect 509302 5818 509334 6374
rect 508714 -3226 509334 5818
rect 508714 -3782 508746 -3226
rect 509302 -3782 509334 -3226
rect 508714 -7654 509334 -3782
rect 509954 708678 510574 711590
rect 509954 708122 509986 708678
rect 510542 708122 510574 708678
rect 509954 691614 510574 708122
rect 509954 691058 509986 691614
rect 510542 691058 510574 691614
rect 509954 655614 510574 691058
rect 509954 655058 509986 655614
rect 510542 655058 510574 655614
rect 509954 619614 510574 655058
rect 509954 619058 509986 619614
rect 510542 619058 510574 619614
rect 509954 583614 510574 619058
rect 509954 583058 509986 583614
rect 510542 583058 510574 583614
rect 509954 547614 510574 583058
rect 509954 547058 509986 547614
rect 510542 547058 510574 547614
rect 509954 511614 510574 547058
rect 509954 511058 509986 511614
rect 510542 511058 510574 511614
rect 509954 475614 510574 511058
rect 509954 475058 509986 475614
rect 510542 475058 510574 475614
rect 509954 439614 510574 475058
rect 509954 439058 509986 439614
rect 510542 439058 510574 439614
rect 509954 403614 510574 439058
rect 509954 403058 509986 403614
rect 510542 403058 510574 403614
rect 509954 367614 510574 403058
rect 509954 367058 509986 367614
rect 510542 367058 510574 367614
rect 509954 331614 510574 367058
rect 509954 331058 509986 331614
rect 510542 331058 510574 331614
rect 509954 295614 510574 331058
rect 509954 295058 509986 295614
rect 510542 295058 510574 295614
rect 509954 259614 510574 295058
rect 509954 259058 509986 259614
rect 510542 259058 510574 259614
rect 509954 223614 510574 259058
rect 509954 223058 509986 223614
rect 510542 223058 510574 223614
rect 509954 187614 510574 223058
rect 509954 187058 509986 187614
rect 510542 187058 510574 187614
rect 509954 151614 510574 187058
rect 509954 151058 509986 151614
rect 510542 151058 510574 151614
rect 509954 115614 510574 151058
rect 509954 115058 509986 115614
rect 510542 115058 510574 115614
rect 509954 79614 510574 115058
rect 509954 79058 509986 79614
rect 510542 79058 510574 79614
rect 509954 43614 510574 79058
rect 509954 43058 509986 43614
rect 510542 43058 510574 43614
rect 509954 7614 510574 43058
rect 509954 7058 509986 7614
rect 510542 7058 510574 7614
rect 509954 -4186 510574 7058
rect 509954 -4742 509986 -4186
rect 510542 -4742 510574 -4186
rect 509954 -7654 510574 -4742
rect 511194 709638 511814 711590
rect 511194 709082 511226 709638
rect 511782 709082 511814 709638
rect 511194 692854 511814 709082
rect 511194 692298 511226 692854
rect 511782 692298 511814 692854
rect 511194 656854 511814 692298
rect 511194 656298 511226 656854
rect 511782 656298 511814 656854
rect 511194 620854 511814 656298
rect 511194 620298 511226 620854
rect 511782 620298 511814 620854
rect 511194 584854 511814 620298
rect 511194 584298 511226 584854
rect 511782 584298 511814 584854
rect 511194 548854 511814 584298
rect 511194 548298 511226 548854
rect 511782 548298 511814 548854
rect 511194 512854 511814 548298
rect 511194 512298 511226 512854
rect 511782 512298 511814 512854
rect 511194 476854 511814 512298
rect 511194 476298 511226 476854
rect 511782 476298 511814 476854
rect 511194 440854 511814 476298
rect 511194 440298 511226 440854
rect 511782 440298 511814 440854
rect 511194 404854 511814 440298
rect 511194 404298 511226 404854
rect 511782 404298 511814 404854
rect 511194 368854 511814 404298
rect 511194 368298 511226 368854
rect 511782 368298 511814 368854
rect 511194 332854 511814 368298
rect 511194 332298 511226 332854
rect 511782 332298 511814 332854
rect 511194 296854 511814 332298
rect 511194 296298 511226 296854
rect 511782 296298 511814 296854
rect 511194 260854 511814 296298
rect 511194 260298 511226 260854
rect 511782 260298 511814 260854
rect 511194 224854 511814 260298
rect 511194 224298 511226 224854
rect 511782 224298 511814 224854
rect 511194 188854 511814 224298
rect 511194 188298 511226 188854
rect 511782 188298 511814 188854
rect 511194 152854 511814 188298
rect 511194 152298 511226 152854
rect 511782 152298 511814 152854
rect 511194 116854 511814 152298
rect 511194 116298 511226 116854
rect 511782 116298 511814 116854
rect 511194 80854 511814 116298
rect 511194 80298 511226 80854
rect 511782 80298 511814 80854
rect 511194 44854 511814 80298
rect 511194 44298 511226 44854
rect 511782 44298 511814 44854
rect 511194 8854 511814 44298
rect 511194 8298 511226 8854
rect 511782 8298 511814 8854
rect 511194 -5146 511814 8298
rect 511194 -5702 511226 -5146
rect 511782 -5702 511814 -5146
rect 511194 -7654 511814 -5702
rect 512434 710598 513054 711590
rect 512434 710042 512466 710598
rect 513022 710042 513054 710598
rect 512434 694094 513054 710042
rect 512434 693538 512466 694094
rect 513022 693538 513054 694094
rect 512434 658094 513054 693538
rect 512434 657538 512466 658094
rect 513022 657538 513054 658094
rect 512434 622094 513054 657538
rect 512434 621538 512466 622094
rect 513022 621538 513054 622094
rect 512434 586094 513054 621538
rect 512434 585538 512466 586094
rect 513022 585538 513054 586094
rect 512434 550094 513054 585538
rect 512434 549538 512466 550094
rect 513022 549538 513054 550094
rect 512434 514094 513054 549538
rect 512434 513538 512466 514094
rect 513022 513538 513054 514094
rect 512434 478094 513054 513538
rect 512434 477538 512466 478094
rect 513022 477538 513054 478094
rect 512434 442094 513054 477538
rect 512434 441538 512466 442094
rect 513022 441538 513054 442094
rect 512434 406094 513054 441538
rect 512434 405538 512466 406094
rect 513022 405538 513054 406094
rect 512434 370094 513054 405538
rect 512434 369538 512466 370094
rect 513022 369538 513054 370094
rect 512434 334094 513054 369538
rect 512434 333538 512466 334094
rect 513022 333538 513054 334094
rect 512434 298094 513054 333538
rect 512434 297538 512466 298094
rect 513022 297538 513054 298094
rect 512434 262094 513054 297538
rect 512434 261538 512466 262094
rect 513022 261538 513054 262094
rect 512434 226094 513054 261538
rect 512434 225538 512466 226094
rect 513022 225538 513054 226094
rect 512434 190094 513054 225538
rect 512434 189538 512466 190094
rect 513022 189538 513054 190094
rect 512434 154094 513054 189538
rect 512434 153538 512466 154094
rect 513022 153538 513054 154094
rect 512434 118094 513054 153538
rect 512434 117538 512466 118094
rect 513022 117538 513054 118094
rect 512434 82094 513054 117538
rect 512434 81538 512466 82094
rect 513022 81538 513054 82094
rect 512434 46094 513054 81538
rect 512434 45538 512466 46094
rect 513022 45538 513054 46094
rect 512434 10094 513054 45538
rect 512434 9538 512466 10094
rect 513022 9538 513054 10094
rect 512434 -6106 513054 9538
rect 512434 -6662 512466 -6106
rect 513022 -6662 513054 -6106
rect 512434 -7654 513054 -6662
rect 513674 711558 514294 711590
rect 513674 711002 513706 711558
rect 514262 711002 514294 711558
rect 513674 695334 514294 711002
rect 513674 694778 513706 695334
rect 514262 694778 514294 695334
rect 513674 659334 514294 694778
rect 513674 658778 513706 659334
rect 514262 658778 514294 659334
rect 513674 623334 514294 658778
rect 513674 622778 513706 623334
rect 514262 622778 514294 623334
rect 513674 587334 514294 622778
rect 513674 586778 513706 587334
rect 514262 586778 514294 587334
rect 513674 551334 514294 586778
rect 513674 550778 513706 551334
rect 514262 550778 514294 551334
rect 513674 515334 514294 550778
rect 513674 514778 513706 515334
rect 514262 514778 514294 515334
rect 513674 479334 514294 514778
rect 513674 478778 513706 479334
rect 514262 478778 514294 479334
rect 513674 443334 514294 478778
rect 540994 704838 541614 711590
rect 540994 704282 541026 704838
rect 541582 704282 541614 704838
rect 540994 686654 541614 704282
rect 540994 686098 541026 686654
rect 541582 686098 541614 686654
rect 540994 650654 541614 686098
rect 540994 650098 541026 650654
rect 541582 650098 541614 650654
rect 540994 614654 541614 650098
rect 540994 614098 541026 614654
rect 541582 614098 541614 614654
rect 540994 578654 541614 614098
rect 540994 578098 541026 578654
rect 541582 578098 541614 578654
rect 540994 542654 541614 578098
rect 540994 542098 541026 542654
rect 541582 542098 541614 542654
rect 540994 506654 541614 542098
rect 540994 506098 541026 506654
rect 541582 506098 541614 506654
rect 540994 470654 541614 506098
rect 540994 470098 541026 470654
rect 541582 470098 541614 470654
rect 540994 445572 541614 470098
rect 542234 705798 542854 711590
rect 542234 705242 542266 705798
rect 542822 705242 542854 705798
rect 542234 687894 542854 705242
rect 542234 687338 542266 687894
rect 542822 687338 542854 687894
rect 542234 651894 542854 687338
rect 542234 651338 542266 651894
rect 542822 651338 542854 651894
rect 542234 615894 542854 651338
rect 542234 615338 542266 615894
rect 542822 615338 542854 615894
rect 542234 579894 542854 615338
rect 542234 579338 542266 579894
rect 542822 579338 542854 579894
rect 542234 543894 542854 579338
rect 542234 543338 542266 543894
rect 542822 543338 542854 543894
rect 542234 507894 542854 543338
rect 542234 507338 542266 507894
rect 542822 507338 542854 507894
rect 542234 471894 542854 507338
rect 542234 471338 542266 471894
rect 542822 471338 542854 471894
rect 542234 445572 542854 471338
rect 543474 706758 544094 711590
rect 543474 706202 543506 706758
rect 544062 706202 544094 706758
rect 543474 689134 544094 706202
rect 543474 688578 543506 689134
rect 544062 688578 544094 689134
rect 543474 653134 544094 688578
rect 543474 652578 543506 653134
rect 544062 652578 544094 653134
rect 543474 617134 544094 652578
rect 543474 616578 543506 617134
rect 544062 616578 544094 617134
rect 543474 581134 544094 616578
rect 543474 580578 543506 581134
rect 544062 580578 544094 581134
rect 543474 545134 544094 580578
rect 543474 544578 543506 545134
rect 544062 544578 544094 545134
rect 543474 509134 544094 544578
rect 543474 508578 543506 509134
rect 544062 508578 544094 509134
rect 543474 473134 544094 508578
rect 543474 472578 543506 473134
rect 544062 472578 544094 473134
rect 543474 445572 544094 472578
rect 544714 707718 545334 711590
rect 544714 707162 544746 707718
rect 545302 707162 545334 707718
rect 544714 690374 545334 707162
rect 544714 689818 544746 690374
rect 545302 689818 545334 690374
rect 544714 654374 545334 689818
rect 544714 653818 544746 654374
rect 545302 653818 545334 654374
rect 544714 618374 545334 653818
rect 544714 617818 544746 618374
rect 545302 617818 545334 618374
rect 544714 582374 545334 617818
rect 544714 581818 544746 582374
rect 545302 581818 545334 582374
rect 544714 546374 545334 581818
rect 544714 545818 544746 546374
rect 545302 545818 545334 546374
rect 544714 510374 545334 545818
rect 544714 509818 544746 510374
rect 545302 509818 545334 510374
rect 544714 474374 545334 509818
rect 544714 473818 544746 474374
rect 545302 473818 545334 474374
rect 544714 445572 545334 473818
rect 545954 708678 546574 711590
rect 545954 708122 545986 708678
rect 546542 708122 546574 708678
rect 545954 691614 546574 708122
rect 545954 691058 545986 691614
rect 546542 691058 546574 691614
rect 545954 655614 546574 691058
rect 545954 655058 545986 655614
rect 546542 655058 546574 655614
rect 545954 619614 546574 655058
rect 545954 619058 545986 619614
rect 546542 619058 546574 619614
rect 545954 583614 546574 619058
rect 545954 583058 545986 583614
rect 546542 583058 546574 583614
rect 545954 547614 546574 583058
rect 545954 547058 545986 547614
rect 546542 547058 546574 547614
rect 545954 511614 546574 547058
rect 545954 511058 545986 511614
rect 546542 511058 546574 511614
rect 545954 475614 546574 511058
rect 545954 475058 545986 475614
rect 546542 475058 546574 475614
rect 545954 445572 546574 475058
rect 547194 709638 547814 711590
rect 547194 709082 547226 709638
rect 547782 709082 547814 709638
rect 547194 692854 547814 709082
rect 547194 692298 547226 692854
rect 547782 692298 547814 692854
rect 547194 656854 547814 692298
rect 547194 656298 547226 656854
rect 547782 656298 547814 656854
rect 547194 620854 547814 656298
rect 547194 620298 547226 620854
rect 547782 620298 547814 620854
rect 547194 584854 547814 620298
rect 547194 584298 547226 584854
rect 547782 584298 547814 584854
rect 547194 548854 547814 584298
rect 547194 548298 547226 548854
rect 547782 548298 547814 548854
rect 547194 512854 547814 548298
rect 547194 512298 547226 512854
rect 547782 512298 547814 512854
rect 547194 476854 547814 512298
rect 547194 476298 547226 476854
rect 547782 476298 547814 476854
rect 541571 445092 541637 445093
rect 541571 445028 541572 445092
rect 541636 445028 541637 445092
rect 541571 445027 541637 445028
rect 544331 445092 544397 445093
rect 544331 445028 544332 445092
rect 544396 445028 544397 445092
rect 544331 445027 544397 445028
rect 513674 442778 513706 443334
rect 514262 442778 514294 443334
rect 513674 407334 514294 442778
rect 540876 435894 541196 435926
rect 540876 435658 540918 435894
rect 541154 435658 541196 435894
rect 540876 435574 541196 435658
rect 540876 435338 540918 435574
rect 541154 435338 541196 435574
rect 540876 435306 541196 435338
rect 539910 434654 540230 434686
rect 539910 434418 539952 434654
rect 540188 434418 540230 434654
rect 539910 434334 540230 434418
rect 539910 434098 539952 434334
rect 540188 434098 540230 434334
rect 539910 434066 540230 434098
rect 541574 409325 541634 445027
rect 542808 435894 543128 435926
rect 542808 435658 542850 435894
rect 543086 435658 543128 435894
rect 542808 435574 543128 435658
rect 542808 435338 542850 435574
rect 543086 435338 543128 435574
rect 542808 435306 543128 435338
rect 541842 434654 542162 434686
rect 541842 434418 541884 434654
rect 542120 434418 542162 434654
rect 541842 434334 542162 434418
rect 541842 434098 541884 434334
rect 542120 434098 542162 434334
rect 541842 434066 542162 434098
rect 543774 434654 544094 434686
rect 543774 434418 543816 434654
rect 544052 434418 544094 434654
rect 543774 434334 544094 434418
rect 543774 434098 543816 434334
rect 544052 434098 544094 434334
rect 543774 434066 544094 434098
rect 544334 409325 544394 445027
rect 547194 440854 547814 476298
rect 547194 440298 547226 440854
rect 547782 440298 547814 440854
rect 544740 435894 545060 435926
rect 544740 435658 544782 435894
rect 545018 435658 545060 435894
rect 544740 435574 545060 435658
rect 544740 435338 544782 435574
rect 545018 435338 545060 435574
rect 544740 435306 545060 435338
rect 546672 435894 546992 435926
rect 546672 435658 546714 435894
rect 546950 435658 546992 435894
rect 546672 435574 546992 435658
rect 546672 435338 546714 435574
rect 546950 435338 546992 435574
rect 546672 435306 546992 435338
rect 545706 434654 546026 434686
rect 545706 434418 545748 434654
rect 545984 434418 546026 434654
rect 545706 434334 546026 434418
rect 545706 434098 545748 434334
rect 545984 434098 546026 434334
rect 545706 434066 546026 434098
rect 541571 409324 541637 409325
rect 541571 409260 541572 409324
rect 541636 409260 541637 409324
rect 541571 409259 541637 409260
rect 544331 409324 544397 409325
rect 544331 409260 544332 409324
rect 544396 409260 544397 409324
rect 544331 409259 544397 409260
rect 513674 406778 513706 407334
rect 514262 406778 514294 407334
rect 513674 371334 514294 406778
rect 540876 399894 541196 399926
rect 540876 399658 540918 399894
rect 541154 399658 541196 399894
rect 540876 399574 541196 399658
rect 540876 399338 540918 399574
rect 541154 399338 541196 399574
rect 540876 399306 541196 399338
rect 539910 398654 540230 398686
rect 539910 398418 539952 398654
rect 540188 398418 540230 398654
rect 539910 398334 540230 398418
rect 539910 398098 539952 398334
rect 540188 398098 540230 398334
rect 539910 398066 540230 398098
rect 541574 373149 541634 409259
rect 542808 399894 543128 399926
rect 542808 399658 542850 399894
rect 543086 399658 543128 399894
rect 542808 399574 543128 399658
rect 542808 399338 542850 399574
rect 543086 399338 543128 399574
rect 542808 399306 543128 399338
rect 541842 398654 542162 398686
rect 541842 398418 541884 398654
rect 542120 398418 542162 398654
rect 541842 398334 542162 398418
rect 541842 398098 541884 398334
rect 542120 398098 542162 398334
rect 541842 398066 542162 398098
rect 543774 398654 544094 398686
rect 543774 398418 543816 398654
rect 544052 398418 544094 398654
rect 543774 398334 544094 398418
rect 543774 398098 543816 398334
rect 544052 398098 544094 398334
rect 543774 398066 544094 398098
rect 544334 383670 544394 409259
rect 547194 404854 547814 440298
rect 547194 404298 547226 404854
rect 547782 404298 547814 404854
rect 544740 399894 545060 399926
rect 544740 399658 544782 399894
rect 545018 399658 545060 399894
rect 544740 399574 545060 399658
rect 544740 399338 544782 399574
rect 545018 399338 545060 399574
rect 544740 399306 545060 399338
rect 546672 399894 546992 399926
rect 546672 399658 546714 399894
rect 546950 399658 546992 399894
rect 546672 399574 546992 399658
rect 546672 399338 546714 399574
rect 546950 399338 546992 399574
rect 546672 399306 546992 399338
rect 545706 398654 546026 398686
rect 545706 398418 545748 398654
rect 545984 398418 546026 398654
rect 545706 398334 546026 398418
rect 545706 398098 545748 398334
rect 545984 398098 546026 398334
rect 545706 398066 546026 398098
rect 544334 383610 544578 383670
rect 544518 373421 544578 383610
rect 544515 373420 544581 373421
rect 544515 373356 544516 373420
rect 544580 373356 544581 373420
rect 544515 373355 544581 373356
rect 541571 373148 541637 373149
rect 541571 373084 541572 373148
rect 541636 373084 541637 373148
rect 541571 373083 541637 373084
rect 513674 370778 513706 371334
rect 514262 370778 514294 371334
rect 513674 335334 514294 370778
rect 540876 363894 541196 363926
rect 540876 363658 540918 363894
rect 541154 363658 541196 363894
rect 540876 363574 541196 363658
rect 540876 363338 540918 363574
rect 541154 363338 541196 363574
rect 540876 363306 541196 363338
rect 539910 362654 540230 362686
rect 539910 362418 539952 362654
rect 540188 362418 540230 362654
rect 539910 362334 540230 362418
rect 539910 362098 539952 362334
rect 540188 362098 540230 362334
rect 539910 362066 540230 362098
rect 541574 339557 541634 373083
rect 542808 363894 543128 363926
rect 542808 363658 542850 363894
rect 543086 363658 543128 363894
rect 542808 363574 543128 363658
rect 542808 363338 542850 363574
rect 543086 363338 543128 363574
rect 542808 363306 543128 363338
rect 541842 362654 542162 362686
rect 541842 362418 541884 362654
rect 542120 362418 542162 362654
rect 541842 362334 542162 362418
rect 541842 362098 541884 362334
rect 542120 362098 542162 362334
rect 541842 362066 542162 362098
rect 543774 362654 544094 362686
rect 543774 362418 543816 362654
rect 544052 362418 544094 362654
rect 543774 362334 544094 362418
rect 543774 362098 543816 362334
rect 544052 362098 544094 362334
rect 543774 362066 544094 362098
rect 544518 354690 544578 373355
rect 547194 368854 547814 404298
rect 547194 368298 547226 368854
rect 547782 368298 547814 368854
rect 544740 363894 545060 363926
rect 544740 363658 544782 363894
rect 545018 363658 545060 363894
rect 544740 363574 545060 363658
rect 544740 363338 544782 363574
rect 545018 363338 545060 363574
rect 544740 363306 545060 363338
rect 546672 363894 546992 363926
rect 546672 363658 546714 363894
rect 546950 363658 546992 363894
rect 546672 363574 546992 363658
rect 546672 363338 546714 363574
rect 546950 363338 546992 363574
rect 546672 363306 546992 363338
rect 545706 362654 546026 362686
rect 545706 362418 545748 362654
rect 545984 362418 546026 362654
rect 545706 362334 546026 362418
rect 545706 362098 545748 362334
rect 545984 362098 546026 362334
rect 545706 362066 546026 362098
rect 544334 354630 544578 354690
rect 544334 351933 544394 354630
rect 544331 351932 544397 351933
rect 544331 351868 544332 351932
rect 544396 351868 544397 351932
rect 544331 351867 544397 351868
rect 544334 339557 544394 351867
rect 541571 339556 541637 339557
rect 541571 339492 541572 339556
rect 541636 339492 541637 339556
rect 541571 339491 541637 339492
rect 544331 339556 544397 339557
rect 544331 339492 544332 339556
rect 544396 339492 544397 339556
rect 544331 339491 544397 339492
rect 513674 334778 513706 335334
rect 514262 334778 514294 335334
rect 513674 299334 514294 334778
rect 540876 327894 541196 327926
rect 540876 327658 540918 327894
rect 541154 327658 541196 327894
rect 540876 327574 541196 327658
rect 540876 327338 540918 327574
rect 541154 327338 541196 327574
rect 540876 327306 541196 327338
rect 539910 326654 540230 326686
rect 539910 326418 539952 326654
rect 540188 326418 540230 326654
rect 539910 326334 540230 326418
rect 539910 326098 539952 326334
rect 540188 326098 540230 326334
rect 539910 326066 540230 326098
rect 541574 303653 541634 339491
rect 542808 327894 543128 327926
rect 542808 327658 542850 327894
rect 543086 327658 543128 327894
rect 542808 327574 543128 327658
rect 542808 327338 542850 327574
rect 543086 327338 543128 327574
rect 542808 327306 543128 327338
rect 541842 326654 542162 326686
rect 541842 326418 541884 326654
rect 542120 326418 542162 326654
rect 541842 326334 542162 326418
rect 541842 326098 541884 326334
rect 542120 326098 542162 326334
rect 541842 326066 542162 326098
rect 543774 326654 544094 326686
rect 543774 326418 543816 326654
rect 544052 326418 544094 326654
rect 543774 326334 544094 326418
rect 543774 326098 543816 326334
rect 544052 326098 544094 326334
rect 543774 326066 544094 326098
rect 544334 303789 544394 339491
rect 547194 332854 547814 368298
rect 547194 332298 547226 332854
rect 547782 332298 547814 332854
rect 544740 327894 545060 327926
rect 544740 327658 544782 327894
rect 545018 327658 545060 327894
rect 544740 327574 545060 327658
rect 544740 327338 544782 327574
rect 545018 327338 545060 327574
rect 544740 327306 545060 327338
rect 546672 327894 546992 327926
rect 546672 327658 546714 327894
rect 546950 327658 546992 327894
rect 546672 327574 546992 327658
rect 546672 327338 546714 327574
rect 546950 327338 546992 327574
rect 546672 327306 546992 327338
rect 545706 326654 546026 326686
rect 545706 326418 545748 326654
rect 545984 326418 546026 326654
rect 545706 326334 546026 326418
rect 545706 326098 545748 326334
rect 545984 326098 546026 326334
rect 545706 326066 546026 326098
rect 544331 303788 544397 303789
rect 544331 303724 544332 303788
rect 544396 303724 544397 303788
rect 544331 303723 544397 303724
rect 541571 303652 541637 303653
rect 541571 303588 541572 303652
rect 541636 303588 541637 303652
rect 541571 303587 541637 303588
rect 513674 298778 513706 299334
rect 514262 298778 514294 299334
rect 513674 263334 514294 298778
rect 547194 296854 547814 332298
rect 547194 296298 547226 296854
rect 547782 296298 547814 296854
rect 540876 291894 541196 291926
rect 540876 291658 540918 291894
rect 541154 291658 541196 291894
rect 540876 291574 541196 291658
rect 540876 291338 540918 291574
rect 541154 291338 541196 291574
rect 540876 291306 541196 291338
rect 542808 291894 543128 291926
rect 542808 291658 542850 291894
rect 543086 291658 543128 291894
rect 542808 291574 543128 291658
rect 542808 291338 542850 291574
rect 543086 291338 543128 291574
rect 542808 291306 543128 291338
rect 544740 291894 545060 291926
rect 544740 291658 544782 291894
rect 545018 291658 545060 291894
rect 544740 291574 545060 291658
rect 544740 291338 544782 291574
rect 545018 291338 545060 291574
rect 544740 291306 545060 291338
rect 546672 291894 546992 291926
rect 546672 291658 546714 291894
rect 546950 291658 546992 291894
rect 546672 291574 546992 291658
rect 546672 291338 546714 291574
rect 546950 291338 546992 291574
rect 546672 291306 546992 291338
rect 539910 290654 540230 290686
rect 539910 290418 539952 290654
rect 540188 290418 540230 290654
rect 539910 290334 540230 290418
rect 539910 290098 539952 290334
rect 540188 290098 540230 290334
rect 539910 290066 540230 290098
rect 541842 290654 542162 290686
rect 541842 290418 541884 290654
rect 542120 290418 542162 290654
rect 541842 290334 542162 290418
rect 541842 290098 541884 290334
rect 542120 290098 542162 290334
rect 541842 290066 542162 290098
rect 543774 290654 544094 290686
rect 543774 290418 543816 290654
rect 544052 290418 544094 290654
rect 543774 290334 544094 290418
rect 543774 290098 543816 290334
rect 544052 290098 544094 290334
rect 543774 290066 544094 290098
rect 545706 290654 546026 290686
rect 545706 290418 545748 290654
rect 545984 290418 546026 290654
rect 545706 290334 546026 290418
rect 545706 290098 545748 290334
rect 545984 290098 546026 290334
rect 545706 290066 546026 290098
rect 513674 262778 513706 263334
rect 514262 262778 514294 263334
rect 513674 227334 514294 262778
rect 513674 226778 513706 227334
rect 514262 226778 514294 227334
rect 513674 191334 514294 226778
rect 513674 190778 513706 191334
rect 514262 190778 514294 191334
rect 513674 155334 514294 190778
rect 513674 154778 513706 155334
rect 514262 154778 514294 155334
rect 513674 119334 514294 154778
rect 513674 118778 513706 119334
rect 514262 118778 514294 119334
rect 513674 83334 514294 118778
rect 513674 82778 513706 83334
rect 514262 82778 514294 83334
rect 513674 47334 514294 82778
rect 513674 46778 513706 47334
rect 514262 46778 514294 47334
rect 513674 11334 514294 46778
rect 513674 10778 513706 11334
rect 514262 10778 514294 11334
rect 513674 -7066 514294 10778
rect 513674 -7622 513706 -7066
rect 514262 -7622 514294 -7066
rect 513674 -7654 514294 -7622
rect 540994 254654 541614 279788
rect 540994 254098 541026 254654
rect 541582 254098 541614 254654
rect 540994 218654 541614 254098
rect 540994 218098 541026 218654
rect 541582 218098 541614 218654
rect 540994 182654 541614 218098
rect 540994 182098 541026 182654
rect 541582 182098 541614 182654
rect 540994 146654 541614 182098
rect 540994 146098 541026 146654
rect 541582 146098 541614 146654
rect 540994 110654 541614 146098
rect 540994 110098 541026 110654
rect 541582 110098 541614 110654
rect 540994 74654 541614 110098
rect 540994 74098 541026 74654
rect 541582 74098 541614 74654
rect 540994 38654 541614 74098
rect 540994 38098 541026 38654
rect 541582 38098 541614 38654
rect 540994 2654 541614 38098
rect 540994 2098 541026 2654
rect 541582 2098 541614 2654
rect 540994 -346 541614 2098
rect 540994 -902 541026 -346
rect 541582 -902 541614 -346
rect 540994 -7654 541614 -902
rect 542234 255894 542854 279788
rect 542234 255338 542266 255894
rect 542822 255338 542854 255894
rect 542234 219894 542854 255338
rect 542234 219338 542266 219894
rect 542822 219338 542854 219894
rect 542234 183894 542854 219338
rect 542234 183338 542266 183894
rect 542822 183338 542854 183894
rect 542234 147894 542854 183338
rect 542234 147338 542266 147894
rect 542822 147338 542854 147894
rect 542234 111894 542854 147338
rect 542234 111338 542266 111894
rect 542822 111338 542854 111894
rect 542234 75894 542854 111338
rect 542234 75338 542266 75894
rect 542822 75338 542854 75894
rect 542234 39894 542854 75338
rect 542234 39338 542266 39894
rect 542822 39338 542854 39894
rect 542234 3894 542854 39338
rect 542234 3338 542266 3894
rect 542822 3338 542854 3894
rect 542234 -1306 542854 3338
rect 542234 -1862 542266 -1306
rect 542822 -1862 542854 -1306
rect 542234 -7654 542854 -1862
rect 543474 257134 544094 279788
rect 543474 256578 543506 257134
rect 544062 256578 544094 257134
rect 543474 221134 544094 256578
rect 543474 220578 543506 221134
rect 544062 220578 544094 221134
rect 543474 185134 544094 220578
rect 543474 184578 543506 185134
rect 544062 184578 544094 185134
rect 543474 149134 544094 184578
rect 543474 148578 543506 149134
rect 544062 148578 544094 149134
rect 543474 113134 544094 148578
rect 543474 112578 543506 113134
rect 544062 112578 544094 113134
rect 543474 77134 544094 112578
rect 543474 76578 543506 77134
rect 544062 76578 544094 77134
rect 543474 41134 544094 76578
rect 543474 40578 543506 41134
rect 544062 40578 544094 41134
rect 543474 5134 544094 40578
rect 543474 4578 543506 5134
rect 544062 4578 544094 5134
rect 543474 -2266 544094 4578
rect 543474 -2822 543506 -2266
rect 544062 -2822 544094 -2266
rect 543474 -7654 544094 -2822
rect 544714 258374 545334 279788
rect 544714 257818 544746 258374
rect 545302 257818 545334 258374
rect 544714 222374 545334 257818
rect 544714 221818 544746 222374
rect 545302 221818 545334 222374
rect 544714 186374 545334 221818
rect 544714 185818 544746 186374
rect 545302 185818 545334 186374
rect 544714 150374 545334 185818
rect 544714 149818 544746 150374
rect 545302 149818 545334 150374
rect 544714 114374 545334 149818
rect 544714 113818 544746 114374
rect 545302 113818 545334 114374
rect 544714 78374 545334 113818
rect 544714 77818 544746 78374
rect 545302 77818 545334 78374
rect 544714 42374 545334 77818
rect 544714 41818 544746 42374
rect 545302 41818 545334 42374
rect 544714 6374 545334 41818
rect 544714 5818 544746 6374
rect 545302 5818 545334 6374
rect 544714 -3226 545334 5818
rect 544714 -3782 544746 -3226
rect 545302 -3782 545334 -3226
rect 544714 -7654 545334 -3782
rect 545954 259614 546574 279788
rect 545954 259058 545986 259614
rect 546542 259058 546574 259614
rect 545954 223614 546574 259058
rect 545954 223058 545986 223614
rect 546542 223058 546574 223614
rect 545954 187614 546574 223058
rect 545954 187058 545986 187614
rect 546542 187058 546574 187614
rect 545954 151614 546574 187058
rect 545954 151058 545986 151614
rect 546542 151058 546574 151614
rect 545954 115614 546574 151058
rect 545954 115058 545986 115614
rect 546542 115058 546574 115614
rect 545954 79614 546574 115058
rect 545954 79058 545986 79614
rect 546542 79058 546574 79614
rect 545954 43614 546574 79058
rect 545954 43058 545986 43614
rect 546542 43058 546574 43614
rect 545954 7614 546574 43058
rect 545954 7058 545986 7614
rect 546542 7058 546574 7614
rect 545954 -4186 546574 7058
rect 545954 -4742 545986 -4186
rect 546542 -4742 546574 -4186
rect 545954 -7654 546574 -4742
rect 547194 260854 547814 296298
rect 547194 260298 547226 260854
rect 547782 260298 547814 260854
rect 547194 224854 547814 260298
rect 547194 224298 547226 224854
rect 547782 224298 547814 224854
rect 547194 188854 547814 224298
rect 547194 188298 547226 188854
rect 547782 188298 547814 188854
rect 547194 152854 547814 188298
rect 547194 152298 547226 152854
rect 547782 152298 547814 152854
rect 547194 116854 547814 152298
rect 547194 116298 547226 116854
rect 547782 116298 547814 116854
rect 547194 80854 547814 116298
rect 547194 80298 547226 80854
rect 547782 80298 547814 80854
rect 547194 44854 547814 80298
rect 547194 44298 547226 44854
rect 547782 44298 547814 44854
rect 547194 8854 547814 44298
rect 547194 8298 547226 8854
rect 547782 8298 547814 8854
rect 547194 -5146 547814 8298
rect 547194 -5702 547226 -5146
rect 547782 -5702 547814 -5146
rect 547194 -7654 547814 -5702
rect 548434 710598 549054 711590
rect 548434 710042 548466 710598
rect 549022 710042 549054 710598
rect 548434 694094 549054 710042
rect 548434 693538 548466 694094
rect 549022 693538 549054 694094
rect 548434 658094 549054 693538
rect 548434 657538 548466 658094
rect 549022 657538 549054 658094
rect 548434 622094 549054 657538
rect 548434 621538 548466 622094
rect 549022 621538 549054 622094
rect 548434 586094 549054 621538
rect 548434 585538 548466 586094
rect 549022 585538 549054 586094
rect 548434 550094 549054 585538
rect 548434 549538 548466 550094
rect 549022 549538 549054 550094
rect 548434 514094 549054 549538
rect 548434 513538 548466 514094
rect 549022 513538 549054 514094
rect 548434 478094 549054 513538
rect 548434 477538 548466 478094
rect 549022 477538 549054 478094
rect 548434 442094 549054 477538
rect 548434 441538 548466 442094
rect 549022 441538 549054 442094
rect 548434 406094 549054 441538
rect 549674 711558 550294 711590
rect 549674 711002 549706 711558
rect 550262 711002 550294 711558
rect 549674 695334 550294 711002
rect 549674 694778 549706 695334
rect 550262 694778 550294 695334
rect 549674 659334 550294 694778
rect 549674 658778 549706 659334
rect 550262 658778 550294 659334
rect 549674 623334 550294 658778
rect 549674 622778 549706 623334
rect 550262 622778 550294 623334
rect 549674 587334 550294 622778
rect 549674 586778 549706 587334
rect 550262 586778 550294 587334
rect 549674 551334 550294 586778
rect 549674 550778 549706 551334
rect 550262 550778 550294 551334
rect 549674 515334 550294 550778
rect 549674 514778 549706 515334
rect 550262 514778 550294 515334
rect 549674 479334 550294 514778
rect 549674 478778 549706 479334
rect 550262 478778 550294 479334
rect 549674 443334 550294 478778
rect 549674 442778 549706 443334
rect 550262 442778 550294 443334
rect 549299 434756 549365 434757
rect 549299 434692 549300 434756
rect 549364 434692 549365 434756
rect 549299 434691 549365 434692
rect 548434 405538 548466 406094
rect 549022 405538 549054 406094
rect 548434 370094 549054 405538
rect 549302 398309 549362 434691
rect 549674 407334 550294 442778
rect 549674 406778 549706 407334
rect 550262 406778 550294 407334
rect 549299 398308 549365 398309
rect 549299 398244 549300 398308
rect 549364 398244 549365 398308
rect 549299 398243 549365 398244
rect 548434 369538 548466 370094
rect 549022 369538 549054 370094
rect 548434 334094 549054 369538
rect 549302 362813 549362 398243
rect 549674 371334 550294 406778
rect 549674 370778 549706 371334
rect 550262 370778 550294 371334
rect 549299 362812 549365 362813
rect 549299 362748 549300 362812
rect 549364 362748 549365 362812
rect 549299 362747 549365 362748
rect 548434 333538 548466 334094
rect 549022 333538 549054 334094
rect 548434 298094 549054 333538
rect 549302 326773 549362 362747
rect 549674 335334 550294 370778
rect 549674 334778 549706 335334
rect 550262 334778 550294 335334
rect 549299 326772 549365 326773
rect 549299 326708 549300 326772
rect 549364 326708 549365 326772
rect 549299 326707 549365 326708
rect 548434 297538 548466 298094
rect 549022 297538 549054 298094
rect 548434 262094 549054 297538
rect 549302 290733 549362 326707
rect 549674 299334 550294 334778
rect 549674 298778 549706 299334
rect 550262 298778 550294 299334
rect 549299 290732 549365 290733
rect 549299 290668 549300 290732
rect 549364 290668 549365 290732
rect 549299 290667 549365 290668
rect 548434 261538 548466 262094
rect 549022 261538 549054 262094
rect 548434 226094 549054 261538
rect 548434 225538 548466 226094
rect 549022 225538 549054 226094
rect 548434 190094 549054 225538
rect 548434 189538 548466 190094
rect 549022 189538 549054 190094
rect 548434 154094 549054 189538
rect 548434 153538 548466 154094
rect 549022 153538 549054 154094
rect 548434 118094 549054 153538
rect 548434 117538 548466 118094
rect 549022 117538 549054 118094
rect 548434 82094 549054 117538
rect 548434 81538 548466 82094
rect 549022 81538 549054 82094
rect 548434 46094 549054 81538
rect 548434 45538 548466 46094
rect 549022 45538 549054 46094
rect 548434 10094 549054 45538
rect 549302 19821 549362 290667
rect 549674 263334 550294 298778
rect 549674 262778 549706 263334
rect 550262 262778 550294 263334
rect 549674 227334 550294 262778
rect 549674 226778 549706 227334
rect 550262 226778 550294 227334
rect 549674 191334 550294 226778
rect 549674 190778 549706 191334
rect 550262 190778 550294 191334
rect 549674 155334 550294 190778
rect 549674 154778 549706 155334
rect 550262 154778 550294 155334
rect 549674 119334 550294 154778
rect 549674 118778 549706 119334
rect 550262 118778 550294 119334
rect 549674 83334 550294 118778
rect 549674 82778 549706 83334
rect 550262 82778 550294 83334
rect 549674 47334 550294 82778
rect 549674 46778 549706 47334
rect 550262 46778 550294 47334
rect 549299 19820 549365 19821
rect 549299 19756 549300 19820
rect 549364 19756 549365 19820
rect 549299 19755 549365 19756
rect 548434 9538 548466 10094
rect 549022 9538 549054 10094
rect 548434 -6106 549054 9538
rect 548434 -6662 548466 -6106
rect 549022 -6662 549054 -6106
rect 548434 -7654 549054 -6662
rect 549674 11334 550294 46778
rect 549674 10778 549706 11334
rect 550262 10778 550294 11334
rect 549674 -7066 550294 10778
rect 549674 -7622 549706 -7066
rect 550262 -7622 550294 -7066
rect 549674 -7654 550294 -7622
rect 576994 704838 577614 711590
rect 576994 704282 577026 704838
rect 577582 704282 577614 704838
rect 576994 686654 577614 704282
rect 576994 686098 577026 686654
rect 577582 686098 577614 686654
rect 576994 650654 577614 686098
rect 576994 650098 577026 650654
rect 577582 650098 577614 650654
rect 576994 614654 577614 650098
rect 576994 614098 577026 614654
rect 577582 614098 577614 614654
rect 576994 578654 577614 614098
rect 576994 578098 577026 578654
rect 577582 578098 577614 578654
rect 576994 542654 577614 578098
rect 576994 542098 577026 542654
rect 577582 542098 577614 542654
rect 576994 506654 577614 542098
rect 576994 506098 577026 506654
rect 577582 506098 577614 506654
rect 576994 470654 577614 506098
rect 576994 470098 577026 470654
rect 577582 470098 577614 470654
rect 576994 434654 577614 470098
rect 576994 434098 577026 434654
rect 577582 434098 577614 434654
rect 576994 398654 577614 434098
rect 576994 398098 577026 398654
rect 577582 398098 577614 398654
rect 576994 362654 577614 398098
rect 576994 362098 577026 362654
rect 577582 362098 577614 362654
rect 576994 326654 577614 362098
rect 576994 326098 577026 326654
rect 577582 326098 577614 326654
rect 576994 290654 577614 326098
rect 576994 290098 577026 290654
rect 577582 290098 577614 290654
rect 576994 254654 577614 290098
rect 576994 254098 577026 254654
rect 577582 254098 577614 254654
rect 576994 218654 577614 254098
rect 576994 218098 577026 218654
rect 577582 218098 577614 218654
rect 576994 182654 577614 218098
rect 576994 182098 577026 182654
rect 577582 182098 577614 182654
rect 576994 146654 577614 182098
rect 576994 146098 577026 146654
rect 577582 146098 577614 146654
rect 576994 110654 577614 146098
rect 576994 110098 577026 110654
rect 577582 110098 577614 110654
rect 576994 74654 577614 110098
rect 576994 74098 577026 74654
rect 577582 74098 577614 74654
rect 576994 38654 577614 74098
rect 576994 38098 577026 38654
rect 577582 38098 577614 38654
rect 576994 2654 577614 38098
rect 576994 2098 577026 2654
rect 577582 2098 577614 2654
rect 576994 -346 577614 2098
rect 576994 -902 577026 -346
rect 577582 -902 577614 -346
rect 576994 -7654 577614 -902
rect 578234 705798 578854 711590
rect 578234 705242 578266 705798
rect 578822 705242 578854 705798
rect 578234 687894 578854 705242
rect 578234 687338 578266 687894
rect 578822 687338 578854 687894
rect 578234 651894 578854 687338
rect 578234 651338 578266 651894
rect 578822 651338 578854 651894
rect 578234 615894 578854 651338
rect 578234 615338 578266 615894
rect 578822 615338 578854 615894
rect 578234 579894 578854 615338
rect 578234 579338 578266 579894
rect 578822 579338 578854 579894
rect 578234 543894 578854 579338
rect 578234 543338 578266 543894
rect 578822 543338 578854 543894
rect 578234 507894 578854 543338
rect 578234 507338 578266 507894
rect 578822 507338 578854 507894
rect 578234 471894 578854 507338
rect 578234 471338 578266 471894
rect 578822 471338 578854 471894
rect 578234 435894 578854 471338
rect 578234 435338 578266 435894
rect 578822 435338 578854 435894
rect 578234 399894 578854 435338
rect 578234 399338 578266 399894
rect 578822 399338 578854 399894
rect 578234 363894 578854 399338
rect 578234 363338 578266 363894
rect 578822 363338 578854 363894
rect 578234 327894 578854 363338
rect 578234 327338 578266 327894
rect 578822 327338 578854 327894
rect 578234 291894 578854 327338
rect 578234 291338 578266 291894
rect 578822 291338 578854 291894
rect 578234 255894 578854 291338
rect 578234 255338 578266 255894
rect 578822 255338 578854 255894
rect 578234 219894 578854 255338
rect 578234 219338 578266 219894
rect 578822 219338 578854 219894
rect 578234 183894 578854 219338
rect 578234 183338 578266 183894
rect 578822 183338 578854 183894
rect 578234 147894 578854 183338
rect 578234 147338 578266 147894
rect 578822 147338 578854 147894
rect 578234 111894 578854 147338
rect 578234 111338 578266 111894
rect 578822 111338 578854 111894
rect 578234 75894 578854 111338
rect 578234 75338 578266 75894
rect 578822 75338 578854 75894
rect 578234 39894 578854 75338
rect 578234 39338 578266 39894
rect 578822 39338 578854 39894
rect 578234 3894 578854 39338
rect 578234 3338 578266 3894
rect 578822 3338 578854 3894
rect 578234 -1306 578854 3338
rect 578234 -1862 578266 -1306
rect 578822 -1862 578854 -1306
rect 578234 -7654 578854 -1862
rect 579474 706758 580094 711590
rect 579474 706202 579506 706758
rect 580062 706202 580094 706758
rect 579474 689134 580094 706202
rect 579474 688578 579506 689134
rect 580062 688578 580094 689134
rect 579474 653134 580094 688578
rect 579474 652578 579506 653134
rect 580062 652578 580094 653134
rect 579474 617134 580094 652578
rect 579474 616578 579506 617134
rect 580062 616578 580094 617134
rect 579474 581134 580094 616578
rect 579474 580578 579506 581134
rect 580062 580578 580094 581134
rect 579474 545134 580094 580578
rect 579474 544578 579506 545134
rect 580062 544578 580094 545134
rect 579474 509134 580094 544578
rect 579474 508578 579506 509134
rect 580062 508578 580094 509134
rect 579474 473134 580094 508578
rect 579474 472578 579506 473134
rect 580062 472578 580094 473134
rect 579474 437134 580094 472578
rect 579474 436578 579506 437134
rect 580062 436578 580094 437134
rect 579474 401134 580094 436578
rect 579474 400578 579506 401134
rect 580062 400578 580094 401134
rect 579474 365134 580094 400578
rect 579474 364578 579506 365134
rect 580062 364578 580094 365134
rect 579474 329134 580094 364578
rect 579474 328578 579506 329134
rect 580062 328578 580094 329134
rect 579474 293134 580094 328578
rect 579474 292578 579506 293134
rect 580062 292578 580094 293134
rect 579474 257134 580094 292578
rect 579474 256578 579506 257134
rect 580062 256578 580094 257134
rect 579474 221134 580094 256578
rect 579474 220578 579506 221134
rect 580062 220578 580094 221134
rect 579474 185134 580094 220578
rect 579474 184578 579506 185134
rect 580062 184578 580094 185134
rect 579474 149134 580094 184578
rect 579474 148578 579506 149134
rect 580062 148578 580094 149134
rect 579474 113134 580094 148578
rect 579474 112578 579506 113134
rect 580062 112578 580094 113134
rect 579474 77134 580094 112578
rect 579474 76578 579506 77134
rect 580062 76578 580094 77134
rect 579474 41134 580094 76578
rect 579474 40578 579506 41134
rect 580062 40578 580094 41134
rect 579474 5134 580094 40578
rect 579474 4578 579506 5134
rect 580062 4578 580094 5134
rect 579474 -2266 580094 4578
rect 579474 -2822 579506 -2266
rect 580062 -2822 580094 -2266
rect 579474 -7654 580094 -2822
rect 580714 707718 581334 711590
rect 580714 707162 580746 707718
rect 581302 707162 581334 707718
rect 580714 690374 581334 707162
rect 580714 689818 580746 690374
rect 581302 689818 581334 690374
rect 580714 654374 581334 689818
rect 580714 653818 580746 654374
rect 581302 653818 581334 654374
rect 580714 618374 581334 653818
rect 580714 617818 580746 618374
rect 581302 617818 581334 618374
rect 580714 582374 581334 617818
rect 580714 581818 580746 582374
rect 581302 581818 581334 582374
rect 580714 546374 581334 581818
rect 580714 545818 580746 546374
rect 581302 545818 581334 546374
rect 580714 510374 581334 545818
rect 580714 509818 580746 510374
rect 581302 509818 581334 510374
rect 580714 474374 581334 509818
rect 580714 473818 580746 474374
rect 581302 473818 581334 474374
rect 580714 438374 581334 473818
rect 580714 437818 580746 438374
rect 581302 437818 581334 438374
rect 580714 402374 581334 437818
rect 580714 401818 580746 402374
rect 581302 401818 581334 402374
rect 580714 366374 581334 401818
rect 580714 365818 580746 366374
rect 581302 365818 581334 366374
rect 580714 330374 581334 365818
rect 580714 329818 580746 330374
rect 581302 329818 581334 330374
rect 580714 294374 581334 329818
rect 580714 293818 580746 294374
rect 581302 293818 581334 294374
rect 580714 258374 581334 293818
rect 580714 257818 580746 258374
rect 581302 257818 581334 258374
rect 580714 222374 581334 257818
rect 580714 221818 580746 222374
rect 581302 221818 581334 222374
rect 580714 186374 581334 221818
rect 580714 185818 580746 186374
rect 581302 185818 581334 186374
rect 580714 150374 581334 185818
rect 580714 149818 580746 150374
rect 581302 149818 581334 150374
rect 580714 114374 581334 149818
rect 580714 113818 580746 114374
rect 581302 113818 581334 114374
rect 580714 78374 581334 113818
rect 580714 77818 580746 78374
rect 581302 77818 581334 78374
rect 580714 42374 581334 77818
rect 580714 41818 580746 42374
rect 581302 41818 581334 42374
rect 580714 6374 581334 41818
rect 580714 5818 580746 6374
rect 581302 5818 581334 6374
rect 580714 -3226 581334 5818
rect 580714 -3782 580746 -3226
rect 581302 -3782 581334 -3226
rect 580714 -7654 581334 -3782
rect 581954 708678 582574 711590
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 581954 708122 581986 708678
rect 582542 708122 582574 708678
rect 581954 691614 582574 708122
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581954 691058 581986 691614
rect 582542 691058 582574 691614
rect 581954 655614 582574 691058
rect 581954 655058 581986 655614
rect 582542 655058 582574 655614
rect 581954 619614 582574 655058
rect 581954 619058 581986 619614
rect 582542 619058 582574 619614
rect 581954 583614 582574 619058
rect 581954 583058 581986 583614
rect 582542 583058 582574 583614
rect 581954 547614 582574 583058
rect 581954 547058 581986 547614
rect 582542 547058 582574 547614
rect 581954 511614 582574 547058
rect 581954 511058 581986 511614
rect 582542 511058 582574 511614
rect 581954 475614 582574 511058
rect 581954 475058 581986 475614
rect 582542 475058 582574 475614
rect 581954 439614 582574 475058
rect 581954 439058 581986 439614
rect 582542 439058 582574 439614
rect 581954 403614 582574 439058
rect 581954 403058 581986 403614
rect 582542 403058 582574 403614
rect 581954 367614 582574 403058
rect 581954 367058 581986 367614
rect 582542 367058 582574 367614
rect 581954 331614 582574 367058
rect 581954 331058 581986 331614
rect 582542 331058 582574 331614
rect 581954 295614 582574 331058
rect 581954 295058 581986 295614
rect 582542 295058 582574 295614
rect 581954 259614 582574 295058
rect 581954 259058 581986 259614
rect 582542 259058 582574 259614
rect 581954 223614 582574 259058
rect 581954 223058 581986 223614
rect 582542 223058 582574 223614
rect 581954 187614 582574 223058
rect 581954 187058 581986 187614
rect 582542 187058 582574 187614
rect 581954 151614 582574 187058
rect 581954 151058 581986 151614
rect 582542 151058 582574 151614
rect 581954 115614 582574 151058
rect 581954 115058 581986 115614
rect 582542 115058 582574 115614
rect 581954 79614 582574 115058
rect 581954 79058 581986 79614
rect 582542 79058 582574 79614
rect 581954 43614 582574 79058
rect 581954 43058 581986 43614
rect 582542 43058 582574 43614
rect 581954 7614 582574 43058
rect 581954 7058 581986 7614
rect 582542 7058 582574 7614
rect 581954 -4186 582574 7058
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 686654 585930 704282
rect 585310 686098 585342 686654
rect 585898 686098 585930 686654
rect 585310 650654 585930 686098
rect 585310 650098 585342 650654
rect 585898 650098 585930 650654
rect 585310 614654 585930 650098
rect 585310 614098 585342 614654
rect 585898 614098 585930 614654
rect 585310 578654 585930 614098
rect 585310 578098 585342 578654
rect 585898 578098 585930 578654
rect 585310 542654 585930 578098
rect 585310 542098 585342 542654
rect 585898 542098 585930 542654
rect 585310 506654 585930 542098
rect 585310 506098 585342 506654
rect 585898 506098 585930 506654
rect 585310 470654 585930 506098
rect 585310 470098 585342 470654
rect 585898 470098 585930 470654
rect 585310 434654 585930 470098
rect 585310 434098 585342 434654
rect 585898 434098 585930 434654
rect 585310 398654 585930 434098
rect 585310 398098 585342 398654
rect 585898 398098 585930 398654
rect 585310 362654 585930 398098
rect 585310 362098 585342 362654
rect 585898 362098 585930 362654
rect 585310 326654 585930 362098
rect 585310 326098 585342 326654
rect 585898 326098 585930 326654
rect 585310 290654 585930 326098
rect 585310 290098 585342 290654
rect 585898 290098 585930 290654
rect 585310 254654 585930 290098
rect 585310 254098 585342 254654
rect 585898 254098 585930 254654
rect 585310 218654 585930 254098
rect 585310 218098 585342 218654
rect 585898 218098 585930 218654
rect 585310 182654 585930 218098
rect 585310 182098 585342 182654
rect 585898 182098 585930 182654
rect 585310 146654 585930 182098
rect 585310 146098 585342 146654
rect 585898 146098 585930 146654
rect 585310 110654 585930 146098
rect 585310 110098 585342 110654
rect 585898 110098 585930 110654
rect 585310 74654 585930 110098
rect 585310 74098 585342 74654
rect 585898 74098 585930 74654
rect 585310 38654 585930 74098
rect 585310 38098 585342 38654
rect 585898 38098 585930 38654
rect 585310 2654 585930 38098
rect 585310 2098 585342 2654
rect 585898 2098 585930 2654
rect 585310 -346 585930 2098
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 687894 586890 705242
rect 586270 687338 586302 687894
rect 586858 687338 586890 687894
rect 586270 651894 586890 687338
rect 586270 651338 586302 651894
rect 586858 651338 586890 651894
rect 586270 615894 586890 651338
rect 586270 615338 586302 615894
rect 586858 615338 586890 615894
rect 586270 579894 586890 615338
rect 586270 579338 586302 579894
rect 586858 579338 586890 579894
rect 586270 543894 586890 579338
rect 586270 543338 586302 543894
rect 586858 543338 586890 543894
rect 586270 507894 586890 543338
rect 586270 507338 586302 507894
rect 586858 507338 586890 507894
rect 586270 471894 586890 507338
rect 586270 471338 586302 471894
rect 586858 471338 586890 471894
rect 586270 435894 586890 471338
rect 586270 435338 586302 435894
rect 586858 435338 586890 435894
rect 586270 399894 586890 435338
rect 586270 399338 586302 399894
rect 586858 399338 586890 399894
rect 586270 363894 586890 399338
rect 586270 363338 586302 363894
rect 586858 363338 586890 363894
rect 586270 327894 586890 363338
rect 586270 327338 586302 327894
rect 586858 327338 586890 327894
rect 586270 291894 586890 327338
rect 586270 291338 586302 291894
rect 586858 291338 586890 291894
rect 586270 255894 586890 291338
rect 586270 255338 586302 255894
rect 586858 255338 586890 255894
rect 586270 219894 586890 255338
rect 586270 219338 586302 219894
rect 586858 219338 586890 219894
rect 586270 183894 586890 219338
rect 586270 183338 586302 183894
rect 586858 183338 586890 183894
rect 586270 147894 586890 183338
rect 586270 147338 586302 147894
rect 586858 147338 586890 147894
rect 586270 111894 586890 147338
rect 586270 111338 586302 111894
rect 586858 111338 586890 111894
rect 586270 75894 586890 111338
rect 586270 75338 586302 75894
rect 586858 75338 586890 75894
rect 586270 39894 586890 75338
rect 586270 39338 586302 39894
rect 586858 39338 586890 39894
rect 586270 3894 586890 39338
rect 586270 3338 586302 3894
rect 586858 3338 586890 3894
rect 586270 -1306 586890 3338
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 689134 587850 706202
rect 587230 688578 587262 689134
rect 587818 688578 587850 689134
rect 587230 653134 587850 688578
rect 587230 652578 587262 653134
rect 587818 652578 587850 653134
rect 587230 617134 587850 652578
rect 587230 616578 587262 617134
rect 587818 616578 587850 617134
rect 587230 581134 587850 616578
rect 587230 580578 587262 581134
rect 587818 580578 587850 581134
rect 587230 545134 587850 580578
rect 587230 544578 587262 545134
rect 587818 544578 587850 545134
rect 587230 509134 587850 544578
rect 587230 508578 587262 509134
rect 587818 508578 587850 509134
rect 587230 473134 587850 508578
rect 587230 472578 587262 473134
rect 587818 472578 587850 473134
rect 587230 437134 587850 472578
rect 587230 436578 587262 437134
rect 587818 436578 587850 437134
rect 587230 401134 587850 436578
rect 587230 400578 587262 401134
rect 587818 400578 587850 401134
rect 587230 365134 587850 400578
rect 587230 364578 587262 365134
rect 587818 364578 587850 365134
rect 587230 329134 587850 364578
rect 587230 328578 587262 329134
rect 587818 328578 587850 329134
rect 587230 293134 587850 328578
rect 587230 292578 587262 293134
rect 587818 292578 587850 293134
rect 587230 257134 587850 292578
rect 587230 256578 587262 257134
rect 587818 256578 587850 257134
rect 587230 221134 587850 256578
rect 587230 220578 587262 221134
rect 587818 220578 587850 221134
rect 587230 185134 587850 220578
rect 587230 184578 587262 185134
rect 587818 184578 587850 185134
rect 587230 149134 587850 184578
rect 587230 148578 587262 149134
rect 587818 148578 587850 149134
rect 587230 113134 587850 148578
rect 587230 112578 587262 113134
rect 587818 112578 587850 113134
rect 587230 77134 587850 112578
rect 587230 76578 587262 77134
rect 587818 76578 587850 77134
rect 587230 41134 587850 76578
rect 587230 40578 587262 41134
rect 587818 40578 587850 41134
rect 587230 5134 587850 40578
rect 587230 4578 587262 5134
rect 587818 4578 587850 5134
rect 587230 -2266 587850 4578
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 690374 588810 707162
rect 588190 689818 588222 690374
rect 588778 689818 588810 690374
rect 588190 654374 588810 689818
rect 588190 653818 588222 654374
rect 588778 653818 588810 654374
rect 588190 618374 588810 653818
rect 588190 617818 588222 618374
rect 588778 617818 588810 618374
rect 588190 582374 588810 617818
rect 588190 581818 588222 582374
rect 588778 581818 588810 582374
rect 588190 546374 588810 581818
rect 588190 545818 588222 546374
rect 588778 545818 588810 546374
rect 588190 510374 588810 545818
rect 588190 509818 588222 510374
rect 588778 509818 588810 510374
rect 588190 474374 588810 509818
rect 588190 473818 588222 474374
rect 588778 473818 588810 474374
rect 588190 438374 588810 473818
rect 588190 437818 588222 438374
rect 588778 437818 588810 438374
rect 588190 402374 588810 437818
rect 588190 401818 588222 402374
rect 588778 401818 588810 402374
rect 588190 366374 588810 401818
rect 588190 365818 588222 366374
rect 588778 365818 588810 366374
rect 588190 330374 588810 365818
rect 588190 329818 588222 330374
rect 588778 329818 588810 330374
rect 588190 294374 588810 329818
rect 588190 293818 588222 294374
rect 588778 293818 588810 294374
rect 588190 258374 588810 293818
rect 588190 257818 588222 258374
rect 588778 257818 588810 258374
rect 588190 222374 588810 257818
rect 588190 221818 588222 222374
rect 588778 221818 588810 222374
rect 588190 186374 588810 221818
rect 588190 185818 588222 186374
rect 588778 185818 588810 186374
rect 588190 150374 588810 185818
rect 588190 149818 588222 150374
rect 588778 149818 588810 150374
rect 588190 114374 588810 149818
rect 588190 113818 588222 114374
rect 588778 113818 588810 114374
rect 588190 78374 588810 113818
rect 588190 77818 588222 78374
rect 588778 77818 588810 78374
rect 588190 42374 588810 77818
rect 588190 41818 588222 42374
rect 588778 41818 588810 42374
rect 588190 6374 588810 41818
rect 588190 5818 588222 6374
rect 588778 5818 588810 6374
rect 588190 -3226 588810 5818
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 691614 589770 708122
rect 589150 691058 589182 691614
rect 589738 691058 589770 691614
rect 589150 655614 589770 691058
rect 589150 655058 589182 655614
rect 589738 655058 589770 655614
rect 589150 619614 589770 655058
rect 589150 619058 589182 619614
rect 589738 619058 589770 619614
rect 589150 583614 589770 619058
rect 589150 583058 589182 583614
rect 589738 583058 589770 583614
rect 589150 547614 589770 583058
rect 589150 547058 589182 547614
rect 589738 547058 589770 547614
rect 589150 511614 589770 547058
rect 589150 511058 589182 511614
rect 589738 511058 589770 511614
rect 589150 475614 589770 511058
rect 589150 475058 589182 475614
rect 589738 475058 589770 475614
rect 589150 439614 589770 475058
rect 589150 439058 589182 439614
rect 589738 439058 589770 439614
rect 589150 403614 589770 439058
rect 589150 403058 589182 403614
rect 589738 403058 589770 403614
rect 589150 367614 589770 403058
rect 589150 367058 589182 367614
rect 589738 367058 589770 367614
rect 589150 331614 589770 367058
rect 589150 331058 589182 331614
rect 589738 331058 589770 331614
rect 589150 295614 589770 331058
rect 589150 295058 589182 295614
rect 589738 295058 589770 295614
rect 589150 259614 589770 295058
rect 589150 259058 589182 259614
rect 589738 259058 589770 259614
rect 589150 223614 589770 259058
rect 589150 223058 589182 223614
rect 589738 223058 589770 223614
rect 589150 187614 589770 223058
rect 589150 187058 589182 187614
rect 589738 187058 589770 187614
rect 589150 151614 589770 187058
rect 589150 151058 589182 151614
rect 589738 151058 589770 151614
rect 589150 115614 589770 151058
rect 589150 115058 589182 115614
rect 589738 115058 589770 115614
rect 589150 79614 589770 115058
rect 589150 79058 589182 79614
rect 589738 79058 589770 79614
rect 589150 43614 589770 79058
rect 589150 43058 589182 43614
rect 589738 43058 589770 43614
rect 589150 7614 589770 43058
rect 589150 7058 589182 7614
rect 589738 7058 589770 7614
rect 581954 -4742 581986 -4186
rect 582542 -4742 582574 -4186
rect 581954 -7654 582574 -4742
rect 589150 -4186 589770 7058
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 692854 590730 709082
rect 590110 692298 590142 692854
rect 590698 692298 590730 692854
rect 590110 656854 590730 692298
rect 590110 656298 590142 656854
rect 590698 656298 590730 656854
rect 590110 620854 590730 656298
rect 590110 620298 590142 620854
rect 590698 620298 590730 620854
rect 590110 584854 590730 620298
rect 590110 584298 590142 584854
rect 590698 584298 590730 584854
rect 590110 548854 590730 584298
rect 590110 548298 590142 548854
rect 590698 548298 590730 548854
rect 590110 512854 590730 548298
rect 590110 512298 590142 512854
rect 590698 512298 590730 512854
rect 590110 476854 590730 512298
rect 590110 476298 590142 476854
rect 590698 476298 590730 476854
rect 590110 440854 590730 476298
rect 590110 440298 590142 440854
rect 590698 440298 590730 440854
rect 590110 404854 590730 440298
rect 590110 404298 590142 404854
rect 590698 404298 590730 404854
rect 590110 368854 590730 404298
rect 590110 368298 590142 368854
rect 590698 368298 590730 368854
rect 590110 332854 590730 368298
rect 590110 332298 590142 332854
rect 590698 332298 590730 332854
rect 590110 296854 590730 332298
rect 590110 296298 590142 296854
rect 590698 296298 590730 296854
rect 590110 260854 590730 296298
rect 590110 260298 590142 260854
rect 590698 260298 590730 260854
rect 590110 224854 590730 260298
rect 590110 224298 590142 224854
rect 590698 224298 590730 224854
rect 590110 188854 590730 224298
rect 590110 188298 590142 188854
rect 590698 188298 590730 188854
rect 590110 152854 590730 188298
rect 590110 152298 590142 152854
rect 590698 152298 590730 152854
rect 590110 116854 590730 152298
rect 590110 116298 590142 116854
rect 590698 116298 590730 116854
rect 590110 80854 590730 116298
rect 590110 80298 590142 80854
rect 590698 80298 590730 80854
rect 590110 44854 590730 80298
rect 590110 44298 590142 44854
rect 590698 44298 590730 44854
rect 590110 8854 590730 44298
rect 590110 8298 590142 8854
rect 590698 8298 590730 8854
rect 590110 -5146 590730 8298
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 694094 591690 710042
rect 591070 693538 591102 694094
rect 591658 693538 591690 694094
rect 591070 658094 591690 693538
rect 591070 657538 591102 658094
rect 591658 657538 591690 658094
rect 591070 622094 591690 657538
rect 591070 621538 591102 622094
rect 591658 621538 591690 622094
rect 591070 586094 591690 621538
rect 591070 585538 591102 586094
rect 591658 585538 591690 586094
rect 591070 550094 591690 585538
rect 591070 549538 591102 550094
rect 591658 549538 591690 550094
rect 591070 514094 591690 549538
rect 591070 513538 591102 514094
rect 591658 513538 591690 514094
rect 591070 478094 591690 513538
rect 591070 477538 591102 478094
rect 591658 477538 591690 478094
rect 591070 442094 591690 477538
rect 591070 441538 591102 442094
rect 591658 441538 591690 442094
rect 591070 406094 591690 441538
rect 591070 405538 591102 406094
rect 591658 405538 591690 406094
rect 591070 370094 591690 405538
rect 591070 369538 591102 370094
rect 591658 369538 591690 370094
rect 591070 334094 591690 369538
rect 591070 333538 591102 334094
rect 591658 333538 591690 334094
rect 591070 298094 591690 333538
rect 591070 297538 591102 298094
rect 591658 297538 591690 298094
rect 591070 262094 591690 297538
rect 591070 261538 591102 262094
rect 591658 261538 591690 262094
rect 591070 226094 591690 261538
rect 591070 225538 591102 226094
rect 591658 225538 591690 226094
rect 591070 190094 591690 225538
rect 591070 189538 591102 190094
rect 591658 189538 591690 190094
rect 591070 154094 591690 189538
rect 591070 153538 591102 154094
rect 591658 153538 591690 154094
rect 591070 118094 591690 153538
rect 591070 117538 591102 118094
rect 591658 117538 591690 118094
rect 591070 82094 591690 117538
rect 591070 81538 591102 82094
rect 591658 81538 591690 82094
rect 591070 46094 591690 81538
rect 591070 45538 591102 46094
rect 591658 45538 591690 46094
rect 591070 10094 591690 45538
rect 591070 9538 591102 10094
rect 591658 9538 591690 10094
rect 591070 -6106 591690 9538
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 695334 592650 711002
rect 592030 694778 592062 695334
rect 592618 694778 592650 695334
rect 592030 659334 592650 694778
rect 592030 658778 592062 659334
rect 592618 658778 592650 659334
rect 592030 623334 592650 658778
rect 592030 622778 592062 623334
rect 592618 622778 592650 623334
rect 592030 587334 592650 622778
rect 592030 586778 592062 587334
rect 592618 586778 592650 587334
rect 592030 551334 592650 586778
rect 592030 550778 592062 551334
rect 592618 550778 592650 551334
rect 592030 515334 592650 550778
rect 592030 514778 592062 515334
rect 592618 514778 592650 515334
rect 592030 479334 592650 514778
rect 592030 478778 592062 479334
rect 592618 478778 592650 479334
rect 592030 443334 592650 478778
rect 592030 442778 592062 443334
rect 592618 442778 592650 443334
rect 592030 407334 592650 442778
rect 592030 406778 592062 407334
rect 592618 406778 592650 407334
rect 592030 371334 592650 406778
rect 592030 370778 592062 371334
rect 592618 370778 592650 371334
rect 592030 335334 592650 370778
rect 592030 334778 592062 335334
rect 592618 334778 592650 335334
rect 592030 299334 592650 334778
rect 592030 298778 592062 299334
rect 592618 298778 592650 299334
rect 592030 263334 592650 298778
rect 592030 262778 592062 263334
rect 592618 262778 592650 263334
rect 592030 227334 592650 262778
rect 592030 226778 592062 227334
rect 592618 226778 592650 227334
rect 592030 191334 592650 226778
rect 592030 190778 592062 191334
rect 592618 190778 592650 191334
rect 592030 155334 592650 190778
rect 592030 154778 592062 155334
rect 592618 154778 592650 155334
rect 592030 119334 592650 154778
rect 592030 118778 592062 119334
rect 592618 118778 592650 119334
rect 592030 83334 592650 118778
rect 592030 82778 592062 83334
rect 592618 82778 592650 83334
rect 592030 47334 592650 82778
rect 592030 46778 592062 47334
rect 592618 46778 592650 47334
rect 592030 11334 592650 46778
rect 592030 10778 592062 11334
rect 592618 10778 592650 11334
rect 592030 -7066 592650 10778
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 694778 -8138 695334
rect -8694 658778 -8138 659334
rect -8694 622778 -8138 623334
rect -8694 586778 -8138 587334
rect -8694 550778 -8138 551334
rect -8694 514778 -8138 515334
rect -8694 478778 -8138 479334
rect -8694 442778 -8138 443334
rect -8694 406778 -8138 407334
rect -8694 370778 -8138 371334
rect -8694 334778 -8138 335334
rect -8694 298778 -8138 299334
rect -8694 262778 -8138 263334
rect -8694 226778 -8138 227334
rect -8694 190778 -8138 191334
rect -8694 154778 -8138 155334
rect -8694 118778 -8138 119334
rect -8694 82778 -8138 83334
rect -8694 46778 -8138 47334
rect -8694 10778 -8138 11334
rect -7734 710042 -7178 710598
rect -7734 693538 -7178 694094
rect -7734 657538 -7178 658094
rect -7734 621538 -7178 622094
rect -7734 585538 -7178 586094
rect -7734 549538 -7178 550094
rect -7734 513538 -7178 514094
rect -7734 477538 -7178 478094
rect -7734 441538 -7178 442094
rect -7734 405538 -7178 406094
rect -7734 369538 -7178 370094
rect -7734 333538 -7178 334094
rect -7734 297538 -7178 298094
rect -7734 261538 -7178 262094
rect -7734 225538 -7178 226094
rect -7734 189538 -7178 190094
rect -7734 153538 -7178 154094
rect -7734 117538 -7178 118094
rect -7734 81538 -7178 82094
rect -7734 45538 -7178 46094
rect -7734 9538 -7178 10094
rect -6774 709082 -6218 709638
rect -6774 692298 -6218 692854
rect -6774 656298 -6218 656854
rect -6774 620298 -6218 620854
rect -6774 584298 -6218 584854
rect -6774 548298 -6218 548854
rect -6774 512298 -6218 512854
rect -6774 476298 -6218 476854
rect -6774 440298 -6218 440854
rect -6774 404298 -6218 404854
rect -6774 368298 -6218 368854
rect -6774 332298 -6218 332854
rect -6774 296298 -6218 296854
rect -6774 260298 -6218 260854
rect -6774 224298 -6218 224854
rect -6774 188298 -6218 188854
rect -6774 152298 -6218 152854
rect -6774 116298 -6218 116854
rect -6774 80298 -6218 80854
rect -6774 44298 -6218 44854
rect -6774 8298 -6218 8854
rect -5814 708122 -5258 708678
rect -5814 691058 -5258 691614
rect -5814 655058 -5258 655614
rect -5814 619058 -5258 619614
rect -5814 583058 -5258 583614
rect -5814 547058 -5258 547614
rect -5814 511058 -5258 511614
rect -5814 475058 -5258 475614
rect -5814 439058 -5258 439614
rect -5814 403058 -5258 403614
rect -5814 367058 -5258 367614
rect -5814 331058 -5258 331614
rect -5814 295058 -5258 295614
rect -5814 259058 -5258 259614
rect -5814 223058 -5258 223614
rect -5814 187058 -5258 187614
rect -5814 151058 -5258 151614
rect -5814 115058 -5258 115614
rect -5814 79058 -5258 79614
rect -5814 43058 -5258 43614
rect -5814 7058 -5258 7614
rect -4854 707162 -4298 707718
rect -4854 689818 -4298 690374
rect -4854 653818 -4298 654374
rect -4854 617818 -4298 618374
rect -4854 581818 -4298 582374
rect -4854 545818 -4298 546374
rect -4854 509818 -4298 510374
rect -4854 473818 -4298 474374
rect -4854 437818 -4298 438374
rect -4854 401818 -4298 402374
rect -4854 365818 -4298 366374
rect -4854 329818 -4298 330374
rect -4854 293818 -4298 294374
rect -4854 257818 -4298 258374
rect -4854 221818 -4298 222374
rect -4854 185818 -4298 186374
rect -4854 149818 -4298 150374
rect -4854 113818 -4298 114374
rect -4854 77818 -4298 78374
rect -4854 41818 -4298 42374
rect -4854 5818 -4298 6374
rect -3894 706202 -3338 706758
rect -3894 688578 -3338 689134
rect -3894 652578 -3338 653134
rect -3894 616578 -3338 617134
rect -3894 580578 -3338 581134
rect -3894 544578 -3338 545134
rect -3894 508578 -3338 509134
rect -3894 472578 -3338 473134
rect -3894 436578 -3338 437134
rect -3894 400578 -3338 401134
rect -3894 364578 -3338 365134
rect -3894 328578 -3338 329134
rect -3894 292578 -3338 293134
rect -3894 256578 -3338 257134
rect -3894 220578 -3338 221134
rect -3894 184578 -3338 185134
rect -3894 148578 -3338 149134
rect -3894 112578 -3338 113134
rect -3894 76578 -3338 77134
rect -3894 40578 -3338 41134
rect -3894 4578 -3338 5134
rect -2934 705242 -2378 705798
rect -2934 687338 -2378 687894
rect -2934 651338 -2378 651894
rect -2934 615338 -2378 615894
rect -2934 579338 -2378 579894
rect -2934 543338 -2378 543894
rect -2934 507338 -2378 507894
rect -2934 471338 -2378 471894
rect -2934 435338 -2378 435894
rect -2934 399338 -2378 399894
rect -2934 363338 -2378 363894
rect -2934 327338 -2378 327894
rect -2934 291338 -2378 291894
rect -2934 255338 -2378 255894
rect -2934 219338 -2378 219894
rect -2934 183338 -2378 183894
rect -2934 147338 -2378 147894
rect -2934 111338 -2378 111894
rect -2934 75338 -2378 75894
rect -2934 39338 -2378 39894
rect -2934 3338 -2378 3894
rect -1974 704282 -1418 704838
rect -1974 686098 -1418 686654
rect -1974 650098 -1418 650654
rect -1974 614098 -1418 614654
rect -1974 578098 -1418 578654
rect -1974 542098 -1418 542654
rect -1974 506098 -1418 506654
rect -1974 470098 -1418 470654
rect -1974 434098 -1418 434654
rect -1974 398098 -1418 398654
rect -1974 362098 -1418 362654
rect -1974 326098 -1418 326654
rect -1974 290098 -1418 290654
rect -1974 254098 -1418 254654
rect -1974 218098 -1418 218654
rect -1974 182098 -1418 182654
rect -1974 146098 -1418 146654
rect -1974 110098 -1418 110654
rect -1974 74098 -1418 74654
rect -1974 38098 -1418 38654
rect -1974 2098 -1418 2654
rect -1974 -902 -1418 -346
rect 1026 704282 1582 704838
rect 1026 686098 1582 686654
rect 1026 650098 1582 650654
rect 1026 614098 1582 614654
rect 1026 578098 1582 578654
rect 1026 542098 1582 542654
rect 1026 506098 1582 506654
rect 1026 470098 1582 470654
rect 1026 434098 1582 434654
rect 1026 398098 1582 398654
rect 1026 362098 1582 362654
rect 1026 326098 1582 326654
rect 1026 290098 1582 290654
rect 1026 254098 1582 254654
rect 1026 218098 1582 218654
rect 1026 182098 1582 182654
rect 1026 146098 1582 146654
rect 1026 110098 1582 110654
rect 1026 74098 1582 74654
rect 1026 38098 1582 38654
rect 1026 2098 1582 2654
rect 1026 -902 1582 -346
rect -2934 -1862 -2378 -1306
rect -3894 -2822 -3338 -2266
rect -4854 -3782 -4298 -3226
rect -5814 -4742 -5258 -4186
rect -6774 -5702 -6218 -5146
rect -7734 -6662 -7178 -6106
rect -8694 -7622 -8138 -7066
rect 2266 705242 2822 705798
rect 2266 687338 2822 687894
rect 2266 651338 2822 651894
rect 2266 615338 2822 615894
rect 2266 579338 2822 579894
rect 2266 543338 2822 543894
rect 2266 507338 2822 507894
rect 2266 471338 2822 471894
rect 2266 435338 2822 435894
rect 2266 399338 2822 399894
rect 2266 363338 2822 363894
rect 2266 327338 2822 327894
rect 2266 291338 2822 291894
rect 2266 255338 2822 255894
rect 2266 219338 2822 219894
rect 2266 183338 2822 183894
rect 2266 147338 2822 147894
rect 2266 111338 2822 111894
rect 2266 75338 2822 75894
rect 2266 39338 2822 39894
rect 2266 3338 2822 3894
rect 2266 -1862 2822 -1306
rect 3506 706202 4062 706758
rect 3506 688578 4062 689134
rect 3506 652578 4062 653134
rect 3506 616578 4062 617134
rect 3506 580578 4062 581134
rect 3506 544578 4062 545134
rect 3506 508578 4062 509134
rect 3506 472578 4062 473134
rect 3506 436578 4062 437134
rect 3506 400578 4062 401134
rect 3506 364578 4062 365134
rect 3506 328578 4062 329134
rect 3506 292578 4062 293134
rect 3506 256578 4062 257134
rect 3506 220578 4062 221134
rect 3506 184578 4062 185134
rect 3506 148578 4062 149134
rect 3506 112578 4062 113134
rect 3506 76578 4062 77134
rect 3506 40578 4062 41134
rect 3506 4578 4062 5134
rect 3506 -2822 4062 -2266
rect 4746 707162 5302 707718
rect 4746 689818 5302 690374
rect 4746 653818 5302 654374
rect 4746 617818 5302 618374
rect 4746 581818 5302 582374
rect 4746 545818 5302 546374
rect 4746 509818 5302 510374
rect 4746 473818 5302 474374
rect 4746 437818 5302 438374
rect 4746 401818 5302 402374
rect 4746 365818 5302 366374
rect 4746 329818 5302 330374
rect 4746 293818 5302 294374
rect 4746 257818 5302 258374
rect 4746 221818 5302 222374
rect 4746 185818 5302 186374
rect 4746 149818 5302 150374
rect 4746 113818 5302 114374
rect 4746 77818 5302 78374
rect 4746 41818 5302 42374
rect 4746 5818 5302 6374
rect 4746 -3782 5302 -3226
rect 5986 708122 6542 708678
rect 5986 691058 6542 691614
rect 5986 655058 6542 655614
rect 5986 619058 6542 619614
rect 5986 583058 6542 583614
rect 5986 547058 6542 547614
rect 5986 511058 6542 511614
rect 5986 475058 6542 475614
rect 5986 439058 6542 439614
rect 5986 403058 6542 403614
rect 5986 367058 6542 367614
rect 5986 331058 6542 331614
rect 5986 295058 6542 295614
rect 5986 259058 6542 259614
rect 5986 223058 6542 223614
rect 5986 187058 6542 187614
rect 5986 151058 6542 151614
rect 5986 115058 6542 115614
rect 5986 79058 6542 79614
rect 5986 43058 6542 43614
rect 5986 7058 6542 7614
rect 5986 -4742 6542 -4186
rect 7226 709082 7782 709638
rect 7226 692298 7782 692854
rect 7226 656298 7782 656854
rect 7226 620298 7782 620854
rect 7226 584298 7782 584854
rect 7226 548298 7782 548854
rect 7226 512298 7782 512854
rect 7226 476298 7782 476854
rect 7226 440298 7782 440854
rect 7226 404298 7782 404854
rect 7226 368298 7782 368854
rect 7226 332298 7782 332854
rect 7226 296298 7782 296854
rect 7226 260298 7782 260854
rect 7226 224298 7782 224854
rect 7226 188298 7782 188854
rect 7226 152298 7782 152854
rect 7226 116298 7782 116854
rect 7226 80298 7782 80854
rect 7226 44298 7782 44854
rect 7226 8298 7782 8854
rect 7226 -5702 7782 -5146
rect 8466 710042 9022 710598
rect 8466 693538 9022 694094
rect 8466 657538 9022 658094
rect 8466 621538 9022 622094
rect 8466 585538 9022 586094
rect 8466 549538 9022 550094
rect 8466 513538 9022 514094
rect 8466 477538 9022 478094
rect 8466 441538 9022 442094
rect 8466 405538 9022 406094
rect 8466 369538 9022 370094
rect 8466 333538 9022 334094
rect 8466 297538 9022 298094
rect 8466 261538 9022 262094
rect 8466 225538 9022 226094
rect 8466 189538 9022 190094
rect 8466 153538 9022 154094
rect 8466 117538 9022 118094
rect 8466 81538 9022 82094
rect 8466 45538 9022 46094
rect 8466 9538 9022 10094
rect 8466 -6662 9022 -6106
rect 9706 711002 10262 711558
rect 9706 694778 10262 695334
rect 9706 658778 10262 659334
rect 9706 622778 10262 623334
rect 9706 586778 10262 587334
rect 9706 550778 10262 551334
rect 9706 514778 10262 515334
rect 9706 478778 10262 479334
rect 9706 442778 10262 443334
rect 9706 406778 10262 407334
rect 9706 370778 10262 371334
rect 9706 334778 10262 335334
rect 9706 298778 10262 299334
rect 9706 262778 10262 263334
rect 9706 226778 10262 227334
rect 9706 190778 10262 191334
rect 9706 154778 10262 155334
rect 9706 118778 10262 119334
rect 9706 82778 10262 83334
rect 9706 46778 10262 47334
rect 9706 10778 10262 11334
rect 9706 -7622 10262 -7066
rect 37026 704282 37582 704838
rect 37026 686098 37582 686654
rect 37026 650098 37582 650654
rect 37026 614098 37582 614654
rect 37026 578098 37582 578654
rect 37026 542098 37582 542654
rect 37026 506098 37582 506654
rect 37026 470098 37582 470654
rect 37026 434098 37582 434654
rect 37026 398098 37582 398654
rect 37026 362098 37582 362654
rect 37026 326098 37582 326654
rect 37026 290098 37582 290654
rect 37026 254098 37582 254654
rect 37026 218098 37582 218654
rect 37026 182098 37582 182654
rect 37026 146098 37582 146654
rect 37026 110098 37582 110654
rect 37026 74098 37582 74654
rect 37026 38098 37582 38654
rect 37026 2098 37582 2654
rect 37026 -902 37582 -346
rect 38266 705242 38822 705798
rect 38266 687338 38822 687894
rect 38266 651338 38822 651894
rect 38266 615338 38822 615894
rect 38266 579338 38822 579894
rect 38266 543338 38822 543894
rect 38266 507338 38822 507894
rect 38266 471338 38822 471894
rect 38266 435338 38822 435894
rect 38266 399338 38822 399894
rect 38266 363338 38822 363894
rect 38266 327338 38822 327894
rect 38266 291338 38822 291894
rect 38266 255338 38822 255894
rect 38266 219338 38822 219894
rect 38266 183338 38822 183894
rect 38266 147338 38822 147894
rect 38266 111338 38822 111894
rect 38266 75338 38822 75894
rect 38266 39338 38822 39894
rect 38266 3338 38822 3894
rect 38266 -1862 38822 -1306
rect 39506 706202 40062 706758
rect 39506 688578 40062 689134
rect 39506 652578 40062 653134
rect 39506 616578 40062 617134
rect 39506 580578 40062 581134
rect 39506 544578 40062 545134
rect 39506 508578 40062 509134
rect 39506 472578 40062 473134
rect 39506 436578 40062 437134
rect 39506 400578 40062 401134
rect 39506 364578 40062 365134
rect 39506 328578 40062 329134
rect 39506 292578 40062 293134
rect 39506 256578 40062 257134
rect 39506 220578 40062 221134
rect 39506 184578 40062 185134
rect 39506 148578 40062 149134
rect 39506 112578 40062 113134
rect 39506 76578 40062 77134
rect 39506 40578 40062 41134
rect 39506 4578 40062 5134
rect 39506 -2822 40062 -2266
rect 40746 707162 41302 707718
rect 40746 689818 41302 690374
rect 40746 653818 41302 654374
rect 40746 617818 41302 618374
rect 40746 581818 41302 582374
rect 40746 545818 41302 546374
rect 40746 509818 41302 510374
rect 40746 473818 41302 474374
rect 40746 437818 41302 438374
rect 40746 401818 41302 402374
rect 40746 365818 41302 366374
rect 40746 329818 41302 330374
rect 40746 293818 41302 294374
rect 40746 257818 41302 258374
rect 40746 221818 41302 222374
rect 40746 185818 41302 186374
rect 40746 149818 41302 150374
rect 40746 113818 41302 114374
rect 40746 77818 41302 78374
rect 40746 41818 41302 42374
rect 40746 5818 41302 6374
rect 40746 -3782 41302 -3226
rect 41986 708122 42542 708678
rect 41986 691058 42542 691614
rect 41986 655058 42542 655614
rect 41986 619058 42542 619614
rect 41986 583058 42542 583614
rect 41986 547058 42542 547614
rect 41986 511058 42542 511614
rect 41986 475058 42542 475614
rect 41986 439058 42542 439614
rect 41986 403058 42542 403614
rect 41986 367058 42542 367614
rect 41986 331058 42542 331614
rect 41986 295058 42542 295614
rect 41986 259058 42542 259614
rect 41986 223058 42542 223614
rect 41986 187058 42542 187614
rect 41986 151058 42542 151614
rect 41986 115058 42542 115614
rect 41986 79058 42542 79614
rect 41986 43058 42542 43614
rect 41986 7058 42542 7614
rect 41986 -4742 42542 -4186
rect 43226 709082 43782 709638
rect 43226 692298 43782 692854
rect 43226 656298 43782 656854
rect 43226 620298 43782 620854
rect 43226 584298 43782 584854
rect 43226 548298 43782 548854
rect 43226 512298 43782 512854
rect 43226 476298 43782 476854
rect 43226 440298 43782 440854
rect 43226 404298 43782 404854
rect 43226 368298 43782 368854
rect 43226 332298 43782 332854
rect 43226 296298 43782 296854
rect 43226 260298 43782 260854
rect 43226 224298 43782 224854
rect 43226 188298 43782 188854
rect 43226 152298 43782 152854
rect 43226 116298 43782 116854
rect 43226 80298 43782 80854
rect 43226 44298 43782 44854
rect 43226 8298 43782 8854
rect 43226 -5702 43782 -5146
rect 44466 710042 45022 710598
rect 44466 693538 45022 694094
rect 44466 657538 45022 658094
rect 44466 621538 45022 622094
rect 44466 585538 45022 586094
rect 44466 549538 45022 550094
rect 44466 513538 45022 514094
rect 44466 477538 45022 478094
rect 44466 441538 45022 442094
rect 44466 405538 45022 406094
rect 44466 369538 45022 370094
rect 44466 333538 45022 334094
rect 44466 297538 45022 298094
rect 44466 261538 45022 262094
rect 44466 225538 45022 226094
rect 44466 189538 45022 190094
rect 44466 153538 45022 154094
rect 44466 117538 45022 118094
rect 44466 81538 45022 82094
rect 44466 45538 45022 46094
rect 44466 9538 45022 10094
rect 44466 -6662 45022 -6106
rect 45706 711002 46262 711558
rect 45706 694778 46262 695334
rect 45706 658778 46262 659334
rect 45706 622778 46262 623334
rect 45706 586778 46262 587334
rect 45706 550778 46262 551334
rect 45706 514778 46262 515334
rect 45706 478778 46262 479334
rect 45706 442778 46262 443334
rect 45706 406778 46262 407334
rect 45706 370778 46262 371334
rect 45706 334778 46262 335334
rect 45706 298778 46262 299334
rect 45706 262778 46262 263334
rect 45706 226778 46262 227334
rect 45706 190778 46262 191334
rect 45706 154778 46262 155334
rect 45706 118778 46262 119334
rect 45706 82778 46262 83334
rect 45706 46778 46262 47334
rect 45706 10778 46262 11334
rect 45706 -7622 46262 -7066
rect 73026 704282 73582 704838
rect 73026 686098 73582 686654
rect 73026 650098 73582 650654
rect 73026 614098 73582 614654
rect 73026 578098 73582 578654
rect 73026 542098 73582 542654
rect 73026 506098 73582 506654
rect 73026 470098 73582 470654
rect 73026 434098 73582 434654
rect 73026 398098 73582 398654
rect 73026 362098 73582 362654
rect 73026 326098 73582 326654
rect 73026 290098 73582 290654
rect 73026 254098 73582 254654
rect 73026 218098 73582 218654
rect 73026 182098 73582 182654
rect 73026 146098 73582 146654
rect 73026 110098 73582 110654
rect 73026 74098 73582 74654
rect 73026 38098 73582 38654
rect 73026 2098 73582 2654
rect 73026 -902 73582 -346
rect 74266 705242 74822 705798
rect 74266 687338 74822 687894
rect 74266 651338 74822 651894
rect 74266 615338 74822 615894
rect 74266 579338 74822 579894
rect 74266 543338 74822 543894
rect 74266 507338 74822 507894
rect 74266 471338 74822 471894
rect 74266 435338 74822 435894
rect 74266 399338 74822 399894
rect 74266 363338 74822 363894
rect 74266 327338 74822 327894
rect 74266 291338 74822 291894
rect 74266 255338 74822 255894
rect 74266 219338 74822 219894
rect 74266 183338 74822 183894
rect 74266 147338 74822 147894
rect 74266 111338 74822 111894
rect 74266 75338 74822 75894
rect 74266 39338 74822 39894
rect 74266 3338 74822 3894
rect 74266 -1862 74822 -1306
rect 75506 706202 76062 706758
rect 75506 688578 76062 689134
rect 75506 652578 76062 653134
rect 75506 616578 76062 617134
rect 75506 580578 76062 581134
rect 75506 544578 76062 545134
rect 75506 508578 76062 509134
rect 75506 472578 76062 473134
rect 75506 436578 76062 437134
rect 75506 400578 76062 401134
rect 75506 364578 76062 365134
rect 75506 328578 76062 329134
rect 75506 292578 76062 293134
rect 75506 256578 76062 257134
rect 75506 220578 76062 221134
rect 75506 184578 76062 185134
rect 75506 148578 76062 149134
rect 75506 112578 76062 113134
rect 75506 76578 76062 77134
rect 75506 40578 76062 41134
rect 75506 4578 76062 5134
rect 75506 -2822 76062 -2266
rect 76746 707162 77302 707718
rect 76746 689818 77302 690374
rect 76746 653818 77302 654374
rect 76746 617818 77302 618374
rect 76746 581818 77302 582374
rect 76746 545818 77302 546374
rect 76746 509818 77302 510374
rect 76746 473818 77302 474374
rect 76746 437818 77302 438374
rect 76746 401818 77302 402374
rect 76746 365818 77302 366374
rect 76746 329818 77302 330374
rect 76746 293818 77302 294374
rect 76746 257818 77302 258374
rect 76746 221818 77302 222374
rect 76746 185818 77302 186374
rect 76746 149818 77302 150374
rect 76746 113818 77302 114374
rect 76746 77818 77302 78374
rect 76746 41818 77302 42374
rect 76746 5818 77302 6374
rect 76746 -3782 77302 -3226
rect 77986 708122 78542 708678
rect 77986 691058 78542 691614
rect 77986 655058 78542 655614
rect 77986 619058 78542 619614
rect 77986 583058 78542 583614
rect 77986 547058 78542 547614
rect 77986 511058 78542 511614
rect 77986 475058 78542 475614
rect 77986 439058 78542 439614
rect 77986 403058 78542 403614
rect 77986 367058 78542 367614
rect 77986 331058 78542 331614
rect 77986 295058 78542 295614
rect 77986 259058 78542 259614
rect 77986 223058 78542 223614
rect 77986 187058 78542 187614
rect 77986 151058 78542 151614
rect 77986 115058 78542 115614
rect 77986 79058 78542 79614
rect 77986 43058 78542 43614
rect 77986 7058 78542 7614
rect 77986 -4742 78542 -4186
rect 79226 709082 79782 709638
rect 79226 692298 79782 692854
rect 79226 656298 79782 656854
rect 79226 620298 79782 620854
rect 79226 584298 79782 584854
rect 79226 548298 79782 548854
rect 79226 512298 79782 512854
rect 79226 476298 79782 476854
rect 79226 440298 79782 440854
rect 79226 404298 79782 404854
rect 79226 368298 79782 368854
rect 79226 332298 79782 332854
rect 79226 296298 79782 296854
rect 79226 260298 79782 260854
rect 79226 224298 79782 224854
rect 79226 188298 79782 188854
rect 79226 152298 79782 152854
rect 79226 116298 79782 116854
rect 79226 80298 79782 80854
rect 79226 44298 79782 44854
rect 79226 8298 79782 8854
rect 79226 -5702 79782 -5146
rect 80466 710042 81022 710598
rect 80466 693538 81022 694094
rect 80466 657538 81022 658094
rect 80466 621538 81022 622094
rect 80466 585538 81022 586094
rect 80466 549538 81022 550094
rect 80466 513538 81022 514094
rect 80466 477538 81022 478094
rect 80466 441538 81022 442094
rect 80466 405538 81022 406094
rect 80466 369538 81022 370094
rect 80466 333538 81022 334094
rect 80466 297538 81022 298094
rect 80466 261538 81022 262094
rect 80466 225538 81022 226094
rect 80466 189538 81022 190094
rect 80466 153538 81022 154094
rect 80466 117538 81022 118094
rect 80466 81538 81022 82094
rect 80466 45538 81022 46094
rect 80466 9538 81022 10094
rect 80466 -6662 81022 -6106
rect 81706 711002 82262 711558
rect 81706 694778 82262 695334
rect 81706 658778 82262 659334
rect 81706 622778 82262 623334
rect 81706 586778 82262 587334
rect 81706 550778 82262 551334
rect 81706 514778 82262 515334
rect 81706 478778 82262 479334
rect 81706 442778 82262 443334
rect 81706 406778 82262 407334
rect 81706 370778 82262 371334
rect 81706 334778 82262 335334
rect 81706 298778 82262 299334
rect 81706 262778 82262 263334
rect 81706 226778 82262 227334
rect 81706 190778 82262 191334
rect 81706 154778 82262 155334
rect 81706 118778 82262 119334
rect 81706 82778 82262 83334
rect 81706 46778 82262 47334
rect 81706 10778 82262 11334
rect 81706 -7622 82262 -7066
rect 109026 704282 109582 704838
rect 109026 686098 109582 686654
rect 109026 650098 109582 650654
rect 109026 614098 109582 614654
rect 109026 578098 109582 578654
rect 109026 542098 109582 542654
rect 109026 506098 109582 506654
rect 109026 470098 109582 470654
rect 109026 434098 109582 434654
rect 109026 398098 109582 398654
rect 109026 362098 109582 362654
rect 109026 326098 109582 326654
rect 109026 290098 109582 290654
rect 109026 254098 109582 254654
rect 109026 218098 109582 218654
rect 109026 182098 109582 182654
rect 109026 146098 109582 146654
rect 109026 110098 109582 110654
rect 109026 74098 109582 74654
rect 109026 38098 109582 38654
rect 109026 2098 109582 2654
rect 109026 -902 109582 -346
rect 110266 705242 110822 705798
rect 110266 687338 110822 687894
rect 110266 651338 110822 651894
rect 110266 615338 110822 615894
rect 110266 579338 110822 579894
rect 110266 543338 110822 543894
rect 110266 507338 110822 507894
rect 110266 471338 110822 471894
rect 110266 435338 110822 435894
rect 110266 399338 110822 399894
rect 110266 363338 110822 363894
rect 110266 327338 110822 327894
rect 110266 291338 110822 291894
rect 110266 255338 110822 255894
rect 110266 219338 110822 219894
rect 110266 183338 110822 183894
rect 110266 147338 110822 147894
rect 110266 111338 110822 111894
rect 110266 75338 110822 75894
rect 110266 39338 110822 39894
rect 110266 3338 110822 3894
rect 110266 -1862 110822 -1306
rect 111506 706202 112062 706758
rect 111506 688578 112062 689134
rect 111506 652578 112062 653134
rect 111506 616578 112062 617134
rect 111506 580578 112062 581134
rect 111506 544578 112062 545134
rect 111506 508578 112062 509134
rect 111506 472578 112062 473134
rect 111506 436578 112062 437134
rect 111506 400578 112062 401134
rect 111506 364578 112062 365134
rect 111506 328578 112062 329134
rect 111506 292578 112062 293134
rect 111506 256578 112062 257134
rect 111506 220578 112062 221134
rect 111506 184578 112062 185134
rect 111506 148578 112062 149134
rect 111506 112578 112062 113134
rect 111506 76578 112062 77134
rect 111506 40578 112062 41134
rect 111506 4578 112062 5134
rect 111506 -2822 112062 -2266
rect 112746 707162 113302 707718
rect 112746 689818 113302 690374
rect 112746 653818 113302 654374
rect 112746 617818 113302 618374
rect 112746 581818 113302 582374
rect 112746 545818 113302 546374
rect 112746 509818 113302 510374
rect 112746 473818 113302 474374
rect 112746 437818 113302 438374
rect 112746 401818 113302 402374
rect 112746 365818 113302 366374
rect 112746 329818 113302 330374
rect 112746 293818 113302 294374
rect 112746 257818 113302 258374
rect 112746 221818 113302 222374
rect 112746 185818 113302 186374
rect 112746 149818 113302 150374
rect 112746 113818 113302 114374
rect 112746 77818 113302 78374
rect 112746 41818 113302 42374
rect 112746 5818 113302 6374
rect 112746 -3782 113302 -3226
rect 113986 708122 114542 708678
rect 113986 691058 114542 691614
rect 113986 655058 114542 655614
rect 113986 619058 114542 619614
rect 113986 583058 114542 583614
rect 113986 547058 114542 547614
rect 113986 511058 114542 511614
rect 113986 475058 114542 475614
rect 113986 439058 114542 439614
rect 113986 403058 114542 403614
rect 113986 367058 114542 367614
rect 113986 331058 114542 331614
rect 113986 295058 114542 295614
rect 113986 259058 114542 259614
rect 113986 223058 114542 223614
rect 113986 187058 114542 187614
rect 113986 151058 114542 151614
rect 113986 115058 114542 115614
rect 113986 79058 114542 79614
rect 113986 43058 114542 43614
rect 113986 7058 114542 7614
rect 113986 -4742 114542 -4186
rect 115226 709082 115782 709638
rect 115226 692298 115782 692854
rect 115226 656298 115782 656854
rect 115226 620298 115782 620854
rect 115226 584298 115782 584854
rect 115226 548298 115782 548854
rect 115226 512298 115782 512854
rect 115226 476298 115782 476854
rect 115226 440298 115782 440854
rect 115226 404298 115782 404854
rect 115226 368298 115782 368854
rect 115226 332298 115782 332854
rect 115226 296298 115782 296854
rect 115226 260298 115782 260854
rect 115226 224298 115782 224854
rect 115226 188298 115782 188854
rect 115226 152298 115782 152854
rect 115226 116298 115782 116854
rect 115226 80298 115782 80854
rect 115226 44298 115782 44854
rect 115226 8298 115782 8854
rect 115226 -5702 115782 -5146
rect 116466 710042 117022 710598
rect 116466 693538 117022 694094
rect 116466 657538 117022 658094
rect 116466 621538 117022 622094
rect 116466 585538 117022 586094
rect 116466 549538 117022 550094
rect 116466 513538 117022 514094
rect 116466 477538 117022 478094
rect 116466 441538 117022 442094
rect 116466 405538 117022 406094
rect 116466 369538 117022 370094
rect 116466 333538 117022 334094
rect 116466 297538 117022 298094
rect 116466 261538 117022 262094
rect 116466 225538 117022 226094
rect 116466 189538 117022 190094
rect 116466 153538 117022 154094
rect 116466 117538 117022 118094
rect 116466 81538 117022 82094
rect 116466 45538 117022 46094
rect 116466 9538 117022 10094
rect 116466 -6662 117022 -6106
rect 117706 711002 118262 711558
rect 117706 694778 118262 695334
rect 117706 658778 118262 659334
rect 117706 622778 118262 623334
rect 117706 586778 118262 587334
rect 117706 550778 118262 551334
rect 117706 514778 118262 515334
rect 117706 478778 118262 479334
rect 117706 442778 118262 443334
rect 117706 406778 118262 407334
rect 117706 370778 118262 371334
rect 117706 334778 118262 335334
rect 117706 298778 118262 299334
rect 117706 262778 118262 263334
rect 117706 226778 118262 227334
rect 117706 190778 118262 191334
rect 117706 154778 118262 155334
rect 117706 118778 118262 119334
rect 117706 82778 118262 83334
rect 117706 46778 118262 47334
rect 117706 10778 118262 11334
rect 117706 -7622 118262 -7066
rect 145026 704282 145582 704838
rect 145026 686098 145582 686654
rect 145026 650098 145582 650654
rect 145026 614098 145582 614654
rect 145026 578098 145582 578654
rect 145026 542098 145582 542654
rect 145026 506098 145582 506654
rect 145026 470098 145582 470654
rect 145026 434098 145582 434654
rect 145026 398098 145582 398654
rect 145026 362098 145582 362654
rect 145026 326098 145582 326654
rect 145026 290098 145582 290654
rect 145026 254098 145582 254654
rect 145026 218098 145582 218654
rect 145026 182098 145582 182654
rect 145026 146098 145582 146654
rect 145026 110098 145582 110654
rect 145026 74098 145582 74654
rect 145026 38098 145582 38654
rect 145026 2098 145582 2654
rect 145026 -902 145582 -346
rect 146266 705242 146822 705798
rect 146266 687338 146822 687894
rect 146266 651338 146822 651894
rect 146266 615338 146822 615894
rect 146266 579338 146822 579894
rect 146266 543338 146822 543894
rect 146266 507338 146822 507894
rect 146266 471338 146822 471894
rect 146266 435338 146822 435894
rect 146266 399338 146822 399894
rect 146266 363338 146822 363894
rect 146266 327338 146822 327894
rect 146266 291338 146822 291894
rect 146266 255338 146822 255894
rect 146266 219338 146822 219894
rect 146266 183338 146822 183894
rect 146266 147338 146822 147894
rect 146266 111338 146822 111894
rect 146266 75338 146822 75894
rect 146266 39338 146822 39894
rect 146266 3338 146822 3894
rect 146266 -1862 146822 -1306
rect 147506 706202 148062 706758
rect 147506 688578 148062 689134
rect 147506 652578 148062 653134
rect 147506 616578 148062 617134
rect 147506 580578 148062 581134
rect 147506 544578 148062 545134
rect 147506 508578 148062 509134
rect 147506 472578 148062 473134
rect 147506 436578 148062 437134
rect 147506 400578 148062 401134
rect 147506 364578 148062 365134
rect 147506 328578 148062 329134
rect 147506 292578 148062 293134
rect 147506 256578 148062 257134
rect 147506 220578 148062 221134
rect 147506 184578 148062 185134
rect 147506 148578 148062 149134
rect 147506 112578 148062 113134
rect 147506 76578 148062 77134
rect 147506 40578 148062 41134
rect 147506 4578 148062 5134
rect 147506 -2822 148062 -2266
rect 148746 707162 149302 707718
rect 148746 689818 149302 690374
rect 148746 653818 149302 654374
rect 148746 617818 149302 618374
rect 148746 581818 149302 582374
rect 148746 545818 149302 546374
rect 148746 509818 149302 510374
rect 148746 473818 149302 474374
rect 148746 437818 149302 438374
rect 148746 401818 149302 402374
rect 148746 365818 149302 366374
rect 148746 329818 149302 330374
rect 148746 293818 149302 294374
rect 148746 257818 149302 258374
rect 148746 221818 149302 222374
rect 148746 185818 149302 186374
rect 148746 149818 149302 150374
rect 148746 113818 149302 114374
rect 148746 77818 149302 78374
rect 148746 41818 149302 42374
rect 148746 5818 149302 6374
rect 148746 -3782 149302 -3226
rect 149986 708122 150542 708678
rect 149986 691058 150542 691614
rect 149986 655058 150542 655614
rect 149986 619058 150542 619614
rect 149986 583058 150542 583614
rect 149986 547058 150542 547614
rect 149986 511058 150542 511614
rect 149986 475058 150542 475614
rect 149986 439058 150542 439614
rect 149986 403058 150542 403614
rect 149986 367058 150542 367614
rect 149986 331058 150542 331614
rect 149986 295058 150542 295614
rect 149986 259058 150542 259614
rect 149986 223058 150542 223614
rect 149986 187058 150542 187614
rect 149986 151058 150542 151614
rect 149986 115058 150542 115614
rect 149986 79058 150542 79614
rect 149986 43058 150542 43614
rect 149986 7058 150542 7614
rect 149986 -4742 150542 -4186
rect 151226 709082 151782 709638
rect 151226 692298 151782 692854
rect 151226 656298 151782 656854
rect 151226 620298 151782 620854
rect 151226 584298 151782 584854
rect 151226 548298 151782 548854
rect 151226 512298 151782 512854
rect 151226 476298 151782 476854
rect 151226 440298 151782 440854
rect 151226 404298 151782 404854
rect 151226 368298 151782 368854
rect 151226 332298 151782 332854
rect 151226 296298 151782 296854
rect 151226 260298 151782 260854
rect 151226 224298 151782 224854
rect 151226 188298 151782 188854
rect 151226 152298 151782 152854
rect 151226 116298 151782 116854
rect 151226 80298 151782 80854
rect 151226 44298 151782 44854
rect 151226 8298 151782 8854
rect 151226 -5702 151782 -5146
rect 152466 710042 153022 710598
rect 152466 693538 153022 694094
rect 152466 657538 153022 658094
rect 152466 621538 153022 622094
rect 152466 585538 153022 586094
rect 152466 549538 153022 550094
rect 152466 513538 153022 514094
rect 152466 477538 153022 478094
rect 152466 441538 153022 442094
rect 152466 405538 153022 406094
rect 152466 369538 153022 370094
rect 152466 333538 153022 334094
rect 152466 297538 153022 298094
rect 152466 261538 153022 262094
rect 152466 225538 153022 226094
rect 152466 189538 153022 190094
rect 152466 153538 153022 154094
rect 152466 117538 153022 118094
rect 152466 81538 153022 82094
rect 152466 45538 153022 46094
rect 152466 9538 153022 10094
rect 152466 -6662 153022 -6106
rect 153706 711002 154262 711558
rect 153706 694778 154262 695334
rect 153706 658778 154262 659334
rect 153706 622778 154262 623334
rect 153706 586778 154262 587334
rect 153706 550778 154262 551334
rect 153706 514778 154262 515334
rect 153706 478778 154262 479334
rect 153706 442778 154262 443334
rect 153706 406778 154262 407334
rect 153706 370778 154262 371334
rect 153706 334778 154262 335334
rect 153706 298778 154262 299334
rect 153706 262778 154262 263334
rect 153706 226778 154262 227334
rect 153706 190778 154262 191334
rect 153706 154778 154262 155334
rect 153706 118778 154262 119334
rect 153706 82778 154262 83334
rect 153706 46778 154262 47334
rect 153706 10778 154262 11334
rect 153706 -7622 154262 -7066
rect 181026 704282 181582 704838
rect 181026 686098 181582 686654
rect 181026 650098 181582 650654
rect 181026 614098 181582 614654
rect 181026 578098 181582 578654
rect 181026 542098 181582 542654
rect 181026 506098 181582 506654
rect 181026 470098 181582 470654
rect 181026 434098 181582 434654
rect 181026 398098 181582 398654
rect 181026 362098 181582 362654
rect 181026 326098 181582 326654
rect 181026 290098 181582 290654
rect 181026 254098 181582 254654
rect 181026 218098 181582 218654
rect 181026 182098 181582 182654
rect 181026 146098 181582 146654
rect 181026 110098 181582 110654
rect 181026 74098 181582 74654
rect 181026 38098 181582 38654
rect 181026 2098 181582 2654
rect 181026 -902 181582 -346
rect 182266 705242 182822 705798
rect 182266 687338 182822 687894
rect 182266 651338 182822 651894
rect 182266 615338 182822 615894
rect 182266 579338 182822 579894
rect 182266 543338 182822 543894
rect 182266 507338 182822 507894
rect 182266 471338 182822 471894
rect 182266 435338 182822 435894
rect 182266 399338 182822 399894
rect 182266 363338 182822 363894
rect 182266 327338 182822 327894
rect 182266 291338 182822 291894
rect 182266 255338 182822 255894
rect 182266 219338 182822 219894
rect 182266 183338 182822 183894
rect 182266 147338 182822 147894
rect 182266 111338 182822 111894
rect 182266 75338 182822 75894
rect 182266 39338 182822 39894
rect 182266 3338 182822 3894
rect 182266 -1862 182822 -1306
rect 183506 706202 184062 706758
rect 183506 688578 184062 689134
rect 183506 652578 184062 653134
rect 183506 616578 184062 617134
rect 183506 580578 184062 581134
rect 183506 544578 184062 545134
rect 183506 508578 184062 509134
rect 183506 472578 184062 473134
rect 183506 436578 184062 437134
rect 183506 400578 184062 401134
rect 183506 364578 184062 365134
rect 183506 328578 184062 329134
rect 183506 292578 184062 293134
rect 183506 256578 184062 257134
rect 183506 220578 184062 221134
rect 183506 184578 184062 185134
rect 183506 148578 184062 149134
rect 183506 112578 184062 113134
rect 183506 76578 184062 77134
rect 183506 40578 184062 41134
rect 183506 4578 184062 5134
rect 183506 -2822 184062 -2266
rect 184746 707162 185302 707718
rect 184746 689818 185302 690374
rect 184746 653818 185302 654374
rect 184746 617818 185302 618374
rect 184746 581818 185302 582374
rect 184746 545818 185302 546374
rect 184746 509818 185302 510374
rect 184746 473818 185302 474374
rect 184746 437818 185302 438374
rect 184746 401818 185302 402374
rect 184746 365818 185302 366374
rect 184746 329818 185302 330374
rect 184746 293818 185302 294374
rect 184746 257818 185302 258374
rect 184746 221818 185302 222374
rect 184746 185818 185302 186374
rect 184746 149818 185302 150374
rect 184746 113818 185302 114374
rect 184746 77818 185302 78374
rect 184746 41818 185302 42374
rect 184746 5818 185302 6374
rect 184746 -3782 185302 -3226
rect 185986 708122 186542 708678
rect 185986 691058 186542 691614
rect 185986 655058 186542 655614
rect 185986 619058 186542 619614
rect 185986 583058 186542 583614
rect 185986 547058 186542 547614
rect 185986 511058 186542 511614
rect 185986 475058 186542 475614
rect 185986 439058 186542 439614
rect 185986 403058 186542 403614
rect 185986 367058 186542 367614
rect 185986 331058 186542 331614
rect 185986 295058 186542 295614
rect 185986 259058 186542 259614
rect 185986 223058 186542 223614
rect 185986 187058 186542 187614
rect 185986 151058 186542 151614
rect 185986 115058 186542 115614
rect 185986 79058 186542 79614
rect 185986 43058 186542 43614
rect 185986 7058 186542 7614
rect 185986 -4742 186542 -4186
rect 187226 709082 187782 709638
rect 187226 692298 187782 692854
rect 187226 656298 187782 656854
rect 187226 620298 187782 620854
rect 187226 584298 187782 584854
rect 187226 548298 187782 548854
rect 187226 512298 187782 512854
rect 187226 476298 187782 476854
rect 187226 440298 187782 440854
rect 187226 404298 187782 404854
rect 187226 368298 187782 368854
rect 187226 332298 187782 332854
rect 187226 296298 187782 296854
rect 187226 260298 187782 260854
rect 187226 224298 187782 224854
rect 187226 188298 187782 188854
rect 187226 152298 187782 152854
rect 187226 116298 187782 116854
rect 187226 80298 187782 80854
rect 187226 44298 187782 44854
rect 187226 8298 187782 8854
rect 187226 -5702 187782 -5146
rect 188466 710042 189022 710598
rect 188466 693538 189022 694094
rect 188466 657538 189022 658094
rect 188466 621538 189022 622094
rect 188466 585538 189022 586094
rect 188466 549538 189022 550094
rect 188466 513538 189022 514094
rect 188466 477538 189022 478094
rect 188466 441538 189022 442094
rect 188466 405538 189022 406094
rect 188466 369538 189022 370094
rect 188466 333538 189022 334094
rect 188466 297538 189022 298094
rect 188466 261538 189022 262094
rect 188466 225538 189022 226094
rect 188466 189538 189022 190094
rect 188466 153538 189022 154094
rect 188466 117538 189022 118094
rect 188466 81538 189022 82094
rect 188466 45538 189022 46094
rect 188466 9538 189022 10094
rect 188466 -6662 189022 -6106
rect 189706 711002 190262 711558
rect 189706 694778 190262 695334
rect 189706 658778 190262 659334
rect 189706 622778 190262 623334
rect 189706 586778 190262 587334
rect 189706 550778 190262 551334
rect 189706 514778 190262 515334
rect 189706 478778 190262 479334
rect 189706 442778 190262 443334
rect 189706 406778 190262 407334
rect 189706 370778 190262 371334
rect 189706 334778 190262 335334
rect 189706 298778 190262 299334
rect 189706 262778 190262 263334
rect 189706 226778 190262 227334
rect 189706 190778 190262 191334
rect 189706 154778 190262 155334
rect 189706 118778 190262 119334
rect 189706 82778 190262 83334
rect 189706 46778 190262 47334
rect 189706 10778 190262 11334
rect 189706 -7622 190262 -7066
rect 217026 704282 217582 704838
rect 217026 686098 217582 686654
rect 217026 650098 217582 650654
rect 217026 614098 217582 614654
rect 217026 578098 217582 578654
rect 217026 542098 217582 542654
rect 217026 506098 217582 506654
rect 217026 470098 217582 470654
rect 217026 434098 217582 434654
rect 217026 398098 217582 398654
rect 217026 362098 217582 362654
rect 217026 326098 217582 326654
rect 217026 290098 217582 290654
rect 217026 254098 217582 254654
rect 217026 218098 217582 218654
rect 217026 182098 217582 182654
rect 217026 146098 217582 146654
rect 217026 110098 217582 110654
rect 217026 74098 217582 74654
rect 217026 38098 217582 38654
rect 217026 2098 217582 2654
rect 217026 -902 217582 -346
rect 218266 705242 218822 705798
rect 218266 687338 218822 687894
rect 218266 651338 218822 651894
rect 218266 615338 218822 615894
rect 218266 579338 218822 579894
rect 218266 543338 218822 543894
rect 218266 507338 218822 507894
rect 218266 471338 218822 471894
rect 218266 435338 218822 435894
rect 218266 399338 218822 399894
rect 218266 363338 218822 363894
rect 218266 327338 218822 327894
rect 218266 291338 218822 291894
rect 218266 255338 218822 255894
rect 218266 219338 218822 219894
rect 218266 183338 218822 183894
rect 218266 147338 218822 147894
rect 218266 111338 218822 111894
rect 218266 75338 218822 75894
rect 218266 39338 218822 39894
rect 218266 3338 218822 3894
rect 218266 -1862 218822 -1306
rect 219506 706202 220062 706758
rect 219506 688578 220062 689134
rect 219506 652578 220062 653134
rect 219506 616578 220062 617134
rect 219506 580578 220062 581134
rect 219506 544578 220062 545134
rect 219506 508578 220062 509134
rect 219506 472578 220062 473134
rect 219506 436578 220062 437134
rect 219506 400578 220062 401134
rect 219506 364578 220062 365134
rect 219506 328578 220062 329134
rect 219506 292578 220062 293134
rect 219506 256578 220062 257134
rect 219506 220578 220062 221134
rect 219506 184578 220062 185134
rect 219506 148578 220062 149134
rect 219506 112578 220062 113134
rect 219506 76578 220062 77134
rect 219506 40578 220062 41134
rect 219506 4578 220062 5134
rect 219506 -2822 220062 -2266
rect 220746 707162 221302 707718
rect 220746 689818 221302 690374
rect 220746 653818 221302 654374
rect 220746 617818 221302 618374
rect 220746 581818 221302 582374
rect 220746 545818 221302 546374
rect 220746 509818 221302 510374
rect 220746 473818 221302 474374
rect 220746 437818 221302 438374
rect 220746 401818 221302 402374
rect 220746 365818 221302 366374
rect 220746 329818 221302 330374
rect 220746 293818 221302 294374
rect 220746 257818 221302 258374
rect 220746 221818 221302 222374
rect 220746 185818 221302 186374
rect 220746 149818 221302 150374
rect 220746 113818 221302 114374
rect 220746 77818 221302 78374
rect 220746 41818 221302 42374
rect 220746 5818 221302 6374
rect 220746 -3782 221302 -3226
rect 221986 708122 222542 708678
rect 221986 691058 222542 691614
rect 221986 655058 222542 655614
rect 221986 619058 222542 619614
rect 221986 583058 222542 583614
rect 221986 547058 222542 547614
rect 221986 511058 222542 511614
rect 221986 475058 222542 475614
rect 221986 439058 222542 439614
rect 221986 403058 222542 403614
rect 221986 367058 222542 367614
rect 221986 331058 222542 331614
rect 221986 295058 222542 295614
rect 221986 259058 222542 259614
rect 221986 223058 222542 223614
rect 221986 187058 222542 187614
rect 221986 151058 222542 151614
rect 221986 115058 222542 115614
rect 221986 79058 222542 79614
rect 221986 43058 222542 43614
rect 221986 7058 222542 7614
rect 221986 -4742 222542 -4186
rect 223226 709082 223782 709638
rect 223226 692298 223782 692854
rect 223226 656298 223782 656854
rect 223226 620298 223782 620854
rect 223226 584298 223782 584854
rect 223226 548298 223782 548854
rect 223226 512298 223782 512854
rect 223226 476298 223782 476854
rect 223226 440298 223782 440854
rect 223226 404298 223782 404854
rect 223226 368298 223782 368854
rect 223226 332298 223782 332854
rect 223226 296298 223782 296854
rect 223226 260298 223782 260854
rect 223226 224298 223782 224854
rect 223226 188298 223782 188854
rect 223226 152298 223782 152854
rect 223226 116298 223782 116854
rect 223226 80298 223782 80854
rect 223226 44298 223782 44854
rect 223226 8298 223782 8854
rect 223226 -5702 223782 -5146
rect 224466 710042 225022 710598
rect 224466 693538 225022 694094
rect 224466 657538 225022 658094
rect 224466 621538 225022 622094
rect 224466 585538 225022 586094
rect 224466 549538 225022 550094
rect 224466 513538 225022 514094
rect 224466 477538 225022 478094
rect 224466 441538 225022 442094
rect 224466 405538 225022 406094
rect 224466 369538 225022 370094
rect 224466 333538 225022 334094
rect 224466 297538 225022 298094
rect 224466 261538 225022 262094
rect 224466 225538 225022 226094
rect 224466 189538 225022 190094
rect 224466 153538 225022 154094
rect 224466 117538 225022 118094
rect 224466 81538 225022 82094
rect 224466 45538 225022 46094
rect 224466 9538 225022 10094
rect 224466 -6662 225022 -6106
rect 225706 711002 226262 711558
rect 225706 694778 226262 695334
rect 225706 658778 226262 659334
rect 225706 622778 226262 623334
rect 225706 586778 226262 587334
rect 225706 550778 226262 551334
rect 225706 514778 226262 515334
rect 225706 478778 226262 479334
rect 225706 442778 226262 443334
rect 225706 406778 226262 407334
rect 225706 370778 226262 371334
rect 225706 334778 226262 335334
rect 225706 298778 226262 299334
rect 225706 262778 226262 263334
rect 225706 226778 226262 227334
rect 225706 190778 226262 191334
rect 225706 154778 226262 155334
rect 225706 118778 226262 119334
rect 225706 82778 226262 83334
rect 225706 46778 226262 47334
rect 225706 10778 226262 11334
rect 225706 -7622 226262 -7066
rect 253026 704282 253582 704838
rect 253026 686098 253582 686654
rect 253026 650098 253582 650654
rect 253026 614098 253582 614654
rect 253026 578098 253582 578654
rect 253026 542098 253582 542654
rect 253026 506098 253582 506654
rect 253026 470098 253582 470654
rect 253026 434098 253582 434654
rect 253026 398098 253582 398654
rect 253026 362098 253582 362654
rect 253026 326098 253582 326654
rect 253026 290098 253582 290654
rect 253026 254098 253582 254654
rect 253026 218098 253582 218654
rect 253026 182098 253582 182654
rect 253026 146098 253582 146654
rect 253026 110098 253582 110654
rect 253026 74098 253582 74654
rect 253026 38098 253582 38654
rect 253026 2098 253582 2654
rect 253026 -902 253582 -346
rect 254266 705242 254822 705798
rect 254266 687338 254822 687894
rect 254266 651338 254822 651894
rect 254266 615338 254822 615894
rect 254266 579338 254822 579894
rect 254266 543338 254822 543894
rect 254266 507338 254822 507894
rect 254266 471338 254822 471894
rect 254266 435338 254822 435894
rect 254266 399338 254822 399894
rect 254266 363338 254822 363894
rect 254266 327338 254822 327894
rect 254266 291338 254822 291894
rect 254266 255338 254822 255894
rect 254266 219338 254822 219894
rect 254266 183338 254822 183894
rect 254266 147338 254822 147894
rect 254266 111338 254822 111894
rect 254266 75338 254822 75894
rect 254266 39338 254822 39894
rect 254266 3338 254822 3894
rect 254266 -1862 254822 -1306
rect 255506 706202 256062 706758
rect 255506 688578 256062 689134
rect 255506 652578 256062 653134
rect 255506 616578 256062 617134
rect 255506 580578 256062 581134
rect 255506 544578 256062 545134
rect 255506 508578 256062 509134
rect 255506 472578 256062 473134
rect 255506 436578 256062 437134
rect 255506 400578 256062 401134
rect 255506 364578 256062 365134
rect 255506 328578 256062 329134
rect 255506 292578 256062 293134
rect 255506 256578 256062 257134
rect 255506 220578 256062 221134
rect 255506 184578 256062 185134
rect 255506 148578 256062 149134
rect 255506 112578 256062 113134
rect 255506 76578 256062 77134
rect 255506 40578 256062 41134
rect 255506 4578 256062 5134
rect 255506 -2822 256062 -2266
rect 256746 707162 257302 707718
rect 256746 689818 257302 690374
rect 256746 653818 257302 654374
rect 256746 617818 257302 618374
rect 256746 581818 257302 582374
rect 256746 545818 257302 546374
rect 256746 509818 257302 510374
rect 256746 473818 257302 474374
rect 256746 437818 257302 438374
rect 256746 401818 257302 402374
rect 256746 365818 257302 366374
rect 256746 329818 257302 330374
rect 256746 293818 257302 294374
rect 256746 257818 257302 258374
rect 256746 221818 257302 222374
rect 256746 185818 257302 186374
rect 256746 149818 257302 150374
rect 256746 113818 257302 114374
rect 256746 77818 257302 78374
rect 256746 41818 257302 42374
rect 256746 5818 257302 6374
rect 256746 -3782 257302 -3226
rect 257986 708122 258542 708678
rect 257986 691058 258542 691614
rect 257986 655058 258542 655614
rect 257986 619058 258542 619614
rect 257986 583058 258542 583614
rect 257986 547058 258542 547614
rect 257986 511058 258542 511614
rect 257986 475058 258542 475614
rect 257986 439058 258542 439614
rect 257986 403058 258542 403614
rect 257986 367058 258542 367614
rect 257986 331058 258542 331614
rect 257986 295058 258542 295614
rect 257986 259058 258542 259614
rect 257986 223058 258542 223614
rect 257986 187058 258542 187614
rect 257986 151058 258542 151614
rect 257986 115058 258542 115614
rect 257986 79058 258542 79614
rect 257986 43058 258542 43614
rect 257986 7058 258542 7614
rect 257986 -4742 258542 -4186
rect 259226 709082 259782 709638
rect 259226 692298 259782 692854
rect 259226 656298 259782 656854
rect 259226 620298 259782 620854
rect 259226 584298 259782 584854
rect 259226 548298 259782 548854
rect 259226 512298 259782 512854
rect 259226 476298 259782 476854
rect 259226 440298 259782 440854
rect 259226 404298 259782 404854
rect 259226 368298 259782 368854
rect 259226 332298 259782 332854
rect 259226 296298 259782 296854
rect 259226 260298 259782 260854
rect 259226 224298 259782 224854
rect 259226 188298 259782 188854
rect 259226 152298 259782 152854
rect 259226 116298 259782 116854
rect 259226 80298 259782 80854
rect 259226 44298 259782 44854
rect 259226 8298 259782 8854
rect 259226 -5702 259782 -5146
rect 260466 710042 261022 710598
rect 260466 693538 261022 694094
rect 260466 657538 261022 658094
rect 260466 621538 261022 622094
rect 260466 585538 261022 586094
rect 260466 549538 261022 550094
rect 260466 513538 261022 514094
rect 260466 477538 261022 478094
rect 260466 441538 261022 442094
rect 260466 405538 261022 406094
rect 260466 369538 261022 370094
rect 260466 333538 261022 334094
rect 260466 297538 261022 298094
rect 260466 261538 261022 262094
rect 260466 225538 261022 226094
rect 260466 189538 261022 190094
rect 260466 153538 261022 154094
rect 260466 117538 261022 118094
rect 260466 81538 261022 82094
rect 260466 45538 261022 46094
rect 260466 9538 261022 10094
rect 260466 -6662 261022 -6106
rect 261706 711002 262262 711558
rect 261706 694778 262262 695334
rect 261706 658778 262262 659334
rect 261706 622778 262262 623334
rect 261706 586778 262262 587334
rect 261706 550778 262262 551334
rect 261706 514778 262262 515334
rect 261706 478778 262262 479334
rect 261706 442778 262262 443334
rect 261706 406778 262262 407334
rect 261706 370778 262262 371334
rect 261706 334778 262262 335334
rect 261706 298778 262262 299334
rect 261706 262778 262262 263334
rect 261706 226778 262262 227334
rect 261706 190778 262262 191334
rect 261706 154778 262262 155334
rect 261706 118778 262262 119334
rect 261706 82778 262262 83334
rect 261706 46778 262262 47334
rect 261706 10778 262262 11334
rect 261706 -7622 262262 -7066
rect 289026 704282 289582 704838
rect 289026 686098 289582 686654
rect 289026 650098 289582 650654
rect 289026 614098 289582 614654
rect 289026 578098 289582 578654
rect 289026 542098 289582 542654
rect 289026 506098 289582 506654
rect 289026 470098 289582 470654
rect 289026 434098 289582 434654
rect 289026 398098 289582 398654
rect 289026 362098 289582 362654
rect 289026 326098 289582 326654
rect 289026 290098 289582 290654
rect 289026 254098 289582 254654
rect 289026 218098 289582 218654
rect 289026 182098 289582 182654
rect 289026 146098 289582 146654
rect 289026 110098 289582 110654
rect 289026 74098 289582 74654
rect 289026 38098 289582 38654
rect 289026 2098 289582 2654
rect 289026 -902 289582 -346
rect 290266 705242 290822 705798
rect 290266 687338 290822 687894
rect 290266 651338 290822 651894
rect 290266 615338 290822 615894
rect 290266 579338 290822 579894
rect 290266 543338 290822 543894
rect 290266 507338 290822 507894
rect 290266 471338 290822 471894
rect 290266 435338 290822 435894
rect 290266 399338 290822 399894
rect 290266 363338 290822 363894
rect 290266 327338 290822 327894
rect 290266 291338 290822 291894
rect 290266 255338 290822 255894
rect 290266 219338 290822 219894
rect 290266 183338 290822 183894
rect 290266 147338 290822 147894
rect 290266 111338 290822 111894
rect 290266 75338 290822 75894
rect 290266 39338 290822 39894
rect 290266 3338 290822 3894
rect 290266 -1862 290822 -1306
rect 291506 706202 292062 706758
rect 291506 688578 292062 689134
rect 291506 652578 292062 653134
rect 291506 616578 292062 617134
rect 291506 580578 292062 581134
rect 291506 544578 292062 545134
rect 291506 508578 292062 509134
rect 291506 472578 292062 473134
rect 291506 436578 292062 437134
rect 291506 400578 292062 401134
rect 291506 364578 292062 365134
rect 291506 328578 292062 329134
rect 291506 292578 292062 293134
rect 291506 256578 292062 257134
rect 291506 220578 292062 221134
rect 291506 184578 292062 185134
rect 291506 148578 292062 149134
rect 291506 112578 292062 113134
rect 291506 76578 292062 77134
rect 291506 40578 292062 41134
rect 291506 4578 292062 5134
rect 291506 -2822 292062 -2266
rect 292746 707162 293302 707718
rect 292746 689818 293302 690374
rect 292746 653818 293302 654374
rect 292746 617818 293302 618374
rect 292746 581818 293302 582374
rect 292746 545818 293302 546374
rect 292746 509818 293302 510374
rect 292746 473818 293302 474374
rect 292746 437818 293302 438374
rect 292746 401818 293302 402374
rect 292746 365818 293302 366374
rect 292746 329818 293302 330374
rect 292746 293818 293302 294374
rect 292746 257818 293302 258374
rect 292746 221818 293302 222374
rect 292746 185818 293302 186374
rect 292746 149818 293302 150374
rect 292746 113818 293302 114374
rect 292746 77818 293302 78374
rect 292746 41818 293302 42374
rect 292746 5818 293302 6374
rect 292746 -3782 293302 -3226
rect 293986 708122 294542 708678
rect 293986 691058 294542 691614
rect 293986 655058 294542 655614
rect 293986 619058 294542 619614
rect 293986 583058 294542 583614
rect 293986 547058 294542 547614
rect 293986 511058 294542 511614
rect 293986 475058 294542 475614
rect 293986 439058 294542 439614
rect 293986 403058 294542 403614
rect 293986 367058 294542 367614
rect 293986 331058 294542 331614
rect 293986 295058 294542 295614
rect 293986 259058 294542 259614
rect 293986 223058 294542 223614
rect 293986 187058 294542 187614
rect 293986 151058 294542 151614
rect 293986 115058 294542 115614
rect 293986 79058 294542 79614
rect 293986 43058 294542 43614
rect 293986 7058 294542 7614
rect 293986 -4742 294542 -4186
rect 295226 709082 295782 709638
rect 295226 692298 295782 692854
rect 295226 656298 295782 656854
rect 295226 620298 295782 620854
rect 295226 584298 295782 584854
rect 295226 548298 295782 548854
rect 295226 512298 295782 512854
rect 295226 476298 295782 476854
rect 295226 440298 295782 440854
rect 295226 404298 295782 404854
rect 295226 368298 295782 368854
rect 295226 332298 295782 332854
rect 295226 296298 295782 296854
rect 295226 260298 295782 260854
rect 295226 224298 295782 224854
rect 295226 188298 295782 188854
rect 295226 152298 295782 152854
rect 295226 116298 295782 116854
rect 295226 80298 295782 80854
rect 295226 44298 295782 44854
rect 295226 8298 295782 8854
rect 295226 -5702 295782 -5146
rect 296466 710042 297022 710598
rect 296466 693538 297022 694094
rect 296466 657538 297022 658094
rect 296466 621538 297022 622094
rect 296466 585538 297022 586094
rect 296466 549538 297022 550094
rect 296466 513538 297022 514094
rect 296466 477538 297022 478094
rect 296466 441538 297022 442094
rect 296466 405538 297022 406094
rect 296466 369538 297022 370094
rect 296466 333538 297022 334094
rect 296466 297538 297022 298094
rect 296466 261538 297022 262094
rect 296466 225538 297022 226094
rect 296466 189538 297022 190094
rect 296466 153538 297022 154094
rect 296466 117538 297022 118094
rect 296466 81538 297022 82094
rect 296466 45538 297022 46094
rect 296466 9538 297022 10094
rect 296466 -6662 297022 -6106
rect 297706 711002 298262 711558
rect 297706 694778 298262 695334
rect 297706 658778 298262 659334
rect 297706 622778 298262 623334
rect 297706 586778 298262 587334
rect 297706 550778 298262 551334
rect 297706 514778 298262 515334
rect 297706 478778 298262 479334
rect 297706 442778 298262 443334
rect 297706 406778 298262 407334
rect 297706 370778 298262 371334
rect 297706 334778 298262 335334
rect 297706 298778 298262 299334
rect 297706 262778 298262 263334
rect 297706 226778 298262 227334
rect 297706 190778 298262 191334
rect 297706 154778 298262 155334
rect 297706 118778 298262 119334
rect 297706 82778 298262 83334
rect 297706 46778 298262 47334
rect 297706 10778 298262 11334
rect 297706 -7622 298262 -7066
rect 325026 704282 325582 704838
rect 325026 686098 325582 686654
rect 325026 650098 325582 650654
rect 325026 614098 325582 614654
rect 325026 578098 325582 578654
rect 325026 542098 325582 542654
rect 325026 506098 325582 506654
rect 325026 470098 325582 470654
rect 325026 434098 325582 434654
rect 325026 398098 325582 398654
rect 325026 362098 325582 362654
rect 325026 326098 325582 326654
rect 325026 290098 325582 290654
rect 325026 254098 325582 254654
rect 325026 218098 325582 218654
rect 325026 182098 325582 182654
rect 325026 146098 325582 146654
rect 325026 110098 325582 110654
rect 325026 74098 325582 74654
rect 325026 38098 325582 38654
rect 325026 2098 325582 2654
rect 325026 -902 325582 -346
rect 326266 705242 326822 705798
rect 326266 687338 326822 687894
rect 326266 651338 326822 651894
rect 326266 615338 326822 615894
rect 326266 579338 326822 579894
rect 326266 543338 326822 543894
rect 326266 507338 326822 507894
rect 326266 471338 326822 471894
rect 326266 435338 326822 435894
rect 326266 399338 326822 399894
rect 326266 363338 326822 363894
rect 326266 327338 326822 327894
rect 326266 291338 326822 291894
rect 326266 255338 326822 255894
rect 326266 219338 326822 219894
rect 326266 183338 326822 183894
rect 326266 147338 326822 147894
rect 326266 111338 326822 111894
rect 326266 75338 326822 75894
rect 326266 39338 326822 39894
rect 326266 3338 326822 3894
rect 326266 -1862 326822 -1306
rect 327506 706202 328062 706758
rect 327506 688578 328062 689134
rect 327506 652578 328062 653134
rect 327506 616578 328062 617134
rect 327506 580578 328062 581134
rect 327506 544578 328062 545134
rect 327506 508578 328062 509134
rect 327506 472578 328062 473134
rect 327506 436578 328062 437134
rect 327506 400578 328062 401134
rect 327506 364578 328062 365134
rect 327506 328578 328062 329134
rect 327506 292578 328062 293134
rect 327506 256578 328062 257134
rect 327506 220578 328062 221134
rect 327506 184578 328062 185134
rect 327506 148578 328062 149134
rect 327506 112578 328062 113134
rect 327506 76578 328062 77134
rect 327506 40578 328062 41134
rect 327506 4578 328062 5134
rect 327506 -2822 328062 -2266
rect 328746 707162 329302 707718
rect 328746 689818 329302 690374
rect 328746 653818 329302 654374
rect 328746 617818 329302 618374
rect 328746 581818 329302 582374
rect 328746 545818 329302 546374
rect 328746 509818 329302 510374
rect 328746 473818 329302 474374
rect 328746 437818 329302 438374
rect 328746 401818 329302 402374
rect 328746 365818 329302 366374
rect 328746 329818 329302 330374
rect 328746 293818 329302 294374
rect 328746 257818 329302 258374
rect 328746 221818 329302 222374
rect 328746 185818 329302 186374
rect 328746 149818 329302 150374
rect 328746 113818 329302 114374
rect 328746 77818 329302 78374
rect 328746 41818 329302 42374
rect 328746 5818 329302 6374
rect 328746 -3782 329302 -3226
rect 329986 708122 330542 708678
rect 329986 691058 330542 691614
rect 329986 655058 330542 655614
rect 329986 619058 330542 619614
rect 329986 583058 330542 583614
rect 329986 547058 330542 547614
rect 329986 511058 330542 511614
rect 329986 475058 330542 475614
rect 329986 439058 330542 439614
rect 329986 403058 330542 403614
rect 329986 367058 330542 367614
rect 329986 331058 330542 331614
rect 329986 295058 330542 295614
rect 329986 259058 330542 259614
rect 329986 223058 330542 223614
rect 329986 187058 330542 187614
rect 329986 151058 330542 151614
rect 329986 115058 330542 115614
rect 329986 79058 330542 79614
rect 329986 43058 330542 43614
rect 329986 7058 330542 7614
rect 329986 -4742 330542 -4186
rect 331226 709082 331782 709638
rect 331226 692298 331782 692854
rect 331226 656298 331782 656854
rect 331226 620298 331782 620854
rect 331226 584298 331782 584854
rect 331226 548298 331782 548854
rect 331226 512298 331782 512854
rect 331226 476298 331782 476854
rect 331226 440298 331782 440854
rect 331226 404298 331782 404854
rect 331226 368298 331782 368854
rect 331226 332298 331782 332854
rect 331226 296298 331782 296854
rect 331226 260298 331782 260854
rect 331226 224298 331782 224854
rect 331226 188298 331782 188854
rect 331226 152298 331782 152854
rect 331226 116298 331782 116854
rect 331226 80298 331782 80854
rect 331226 44298 331782 44854
rect 331226 8298 331782 8854
rect 331226 -5702 331782 -5146
rect 332466 710042 333022 710598
rect 332466 693538 333022 694094
rect 332466 657538 333022 658094
rect 332466 621538 333022 622094
rect 332466 585538 333022 586094
rect 332466 549538 333022 550094
rect 332466 513538 333022 514094
rect 332466 477538 333022 478094
rect 332466 441538 333022 442094
rect 332466 405538 333022 406094
rect 332466 369538 333022 370094
rect 332466 333538 333022 334094
rect 332466 297538 333022 298094
rect 332466 261538 333022 262094
rect 332466 225538 333022 226094
rect 332466 189538 333022 190094
rect 332466 153538 333022 154094
rect 332466 117538 333022 118094
rect 332466 81538 333022 82094
rect 332466 45538 333022 46094
rect 332466 9538 333022 10094
rect 332466 -6662 333022 -6106
rect 333706 711002 334262 711558
rect 333706 694778 334262 695334
rect 333706 658778 334262 659334
rect 333706 622778 334262 623334
rect 333706 586778 334262 587334
rect 333706 550778 334262 551334
rect 333706 514778 334262 515334
rect 333706 478778 334262 479334
rect 333706 442778 334262 443334
rect 333706 406778 334262 407334
rect 333706 370778 334262 371334
rect 333706 334778 334262 335334
rect 333706 298778 334262 299334
rect 333706 262778 334262 263334
rect 333706 226778 334262 227334
rect 333706 190778 334262 191334
rect 333706 154778 334262 155334
rect 333706 118778 334262 119334
rect 333706 82778 334262 83334
rect 333706 46778 334262 47334
rect 333706 10778 334262 11334
rect 333706 -7622 334262 -7066
rect 361026 704282 361582 704838
rect 361026 686098 361582 686654
rect 361026 650098 361582 650654
rect 361026 614098 361582 614654
rect 361026 578098 361582 578654
rect 361026 542098 361582 542654
rect 361026 506098 361582 506654
rect 361026 470098 361582 470654
rect 361026 434098 361582 434654
rect 361026 398098 361582 398654
rect 361026 362098 361582 362654
rect 361026 326098 361582 326654
rect 361026 290098 361582 290654
rect 361026 254098 361582 254654
rect 361026 218098 361582 218654
rect 361026 182098 361582 182654
rect 361026 146098 361582 146654
rect 361026 110098 361582 110654
rect 361026 74098 361582 74654
rect 361026 38098 361582 38654
rect 361026 2098 361582 2654
rect 361026 -902 361582 -346
rect 362266 705242 362822 705798
rect 362266 687338 362822 687894
rect 362266 651338 362822 651894
rect 362266 615338 362822 615894
rect 362266 579338 362822 579894
rect 362266 543338 362822 543894
rect 362266 507338 362822 507894
rect 362266 471338 362822 471894
rect 362266 435338 362822 435894
rect 362266 399338 362822 399894
rect 362266 363338 362822 363894
rect 362266 327338 362822 327894
rect 362266 291338 362822 291894
rect 362266 255338 362822 255894
rect 362266 219338 362822 219894
rect 362266 183338 362822 183894
rect 362266 147338 362822 147894
rect 362266 111338 362822 111894
rect 362266 75338 362822 75894
rect 362266 39338 362822 39894
rect 362266 3338 362822 3894
rect 362266 -1862 362822 -1306
rect 363506 706202 364062 706758
rect 363506 688578 364062 689134
rect 363506 652578 364062 653134
rect 363506 616578 364062 617134
rect 363506 580578 364062 581134
rect 363506 544578 364062 545134
rect 363506 508578 364062 509134
rect 363506 472578 364062 473134
rect 363506 436578 364062 437134
rect 363506 400578 364062 401134
rect 363506 364578 364062 365134
rect 363506 328578 364062 329134
rect 363506 292578 364062 293134
rect 363506 256578 364062 257134
rect 363506 220578 364062 221134
rect 363506 184578 364062 185134
rect 363506 148578 364062 149134
rect 363506 112578 364062 113134
rect 363506 76578 364062 77134
rect 363506 40578 364062 41134
rect 363506 4578 364062 5134
rect 363506 -2822 364062 -2266
rect 364746 707162 365302 707718
rect 364746 689818 365302 690374
rect 364746 653818 365302 654374
rect 364746 617818 365302 618374
rect 364746 581818 365302 582374
rect 364746 545818 365302 546374
rect 364746 509818 365302 510374
rect 364746 473818 365302 474374
rect 364746 437818 365302 438374
rect 364746 401818 365302 402374
rect 364746 365818 365302 366374
rect 364746 329818 365302 330374
rect 364746 293818 365302 294374
rect 364746 257818 365302 258374
rect 364746 221818 365302 222374
rect 364746 185818 365302 186374
rect 364746 149818 365302 150374
rect 364746 113818 365302 114374
rect 364746 77818 365302 78374
rect 364746 41818 365302 42374
rect 364746 5818 365302 6374
rect 364746 -3782 365302 -3226
rect 365986 708122 366542 708678
rect 365986 691058 366542 691614
rect 365986 655058 366542 655614
rect 365986 619058 366542 619614
rect 365986 583058 366542 583614
rect 365986 547058 366542 547614
rect 365986 511058 366542 511614
rect 365986 475058 366542 475614
rect 365986 439058 366542 439614
rect 365986 403058 366542 403614
rect 365986 367058 366542 367614
rect 365986 331058 366542 331614
rect 365986 295058 366542 295614
rect 365986 259058 366542 259614
rect 365986 223058 366542 223614
rect 365986 187058 366542 187614
rect 365986 151058 366542 151614
rect 365986 115058 366542 115614
rect 365986 79058 366542 79614
rect 365986 43058 366542 43614
rect 365986 7058 366542 7614
rect 365986 -4742 366542 -4186
rect 367226 709082 367782 709638
rect 367226 692298 367782 692854
rect 367226 656298 367782 656854
rect 367226 620298 367782 620854
rect 367226 584298 367782 584854
rect 367226 548298 367782 548854
rect 367226 512298 367782 512854
rect 367226 476298 367782 476854
rect 367226 440298 367782 440854
rect 367226 404298 367782 404854
rect 367226 368298 367782 368854
rect 367226 332298 367782 332854
rect 367226 296298 367782 296854
rect 367226 260298 367782 260854
rect 367226 224298 367782 224854
rect 367226 188298 367782 188854
rect 367226 152298 367782 152854
rect 367226 116298 367782 116854
rect 367226 80298 367782 80854
rect 367226 44298 367782 44854
rect 367226 8298 367782 8854
rect 367226 -5702 367782 -5146
rect 368466 710042 369022 710598
rect 368466 693538 369022 694094
rect 368466 657538 369022 658094
rect 368466 621538 369022 622094
rect 368466 585538 369022 586094
rect 368466 549538 369022 550094
rect 368466 513538 369022 514094
rect 368466 477538 369022 478094
rect 368466 441538 369022 442094
rect 368466 405538 369022 406094
rect 368466 369538 369022 370094
rect 368466 333538 369022 334094
rect 368466 297538 369022 298094
rect 368466 261538 369022 262094
rect 368466 225538 369022 226094
rect 368466 189538 369022 190094
rect 368466 153538 369022 154094
rect 368466 117538 369022 118094
rect 368466 81538 369022 82094
rect 368466 45538 369022 46094
rect 368466 9538 369022 10094
rect 368466 -6662 369022 -6106
rect 369706 711002 370262 711558
rect 369706 694778 370262 695334
rect 369706 658778 370262 659334
rect 369706 622778 370262 623334
rect 369706 586778 370262 587334
rect 369706 550778 370262 551334
rect 369706 514778 370262 515334
rect 369706 478778 370262 479334
rect 369706 442778 370262 443334
rect 369706 406778 370262 407334
rect 369706 370778 370262 371334
rect 369706 334778 370262 335334
rect 369706 298778 370262 299334
rect 369706 262778 370262 263334
rect 369706 226778 370262 227334
rect 369706 190778 370262 191334
rect 369706 154778 370262 155334
rect 369706 118778 370262 119334
rect 369706 82778 370262 83334
rect 369706 46778 370262 47334
rect 369706 10778 370262 11334
rect 369706 -7622 370262 -7066
rect 397026 704282 397582 704838
rect 397026 686098 397582 686654
rect 397026 650098 397582 650654
rect 397026 614098 397582 614654
rect 397026 578098 397582 578654
rect 397026 542098 397582 542654
rect 397026 506098 397582 506654
rect 397026 470098 397582 470654
rect 397026 434098 397582 434654
rect 397026 398098 397582 398654
rect 397026 362098 397582 362654
rect 397026 326098 397582 326654
rect 397026 290098 397582 290654
rect 397026 254098 397582 254654
rect 397026 218098 397582 218654
rect 397026 182098 397582 182654
rect 397026 146098 397582 146654
rect 397026 110098 397582 110654
rect 397026 74098 397582 74654
rect 397026 38098 397582 38654
rect 397026 2098 397582 2654
rect 397026 -902 397582 -346
rect 398266 705242 398822 705798
rect 398266 687338 398822 687894
rect 398266 651338 398822 651894
rect 398266 615338 398822 615894
rect 398266 579338 398822 579894
rect 398266 543338 398822 543894
rect 398266 507338 398822 507894
rect 398266 471338 398822 471894
rect 398266 435338 398822 435894
rect 398266 399338 398822 399894
rect 398266 363338 398822 363894
rect 398266 327338 398822 327894
rect 398266 291338 398822 291894
rect 398266 255338 398822 255894
rect 398266 219338 398822 219894
rect 398266 183338 398822 183894
rect 398266 147338 398822 147894
rect 398266 111338 398822 111894
rect 398266 75338 398822 75894
rect 398266 39338 398822 39894
rect 398266 3338 398822 3894
rect 398266 -1862 398822 -1306
rect 399506 706202 400062 706758
rect 399506 688578 400062 689134
rect 399506 652578 400062 653134
rect 399506 616578 400062 617134
rect 399506 580578 400062 581134
rect 399506 544578 400062 545134
rect 399506 508578 400062 509134
rect 399506 472578 400062 473134
rect 399506 436578 400062 437134
rect 399506 400578 400062 401134
rect 399506 364578 400062 365134
rect 399506 328578 400062 329134
rect 399506 292578 400062 293134
rect 399506 256578 400062 257134
rect 399506 220578 400062 221134
rect 399506 184578 400062 185134
rect 399506 148578 400062 149134
rect 399506 112578 400062 113134
rect 399506 76578 400062 77134
rect 399506 40578 400062 41134
rect 399506 4578 400062 5134
rect 399506 -2822 400062 -2266
rect 400746 707162 401302 707718
rect 400746 689818 401302 690374
rect 400746 653818 401302 654374
rect 400746 617818 401302 618374
rect 400746 581818 401302 582374
rect 400746 545818 401302 546374
rect 400746 509818 401302 510374
rect 400746 473818 401302 474374
rect 400746 437818 401302 438374
rect 400746 401818 401302 402374
rect 400746 365818 401302 366374
rect 400746 329818 401302 330374
rect 400746 293818 401302 294374
rect 400746 257818 401302 258374
rect 400746 221818 401302 222374
rect 400746 185818 401302 186374
rect 400746 149818 401302 150374
rect 400746 113818 401302 114374
rect 400746 77818 401302 78374
rect 400746 41818 401302 42374
rect 400746 5818 401302 6374
rect 400746 -3782 401302 -3226
rect 401986 708122 402542 708678
rect 401986 691058 402542 691614
rect 401986 655058 402542 655614
rect 401986 619058 402542 619614
rect 401986 583058 402542 583614
rect 401986 547058 402542 547614
rect 401986 511058 402542 511614
rect 401986 475058 402542 475614
rect 401986 439058 402542 439614
rect 401986 403058 402542 403614
rect 401986 367058 402542 367614
rect 401986 331058 402542 331614
rect 401986 295058 402542 295614
rect 401986 259058 402542 259614
rect 401986 223058 402542 223614
rect 401986 187058 402542 187614
rect 401986 151058 402542 151614
rect 401986 115058 402542 115614
rect 401986 79058 402542 79614
rect 401986 43058 402542 43614
rect 401986 7058 402542 7614
rect 401986 -4742 402542 -4186
rect 403226 709082 403782 709638
rect 403226 692298 403782 692854
rect 403226 656298 403782 656854
rect 403226 620298 403782 620854
rect 403226 584298 403782 584854
rect 403226 548298 403782 548854
rect 403226 512298 403782 512854
rect 403226 476298 403782 476854
rect 403226 440298 403782 440854
rect 403226 404298 403782 404854
rect 403226 368298 403782 368854
rect 403226 332298 403782 332854
rect 403226 296298 403782 296854
rect 403226 260298 403782 260854
rect 403226 224298 403782 224854
rect 403226 188298 403782 188854
rect 403226 152298 403782 152854
rect 403226 116298 403782 116854
rect 403226 80298 403782 80854
rect 403226 44298 403782 44854
rect 403226 8298 403782 8854
rect 403226 -5702 403782 -5146
rect 404466 710042 405022 710598
rect 404466 693538 405022 694094
rect 404466 657538 405022 658094
rect 404466 621538 405022 622094
rect 404466 585538 405022 586094
rect 404466 549538 405022 550094
rect 404466 513538 405022 514094
rect 404466 477538 405022 478094
rect 404466 441538 405022 442094
rect 404466 405538 405022 406094
rect 404466 369538 405022 370094
rect 404466 333538 405022 334094
rect 404466 297538 405022 298094
rect 404466 261538 405022 262094
rect 404466 225538 405022 226094
rect 404466 189538 405022 190094
rect 404466 153538 405022 154094
rect 404466 117538 405022 118094
rect 404466 81538 405022 82094
rect 404466 45538 405022 46094
rect 404466 9538 405022 10094
rect 404466 -6662 405022 -6106
rect 405706 711002 406262 711558
rect 405706 694778 406262 695334
rect 405706 658778 406262 659334
rect 405706 622778 406262 623334
rect 405706 586778 406262 587334
rect 405706 550778 406262 551334
rect 405706 514778 406262 515334
rect 405706 478778 406262 479334
rect 405706 442778 406262 443334
rect 405706 406778 406262 407334
rect 405706 370778 406262 371334
rect 405706 334778 406262 335334
rect 405706 298778 406262 299334
rect 405706 262778 406262 263334
rect 405706 226778 406262 227334
rect 405706 190778 406262 191334
rect 405706 154778 406262 155334
rect 405706 118778 406262 119334
rect 405706 82778 406262 83334
rect 405706 46778 406262 47334
rect 405706 10778 406262 11334
rect 405706 -7622 406262 -7066
rect 433026 704282 433582 704838
rect 433026 686098 433582 686654
rect 433026 650098 433582 650654
rect 433026 614098 433582 614654
rect 433026 578098 433582 578654
rect 433026 542098 433582 542654
rect 433026 506098 433582 506654
rect 433026 470098 433582 470654
rect 433026 434098 433582 434654
rect 433026 398098 433582 398654
rect 433026 362098 433582 362654
rect 433026 326098 433582 326654
rect 433026 290098 433582 290654
rect 433026 254098 433582 254654
rect 433026 218098 433582 218654
rect 433026 182098 433582 182654
rect 433026 146098 433582 146654
rect 433026 110098 433582 110654
rect 433026 74098 433582 74654
rect 433026 38098 433582 38654
rect 433026 2098 433582 2654
rect 433026 -902 433582 -346
rect 434266 705242 434822 705798
rect 434266 687338 434822 687894
rect 434266 651338 434822 651894
rect 434266 615338 434822 615894
rect 434266 579338 434822 579894
rect 434266 543338 434822 543894
rect 434266 507338 434822 507894
rect 434266 471338 434822 471894
rect 434266 435338 434822 435894
rect 434266 399338 434822 399894
rect 434266 363338 434822 363894
rect 434266 327338 434822 327894
rect 434266 291338 434822 291894
rect 434266 255338 434822 255894
rect 434266 219338 434822 219894
rect 434266 183338 434822 183894
rect 434266 147338 434822 147894
rect 434266 111338 434822 111894
rect 434266 75338 434822 75894
rect 434266 39338 434822 39894
rect 434266 3338 434822 3894
rect 434266 -1862 434822 -1306
rect 435506 706202 436062 706758
rect 435506 688578 436062 689134
rect 435506 652578 436062 653134
rect 435506 616578 436062 617134
rect 435506 580578 436062 581134
rect 435506 544578 436062 545134
rect 435506 508578 436062 509134
rect 435506 472578 436062 473134
rect 435506 436578 436062 437134
rect 435506 400578 436062 401134
rect 435506 364578 436062 365134
rect 435506 328578 436062 329134
rect 435506 292578 436062 293134
rect 435506 256578 436062 257134
rect 435506 220578 436062 221134
rect 435506 184578 436062 185134
rect 435506 148578 436062 149134
rect 435506 112578 436062 113134
rect 435506 76578 436062 77134
rect 435506 40578 436062 41134
rect 435506 4578 436062 5134
rect 435506 -2822 436062 -2266
rect 436746 707162 437302 707718
rect 436746 689818 437302 690374
rect 436746 653818 437302 654374
rect 436746 617818 437302 618374
rect 436746 581818 437302 582374
rect 436746 545818 437302 546374
rect 436746 509818 437302 510374
rect 436746 473818 437302 474374
rect 436746 437818 437302 438374
rect 436746 401818 437302 402374
rect 436746 365818 437302 366374
rect 436746 329818 437302 330374
rect 436746 293818 437302 294374
rect 436746 257818 437302 258374
rect 436746 221818 437302 222374
rect 436746 185818 437302 186374
rect 436746 149818 437302 150374
rect 436746 113818 437302 114374
rect 436746 77818 437302 78374
rect 436746 41818 437302 42374
rect 436746 5818 437302 6374
rect 436746 -3782 437302 -3226
rect 437986 708122 438542 708678
rect 437986 691058 438542 691614
rect 437986 655058 438542 655614
rect 437986 619058 438542 619614
rect 437986 583058 438542 583614
rect 437986 547058 438542 547614
rect 437986 511058 438542 511614
rect 437986 475058 438542 475614
rect 437986 439058 438542 439614
rect 437986 403058 438542 403614
rect 437986 367058 438542 367614
rect 437986 331058 438542 331614
rect 437986 295058 438542 295614
rect 437986 259058 438542 259614
rect 437986 223058 438542 223614
rect 437986 187058 438542 187614
rect 437986 151058 438542 151614
rect 437986 115058 438542 115614
rect 437986 79058 438542 79614
rect 437986 43058 438542 43614
rect 437986 7058 438542 7614
rect 437986 -4742 438542 -4186
rect 439226 709082 439782 709638
rect 439226 692298 439782 692854
rect 439226 656298 439782 656854
rect 439226 620298 439782 620854
rect 439226 584298 439782 584854
rect 439226 548298 439782 548854
rect 439226 512298 439782 512854
rect 439226 476298 439782 476854
rect 439226 440298 439782 440854
rect 439226 404298 439782 404854
rect 439226 368298 439782 368854
rect 439226 332298 439782 332854
rect 439226 296298 439782 296854
rect 439226 260298 439782 260854
rect 439226 224298 439782 224854
rect 439226 188298 439782 188854
rect 439226 152298 439782 152854
rect 439226 116298 439782 116854
rect 439226 80298 439782 80854
rect 439226 44298 439782 44854
rect 439226 8298 439782 8854
rect 439226 -5702 439782 -5146
rect 440466 710042 441022 710598
rect 440466 693538 441022 694094
rect 440466 657538 441022 658094
rect 440466 621538 441022 622094
rect 440466 585538 441022 586094
rect 440466 549538 441022 550094
rect 440466 513538 441022 514094
rect 440466 477538 441022 478094
rect 440466 441538 441022 442094
rect 440466 405538 441022 406094
rect 440466 369538 441022 370094
rect 440466 333538 441022 334094
rect 440466 297538 441022 298094
rect 440466 261538 441022 262094
rect 440466 225538 441022 226094
rect 440466 189538 441022 190094
rect 440466 153538 441022 154094
rect 440466 117538 441022 118094
rect 440466 81538 441022 82094
rect 440466 45538 441022 46094
rect 440466 9538 441022 10094
rect 440466 -6662 441022 -6106
rect 441706 711002 442262 711558
rect 441706 694778 442262 695334
rect 441706 658778 442262 659334
rect 441706 622778 442262 623334
rect 441706 586778 442262 587334
rect 441706 550778 442262 551334
rect 441706 514778 442262 515334
rect 441706 478778 442262 479334
rect 441706 442778 442262 443334
rect 441706 406778 442262 407334
rect 441706 370778 442262 371334
rect 441706 334778 442262 335334
rect 441706 298778 442262 299334
rect 441706 262778 442262 263334
rect 441706 226778 442262 227334
rect 441706 190778 442262 191334
rect 441706 154778 442262 155334
rect 441706 118778 442262 119334
rect 441706 82778 442262 83334
rect 441706 46778 442262 47334
rect 441706 10778 442262 11334
rect 441706 -7622 442262 -7066
rect 469026 704282 469582 704838
rect 469026 686098 469582 686654
rect 469026 650098 469582 650654
rect 469026 614098 469582 614654
rect 469026 578098 469582 578654
rect 469026 542098 469582 542654
rect 469026 506098 469582 506654
rect 469026 470098 469582 470654
rect 469026 434098 469582 434654
rect 469026 398098 469582 398654
rect 469026 362098 469582 362654
rect 469026 326098 469582 326654
rect 469026 290098 469582 290654
rect 469026 254098 469582 254654
rect 469026 218098 469582 218654
rect 469026 182098 469582 182654
rect 469026 146098 469582 146654
rect 469026 110098 469582 110654
rect 469026 74098 469582 74654
rect 469026 38098 469582 38654
rect 469026 2098 469582 2654
rect 469026 -902 469582 -346
rect 470266 705242 470822 705798
rect 470266 687338 470822 687894
rect 470266 651338 470822 651894
rect 470266 615338 470822 615894
rect 470266 579338 470822 579894
rect 470266 543338 470822 543894
rect 470266 507338 470822 507894
rect 470266 471338 470822 471894
rect 470266 435338 470822 435894
rect 470266 399338 470822 399894
rect 470266 363338 470822 363894
rect 470266 327338 470822 327894
rect 470266 291338 470822 291894
rect 470266 255338 470822 255894
rect 470266 219338 470822 219894
rect 470266 183338 470822 183894
rect 470266 147338 470822 147894
rect 470266 111338 470822 111894
rect 470266 75338 470822 75894
rect 470266 39338 470822 39894
rect 470266 3338 470822 3894
rect 470266 -1862 470822 -1306
rect 471506 706202 472062 706758
rect 471506 688578 472062 689134
rect 471506 652578 472062 653134
rect 471506 616578 472062 617134
rect 471506 580578 472062 581134
rect 471506 544578 472062 545134
rect 471506 508578 472062 509134
rect 471506 472578 472062 473134
rect 471506 436578 472062 437134
rect 471506 400578 472062 401134
rect 471506 364578 472062 365134
rect 472746 707162 473302 707718
rect 472746 689818 473302 690374
rect 472746 653818 473302 654374
rect 472746 617818 473302 618374
rect 472746 581818 473302 582374
rect 472746 545818 473302 546374
rect 472746 509818 473302 510374
rect 472746 473818 473302 474374
rect 473986 708122 474542 708678
rect 473986 691058 474542 691614
rect 473986 655058 474542 655614
rect 473986 619058 474542 619614
rect 473986 583058 474542 583614
rect 473986 547058 474542 547614
rect 473986 511058 474542 511614
rect 473986 475058 474542 475614
rect 472746 437818 473302 438374
rect 473986 439058 474542 439614
rect 472746 401818 473302 402374
rect 473986 403058 474542 403614
rect 472746 365818 473302 366374
rect 475226 709082 475782 709638
rect 475226 692298 475782 692854
rect 475226 656298 475782 656854
rect 475226 620298 475782 620854
rect 475226 584298 475782 584854
rect 475226 548298 475782 548854
rect 475226 512298 475782 512854
rect 475226 476298 475782 476854
rect 475226 440298 475782 440854
rect 475226 404298 475782 404854
rect 473986 367058 474542 367614
rect 475226 368298 475782 368854
rect 476466 710042 477022 710598
rect 476466 693538 477022 694094
rect 476466 657538 477022 658094
rect 476466 621538 477022 622094
rect 476466 585538 477022 586094
rect 476466 549538 477022 550094
rect 476466 513538 477022 514094
rect 476466 477538 477022 478094
rect 476466 441538 477022 442094
rect 476466 405538 477022 406094
rect 476466 369538 477022 370094
rect 477706 711002 478262 711558
rect 477706 694778 478262 695334
rect 477706 658778 478262 659334
rect 477706 622778 478262 623334
rect 477706 586778 478262 587334
rect 477706 550778 478262 551334
rect 477706 514778 478262 515334
rect 477706 478778 478262 479334
rect 505026 704282 505582 704838
rect 505026 686098 505582 686654
rect 505026 650098 505582 650654
rect 505026 614098 505582 614654
rect 505026 578098 505582 578654
rect 505026 542098 505582 542654
rect 505026 506098 505582 506654
rect 505026 470098 505582 470654
rect 477706 442778 478262 443334
rect 477706 406778 478262 407334
rect 505026 434098 505582 434654
rect 477706 370778 478262 371334
rect 471506 328578 472062 329134
rect 471506 292578 472062 293134
rect 472746 329818 473302 330374
rect 473986 331058 474542 331614
rect 472746 293818 473302 294374
rect 473986 295058 474542 295614
rect 475226 332298 475782 332854
rect 475226 296298 475782 296854
rect 476466 333538 477022 334094
rect 476466 297538 477022 298094
rect 477706 334778 478262 335334
rect 505026 398098 505582 398654
rect 505026 362098 505582 362654
rect 477706 298778 478262 299334
rect 505026 326098 505582 326654
rect 505026 290098 505582 290654
rect 471506 256578 472062 257134
rect 471506 220578 472062 221134
rect 471506 184578 472062 185134
rect 471506 148578 472062 149134
rect 471506 112578 472062 113134
rect 471506 76578 472062 77134
rect 471506 40578 472062 41134
rect 471506 4578 472062 5134
rect 471506 -2822 472062 -2266
rect 472746 257818 473302 258374
rect 472746 221818 473302 222374
rect 472746 185818 473302 186374
rect 472746 149818 473302 150374
rect 472746 113818 473302 114374
rect 472746 77818 473302 78374
rect 472746 41818 473302 42374
rect 472746 5818 473302 6374
rect 472746 -3782 473302 -3226
rect 473986 259058 474542 259614
rect 473986 223058 474542 223614
rect 473986 187058 474542 187614
rect 473986 151058 474542 151614
rect 473986 115058 474542 115614
rect 473986 79058 474542 79614
rect 473986 43058 474542 43614
rect 473986 7058 474542 7614
rect 473986 -4742 474542 -4186
rect 475226 260298 475782 260854
rect 475226 224298 475782 224854
rect 475226 188298 475782 188854
rect 475226 152298 475782 152854
rect 475226 116298 475782 116854
rect 475226 80298 475782 80854
rect 475226 44298 475782 44854
rect 475226 8298 475782 8854
rect 475226 -5702 475782 -5146
rect 476466 261538 477022 262094
rect 476466 225538 477022 226094
rect 476466 189538 477022 190094
rect 476466 153538 477022 154094
rect 476466 117538 477022 118094
rect 476466 81538 477022 82094
rect 476466 45538 477022 46094
rect 476466 9538 477022 10094
rect 477706 262778 478262 263334
rect 477706 226778 478262 227334
rect 477706 190778 478262 191334
rect 477706 154778 478262 155334
rect 477706 118778 478262 119334
rect 477706 82778 478262 83334
rect 477706 46778 478262 47334
rect 505026 254098 505582 254654
rect 505026 218098 505582 218654
rect 505026 182098 505582 182654
rect 505026 146098 505582 146654
rect 505026 110098 505582 110654
rect 505026 74098 505582 74654
rect 477706 10778 478262 11334
rect 476466 -6662 477022 -6106
rect 477706 -7622 478262 -7066
rect 505026 38098 505582 38654
rect 505026 2098 505582 2654
rect 505026 -902 505582 -346
rect 506266 705242 506822 705798
rect 506266 687338 506822 687894
rect 506266 651338 506822 651894
rect 506266 615338 506822 615894
rect 506266 579338 506822 579894
rect 506266 543338 506822 543894
rect 506266 507338 506822 507894
rect 506266 471338 506822 471894
rect 506266 435338 506822 435894
rect 506266 399338 506822 399894
rect 506266 363338 506822 363894
rect 506266 327338 506822 327894
rect 506266 291338 506822 291894
rect 506266 255338 506822 255894
rect 506266 219338 506822 219894
rect 506266 183338 506822 183894
rect 506266 147338 506822 147894
rect 506266 111338 506822 111894
rect 506266 75338 506822 75894
rect 506266 39338 506822 39894
rect 506266 3338 506822 3894
rect 506266 -1862 506822 -1306
rect 507506 706202 508062 706758
rect 507506 688578 508062 689134
rect 507506 652578 508062 653134
rect 507506 616578 508062 617134
rect 507506 580578 508062 581134
rect 507506 544578 508062 545134
rect 507506 508578 508062 509134
rect 507506 472578 508062 473134
rect 507506 436578 508062 437134
rect 507506 400578 508062 401134
rect 507506 364578 508062 365134
rect 507506 328578 508062 329134
rect 507506 292578 508062 293134
rect 507506 256578 508062 257134
rect 507506 220578 508062 221134
rect 507506 184578 508062 185134
rect 507506 148578 508062 149134
rect 507506 112578 508062 113134
rect 507506 76578 508062 77134
rect 507506 40578 508062 41134
rect 507506 4578 508062 5134
rect 507506 -2822 508062 -2266
rect 508746 707162 509302 707718
rect 508746 689818 509302 690374
rect 508746 653818 509302 654374
rect 508746 617818 509302 618374
rect 508746 581818 509302 582374
rect 508746 545818 509302 546374
rect 508746 509818 509302 510374
rect 508746 473818 509302 474374
rect 508746 437818 509302 438374
rect 508746 401818 509302 402374
rect 508746 365818 509302 366374
rect 508746 329818 509302 330374
rect 508746 293818 509302 294374
rect 508746 257818 509302 258374
rect 508746 221818 509302 222374
rect 508746 185818 509302 186374
rect 508746 149818 509302 150374
rect 508746 113818 509302 114374
rect 508746 77818 509302 78374
rect 508746 41818 509302 42374
rect 508746 5818 509302 6374
rect 508746 -3782 509302 -3226
rect 509986 708122 510542 708678
rect 509986 691058 510542 691614
rect 509986 655058 510542 655614
rect 509986 619058 510542 619614
rect 509986 583058 510542 583614
rect 509986 547058 510542 547614
rect 509986 511058 510542 511614
rect 509986 475058 510542 475614
rect 509986 439058 510542 439614
rect 509986 403058 510542 403614
rect 509986 367058 510542 367614
rect 509986 331058 510542 331614
rect 509986 295058 510542 295614
rect 509986 259058 510542 259614
rect 509986 223058 510542 223614
rect 509986 187058 510542 187614
rect 509986 151058 510542 151614
rect 509986 115058 510542 115614
rect 509986 79058 510542 79614
rect 509986 43058 510542 43614
rect 509986 7058 510542 7614
rect 509986 -4742 510542 -4186
rect 511226 709082 511782 709638
rect 511226 692298 511782 692854
rect 511226 656298 511782 656854
rect 511226 620298 511782 620854
rect 511226 584298 511782 584854
rect 511226 548298 511782 548854
rect 511226 512298 511782 512854
rect 511226 476298 511782 476854
rect 511226 440298 511782 440854
rect 511226 404298 511782 404854
rect 511226 368298 511782 368854
rect 511226 332298 511782 332854
rect 511226 296298 511782 296854
rect 511226 260298 511782 260854
rect 511226 224298 511782 224854
rect 511226 188298 511782 188854
rect 511226 152298 511782 152854
rect 511226 116298 511782 116854
rect 511226 80298 511782 80854
rect 511226 44298 511782 44854
rect 511226 8298 511782 8854
rect 511226 -5702 511782 -5146
rect 512466 710042 513022 710598
rect 512466 693538 513022 694094
rect 512466 657538 513022 658094
rect 512466 621538 513022 622094
rect 512466 585538 513022 586094
rect 512466 549538 513022 550094
rect 512466 513538 513022 514094
rect 512466 477538 513022 478094
rect 512466 441538 513022 442094
rect 512466 405538 513022 406094
rect 512466 369538 513022 370094
rect 512466 333538 513022 334094
rect 512466 297538 513022 298094
rect 512466 261538 513022 262094
rect 512466 225538 513022 226094
rect 512466 189538 513022 190094
rect 512466 153538 513022 154094
rect 512466 117538 513022 118094
rect 512466 81538 513022 82094
rect 512466 45538 513022 46094
rect 512466 9538 513022 10094
rect 512466 -6662 513022 -6106
rect 513706 711002 514262 711558
rect 513706 694778 514262 695334
rect 513706 658778 514262 659334
rect 513706 622778 514262 623334
rect 513706 586778 514262 587334
rect 513706 550778 514262 551334
rect 513706 514778 514262 515334
rect 513706 478778 514262 479334
rect 541026 704282 541582 704838
rect 541026 686098 541582 686654
rect 541026 650098 541582 650654
rect 541026 614098 541582 614654
rect 541026 578098 541582 578654
rect 541026 542098 541582 542654
rect 541026 506098 541582 506654
rect 541026 470098 541582 470654
rect 542266 705242 542822 705798
rect 542266 687338 542822 687894
rect 542266 651338 542822 651894
rect 542266 615338 542822 615894
rect 542266 579338 542822 579894
rect 542266 543338 542822 543894
rect 542266 507338 542822 507894
rect 542266 471338 542822 471894
rect 543506 706202 544062 706758
rect 543506 688578 544062 689134
rect 543506 652578 544062 653134
rect 543506 616578 544062 617134
rect 543506 580578 544062 581134
rect 543506 544578 544062 545134
rect 543506 508578 544062 509134
rect 543506 472578 544062 473134
rect 544746 707162 545302 707718
rect 544746 689818 545302 690374
rect 544746 653818 545302 654374
rect 544746 617818 545302 618374
rect 544746 581818 545302 582374
rect 544746 545818 545302 546374
rect 544746 509818 545302 510374
rect 544746 473818 545302 474374
rect 545986 708122 546542 708678
rect 545986 691058 546542 691614
rect 545986 655058 546542 655614
rect 545986 619058 546542 619614
rect 545986 583058 546542 583614
rect 545986 547058 546542 547614
rect 545986 511058 546542 511614
rect 545986 475058 546542 475614
rect 547226 709082 547782 709638
rect 547226 692298 547782 692854
rect 547226 656298 547782 656854
rect 547226 620298 547782 620854
rect 547226 584298 547782 584854
rect 547226 548298 547782 548854
rect 547226 512298 547782 512854
rect 547226 476298 547782 476854
rect 513706 442778 514262 443334
rect 540918 435658 541154 435894
rect 540918 435338 541154 435574
rect 539952 434418 540188 434654
rect 539952 434098 540188 434334
rect 542850 435658 543086 435894
rect 542850 435338 543086 435574
rect 541884 434418 542120 434654
rect 541884 434098 542120 434334
rect 543816 434418 544052 434654
rect 543816 434098 544052 434334
rect 547226 440298 547782 440854
rect 544782 435658 545018 435894
rect 544782 435338 545018 435574
rect 546714 435658 546950 435894
rect 546714 435338 546950 435574
rect 545748 434418 545984 434654
rect 545748 434098 545984 434334
rect 513706 406778 514262 407334
rect 540918 399658 541154 399894
rect 540918 399338 541154 399574
rect 539952 398418 540188 398654
rect 539952 398098 540188 398334
rect 542850 399658 543086 399894
rect 542850 399338 543086 399574
rect 541884 398418 542120 398654
rect 541884 398098 542120 398334
rect 543816 398418 544052 398654
rect 543816 398098 544052 398334
rect 547226 404298 547782 404854
rect 544782 399658 545018 399894
rect 544782 399338 545018 399574
rect 546714 399658 546950 399894
rect 546714 399338 546950 399574
rect 545748 398418 545984 398654
rect 545748 398098 545984 398334
rect 513706 370778 514262 371334
rect 540918 363658 541154 363894
rect 540918 363338 541154 363574
rect 539952 362418 540188 362654
rect 539952 362098 540188 362334
rect 542850 363658 543086 363894
rect 542850 363338 543086 363574
rect 541884 362418 542120 362654
rect 541884 362098 542120 362334
rect 543816 362418 544052 362654
rect 543816 362098 544052 362334
rect 547226 368298 547782 368854
rect 544782 363658 545018 363894
rect 544782 363338 545018 363574
rect 546714 363658 546950 363894
rect 546714 363338 546950 363574
rect 545748 362418 545984 362654
rect 545748 362098 545984 362334
rect 513706 334778 514262 335334
rect 540918 327658 541154 327894
rect 540918 327338 541154 327574
rect 539952 326418 540188 326654
rect 539952 326098 540188 326334
rect 542850 327658 543086 327894
rect 542850 327338 543086 327574
rect 541884 326418 542120 326654
rect 541884 326098 542120 326334
rect 543816 326418 544052 326654
rect 543816 326098 544052 326334
rect 547226 332298 547782 332854
rect 544782 327658 545018 327894
rect 544782 327338 545018 327574
rect 546714 327658 546950 327894
rect 546714 327338 546950 327574
rect 545748 326418 545984 326654
rect 545748 326098 545984 326334
rect 513706 298778 514262 299334
rect 547226 296298 547782 296854
rect 540918 291658 541154 291894
rect 540918 291338 541154 291574
rect 542850 291658 543086 291894
rect 542850 291338 543086 291574
rect 544782 291658 545018 291894
rect 544782 291338 545018 291574
rect 546714 291658 546950 291894
rect 546714 291338 546950 291574
rect 539952 290418 540188 290654
rect 539952 290098 540188 290334
rect 541884 290418 542120 290654
rect 541884 290098 542120 290334
rect 543816 290418 544052 290654
rect 543816 290098 544052 290334
rect 545748 290418 545984 290654
rect 545748 290098 545984 290334
rect 513706 262778 514262 263334
rect 513706 226778 514262 227334
rect 513706 190778 514262 191334
rect 513706 154778 514262 155334
rect 513706 118778 514262 119334
rect 513706 82778 514262 83334
rect 513706 46778 514262 47334
rect 513706 10778 514262 11334
rect 513706 -7622 514262 -7066
rect 541026 254098 541582 254654
rect 541026 218098 541582 218654
rect 541026 182098 541582 182654
rect 541026 146098 541582 146654
rect 541026 110098 541582 110654
rect 541026 74098 541582 74654
rect 541026 38098 541582 38654
rect 541026 2098 541582 2654
rect 541026 -902 541582 -346
rect 542266 255338 542822 255894
rect 542266 219338 542822 219894
rect 542266 183338 542822 183894
rect 542266 147338 542822 147894
rect 542266 111338 542822 111894
rect 542266 75338 542822 75894
rect 542266 39338 542822 39894
rect 542266 3338 542822 3894
rect 542266 -1862 542822 -1306
rect 543506 256578 544062 257134
rect 543506 220578 544062 221134
rect 543506 184578 544062 185134
rect 543506 148578 544062 149134
rect 543506 112578 544062 113134
rect 543506 76578 544062 77134
rect 543506 40578 544062 41134
rect 543506 4578 544062 5134
rect 543506 -2822 544062 -2266
rect 544746 257818 545302 258374
rect 544746 221818 545302 222374
rect 544746 185818 545302 186374
rect 544746 149818 545302 150374
rect 544746 113818 545302 114374
rect 544746 77818 545302 78374
rect 544746 41818 545302 42374
rect 544746 5818 545302 6374
rect 544746 -3782 545302 -3226
rect 545986 259058 546542 259614
rect 545986 223058 546542 223614
rect 545986 187058 546542 187614
rect 545986 151058 546542 151614
rect 545986 115058 546542 115614
rect 545986 79058 546542 79614
rect 545986 43058 546542 43614
rect 545986 7058 546542 7614
rect 545986 -4742 546542 -4186
rect 547226 260298 547782 260854
rect 547226 224298 547782 224854
rect 547226 188298 547782 188854
rect 547226 152298 547782 152854
rect 547226 116298 547782 116854
rect 547226 80298 547782 80854
rect 547226 44298 547782 44854
rect 547226 8298 547782 8854
rect 547226 -5702 547782 -5146
rect 548466 710042 549022 710598
rect 548466 693538 549022 694094
rect 548466 657538 549022 658094
rect 548466 621538 549022 622094
rect 548466 585538 549022 586094
rect 548466 549538 549022 550094
rect 548466 513538 549022 514094
rect 548466 477538 549022 478094
rect 548466 441538 549022 442094
rect 549706 711002 550262 711558
rect 549706 694778 550262 695334
rect 549706 658778 550262 659334
rect 549706 622778 550262 623334
rect 549706 586778 550262 587334
rect 549706 550778 550262 551334
rect 549706 514778 550262 515334
rect 549706 478778 550262 479334
rect 549706 442778 550262 443334
rect 548466 405538 549022 406094
rect 549706 406778 550262 407334
rect 548466 369538 549022 370094
rect 549706 370778 550262 371334
rect 548466 333538 549022 334094
rect 549706 334778 550262 335334
rect 548466 297538 549022 298094
rect 549706 298778 550262 299334
rect 548466 261538 549022 262094
rect 548466 225538 549022 226094
rect 548466 189538 549022 190094
rect 548466 153538 549022 154094
rect 548466 117538 549022 118094
rect 548466 81538 549022 82094
rect 548466 45538 549022 46094
rect 549706 262778 550262 263334
rect 549706 226778 550262 227334
rect 549706 190778 550262 191334
rect 549706 154778 550262 155334
rect 549706 118778 550262 119334
rect 549706 82778 550262 83334
rect 549706 46778 550262 47334
rect 548466 9538 549022 10094
rect 548466 -6662 549022 -6106
rect 549706 10778 550262 11334
rect 549706 -7622 550262 -7066
rect 577026 704282 577582 704838
rect 577026 686098 577582 686654
rect 577026 650098 577582 650654
rect 577026 614098 577582 614654
rect 577026 578098 577582 578654
rect 577026 542098 577582 542654
rect 577026 506098 577582 506654
rect 577026 470098 577582 470654
rect 577026 434098 577582 434654
rect 577026 398098 577582 398654
rect 577026 362098 577582 362654
rect 577026 326098 577582 326654
rect 577026 290098 577582 290654
rect 577026 254098 577582 254654
rect 577026 218098 577582 218654
rect 577026 182098 577582 182654
rect 577026 146098 577582 146654
rect 577026 110098 577582 110654
rect 577026 74098 577582 74654
rect 577026 38098 577582 38654
rect 577026 2098 577582 2654
rect 577026 -902 577582 -346
rect 578266 705242 578822 705798
rect 578266 687338 578822 687894
rect 578266 651338 578822 651894
rect 578266 615338 578822 615894
rect 578266 579338 578822 579894
rect 578266 543338 578822 543894
rect 578266 507338 578822 507894
rect 578266 471338 578822 471894
rect 578266 435338 578822 435894
rect 578266 399338 578822 399894
rect 578266 363338 578822 363894
rect 578266 327338 578822 327894
rect 578266 291338 578822 291894
rect 578266 255338 578822 255894
rect 578266 219338 578822 219894
rect 578266 183338 578822 183894
rect 578266 147338 578822 147894
rect 578266 111338 578822 111894
rect 578266 75338 578822 75894
rect 578266 39338 578822 39894
rect 578266 3338 578822 3894
rect 578266 -1862 578822 -1306
rect 579506 706202 580062 706758
rect 579506 688578 580062 689134
rect 579506 652578 580062 653134
rect 579506 616578 580062 617134
rect 579506 580578 580062 581134
rect 579506 544578 580062 545134
rect 579506 508578 580062 509134
rect 579506 472578 580062 473134
rect 579506 436578 580062 437134
rect 579506 400578 580062 401134
rect 579506 364578 580062 365134
rect 579506 328578 580062 329134
rect 579506 292578 580062 293134
rect 579506 256578 580062 257134
rect 579506 220578 580062 221134
rect 579506 184578 580062 185134
rect 579506 148578 580062 149134
rect 579506 112578 580062 113134
rect 579506 76578 580062 77134
rect 579506 40578 580062 41134
rect 579506 4578 580062 5134
rect 579506 -2822 580062 -2266
rect 580746 707162 581302 707718
rect 580746 689818 581302 690374
rect 580746 653818 581302 654374
rect 580746 617818 581302 618374
rect 580746 581818 581302 582374
rect 580746 545818 581302 546374
rect 580746 509818 581302 510374
rect 580746 473818 581302 474374
rect 580746 437818 581302 438374
rect 580746 401818 581302 402374
rect 580746 365818 581302 366374
rect 580746 329818 581302 330374
rect 580746 293818 581302 294374
rect 580746 257818 581302 258374
rect 580746 221818 581302 222374
rect 580746 185818 581302 186374
rect 580746 149818 581302 150374
rect 580746 113818 581302 114374
rect 580746 77818 581302 78374
rect 580746 41818 581302 42374
rect 580746 5818 581302 6374
rect 580746 -3782 581302 -3226
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 581986 708122 582542 708678
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581986 691058 582542 691614
rect 581986 655058 582542 655614
rect 581986 619058 582542 619614
rect 581986 583058 582542 583614
rect 581986 547058 582542 547614
rect 581986 511058 582542 511614
rect 581986 475058 582542 475614
rect 581986 439058 582542 439614
rect 581986 403058 582542 403614
rect 581986 367058 582542 367614
rect 581986 331058 582542 331614
rect 581986 295058 582542 295614
rect 581986 259058 582542 259614
rect 581986 223058 582542 223614
rect 581986 187058 582542 187614
rect 581986 151058 582542 151614
rect 581986 115058 582542 115614
rect 581986 79058 582542 79614
rect 581986 43058 582542 43614
rect 581986 7058 582542 7614
rect 585342 704282 585898 704838
rect 585342 686098 585898 686654
rect 585342 650098 585898 650654
rect 585342 614098 585898 614654
rect 585342 578098 585898 578654
rect 585342 542098 585898 542654
rect 585342 506098 585898 506654
rect 585342 470098 585898 470654
rect 585342 434098 585898 434654
rect 585342 398098 585898 398654
rect 585342 362098 585898 362654
rect 585342 326098 585898 326654
rect 585342 290098 585898 290654
rect 585342 254098 585898 254654
rect 585342 218098 585898 218654
rect 585342 182098 585898 182654
rect 585342 146098 585898 146654
rect 585342 110098 585898 110654
rect 585342 74098 585898 74654
rect 585342 38098 585898 38654
rect 585342 2098 585898 2654
rect 585342 -902 585898 -346
rect 586302 687338 586858 687894
rect 586302 651338 586858 651894
rect 586302 615338 586858 615894
rect 586302 579338 586858 579894
rect 586302 543338 586858 543894
rect 586302 507338 586858 507894
rect 586302 471338 586858 471894
rect 586302 435338 586858 435894
rect 586302 399338 586858 399894
rect 586302 363338 586858 363894
rect 586302 327338 586858 327894
rect 586302 291338 586858 291894
rect 586302 255338 586858 255894
rect 586302 219338 586858 219894
rect 586302 183338 586858 183894
rect 586302 147338 586858 147894
rect 586302 111338 586858 111894
rect 586302 75338 586858 75894
rect 586302 39338 586858 39894
rect 586302 3338 586858 3894
rect 586302 -1862 586858 -1306
rect 587262 688578 587818 689134
rect 587262 652578 587818 653134
rect 587262 616578 587818 617134
rect 587262 580578 587818 581134
rect 587262 544578 587818 545134
rect 587262 508578 587818 509134
rect 587262 472578 587818 473134
rect 587262 436578 587818 437134
rect 587262 400578 587818 401134
rect 587262 364578 587818 365134
rect 587262 328578 587818 329134
rect 587262 292578 587818 293134
rect 587262 256578 587818 257134
rect 587262 220578 587818 221134
rect 587262 184578 587818 185134
rect 587262 148578 587818 149134
rect 587262 112578 587818 113134
rect 587262 76578 587818 77134
rect 587262 40578 587818 41134
rect 587262 4578 587818 5134
rect 587262 -2822 587818 -2266
rect 588222 689818 588778 690374
rect 588222 653818 588778 654374
rect 588222 617818 588778 618374
rect 588222 581818 588778 582374
rect 588222 545818 588778 546374
rect 588222 509818 588778 510374
rect 588222 473818 588778 474374
rect 588222 437818 588778 438374
rect 588222 401818 588778 402374
rect 588222 365818 588778 366374
rect 588222 329818 588778 330374
rect 588222 293818 588778 294374
rect 588222 257818 588778 258374
rect 588222 221818 588778 222374
rect 588222 185818 588778 186374
rect 588222 149818 588778 150374
rect 588222 113818 588778 114374
rect 588222 77818 588778 78374
rect 588222 41818 588778 42374
rect 588222 5818 588778 6374
rect 588222 -3782 588778 -3226
rect 589182 691058 589738 691614
rect 589182 655058 589738 655614
rect 589182 619058 589738 619614
rect 589182 583058 589738 583614
rect 589182 547058 589738 547614
rect 589182 511058 589738 511614
rect 589182 475058 589738 475614
rect 589182 439058 589738 439614
rect 589182 403058 589738 403614
rect 589182 367058 589738 367614
rect 589182 331058 589738 331614
rect 589182 295058 589738 295614
rect 589182 259058 589738 259614
rect 589182 223058 589738 223614
rect 589182 187058 589738 187614
rect 589182 151058 589738 151614
rect 589182 115058 589738 115614
rect 589182 79058 589738 79614
rect 589182 43058 589738 43614
rect 589182 7058 589738 7614
rect 581986 -4742 582542 -4186
rect 589182 -4742 589738 -4186
rect 590142 692298 590698 692854
rect 590142 656298 590698 656854
rect 590142 620298 590698 620854
rect 590142 584298 590698 584854
rect 590142 548298 590698 548854
rect 590142 512298 590698 512854
rect 590142 476298 590698 476854
rect 590142 440298 590698 440854
rect 590142 404298 590698 404854
rect 590142 368298 590698 368854
rect 590142 332298 590698 332854
rect 590142 296298 590698 296854
rect 590142 260298 590698 260854
rect 590142 224298 590698 224854
rect 590142 188298 590698 188854
rect 590142 152298 590698 152854
rect 590142 116298 590698 116854
rect 590142 80298 590698 80854
rect 590142 44298 590698 44854
rect 590142 8298 590698 8854
rect 590142 -5702 590698 -5146
rect 591102 693538 591658 694094
rect 591102 657538 591658 658094
rect 591102 621538 591658 622094
rect 591102 585538 591658 586094
rect 591102 549538 591658 550094
rect 591102 513538 591658 514094
rect 591102 477538 591658 478094
rect 591102 441538 591658 442094
rect 591102 405538 591658 406094
rect 591102 369538 591658 370094
rect 591102 333538 591658 334094
rect 591102 297538 591658 298094
rect 591102 261538 591658 262094
rect 591102 225538 591658 226094
rect 591102 189538 591658 190094
rect 591102 153538 591658 154094
rect 591102 117538 591658 118094
rect 591102 81538 591658 82094
rect 591102 45538 591658 46094
rect 591102 9538 591658 10094
rect 591102 -6662 591658 -6106
rect 592062 694778 592618 695334
rect 592062 658778 592618 659334
rect 592062 622778 592618 623334
rect 592062 586778 592618 587334
rect 592062 550778 592618 551334
rect 592062 514778 592618 515334
rect 592062 478778 592618 479334
rect 592062 442778 592618 443334
rect 592062 406778 592618 407334
rect 592062 370778 592618 371334
rect 592062 334778 592618 335334
rect 592062 298778 592618 299334
rect 592062 262778 592618 263334
rect 592062 226778 592618 227334
rect 592062 190778 592618 191334
rect 592062 154778 592618 155334
rect 592062 118778 592618 119334
rect 592062 82778 592618 83334
rect 592062 46778 592618 47334
rect 592062 10778 592618 11334
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 9706 711558
rect 10262 711002 45706 711558
rect 46262 711002 81706 711558
rect 82262 711002 117706 711558
rect 118262 711002 153706 711558
rect 154262 711002 189706 711558
rect 190262 711002 225706 711558
rect 226262 711002 261706 711558
rect 262262 711002 297706 711558
rect 298262 711002 333706 711558
rect 334262 711002 369706 711558
rect 370262 711002 405706 711558
rect 406262 711002 441706 711558
rect 442262 711002 477706 711558
rect 478262 711002 513706 711558
rect 514262 711002 549706 711558
rect 550262 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 8466 710598
rect 9022 710042 44466 710598
rect 45022 710042 80466 710598
rect 81022 710042 116466 710598
rect 117022 710042 152466 710598
rect 153022 710042 188466 710598
rect 189022 710042 224466 710598
rect 225022 710042 260466 710598
rect 261022 710042 296466 710598
rect 297022 710042 332466 710598
rect 333022 710042 368466 710598
rect 369022 710042 404466 710598
rect 405022 710042 440466 710598
rect 441022 710042 476466 710598
rect 477022 710042 512466 710598
rect 513022 710042 548466 710598
rect 549022 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 7226 709638
rect 7782 709082 43226 709638
rect 43782 709082 79226 709638
rect 79782 709082 115226 709638
rect 115782 709082 151226 709638
rect 151782 709082 187226 709638
rect 187782 709082 223226 709638
rect 223782 709082 259226 709638
rect 259782 709082 295226 709638
rect 295782 709082 331226 709638
rect 331782 709082 367226 709638
rect 367782 709082 403226 709638
rect 403782 709082 439226 709638
rect 439782 709082 475226 709638
rect 475782 709082 511226 709638
rect 511782 709082 547226 709638
rect 547782 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 5986 708678
rect 6542 708122 41986 708678
rect 42542 708122 77986 708678
rect 78542 708122 113986 708678
rect 114542 708122 149986 708678
rect 150542 708122 185986 708678
rect 186542 708122 221986 708678
rect 222542 708122 257986 708678
rect 258542 708122 293986 708678
rect 294542 708122 329986 708678
rect 330542 708122 365986 708678
rect 366542 708122 401986 708678
rect 402542 708122 437986 708678
rect 438542 708122 473986 708678
rect 474542 708122 509986 708678
rect 510542 708122 545986 708678
rect 546542 708122 581986 708678
rect 582542 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 4746 707718
rect 5302 707162 40746 707718
rect 41302 707162 76746 707718
rect 77302 707162 112746 707718
rect 113302 707162 148746 707718
rect 149302 707162 184746 707718
rect 185302 707162 220746 707718
rect 221302 707162 256746 707718
rect 257302 707162 292746 707718
rect 293302 707162 328746 707718
rect 329302 707162 364746 707718
rect 365302 707162 400746 707718
rect 401302 707162 436746 707718
rect 437302 707162 472746 707718
rect 473302 707162 508746 707718
rect 509302 707162 544746 707718
rect 545302 707162 580746 707718
rect 581302 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 3506 706758
rect 4062 706202 39506 706758
rect 40062 706202 75506 706758
rect 76062 706202 111506 706758
rect 112062 706202 147506 706758
rect 148062 706202 183506 706758
rect 184062 706202 219506 706758
rect 220062 706202 255506 706758
rect 256062 706202 291506 706758
rect 292062 706202 327506 706758
rect 328062 706202 363506 706758
rect 364062 706202 399506 706758
rect 400062 706202 435506 706758
rect 436062 706202 471506 706758
rect 472062 706202 507506 706758
rect 508062 706202 543506 706758
rect 544062 706202 579506 706758
rect 580062 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 2266 705798
rect 2822 705242 38266 705798
rect 38822 705242 74266 705798
rect 74822 705242 110266 705798
rect 110822 705242 146266 705798
rect 146822 705242 182266 705798
rect 182822 705242 218266 705798
rect 218822 705242 254266 705798
rect 254822 705242 290266 705798
rect 290822 705242 326266 705798
rect 326822 705242 362266 705798
rect 362822 705242 398266 705798
rect 398822 705242 434266 705798
rect 434822 705242 470266 705798
rect 470822 705242 506266 705798
rect 506822 705242 542266 705798
rect 542822 705242 578266 705798
rect 578822 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1026 704838
rect 1582 704282 37026 704838
rect 37582 704282 73026 704838
rect 73582 704282 109026 704838
rect 109582 704282 145026 704838
rect 145582 704282 181026 704838
rect 181582 704282 217026 704838
rect 217582 704282 253026 704838
rect 253582 704282 289026 704838
rect 289582 704282 325026 704838
rect 325582 704282 361026 704838
rect 361582 704282 397026 704838
rect 397582 704282 433026 704838
rect 433582 704282 469026 704838
rect 469582 704282 505026 704838
rect 505582 704282 541026 704838
rect 541582 704282 577026 704838
rect 577582 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 695334 592650 695366
rect -8726 694778 -8694 695334
rect -8138 694778 9706 695334
rect 10262 694778 45706 695334
rect 46262 694778 81706 695334
rect 82262 694778 117706 695334
rect 118262 694778 153706 695334
rect 154262 694778 189706 695334
rect 190262 694778 225706 695334
rect 226262 694778 261706 695334
rect 262262 694778 297706 695334
rect 298262 694778 333706 695334
rect 334262 694778 369706 695334
rect 370262 694778 405706 695334
rect 406262 694778 441706 695334
rect 442262 694778 477706 695334
rect 478262 694778 513706 695334
rect 514262 694778 549706 695334
rect 550262 694778 592062 695334
rect 592618 694778 592650 695334
rect -8726 694746 592650 694778
rect -8726 694094 592650 694126
rect -8726 693538 -7734 694094
rect -7178 693538 8466 694094
rect 9022 693538 44466 694094
rect 45022 693538 80466 694094
rect 81022 693538 116466 694094
rect 117022 693538 152466 694094
rect 153022 693538 188466 694094
rect 189022 693538 224466 694094
rect 225022 693538 260466 694094
rect 261022 693538 296466 694094
rect 297022 693538 332466 694094
rect 333022 693538 368466 694094
rect 369022 693538 404466 694094
rect 405022 693538 440466 694094
rect 441022 693538 476466 694094
rect 477022 693538 512466 694094
rect 513022 693538 548466 694094
rect 549022 693538 591102 694094
rect 591658 693538 592650 694094
rect -8726 693506 592650 693538
rect -8726 692854 592650 692886
rect -8726 692298 -6774 692854
rect -6218 692298 7226 692854
rect 7782 692298 43226 692854
rect 43782 692298 79226 692854
rect 79782 692298 115226 692854
rect 115782 692298 151226 692854
rect 151782 692298 187226 692854
rect 187782 692298 223226 692854
rect 223782 692298 259226 692854
rect 259782 692298 295226 692854
rect 295782 692298 331226 692854
rect 331782 692298 367226 692854
rect 367782 692298 403226 692854
rect 403782 692298 439226 692854
rect 439782 692298 475226 692854
rect 475782 692298 511226 692854
rect 511782 692298 547226 692854
rect 547782 692298 590142 692854
rect 590698 692298 592650 692854
rect -8726 692266 592650 692298
rect -8726 691614 592650 691646
rect -8726 691058 -5814 691614
rect -5258 691058 5986 691614
rect 6542 691058 41986 691614
rect 42542 691058 77986 691614
rect 78542 691058 113986 691614
rect 114542 691058 149986 691614
rect 150542 691058 185986 691614
rect 186542 691058 221986 691614
rect 222542 691058 257986 691614
rect 258542 691058 293986 691614
rect 294542 691058 329986 691614
rect 330542 691058 365986 691614
rect 366542 691058 401986 691614
rect 402542 691058 437986 691614
rect 438542 691058 473986 691614
rect 474542 691058 509986 691614
rect 510542 691058 545986 691614
rect 546542 691058 581986 691614
rect 582542 691058 589182 691614
rect 589738 691058 592650 691614
rect -8726 691026 592650 691058
rect -8726 690374 592650 690406
rect -8726 689818 -4854 690374
rect -4298 689818 4746 690374
rect 5302 689818 40746 690374
rect 41302 689818 76746 690374
rect 77302 689818 112746 690374
rect 113302 689818 148746 690374
rect 149302 689818 184746 690374
rect 185302 689818 220746 690374
rect 221302 689818 256746 690374
rect 257302 689818 292746 690374
rect 293302 689818 328746 690374
rect 329302 689818 364746 690374
rect 365302 689818 400746 690374
rect 401302 689818 436746 690374
rect 437302 689818 472746 690374
rect 473302 689818 508746 690374
rect 509302 689818 544746 690374
rect 545302 689818 580746 690374
rect 581302 689818 588222 690374
rect 588778 689818 592650 690374
rect -8726 689786 592650 689818
rect -8726 689134 592650 689166
rect -8726 688578 -3894 689134
rect -3338 688578 3506 689134
rect 4062 688578 39506 689134
rect 40062 688578 75506 689134
rect 76062 688578 111506 689134
rect 112062 688578 147506 689134
rect 148062 688578 183506 689134
rect 184062 688578 219506 689134
rect 220062 688578 255506 689134
rect 256062 688578 291506 689134
rect 292062 688578 327506 689134
rect 328062 688578 363506 689134
rect 364062 688578 399506 689134
rect 400062 688578 435506 689134
rect 436062 688578 471506 689134
rect 472062 688578 507506 689134
rect 508062 688578 543506 689134
rect 544062 688578 579506 689134
rect 580062 688578 587262 689134
rect 587818 688578 592650 689134
rect -8726 688546 592650 688578
rect -8726 687894 592650 687926
rect -8726 687338 -2934 687894
rect -2378 687338 2266 687894
rect 2822 687338 38266 687894
rect 38822 687338 74266 687894
rect 74822 687338 110266 687894
rect 110822 687338 146266 687894
rect 146822 687338 182266 687894
rect 182822 687338 218266 687894
rect 218822 687338 254266 687894
rect 254822 687338 290266 687894
rect 290822 687338 326266 687894
rect 326822 687338 362266 687894
rect 362822 687338 398266 687894
rect 398822 687338 434266 687894
rect 434822 687338 470266 687894
rect 470822 687338 506266 687894
rect 506822 687338 542266 687894
rect 542822 687338 578266 687894
rect 578822 687338 586302 687894
rect 586858 687338 592650 687894
rect -8726 687306 592650 687338
rect -8726 686654 592650 686686
rect -8726 686098 -1974 686654
rect -1418 686098 1026 686654
rect 1582 686098 37026 686654
rect 37582 686098 73026 686654
rect 73582 686098 109026 686654
rect 109582 686098 145026 686654
rect 145582 686098 181026 686654
rect 181582 686098 217026 686654
rect 217582 686098 253026 686654
rect 253582 686098 289026 686654
rect 289582 686098 325026 686654
rect 325582 686098 361026 686654
rect 361582 686098 397026 686654
rect 397582 686098 433026 686654
rect 433582 686098 469026 686654
rect 469582 686098 505026 686654
rect 505582 686098 541026 686654
rect 541582 686098 577026 686654
rect 577582 686098 585342 686654
rect 585898 686098 592650 686654
rect -8726 686066 592650 686098
rect -8726 659334 592650 659366
rect -8726 658778 -8694 659334
rect -8138 658778 9706 659334
rect 10262 658778 45706 659334
rect 46262 658778 81706 659334
rect 82262 658778 117706 659334
rect 118262 658778 153706 659334
rect 154262 658778 189706 659334
rect 190262 658778 225706 659334
rect 226262 658778 261706 659334
rect 262262 658778 297706 659334
rect 298262 658778 333706 659334
rect 334262 658778 369706 659334
rect 370262 658778 405706 659334
rect 406262 658778 441706 659334
rect 442262 658778 477706 659334
rect 478262 658778 513706 659334
rect 514262 658778 549706 659334
rect 550262 658778 592062 659334
rect 592618 658778 592650 659334
rect -8726 658746 592650 658778
rect -8726 658094 592650 658126
rect -8726 657538 -7734 658094
rect -7178 657538 8466 658094
rect 9022 657538 44466 658094
rect 45022 657538 80466 658094
rect 81022 657538 116466 658094
rect 117022 657538 152466 658094
rect 153022 657538 188466 658094
rect 189022 657538 224466 658094
rect 225022 657538 260466 658094
rect 261022 657538 296466 658094
rect 297022 657538 332466 658094
rect 333022 657538 368466 658094
rect 369022 657538 404466 658094
rect 405022 657538 440466 658094
rect 441022 657538 476466 658094
rect 477022 657538 512466 658094
rect 513022 657538 548466 658094
rect 549022 657538 591102 658094
rect 591658 657538 592650 658094
rect -8726 657506 592650 657538
rect -8726 656854 592650 656886
rect -8726 656298 -6774 656854
rect -6218 656298 7226 656854
rect 7782 656298 43226 656854
rect 43782 656298 79226 656854
rect 79782 656298 115226 656854
rect 115782 656298 151226 656854
rect 151782 656298 187226 656854
rect 187782 656298 223226 656854
rect 223782 656298 259226 656854
rect 259782 656298 295226 656854
rect 295782 656298 331226 656854
rect 331782 656298 367226 656854
rect 367782 656298 403226 656854
rect 403782 656298 439226 656854
rect 439782 656298 475226 656854
rect 475782 656298 511226 656854
rect 511782 656298 547226 656854
rect 547782 656298 590142 656854
rect 590698 656298 592650 656854
rect -8726 656266 592650 656298
rect -8726 655614 592650 655646
rect -8726 655058 -5814 655614
rect -5258 655058 5986 655614
rect 6542 655058 41986 655614
rect 42542 655058 77986 655614
rect 78542 655058 113986 655614
rect 114542 655058 149986 655614
rect 150542 655058 185986 655614
rect 186542 655058 221986 655614
rect 222542 655058 257986 655614
rect 258542 655058 293986 655614
rect 294542 655058 329986 655614
rect 330542 655058 365986 655614
rect 366542 655058 401986 655614
rect 402542 655058 437986 655614
rect 438542 655058 473986 655614
rect 474542 655058 509986 655614
rect 510542 655058 545986 655614
rect 546542 655058 581986 655614
rect 582542 655058 589182 655614
rect 589738 655058 592650 655614
rect -8726 655026 592650 655058
rect -8726 654374 592650 654406
rect -8726 653818 -4854 654374
rect -4298 653818 4746 654374
rect 5302 653818 40746 654374
rect 41302 653818 76746 654374
rect 77302 653818 112746 654374
rect 113302 653818 148746 654374
rect 149302 653818 184746 654374
rect 185302 653818 220746 654374
rect 221302 653818 256746 654374
rect 257302 653818 292746 654374
rect 293302 653818 328746 654374
rect 329302 653818 364746 654374
rect 365302 653818 400746 654374
rect 401302 653818 436746 654374
rect 437302 653818 472746 654374
rect 473302 653818 508746 654374
rect 509302 653818 544746 654374
rect 545302 653818 580746 654374
rect 581302 653818 588222 654374
rect 588778 653818 592650 654374
rect -8726 653786 592650 653818
rect -8726 653134 592650 653166
rect -8726 652578 -3894 653134
rect -3338 652578 3506 653134
rect 4062 652578 39506 653134
rect 40062 652578 75506 653134
rect 76062 652578 111506 653134
rect 112062 652578 147506 653134
rect 148062 652578 183506 653134
rect 184062 652578 219506 653134
rect 220062 652578 255506 653134
rect 256062 652578 291506 653134
rect 292062 652578 327506 653134
rect 328062 652578 363506 653134
rect 364062 652578 399506 653134
rect 400062 652578 435506 653134
rect 436062 652578 471506 653134
rect 472062 652578 507506 653134
rect 508062 652578 543506 653134
rect 544062 652578 579506 653134
rect 580062 652578 587262 653134
rect 587818 652578 592650 653134
rect -8726 652546 592650 652578
rect -8726 651894 592650 651926
rect -8726 651338 -2934 651894
rect -2378 651338 2266 651894
rect 2822 651338 38266 651894
rect 38822 651338 74266 651894
rect 74822 651338 110266 651894
rect 110822 651338 146266 651894
rect 146822 651338 182266 651894
rect 182822 651338 218266 651894
rect 218822 651338 254266 651894
rect 254822 651338 290266 651894
rect 290822 651338 326266 651894
rect 326822 651338 362266 651894
rect 362822 651338 398266 651894
rect 398822 651338 434266 651894
rect 434822 651338 470266 651894
rect 470822 651338 506266 651894
rect 506822 651338 542266 651894
rect 542822 651338 578266 651894
rect 578822 651338 586302 651894
rect 586858 651338 592650 651894
rect -8726 651306 592650 651338
rect -8726 650654 592650 650686
rect -8726 650098 -1974 650654
rect -1418 650098 1026 650654
rect 1582 650098 37026 650654
rect 37582 650098 73026 650654
rect 73582 650098 109026 650654
rect 109582 650098 145026 650654
rect 145582 650098 181026 650654
rect 181582 650098 217026 650654
rect 217582 650098 253026 650654
rect 253582 650098 289026 650654
rect 289582 650098 325026 650654
rect 325582 650098 361026 650654
rect 361582 650098 397026 650654
rect 397582 650098 433026 650654
rect 433582 650098 469026 650654
rect 469582 650098 505026 650654
rect 505582 650098 541026 650654
rect 541582 650098 577026 650654
rect 577582 650098 585342 650654
rect 585898 650098 592650 650654
rect -8726 650066 592650 650098
rect -8726 623334 592650 623366
rect -8726 622778 -8694 623334
rect -8138 622778 9706 623334
rect 10262 622778 45706 623334
rect 46262 622778 81706 623334
rect 82262 622778 117706 623334
rect 118262 622778 153706 623334
rect 154262 622778 189706 623334
rect 190262 622778 225706 623334
rect 226262 622778 261706 623334
rect 262262 622778 297706 623334
rect 298262 622778 333706 623334
rect 334262 622778 369706 623334
rect 370262 622778 405706 623334
rect 406262 622778 441706 623334
rect 442262 622778 477706 623334
rect 478262 622778 513706 623334
rect 514262 622778 549706 623334
rect 550262 622778 592062 623334
rect 592618 622778 592650 623334
rect -8726 622746 592650 622778
rect -8726 622094 592650 622126
rect -8726 621538 -7734 622094
rect -7178 621538 8466 622094
rect 9022 621538 44466 622094
rect 45022 621538 80466 622094
rect 81022 621538 116466 622094
rect 117022 621538 152466 622094
rect 153022 621538 188466 622094
rect 189022 621538 224466 622094
rect 225022 621538 260466 622094
rect 261022 621538 296466 622094
rect 297022 621538 332466 622094
rect 333022 621538 368466 622094
rect 369022 621538 404466 622094
rect 405022 621538 440466 622094
rect 441022 621538 476466 622094
rect 477022 621538 512466 622094
rect 513022 621538 548466 622094
rect 549022 621538 591102 622094
rect 591658 621538 592650 622094
rect -8726 621506 592650 621538
rect -8726 620854 592650 620886
rect -8726 620298 -6774 620854
rect -6218 620298 7226 620854
rect 7782 620298 43226 620854
rect 43782 620298 79226 620854
rect 79782 620298 115226 620854
rect 115782 620298 151226 620854
rect 151782 620298 187226 620854
rect 187782 620298 223226 620854
rect 223782 620298 259226 620854
rect 259782 620298 295226 620854
rect 295782 620298 331226 620854
rect 331782 620298 367226 620854
rect 367782 620298 403226 620854
rect 403782 620298 439226 620854
rect 439782 620298 475226 620854
rect 475782 620298 511226 620854
rect 511782 620298 547226 620854
rect 547782 620298 590142 620854
rect 590698 620298 592650 620854
rect -8726 620266 592650 620298
rect -8726 619614 592650 619646
rect -8726 619058 -5814 619614
rect -5258 619058 5986 619614
rect 6542 619058 41986 619614
rect 42542 619058 77986 619614
rect 78542 619058 113986 619614
rect 114542 619058 149986 619614
rect 150542 619058 185986 619614
rect 186542 619058 221986 619614
rect 222542 619058 257986 619614
rect 258542 619058 293986 619614
rect 294542 619058 329986 619614
rect 330542 619058 365986 619614
rect 366542 619058 401986 619614
rect 402542 619058 437986 619614
rect 438542 619058 473986 619614
rect 474542 619058 509986 619614
rect 510542 619058 545986 619614
rect 546542 619058 581986 619614
rect 582542 619058 589182 619614
rect 589738 619058 592650 619614
rect -8726 619026 592650 619058
rect -8726 618374 592650 618406
rect -8726 617818 -4854 618374
rect -4298 617818 4746 618374
rect 5302 617818 40746 618374
rect 41302 617818 76746 618374
rect 77302 617818 112746 618374
rect 113302 617818 148746 618374
rect 149302 617818 184746 618374
rect 185302 617818 220746 618374
rect 221302 617818 256746 618374
rect 257302 617818 292746 618374
rect 293302 617818 328746 618374
rect 329302 617818 364746 618374
rect 365302 617818 400746 618374
rect 401302 617818 436746 618374
rect 437302 617818 472746 618374
rect 473302 617818 508746 618374
rect 509302 617818 544746 618374
rect 545302 617818 580746 618374
rect 581302 617818 588222 618374
rect 588778 617818 592650 618374
rect -8726 617786 592650 617818
rect -8726 617134 592650 617166
rect -8726 616578 -3894 617134
rect -3338 616578 3506 617134
rect 4062 616578 39506 617134
rect 40062 616578 75506 617134
rect 76062 616578 111506 617134
rect 112062 616578 147506 617134
rect 148062 616578 183506 617134
rect 184062 616578 219506 617134
rect 220062 616578 255506 617134
rect 256062 616578 291506 617134
rect 292062 616578 327506 617134
rect 328062 616578 363506 617134
rect 364062 616578 399506 617134
rect 400062 616578 435506 617134
rect 436062 616578 471506 617134
rect 472062 616578 507506 617134
rect 508062 616578 543506 617134
rect 544062 616578 579506 617134
rect 580062 616578 587262 617134
rect 587818 616578 592650 617134
rect -8726 616546 592650 616578
rect -8726 615894 592650 615926
rect -8726 615338 -2934 615894
rect -2378 615338 2266 615894
rect 2822 615338 38266 615894
rect 38822 615338 74266 615894
rect 74822 615338 110266 615894
rect 110822 615338 146266 615894
rect 146822 615338 182266 615894
rect 182822 615338 218266 615894
rect 218822 615338 254266 615894
rect 254822 615338 290266 615894
rect 290822 615338 326266 615894
rect 326822 615338 362266 615894
rect 362822 615338 398266 615894
rect 398822 615338 434266 615894
rect 434822 615338 470266 615894
rect 470822 615338 506266 615894
rect 506822 615338 542266 615894
rect 542822 615338 578266 615894
rect 578822 615338 586302 615894
rect 586858 615338 592650 615894
rect -8726 615306 592650 615338
rect -8726 614654 592650 614686
rect -8726 614098 -1974 614654
rect -1418 614098 1026 614654
rect 1582 614098 37026 614654
rect 37582 614098 73026 614654
rect 73582 614098 109026 614654
rect 109582 614098 145026 614654
rect 145582 614098 181026 614654
rect 181582 614098 217026 614654
rect 217582 614098 253026 614654
rect 253582 614098 289026 614654
rect 289582 614098 325026 614654
rect 325582 614098 361026 614654
rect 361582 614098 397026 614654
rect 397582 614098 433026 614654
rect 433582 614098 469026 614654
rect 469582 614098 505026 614654
rect 505582 614098 541026 614654
rect 541582 614098 577026 614654
rect 577582 614098 585342 614654
rect 585898 614098 592650 614654
rect -8726 614066 592650 614098
rect -8726 587334 592650 587366
rect -8726 586778 -8694 587334
rect -8138 586778 9706 587334
rect 10262 586778 45706 587334
rect 46262 586778 81706 587334
rect 82262 586778 117706 587334
rect 118262 586778 153706 587334
rect 154262 586778 189706 587334
rect 190262 586778 225706 587334
rect 226262 586778 261706 587334
rect 262262 586778 297706 587334
rect 298262 586778 333706 587334
rect 334262 586778 369706 587334
rect 370262 586778 405706 587334
rect 406262 586778 441706 587334
rect 442262 586778 477706 587334
rect 478262 586778 513706 587334
rect 514262 586778 549706 587334
rect 550262 586778 592062 587334
rect 592618 586778 592650 587334
rect -8726 586746 592650 586778
rect -8726 586094 592650 586126
rect -8726 585538 -7734 586094
rect -7178 585538 8466 586094
rect 9022 585538 44466 586094
rect 45022 585538 80466 586094
rect 81022 585538 116466 586094
rect 117022 585538 152466 586094
rect 153022 585538 188466 586094
rect 189022 585538 224466 586094
rect 225022 585538 260466 586094
rect 261022 585538 296466 586094
rect 297022 585538 332466 586094
rect 333022 585538 368466 586094
rect 369022 585538 404466 586094
rect 405022 585538 440466 586094
rect 441022 585538 476466 586094
rect 477022 585538 512466 586094
rect 513022 585538 548466 586094
rect 549022 585538 591102 586094
rect 591658 585538 592650 586094
rect -8726 585506 592650 585538
rect -8726 584854 592650 584886
rect -8726 584298 -6774 584854
rect -6218 584298 7226 584854
rect 7782 584298 43226 584854
rect 43782 584298 79226 584854
rect 79782 584298 115226 584854
rect 115782 584298 151226 584854
rect 151782 584298 187226 584854
rect 187782 584298 223226 584854
rect 223782 584298 259226 584854
rect 259782 584298 295226 584854
rect 295782 584298 331226 584854
rect 331782 584298 367226 584854
rect 367782 584298 403226 584854
rect 403782 584298 439226 584854
rect 439782 584298 475226 584854
rect 475782 584298 511226 584854
rect 511782 584298 547226 584854
rect 547782 584298 590142 584854
rect 590698 584298 592650 584854
rect -8726 584266 592650 584298
rect -8726 583614 592650 583646
rect -8726 583058 -5814 583614
rect -5258 583058 5986 583614
rect 6542 583058 41986 583614
rect 42542 583058 77986 583614
rect 78542 583058 113986 583614
rect 114542 583058 149986 583614
rect 150542 583058 185986 583614
rect 186542 583058 221986 583614
rect 222542 583058 257986 583614
rect 258542 583058 293986 583614
rect 294542 583058 329986 583614
rect 330542 583058 365986 583614
rect 366542 583058 401986 583614
rect 402542 583058 437986 583614
rect 438542 583058 473986 583614
rect 474542 583058 509986 583614
rect 510542 583058 545986 583614
rect 546542 583058 581986 583614
rect 582542 583058 589182 583614
rect 589738 583058 592650 583614
rect -8726 583026 592650 583058
rect -8726 582374 592650 582406
rect -8726 581818 -4854 582374
rect -4298 581818 4746 582374
rect 5302 581818 40746 582374
rect 41302 581818 76746 582374
rect 77302 581818 112746 582374
rect 113302 581818 148746 582374
rect 149302 581818 184746 582374
rect 185302 581818 220746 582374
rect 221302 581818 256746 582374
rect 257302 581818 292746 582374
rect 293302 581818 328746 582374
rect 329302 581818 364746 582374
rect 365302 581818 400746 582374
rect 401302 581818 436746 582374
rect 437302 581818 472746 582374
rect 473302 581818 508746 582374
rect 509302 581818 544746 582374
rect 545302 581818 580746 582374
rect 581302 581818 588222 582374
rect 588778 581818 592650 582374
rect -8726 581786 592650 581818
rect -8726 581134 592650 581166
rect -8726 580578 -3894 581134
rect -3338 580578 3506 581134
rect 4062 580578 39506 581134
rect 40062 580578 75506 581134
rect 76062 580578 111506 581134
rect 112062 580578 147506 581134
rect 148062 580578 183506 581134
rect 184062 580578 219506 581134
rect 220062 580578 255506 581134
rect 256062 580578 291506 581134
rect 292062 580578 327506 581134
rect 328062 580578 363506 581134
rect 364062 580578 399506 581134
rect 400062 580578 435506 581134
rect 436062 580578 471506 581134
rect 472062 580578 507506 581134
rect 508062 580578 543506 581134
rect 544062 580578 579506 581134
rect 580062 580578 587262 581134
rect 587818 580578 592650 581134
rect -8726 580546 592650 580578
rect -8726 579894 592650 579926
rect -8726 579338 -2934 579894
rect -2378 579338 2266 579894
rect 2822 579338 38266 579894
rect 38822 579338 74266 579894
rect 74822 579338 110266 579894
rect 110822 579338 146266 579894
rect 146822 579338 182266 579894
rect 182822 579338 218266 579894
rect 218822 579338 254266 579894
rect 254822 579338 290266 579894
rect 290822 579338 326266 579894
rect 326822 579338 362266 579894
rect 362822 579338 398266 579894
rect 398822 579338 434266 579894
rect 434822 579338 470266 579894
rect 470822 579338 506266 579894
rect 506822 579338 542266 579894
rect 542822 579338 578266 579894
rect 578822 579338 586302 579894
rect 586858 579338 592650 579894
rect -8726 579306 592650 579338
rect -8726 578654 592650 578686
rect -8726 578098 -1974 578654
rect -1418 578098 1026 578654
rect 1582 578098 37026 578654
rect 37582 578098 73026 578654
rect 73582 578098 109026 578654
rect 109582 578098 145026 578654
rect 145582 578098 181026 578654
rect 181582 578098 217026 578654
rect 217582 578098 253026 578654
rect 253582 578098 289026 578654
rect 289582 578098 325026 578654
rect 325582 578098 361026 578654
rect 361582 578098 397026 578654
rect 397582 578098 433026 578654
rect 433582 578098 469026 578654
rect 469582 578098 505026 578654
rect 505582 578098 541026 578654
rect 541582 578098 577026 578654
rect 577582 578098 585342 578654
rect 585898 578098 592650 578654
rect -8726 578066 592650 578098
rect -8726 551334 592650 551366
rect -8726 550778 -8694 551334
rect -8138 550778 9706 551334
rect 10262 550778 45706 551334
rect 46262 550778 81706 551334
rect 82262 550778 117706 551334
rect 118262 550778 153706 551334
rect 154262 550778 189706 551334
rect 190262 550778 225706 551334
rect 226262 550778 261706 551334
rect 262262 550778 297706 551334
rect 298262 550778 333706 551334
rect 334262 550778 369706 551334
rect 370262 550778 405706 551334
rect 406262 550778 441706 551334
rect 442262 550778 477706 551334
rect 478262 550778 513706 551334
rect 514262 550778 549706 551334
rect 550262 550778 592062 551334
rect 592618 550778 592650 551334
rect -8726 550746 592650 550778
rect -8726 550094 592650 550126
rect -8726 549538 -7734 550094
rect -7178 549538 8466 550094
rect 9022 549538 44466 550094
rect 45022 549538 80466 550094
rect 81022 549538 116466 550094
rect 117022 549538 152466 550094
rect 153022 549538 188466 550094
rect 189022 549538 224466 550094
rect 225022 549538 260466 550094
rect 261022 549538 296466 550094
rect 297022 549538 332466 550094
rect 333022 549538 368466 550094
rect 369022 549538 404466 550094
rect 405022 549538 440466 550094
rect 441022 549538 476466 550094
rect 477022 549538 512466 550094
rect 513022 549538 548466 550094
rect 549022 549538 591102 550094
rect 591658 549538 592650 550094
rect -8726 549506 592650 549538
rect -8726 548854 592650 548886
rect -8726 548298 -6774 548854
rect -6218 548298 7226 548854
rect 7782 548298 43226 548854
rect 43782 548298 79226 548854
rect 79782 548298 115226 548854
rect 115782 548298 151226 548854
rect 151782 548298 187226 548854
rect 187782 548298 223226 548854
rect 223782 548298 259226 548854
rect 259782 548298 295226 548854
rect 295782 548298 331226 548854
rect 331782 548298 367226 548854
rect 367782 548298 403226 548854
rect 403782 548298 439226 548854
rect 439782 548298 475226 548854
rect 475782 548298 511226 548854
rect 511782 548298 547226 548854
rect 547782 548298 590142 548854
rect 590698 548298 592650 548854
rect -8726 548266 592650 548298
rect -8726 547614 592650 547646
rect -8726 547058 -5814 547614
rect -5258 547058 5986 547614
rect 6542 547058 41986 547614
rect 42542 547058 77986 547614
rect 78542 547058 113986 547614
rect 114542 547058 149986 547614
rect 150542 547058 185986 547614
rect 186542 547058 221986 547614
rect 222542 547058 257986 547614
rect 258542 547058 293986 547614
rect 294542 547058 329986 547614
rect 330542 547058 365986 547614
rect 366542 547058 401986 547614
rect 402542 547058 437986 547614
rect 438542 547058 473986 547614
rect 474542 547058 509986 547614
rect 510542 547058 545986 547614
rect 546542 547058 581986 547614
rect 582542 547058 589182 547614
rect 589738 547058 592650 547614
rect -8726 547026 592650 547058
rect -8726 546374 592650 546406
rect -8726 545818 -4854 546374
rect -4298 545818 4746 546374
rect 5302 545818 40746 546374
rect 41302 545818 76746 546374
rect 77302 545818 112746 546374
rect 113302 545818 148746 546374
rect 149302 545818 184746 546374
rect 185302 545818 220746 546374
rect 221302 545818 256746 546374
rect 257302 545818 292746 546374
rect 293302 545818 328746 546374
rect 329302 545818 364746 546374
rect 365302 545818 400746 546374
rect 401302 545818 436746 546374
rect 437302 545818 472746 546374
rect 473302 545818 508746 546374
rect 509302 545818 544746 546374
rect 545302 545818 580746 546374
rect 581302 545818 588222 546374
rect 588778 545818 592650 546374
rect -8726 545786 592650 545818
rect -8726 545134 592650 545166
rect -8726 544578 -3894 545134
rect -3338 544578 3506 545134
rect 4062 544578 39506 545134
rect 40062 544578 75506 545134
rect 76062 544578 111506 545134
rect 112062 544578 147506 545134
rect 148062 544578 183506 545134
rect 184062 544578 219506 545134
rect 220062 544578 255506 545134
rect 256062 544578 291506 545134
rect 292062 544578 327506 545134
rect 328062 544578 363506 545134
rect 364062 544578 399506 545134
rect 400062 544578 435506 545134
rect 436062 544578 471506 545134
rect 472062 544578 507506 545134
rect 508062 544578 543506 545134
rect 544062 544578 579506 545134
rect 580062 544578 587262 545134
rect 587818 544578 592650 545134
rect -8726 544546 592650 544578
rect -8726 543894 592650 543926
rect -8726 543338 -2934 543894
rect -2378 543338 2266 543894
rect 2822 543338 38266 543894
rect 38822 543338 74266 543894
rect 74822 543338 110266 543894
rect 110822 543338 146266 543894
rect 146822 543338 182266 543894
rect 182822 543338 218266 543894
rect 218822 543338 254266 543894
rect 254822 543338 290266 543894
rect 290822 543338 326266 543894
rect 326822 543338 362266 543894
rect 362822 543338 398266 543894
rect 398822 543338 434266 543894
rect 434822 543338 470266 543894
rect 470822 543338 506266 543894
rect 506822 543338 542266 543894
rect 542822 543338 578266 543894
rect 578822 543338 586302 543894
rect 586858 543338 592650 543894
rect -8726 543306 592650 543338
rect -8726 542654 592650 542686
rect -8726 542098 -1974 542654
rect -1418 542098 1026 542654
rect 1582 542098 37026 542654
rect 37582 542098 73026 542654
rect 73582 542098 109026 542654
rect 109582 542098 145026 542654
rect 145582 542098 181026 542654
rect 181582 542098 217026 542654
rect 217582 542098 253026 542654
rect 253582 542098 289026 542654
rect 289582 542098 325026 542654
rect 325582 542098 361026 542654
rect 361582 542098 397026 542654
rect 397582 542098 433026 542654
rect 433582 542098 469026 542654
rect 469582 542098 505026 542654
rect 505582 542098 541026 542654
rect 541582 542098 577026 542654
rect 577582 542098 585342 542654
rect 585898 542098 592650 542654
rect -8726 542066 592650 542098
rect -8726 515334 592650 515366
rect -8726 514778 -8694 515334
rect -8138 514778 9706 515334
rect 10262 514778 45706 515334
rect 46262 514778 81706 515334
rect 82262 514778 117706 515334
rect 118262 514778 153706 515334
rect 154262 514778 189706 515334
rect 190262 514778 225706 515334
rect 226262 514778 261706 515334
rect 262262 514778 297706 515334
rect 298262 514778 333706 515334
rect 334262 514778 369706 515334
rect 370262 514778 405706 515334
rect 406262 514778 441706 515334
rect 442262 514778 477706 515334
rect 478262 514778 513706 515334
rect 514262 514778 549706 515334
rect 550262 514778 592062 515334
rect 592618 514778 592650 515334
rect -8726 514746 592650 514778
rect -8726 514094 592650 514126
rect -8726 513538 -7734 514094
rect -7178 513538 8466 514094
rect 9022 513538 44466 514094
rect 45022 513538 80466 514094
rect 81022 513538 116466 514094
rect 117022 513538 152466 514094
rect 153022 513538 188466 514094
rect 189022 513538 224466 514094
rect 225022 513538 260466 514094
rect 261022 513538 296466 514094
rect 297022 513538 332466 514094
rect 333022 513538 368466 514094
rect 369022 513538 404466 514094
rect 405022 513538 440466 514094
rect 441022 513538 476466 514094
rect 477022 513538 512466 514094
rect 513022 513538 548466 514094
rect 549022 513538 591102 514094
rect 591658 513538 592650 514094
rect -8726 513506 592650 513538
rect -8726 512854 592650 512886
rect -8726 512298 -6774 512854
rect -6218 512298 7226 512854
rect 7782 512298 43226 512854
rect 43782 512298 79226 512854
rect 79782 512298 115226 512854
rect 115782 512298 151226 512854
rect 151782 512298 187226 512854
rect 187782 512298 223226 512854
rect 223782 512298 259226 512854
rect 259782 512298 295226 512854
rect 295782 512298 331226 512854
rect 331782 512298 367226 512854
rect 367782 512298 403226 512854
rect 403782 512298 439226 512854
rect 439782 512298 475226 512854
rect 475782 512298 511226 512854
rect 511782 512298 547226 512854
rect 547782 512298 590142 512854
rect 590698 512298 592650 512854
rect -8726 512266 592650 512298
rect -8726 511614 592650 511646
rect -8726 511058 -5814 511614
rect -5258 511058 5986 511614
rect 6542 511058 41986 511614
rect 42542 511058 77986 511614
rect 78542 511058 113986 511614
rect 114542 511058 149986 511614
rect 150542 511058 185986 511614
rect 186542 511058 221986 511614
rect 222542 511058 257986 511614
rect 258542 511058 293986 511614
rect 294542 511058 329986 511614
rect 330542 511058 365986 511614
rect 366542 511058 401986 511614
rect 402542 511058 437986 511614
rect 438542 511058 473986 511614
rect 474542 511058 509986 511614
rect 510542 511058 545986 511614
rect 546542 511058 581986 511614
rect 582542 511058 589182 511614
rect 589738 511058 592650 511614
rect -8726 511026 592650 511058
rect -8726 510374 592650 510406
rect -8726 509818 -4854 510374
rect -4298 509818 4746 510374
rect 5302 509818 40746 510374
rect 41302 509818 76746 510374
rect 77302 509818 112746 510374
rect 113302 509818 148746 510374
rect 149302 509818 184746 510374
rect 185302 509818 220746 510374
rect 221302 509818 256746 510374
rect 257302 509818 292746 510374
rect 293302 509818 328746 510374
rect 329302 509818 364746 510374
rect 365302 509818 400746 510374
rect 401302 509818 436746 510374
rect 437302 509818 472746 510374
rect 473302 509818 508746 510374
rect 509302 509818 544746 510374
rect 545302 509818 580746 510374
rect 581302 509818 588222 510374
rect 588778 509818 592650 510374
rect -8726 509786 592650 509818
rect -8726 509134 592650 509166
rect -8726 508578 -3894 509134
rect -3338 508578 3506 509134
rect 4062 508578 39506 509134
rect 40062 508578 75506 509134
rect 76062 508578 111506 509134
rect 112062 508578 147506 509134
rect 148062 508578 183506 509134
rect 184062 508578 219506 509134
rect 220062 508578 255506 509134
rect 256062 508578 291506 509134
rect 292062 508578 327506 509134
rect 328062 508578 363506 509134
rect 364062 508578 399506 509134
rect 400062 508578 435506 509134
rect 436062 508578 471506 509134
rect 472062 508578 507506 509134
rect 508062 508578 543506 509134
rect 544062 508578 579506 509134
rect 580062 508578 587262 509134
rect 587818 508578 592650 509134
rect -8726 508546 592650 508578
rect -8726 507894 592650 507926
rect -8726 507338 -2934 507894
rect -2378 507338 2266 507894
rect 2822 507338 38266 507894
rect 38822 507338 74266 507894
rect 74822 507338 110266 507894
rect 110822 507338 146266 507894
rect 146822 507338 182266 507894
rect 182822 507338 218266 507894
rect 218822 507338 254266 507894
rect 254822 507338 290266 507894
rect 290822 507338 326266 507894
rect 326822 507338 362266 507894
rect 362822 507338 398266 507894
rect 398822 507338 434266 507894
rect 434822 507338 470266 507894
rect 470822 507338 506266 507894
rect 506822 507338 542266 507894
rect 542822 507338 578266 507894
rect 578822 507338 586302 507894
rect 586858 507338 592650 507894
rect -8726 507306 592650 507338
rect -8726 506654 592650 506686
rect -8726 506098 -1974 506654
rect -1418 506098 1026 506654
rect 1582 506098 37026 506654
rect 37582 506098 73026 506654
rect 73582 506098 109026 506654
rect 109582 506098 145026 506654
rect 145582 506098 181026 506654
rect 181582 506098 217026 506654
rect 217582 506098 253026 506654
rect 253582 506098 289026 506654
rect 289582 506098 325026 506654
rect 325582 506098 361026 506654
rect 361582 506098 397026 506654
rect 397582 506098 433026 506654
rect 433582 506098 469026 506654
rect 469582 506098 505026 506654
rect 505582 506098 541026 506654
rect 541582 506098 577026 506654
rect 577582 506098 585342 506654
rect 585898 506098 592650 506654
rect -8726 506066 592650 506098
rect -8726 479334 592650 479366
rect -8726 478778 -8694 479334
rect -8138 478778 9706 479334
rect 10262 478778 45706 479334
rect 46262 478778 81706 479334
rect 82262 478778 117706 479334
rect 118262 478778 153706 479334
rect 154262 478778 189706 479334
rect 190262 478778 225706 479334
rect 226262 478778 261706 479334
rect 262262 478778 297706 479334
rect 298262 478778 333706 479334
rect 334262 478778 369706 479334
rect 370262 478778 405706 479334
rect 406262 478778 441706 479334
rect 442262 478778 477706 479334
rect 478262 478778 513706 479334
rect 514262 478778 549706 479334
rect 550262 478778 592062 479334
rect 592618 478778 592650 479334
rect -8726 478746 592650 478778
rect -8726 478094 592650 478126
rect -8726 477538 -7734 478094
rect -7178 477538 8466 478094
rect 9022 477538 44466 478094
rect 45022 477538 80466 478094
rect 81022 477538 116466 478094
rect 117022 477538 152466 478094
rect 153022 477538 188466 478094
rect 189022 477538 224466 478094
rect 225022 477538 260466 478094
rect 261022 477538 296466 478094
rect 297022 477538 332466 478094
rect 333022 477538 368466 478094
rect 369022 477538 404466 478094
rect 405022 477538 440466 478094
rect 441022 477538 476466 478094
rect 477022 477538 512466 478094
rect 513022 477538 548466 478094
rect 549022 477538 591102 478094
rect 591658 477538 592650 478094
rect -8726 477506 592650 477538
rect -8726 476854 592650 476886
rect -8726 476298 -6774 476854
rect -6218 476298 7226 476854
rect 7782 476298 43226 476854
rect 43782 476298 79226 476854
rect 79782 476298 115226 476854
rect 115782 476298 151226 476854
rect 151782 476298 187226 476854
rect 187782 476298 223226 476854
rect 223782 476298 259226 476854
rect 259782 476298 295226 476854
rect 295782 476298 331226 476854
rect 331782 476298 367226 476854
rect 367782 476298 403226 476854
rect 403782 476298 439226 476854
rect 439782 476298 475226 476854
rect 475782 476298 511226 476854
rect 511782 476298 547226 476854
rect 547782 476298 590142 476854
rect 590698 476298 592650 476854
rect -8726 476266 592650 476298
rect -8726 475614 592650 475646
rect -8726 475058 -5814 475614
rect -5258 475058 5986 475614
rect 6542 475058 41986 475614
rect 42542 475058 77986 475614
rect 78542 475058 113986 475614
rect 114542 475058 149986 475614
rect 150542 475058 185986 475614
rect 186542 475058 221986 475614
rect 222542 475058 257986 475614
rect 258542 475058 293986 475614
rect 294542 475058 329986 475614
rect 330542 475058 365986 475614
rect 366542 475058 401986 475614
rect 402542 475058 437986 475614
rect 438542 475058 473986 475614
rect 474542 475058 509986 475614
rect 510542 475058 545986 475614
rect 546542 475058 581986 475614
rect 582542 475058 589182 475614
rect 589738 475058 592650 475614
rect -8726 475026 592650 475058
rect -8726 474374 592650 474406
rect -8726 473818 -4854 474374
rect -4298 473818 4746 474374
rect 5302 473818 40746 474374
rect 41302 473818 76746 474374
rect 77302 473818 112746 474374
rect 113302 473818 148746 474374
rect 149302 473818 184746 474374
rect 185302 473818 220746 474374
rect 221302 473818 256746 474374
rect 257302 473818 292746 474374
rect 293302 473818 328746 474374
rect 329302 473818 364746 474374
rect 365302 473818 400746 474374
rect 401302 473818 436746 474374
rect 437302 473818 472746 474374
rect 473302 473818 508746 474374
rect 509302 473818 544746 474374
rect 545302 473818 580746 474374
rect 581302 473818 588222 474374
rect 588778 473818 592650 474374
rect -8726 473786 592650 473818
rect -8726 473134 592650 473166
rect -8726 472578 -3894 473134
rect -3338 472578 3506 473134
rect 4062 472578 39506 473134
rect 40062 472578 75506 473134
rect 76062 472578 111506 473134
rect 112062 472578 147506 473134
rect 148062 472578 183506 473134
rect 184062 472578 219506 473134
rect 220062 472578 255506 473134
rect 256062 472578 291506 473134
rect 292062 472578 327506 473134
rect 328062 472578 363506 473134
rect 364062 472578 399506 473134
rect 400062 472578 435506 473134
rect 436062 472578 471506 473134
rect 472062 472578 507506 473134
rect 508062 472578 543506 473134
rect 544062 472578 579506 473134
rect 580062 472578 587262 473134
rect 587818 472578 592650 473134
rect -8726 472546 592650 472578
rect -8726 471894 592650 471926
rect -8726 471338 -2934 471894
rect -2378 471338 2266 471894
rect 2822 471338 38266 471894
rect 38822 471338 74266 471894
rect 74822 471338 110266 471894
rect 110822 471338 146266 471894
rect 146822 471338 182266 471894
rect 182822 471338 218266 471894
rect 218822 471338 254266 471894
rect 254822 471338 290266 471894
rect 290822 471338 326266 471894
rect 326822 471338 362266 471894
rect 362822 471338 398266 471894
rect 398822 471338 434266 471894
rect 434822 471338 470266 471894
rect 470822 471338 506266 471894
rect 506822 471338 542266 471894
rect 542822 471338 578266 471894
rect 578822 471338 586302 471894
rect 586858 471338 592650 471894
rect -8726 471306 592650 471338
rect -8726 470654 592650 470686
rect -8726 470098 -1974 470654
rect -1418 470098 1026 470654
rect 1582 470098 37026 470654
rect 37582 470098 73026 470654
rect 73582 470098 109026 470654
rect 109582 470098 145026 470654
rect 145582 470098 181026 470654
rect 181582 470098 217026 470654
rect 217582 470098 253026 470654
rect 253582 470098 289026 470654
rect 289582 470098 325026 470654
rect 325582 470098 361026 470654
rect 361582 470098 397026 470654
rect 397582 470098 433026 470654
rect 433582 470098 469026 470654
rect 469582 470098 505026 470654
rect 505582 470098 541026 470654
rect 541582 470098 577026 470654
rect 577582 470098 585342 470654
rect 585898 470098 592650 470654
rect -8726 470066 592650 470098
rect -8726 443334 592650 443366
rect -8726 442778 -8694 443334
rect -8138 442778 9706 443334
rect 10262 442778 45706 443334
rect 46262 442778 81706 443334
rect 82262 442778 117706 443334
rect 118262 442778 153706 443334
rect 154262 442778 189706 443334
rect 190262 442778 225706 443334
rect 226262 442778 261706 443334
rect 262262 442778 297706 443334
rect 298262 442778 333706 443334
rect 334262 442778 369706 443334
rect 370262 442778 405706 443334
rect 406262 442778 441706 443334
rect 442262 442778 477706 443334
rect 478262 442778 513706 443334
rect 514262 442778 549706 443334
rect 550262 442778 592062 443334
rect 592618 442778 592650 443334
rect -8726 442746 592650 442778
rect -8726 442094 592650 442126
rect -8726 441538 -7734 442094
rect -7178 441538 8466 442094
rect 9022 441538 44466 442094
rect 45022 441538 80466 442094
rect 81022 441538 116466 442094
rect 117022 441538 152466 442094
rect 153022 441538 188466 442094
rect 189022 441538 224466 442094
rect 225022 441538 260466 442094
rect 261022 441538 296466 442094
rect 297022 441538 332466 442094
rect 333022 441538 368466 442094
rect 369022 441538 404466 442094
rect 405022 441538 440466 442094
rect 441022 441538 476466 442094
rect 477022 441538 512466 442094
rect 513022 441538 548466 442094
rect 549022 441538 591102 442094
rect 591658 441538 592650 442094
rect -8726 441506 592650 441538
rect -8726 440854 592650 440886
rect -8726 440298 -6774 440854
rect -6218 440298 7226 440854
rect 7782 440298 43226 440854
rect 43782 440298 79226 440854
rect 79782 440298 115226 440854
rect 115782 440298 151226 440854
rect 151782 440298 187226 440854
rect 187782 440298 223226 440854
rect 223782 440298 259226 440854
rect 259782 440298 295226 440854
rect 295782 440298 331226 440854
rect 331782 440298 367226 440854
rect 367782 440298 403226 440854
rect 403782 440298 439226 440854
rect 439782 440298 475226 440854
rect 475782 440298 511226 440854
rect 511782 440298 547226 440854
rect 547782 440298 590142 440854
rect 590698 440298 592650 440854
rect -8726 440266 592650 440298
rect -8726 439614 592650 439646
rect -8726 439058 -5814 439614
rect -5258 439058 5986 439614
rect 6542 439058 41986 439614
rect 42542 439058 77986 439614
rect 78542 439058 113986 439614
rect 114542 439058 149986 439614
rect 150542 439058 185986 439614
rect 186542 439058 221986 439614
rect 222542 439058 257986 439614
rect 258542 439058 293986 439614
rect 294542 439058 329986 439614
rect 330542 439058 365986 439614
rect 366542 439058 401986 439614
rect 402542 439058 437986 439614
rect 438542 439058 473986 439614
rect 474542 439058 509986 439614
rect 510542 439058 581986 439614
rect 582542 439058 589182 439614
rect 589738 439058 592650 439614
rect -8726 439026 592650 439058
rect -8726 438374 592650 438406
rect -8726 437818 -4854 438374
rect -4298 437818 4746 438374
rect 5302 437818 40746 438374
rect 41302 437818 76746 438374
rect 77302 437818 112746 438374
rect 113302 437818 148746 438374
rect 149302 437818 184746 438374
rect 185302 437818 220746 438374
rect 221302 437818 256746 438374
rect 257302 437818 292746 438374
rect 293302 437818 328746 438374
rect 329302 437818 364746 438374
rect 365302 437818 400746 438374
rect 401302 437818 436746 438374
rect 437302 437818 472746 438374
rect 473302 437818 508746 438374
rect 509302 437818 580746 438374
rect 581302 437818 588222 438374
rect 588778 437818 592650 438374
rect -8726 437786 592650 437818
rect -8726 437134 592650 437166
rect -8726 436578 -3894 437134
rect -3338 436578 3506 437134
rect 4062 436578 39506 437134
rect 40062 436578 75506 437134
rect 76062 436578 111506 437134
rect 112062 436578 147506 437134
rect 148062 436578 183506 437134
rect 184062 436578 219506 437134
rect 220062 436578 255506 437134
rect 256062 436578 291506 437134
rect 292062 436578 327506 437134
rect 328062 436578 363506 437134
rect 364062 436578 399506 437134
rect 400062 436578 435506 437134
rect 436062 436578 471506 437134
rect 472062 436578 507506 437134
rect 508062 436578 579506 437134
rect 580062 436578 587262 437134
rect 587818 436578 592650 437134
rect -8726 436546 592650 436578
rect -8726 435894 592650 435926
rect -8726 435338 -2934 435894
rect -2378 435338 2266 435894
rect 2822 435338 38266 435894
rect 38822 435338 74266 435894
rect 74822 435338 110266 435894
rect 110822 435338 146266 435894
rect 146822 435338 182266 435894
rect 182822 435338 218266 435894
rect 218822 435338 254266 435894
rect 254822 435338 290266 435894
rect 290822 435338 326266 435894
rect 326822 435338 362266 435894
rect 362822 435338 398266 435894
rect 398822 435338 434266 435894
rect 434822 435338 470266 435894
rect 470822 435338 506266 435894
rect 506822 435658 540918 435894
rect 541154 435658 542850 435894
rect 543086 435658 544782 435894
rect 545018 435658 546714 435894
rect 546950 435658 578266 435894
rect 506822 435574 578266 435658
rect 506822 435338 540918 435574
rect 541154 435338 542850 435574
rect 543086 435338 544782 435574
rect 545018 435338 546714 435574
rect 546950 435338 578266 435574
rect 578822 435338 586302 435894
rect 586858 435338 592650 435894
rect -8726 435306 592650 435338
rect -8726 434654 592650 434686
rect -8726 434098 -1974 434654
rect -1418 434098 1026 434654
rect 1582 434098 37026 434654
rect 37582 434098 73026 434654
rect 73582 434098 109026 434654
rect 109582 434098 145026 434654
rect 145582 434098 181026 434654
rect 181582 434098 217026 434654
rect 217582 434098 253026 434654
rect 253582 434098 289026 434654
rect 289582 434098 325026 434654
rect 325582 434098 361026 434654
rect 361582 434098 397026 434654
rect 397582 434098 433026 434654
rect 433582 434098 469026 434654
rect 469582 434098 505026 434654
rect 505582 434418 539952 434654
rect 540188 434418 541884 434654
rect 542120 434418 543816 434654
rect 544052 434418 545748 434654
rect 545984 434418 577026 434654
rect 505582 434334 577026 434418
rect 505582 434098 539952 434334
rect 540188 434098 541884 434334
rect 542120 434098 543816 434334
rect 544052 434098 545748 434334
rect 545984 434098 577026 434334
rect 577582 434098 585342 434654
rect 585898 434098 592650 434654
rect -8726 434066 592650 434098
rect -8726 407334 592650 407366
rect -8726 406778 -8694 407334
rect -8138 406778 9706 407334
rect 10262 406778 45706 407334
rect 46262 406778 81706 407334
rect 82262 406778 117706 407334
rect 118262 406778 153706 407334
rect 154262 406778 189706 407334
rect 190262 406778 225706 407334
rect 226262 406778 261706 407334
rect 262262 406778 297706 407334
rect 298262 406778 333706 407334
rect 334262 406778 369706 407334
rect 370262 406778 405706 407334
rect 406262 406778 441706 407334
rect 442262 406778 477706 407334
rect 478262 406778 513706 407334
rect 514262 406778 549706 407334
rect 550262 406778 592062 407334
rect 592618 406778 592650 407334
rect -8726 406746 592650 406778
rect -8726 406094 592650 406126
rect -8726 405538 -7734 406094
rect -7178 405538 8466 406094
rect 9022 405538 44466 406094
rect 45022 405538 80466 406094
rect 81022 405538 116466 406094
rect 117022 405538 152466 406094
rect 153022 405538 188466 406094
rect 189022 405538 224466 406094
rect 225022 405538 260466 406094
rect 261022 405538 296466 406094
rect 297022 405538 332466 406094
rect 333022 405538 368466 406094
rect 369022 405538 404466 406094
rect 405022 405538 440466 406094
rect 441022 405538 476466 406094
rect 477022 405538 512466 406094
rect 513022 405538 548466 406094
rect 549022 405538 591102 406094
rect 591658 405538 592650 406094
rect -8726 405506 592650 405538
rect -8726 404854 592650 404886
rect -8726 404298 -6774 404854
rect -6218 404298 7226 404854
rect 7782 404298 43226 404854
rect 43782 404298 79226 404854
rect 79782 404298 115226 404854
rect 115782 404298 151226 404854
rect 151782 404298 187226 404854
rect 187782 404298 223226 404854
rect 223782 404298 259226 404854
rect 259782 404298 295226 404854
rect 295782 404298 331226 404854
rect 331782 404298 367226 404854
rect 367782 404298 403226 404854
rect 403782 404298 439226 404854
rect 439782 404298 475226 404854
rect 475782 404298 511226 404854
rect 511782 404298 547226 404854
rect 547782 404298 590142 404854
rect 590698 404298 592650 404854
rect -8726 404266 592650 404298
rect -8726 403614 592650 403646
rect -8726 403058 -5814 403614
rect -5258 403058 5986 403614
rect 6542 403058 41986 403614
rect 42542 403058 77986 403614
rect 78542 403058 113986 403614
rect 114542 403058 149986 403614
rect 150542 403058 185986 403614
rect 186542 403058 221986 403614
rect 222542 403058 257986 403614
rect 258542 403058 293986 403614
rect 294542 403058 329986 403614
rect 330542 403058 365986 403614
rect 366542 403058 401986 403614
rect 402542 403058 437986 403614
rect 438542 403058 473986 403614
rect 474542 403058 509986 403614
rect 510542 403058 581986 403614
rect 582542 403058 589182 403614
rect 589738 403058 592650 403614
rect -8726 403026 592650 403058
rect -8726 402374 592650 402406
rect -8726 401818 -4854 402374
rect -4298 401818 4746 402374
rect 5302 401818 40746 402374
rect 41302 401818 76746 402374
rect 77302 401818 112746 402374
rect 113302 401818 148746 402374
rect 149302 401818 184746 402374
rect 185302 401818 220746 402374
rect 221302 401818 256746 402374
rect 257302 401818 292746 402374
rect 293302 401818 328746 402374
rect 329302 401818 364746 402374
rect 365302 401818 400746 402374
rect 401302 401818 436746 402374
rect 437302 401818 472746 402374
rect 473302 401818 508746 402374
rect 509302 401818 580746 402374
rect 581302 401818 588222 402374
rect 588778 401818 592650 402374
rect -8726 401786 592650 401818
rect -8726 401134 592650 401166
rect -8726 400578 -3894 401134
rect -3338 400578 3506 401134
rect 4062 400578 39506 401134
rect 40062 400578 75506 401134
rect 76062 400578 111506 401134
rect 112062 400578 147506 401134
rect 148062 400578 183506 401134
rect 184062 400578 219506 401134
rect 220062 400578 255506 401134
rect 256062 400578 291506 401134
rect 292062 400578 327506 401134
rect 328062 400578 363506 401134
rect 364062 400578 399506 401134
rect 400062 400578 435506 401134
rect 436062 400578 471506 401134
rect 472062 400578 507506 401134
rect 508062 400578 579506 401134
rect 580062 400578 587262 401134
rect 587818 400578 592650 401134
rect -8726 400546 592650 400578
rect -8726 399894 592650 399926
rect -8726 399338 -2934 399894
rect -2378 399338 2266 399894
rect 2822 399338 38266 399894
rect 38822 399338 74266 399894
rect 74822 399338 110266 399894
rect 110822 399338 146266 399894
rect 146822 399338 182266 399894
rect 182822 399338 218266 399894
rect 218822 399338 254266 399894
rect 254822 399338 290266 399894
rect 290822 399338 326266 399894
rect 326822 399338 362266 399894
rect 362822 399338 398266 399894
rect 398822 399338 434266 399894
rect 434822 399338 470266 399894
rect 470822 399338 506266 399894
rect 506822 399658 540918 399894
rect 541154 399658 542850 399894
rect 543086 399658 544782 399894
rect 545018 399658 546714 399894
rect 546950 399658 578266 399894
rect 506822 399574 578266 399658
rect 506822 399338 540918 399574
rect 541154 399338 542850 399574
rect 543086 399338 544782 399574
rect 545018 399338 546714 399574
rect 546950 399338 578266 399574
rect 578822 399338 586302 399894
rect 586858 399338 592650 399894
rect -8726 399306 592650 399338
rect -8726 398654 592650 398686
rect -8726 398098 -1974 398654
rect -1418 398098 1026 398654
rect 1582 398098 37026 398654
rect 37582 398098 73026 398654
rect 73582 398098 109026 398654
rect 109582 398098 145026 398654
rect 145582 398098 181026 398654
rect 181582 398098 217026 398654
rect 217582 398098 253026 398654
rect 253582 398098 289026 398654
rect 289582 398098 325026 398654
rect 325582 398098 361026 398654
rect 361582 398098 397026 398654
rect 397582 398098 433026 398654
rect 433582 398098 469026 398654
rect 469582 398098 505026 398654
rect 505582 398418 539952 398654
rect 540188 398418 541884 398654
rect 542120 398418 543816 398654
rect 544052 398418 545748 398654
rect 545984 398418 577026 398654
rect 505582 398334 577026 398418
rect 505582 398098 539952 398334
rect 540188 398098 541884 398334
rect 542120 398098 543816 398334
rect 544052 398098 545748 398334
rect 545984 398098 577026 398334
rect 577582 398098 585342 398654
rect 585898 398098 592650 398654
rect -8726 398066 592650 398098
rect -8726 371334 592650 371366
rect -8726 370778 -8694 371334
rect -8138 370778 9706 371334
rect 10262 370778 45706 371334
rect 46262 370778 81706 371334
rect 82262 370778 117706 371334
rect 118262 370778 153706 371334
rect 154262 370778 189706 371334
rect 190262 370778 225706 371334
rect 226262 370778 261706 371334
rect 262262 370778 297706 371334
rect 298262 370778 333706 371334
rect 334262 370778 369706 371334
rect 370262 370778 405706 371334
rect 406262 370778 441706 371334
rect 442262 370778 477706 371334
rect 478262 370778 513706 371334
rect 514262 370778 549706 371334
rect 550262 370778 592062 371334
rect 592618 370778 592650 371334
rect -8726 370746 592650 370778
rect -8726 370094 592650 370126
rect -8726 369538 -7734 370094
rect -7178 369538 8466 370094
rect 9022 369538 44466 370094
rect 45022 369538 80466 370094
rect 81022 369538 116466 370094
rect 117022 369538 152466 370094
rect 153022 369538 188466 370094
rect 189022 369538 224466 370094
rect 225022 369538 260466 370094
rect 261022 369538 296466 370094
rect 297022 369538 332466 370094
rect 333022 369538 368466 370094
rect 369022 369538 404466 370094
rect 405022 369538 440466 370094
rect 441022 369538 476466 370094
rect 477022 369538 512466 370094
rect 513022 369538 548466 370094
rect 549022 369538 591102 370094
rect 591658 369538 592650 370094
rect -8726 369506 592650 369538
rect -8726 368854 592650 368886
rect -8726 368298 -6774 368854
rect -6218 368298 7226 368854
rect 7782 368298 43226 368854
rect 43782 368298 79226 368854
rect 79782 368298 115226 368854
rect 115782 368298 151226 368854
rect 151782 368298 187226 368854
rect 187782 368298 223226 368854
rect 223782 368298 259226 368854
rect 259782 368298 295226 368854
rect 295782 368298 331226 368854
rect 331782 368298 367226 368854
rect 367782 368298 403226 368854
rect 403782 368298 439226 368854
rect 439782 368298 475226 368854
rect 475782 368298 511226 368854
rect 511782 368298 547226 368854
rect 547782 368298 590142 368854
rect 590698 368298 592650 368854
rect -8726 368266 592650 368298
rect -8726 367614 592650 367646
rect -8726 367058 -5814 367614
rect -5258 367058 5986 367614
rect 6542 367058 41986 367614
rect 42542 367058 77986 367614
rect 78542 367058 113986 367614
rect 114542 367058 149986 367614
rect 150542 367058 185986 367614
rect 186542 367058 221986 367614
rect 222542 367058 257986 367614
rect 258542 367058 293986 367614
rect 294542 367058 329986 367614
rect 330542 367058 365986 367614
rect 366542 367058 401986 367614
rect 402542 367058 437986 367614
rect 438542 367058 473986 367614
rect 474542 367058 509986 367614
rect 510542 367058 581986 367614
rect 582542 367058 589182 367614
rect 589738 367058 592650 367614
rect -8726 367026 592650 367058
rect -8726 366374 592650 366406
rect -8726 365818 -4854 366374
rect -4298 365818 4746 366374
rect 5302 365818 40746 366374
rect 41302 365818 76746 366374
rect 77302 365818 112746 366374
rect 113302 365818 148746 366374
rect 149302 365818 184746 366374
rect 185302 365818 220746 366374
rect 221302 365818 256746 366374
rect 257302 365818 292746 366374
rect 293302 365818 328746 366374
rect 329302 365818 364746 366374
rect 365302 365818 400746 366374
rect 401302 365818 436746 366374
rect 437302 365818 472746 366374
rect 473302 365818 508746 366374
rect 509302 365818 580746 366374
rect 581302 365818 588222 366374
rect 588778 365818 592650 366374
rect -8726 365786 592650 365818
rect -8726 365134 592650 365166
rect -8726 364578 -3894 365134
rect -3338 364578 3506 365134
rect 4062 364578 39506 365134
rect 40062 364578 75506 365134
rect 76062 364578 111506 365134
rect 112062 364578 147506 365134
rect 148062 364578 183506 365134
rect 184062 364578 219506 365134
rect 220062 364578 255506 365134
rect 256062 364578 291506 365134
rect 292062 364578 327506 365134
rect 328062 364578 363506 365134
rect 364062 364578 399506 365134
rect 400062 364578 435506 365134
rect 436062 364578 471506 365134
rect 472062 364578 507506 365134
rect 508062 364578 579506 365134
rect 580062 364578 587262 365134
rect 587818 364578 592650 365134
rect -8726 364546 592650 364578
rect -8726 363894 592650 363926
rect -8726 363338 -2934 363894
rect -2378 363338 2266 363894
rect 2822 363338 38266 363894
rect 38822 363338 74266 363894
rect 74822 363338 110266 363894
rect 110822 363338 146266 363894
rect 146822 363338 182266 363894
rect 182822 363338 218266 363894
rect 218822 363338 254266 363894
rect 254822 363338 290266 363894
rect 290822 363338 326266 363894
rect 326822 363338 362266 363894
rect 362822 363338 398266 363894
rect 398822 363338 434266 363894
rect 434822 363338 470266 363894
rect 470822 363338 506266 363894
rect 506822 363658 540918 363894
rect 541154 363658 542850 363894
rect 543086 363658 544782 363894
rect 545018 363658 546714 363894
rect 546950 363658 578266 363894
rect 506822 363574 578266 363658
rect 506822 363338 540918 363574
rect 541154 363338 542850 363574
rect 543086 363338 544782 363574
rect 545018 363338 546714 363574
rect 546950 363338 578266 363574
rect 578822 363338 586302 363894
rect 586858 363338 592650 363894
rect -8726 363306 592650 363338
rect -8726 362654 592650 362686
rect -8726 362098 -1974 362654
rect -1418 362098 1026 362654
rect 1582 362098 37026 362654
rect 37582 362098 73026 362654
rect 73582 362098 109026 362654
rect 109582 362098 145026 362654
rect 145582 362098 181026 362654
rect 181582 362098 217026 362654
rect 217582 362098 253026 362654
rect 253582 362098 289026 362654
rect 289582 362098 325026 362654
rect 325582 362098 361026 362654
rect 361582 362098 397026 362654
rect 397582 362098 433026 362654
rect 433582 362098 469026 362654
rect 469582 362098 505026 362654
rect 505582 362418 539952 362654
rect 540188 362418 541884 362654
rect 542120 362418 543816 362654
rect 544052 362418 545748 362654
rect 545984 362418 577026 362654
rect 505582 362334 577026 362418
rect 505582 362098 539952 362334
rect 540188 362098 541884 362334
rect 542120 362098 543816 362334
rect 544052 362098 545748 362334
rect 545984 362098 577026 362334
rect 577582 362098 585342 362654
rect 585898 362098 592650 362654
rect -8726 362066 592650 362098
rect -8726 335334 592650 335366
rect -8726 334778 -8694 335334
rect -8138 334778 9706 335334
rect 10262 334778 45706 335334
rect 46262 334778 81706 335334
rect 82262 334778 117706 335334
rect 118262 334778 153706 335334
rect 154262 334778 189706 335334
rect 190262 334778 225706 335334
rect 226262 334778 261706 335334
rect 262262 334778 297706 335334
rect 298262 334778 333706 335334
rect 334262 334778 369706 335334
rect 370262 334778 405706 335334
rect 406262 334778 441706 335334
rect 442262 334778 477706 335334
rect 478262 334778 513706 335334
rect 514262 334778 549706 335334
rect 550262 334778 592062 335334
rect 592618 334778 592650 335334
rect -8726 334746 592650 334778
rect -8726 334094 592650 334126
rect -8726 333538 -7734 334094
rect -7178 333538 8466 334094
rect 9022 333538 44466 334094
rect 45022 333538 80466 334094
rect 81022 333538 116466 334094
rect 117022 333538 152466 334094
rect 153022 333538 188466 334094
rect 189022 333538 224466 334094
rect 225022 333538 260466 334094
rect 261022 333538 296466 334094
rect 297022 333538 332466 334094
rect 333022 333538 368466 334094
rect 369022 333538 404466 334094
rect 405022 333538 440466 334094
rect 441022 333538 476466 334094
rect 477022 333538 512466 334094
rect 513022 333538 548466 334094
rect 549022 333538 591102 334094
rect 591658 333538 592650 334094
rect -8726 333506 592650 333538
rect -8726 332854 592650 332886
rect -8726 332298 -6774 332854
rect -6218 332298 7226 332854
rect 7782 332298 43226 332854
rect 43782 332298 79226 332854
rect 79782 332298 115226 332854
rect 115782 332298 151226 332854
rect 151782 332298 187226 332854
rect 187782 332298 223226 332854
rect 223782 332298 259226 332854
rect 259782 332298 295226 332854
rect 295782 332298 331226 332854
rect 331782 332298 367226 332854
rect 367782 332298 403226 332854
rect 403782 332298 439226 332854
rect 439782 332298 475226 332854
rect 475782 332298 511226 332854
rect 511782 332298 547226 332854
rect 547782 332298 590142 332854
rect 590698 332298 592650 332854
rect -8726 332266 592650 332298
rect -8726 331614 592650 331646
rect -8726 331058 -5814 331614
rect -5258 331058 5986 331614
rect 6542 331058 41986 331614
rect 42542 331058 77986 331614
rect 78542 331058 113986 331614
rect 114542 331058 149986 331614
rect 150542 331058 185986 331614
rect 186542 331058 221986 331614
rect 222542 331058 257986 331614
rect 258542 331058 293986 331614
rect 294542 331058 329986 331614
rect 330542 331058 365986 331614
rect 366542 331058 401986 331614
rect 402542 331058 437986 331614
rect 438542 331058 473986 331614
rect 474542 331058 509986 331614
rect 510542 331058 581986 331614
rect 582542 331058 589182 331614
rect 589738 331058 592650 331614
rect -8726 331026 592650 331058
rect -8726 330374 592650 330406
rect -8726 329818 -4854 330374
rect -4298 329818 4746 330374
rect 5302 329818 40746 330374
rect 41302 329818 76746 330374
rect 77302 329818 112746 330374
rect 113302 329818 148746 330374
rect 149302 329818 184746 330374
rect 185302 329818 220746 330374
rect 221302 329818 256746 330374
rect 257302 329818 292746 330374
rect 293302 329818 328746 330374
rect 329302 329818 364746 330374
rect 365302 329818 400746 330374
rect 401302 329818 436746 330374
rect 437302 329818 472746 330374
rect 473302 329818 508746 330374
rect 509302 329818 580746 330374
rect 581302 329818 588222 330374
rect 588778 329818 592650 330374
rect -8726 329786 592650 329818
rect -8726 329134 592650 329166
rect -8726 328578 -3894 329134
rect -3338 328578 3506 329134
rect 4062 328578 39506 329134
rect 40062 328578 75506 329134
rect 76062 328578 111506 329134
rect 112062 328578 147506 329134
rect 148062 328578 183506 329134
rect 184062 328578 219506 329134
rect 220062 328578 255506 329134
rect 256062 328578 291506 329134
rect 292062 328578 327506 329134
rect 328062 328578 363506 329134
rect 364062 328578 399506 329134
rect 400062 328578 435506 329134
rect 436062 328578 471506 329134
rect 472062 328578 507506 329134
rect 508062 328578 579506 329134
rect 580062 328578 587262 329134
rect 587818 328578 592650 329134
rect -8726 328546 592650 328578
rect -8726 327894 592650 327926
rect -8726 327338 -2934 327894
rect -2378 327338 2266 327894
rect 2822 327338 38266 327894
rect 38822 327338 74266 327894
rect 74822 327338 110266 327894
rect 110822 327338 146266 327894
rect 146822 327338 182266 327894
rect 182822 327338 218266 327894
rect 218822 327338 254266 327894
rect 254822 327338 290266 327894
rect 290822 327338 326266 327894
rect 326822 327338 362266 327894
rect 362822 327338 398266 327894
rect 398822 327338 434266 327894
rect 434822 327338 470266 327894
rect 470822 327338 506266 327894
rect 506822 327658 540918 327894
rect 541154 327658 542850 327894
rect 543086 327658 544782 327894
rect 545018 327658 546714 327894
rect 546950 327658 578266 327894
rect 506822 327574 578266 327658
rect 506822 327338 540918 327574
rect 541154 327338 542850 327574
rect 543086 327338 544782 327574
rect 545018 327338 546714 327574
rect 546950 327338 578266 327574
rect 578822 327338 586302 327894
rect 586858 327338 592650 327894
rect -8726 327306 592650 327338
rect -8726 326654 592650 326686
rect -8726 326098 -1974 326654
rect -1418 326098 1026 326654
rect 1582 326098 37026 326654
rect 37582 326098 73026 326654
rect 73582 326098 109026 326654
rect 109582 326098 145026 326654
rect 145582 326098 181026 326654
rect 181582 326098 217026 326654
rect 217582 326098 253026 326654
rect 253582 326098 289026 326654
rect 289582 326098 325026 326654
rect 325582 326098 361026 326654
rect 361582 326098 397026 326654
rect 397582 326098 433026 326654
rect 433582 326098 469026 326654
rect 469582 326098 505026 326654
rect 505582 326418 539952 326654
rect 540188 326418 541884 326654
rect 542120 326418 543816 326654
rect 544052 326418 545748 326654
rect 545984 326418 577026 326654
rect 505582 326334 577026 326418
rect 505582 326098 539952 326334
rect 540188 326098 541884 326334
rect 542120 326098 543816 326334
rect 544052 326098 545748 326334
rect 545984 326098 577026 326334
rect 577582 326098 585342 326654
rect 585898 326098 592650 326654
rect -8726 326066 592650 326098
rect -8726 299334 592650 299366
rect -8726 298778 -8694 299334
rect -8138 298778 9706 299334
rect 10262 298778 45706 299334
rect 46262 298778 81706 299334
rect 82262 298778 117706 299334
rect 118262 298778 153706 299334
rect 154262 298778 189706 299334
rect 190262 298778 225706 299334
rect 226262 298778 261706 299334
rect 262262 298778 297706 299334
rect 298262 298778 333706 299334
rect 334262 298778 369706 299334
rect 370262 298778 405706 299334
rect 406262 298778 441706 299334
rect 442262 298778 477706 299334
rect 478262 298778 513706 299334
rect 514262 298778 549706 299334
rect 550262 298778 592062 299334
rect 592618 298778 592650 299334
rect -8726 298746 592650 298778
rect -8726 298094 592650 298126
rect -8726 297538 -7734 298094
rect -7178 297538 8466 298094
rect 9022 297538 44466 298094
rect 45022 297538 80466 298094
rect 81022 297538 116466 298094
rect 117022 297538 152466 298094
rect 153022 297538 188466 298094
rect 189022 297538 224466 298094
rect 225022 297538 260466 298094
rect 261022 297538 296466 298094
rect 297022 297538 332466 298094
rect 333022 297538 368466 298094
rect 369022 297538 404466 298094
rect 405022 297538 440466 298094
rect 441022 297538 476466 298094
rect 477022 297538 512466 298094
rect 513022 297538 548466 298094
rect 549022 297538 591102 298094
rect 591658 297538 592650 298094
rect -8726 297506 592650 297538
rect -8726 296854 592650 296886
rect -8726 296298 -6774 296854
rect -6218 296298 7226 296854
rect 7782 296298 43226 296854
rect 43782 296298 79226 296854
rect 79782 296298 115226 296854
rect 115782 296298 151226 296854
rect 151782 296298 187226 296854
rect 187782 296298 223226 296854
rect 223782 296298 259226 296854
rect 259782 296298 295226 296854
rect 295782 296298 331226 296854
rect 331782 296298 367226 296854
rect 367782 296298 403226 296854
rect 403782 296298 439226 296854
rect 439782 296298 475226 296854
rect 475782 296298 511226 296854
rect 511782 296298 547226 296854
rect 547782 296298 590142 296854
rect 590698 296298 592650 296854
rect -8726 296266 592650 296298
rect -8726 295614 592650 295646
rect -8726 295058 -5814 295614
rect -5258 295058 5986 295614
rect 6542 295058 41986 295614
rect 42542 295058 77986 295614
rect 78542 295058 113986 295614
rect 114542 295058 149986 295614
rect 150542 295058 185986 295614
rect 186542 295058 221986 295614
rect 222542 295058 257986 295614
rect 258542 295058 293986 295614
rect 294542 295058 329986 295614
rect 330542 295058 365986 295614
rect 366542 295058 401986 295614
rect 402542 295058 437986 295614
rect 438542 295058 473986 295614
rect 474542 295058 509986 295614
rect 510542 295058 581986 295614
rect 582542 295058 589182 295614
rect 589738 295058 592650 295614
rect -8726 295026 592650 295058
rect -8726 294374 592650 294406
rect -8726 293818 -4854 294374
rect -4298 293818 4746 294374
rect 5302 293818 40746 294374
rect 41302 293818 76746 294374
rect 77302 293818 112746 294374
rect 113302 293818 148746 294374
rect 149302 293818 184746 294374
rect 185302 293818 220746 294374
rect 221302 293818 256746 294374
rect 257302 293818 292746 294374
rect 293302 293818 328746 294374
rect 329302 293818 364746 294374
rect 365302 293818 400746 294374
rect 401302 293818 436746 294374
rect 437302 293818 472746 294374
rect 473302 293818 508746 294374
rect 509302 293818 580746 294374
rect 581302 293818 588222 294374
rect 588778 293818 592650 294374
rect -8726 293786 592650 293818
rect -8726 293134 592650 293166
rect -8726 292578 -3894 293134
rect -3338 292578 3506 293134
rect 4062 292578 39506 293134
rect 40062 292578 75506 293134
rect 76062 292578 111506 293134
rect 112062 292578 147506 293134
rect 148062 292578 183506 293134
rect 184062 292578 219506 293134
rect 220062 292578 255506 293134
rect 256062 292578 291506 293134
rect 292062 292578 327506 293134
rect 328062 292578 363506 293134
rect 364062 292578 399506 293134
rect 400062 292578 435506 293134
rect 436062 292578 471506 293134
rect 472062 292578 507506 293134
rect 508062 292578 579506 293134
rect 580062 292578 587262 293134
rect 587818 292578 592650 293134
rect -8726 292546 592650 292578
rect -8726 291894 592650 291926
rect -8726 291338 -2934 291894
rect -2378 291338 2266 291894
rect 2822 291338 38266 291894
rect 38822 291338 74266 291894
rect 74822 291338 110266 291894
rect 110822 291338 146266 291894
rect 146822 291338 182266 291894
rect 182822 291338 218266 291894
rect 218822 291338 254266 291894
rect 254822 291338 290266 291894
rect 290822 291338 326266 291894
rect 326822 291338 362266 291894
rect 362822 291338 398266 291894
rect 398822 291338 434266 291894
rect 434822 291338 470266 291894
rect 470822 291338 506266 291894
rect 506822 291658 540918 291894
rect 541154 291658 542850 291894
rect 543086 291658 544782 291894
rect 545018 291658 546714 291894
rect 546950 291658 578266 291894
rect 506822 291574 578266 291658
rect 506822 291338 540918 291574
rect 541154 291338 542850 291574
rect 543086 291338 544782 291574
rect 545018 291338 546714 291574
rect 546950 291338 578266 291574
rect 578822 291338 586302 291894
rect 586858 291338 592650 291894
rect -8726 291306 592650 291338
rect -8726 290654 592650 290686
rect -8726 290098 -1974 290654
rect -1418 290098 1026 290654
rect 1582 290098 37026 290654
rect 37582 290098 73026 290654
rect 73582 290098 109026 290654
rect 109582 290098 145026 290654
rect 145582 290098 181026 290654
rect 181582 290098 217026 290654
rect 217582 290098 253026 290654
rect 253582 290098 289026 290654
rect 289582 290098 325026 290654
rect 325582 290098 361026 290654
rect 361582 290098 397026 290654
rect 397582 290098 433026 290654
rect 433582 290098 469026 290654
rect 469582 290098 505026 290654
rect 505582 290418 539952 290654
rect 540188 290418 541884 290654
rect 542120 290418 543816 290654
rect 544052 290418 545748 290654
rect 545984 290418 577026 290654
rect 505582 290334 577026 290418
rect 505582 290098 539952 290334
rect 540188 290098 541884 290334
rect 542120 290098 543816 290334
rect 544052 290098 545748 290334
rect 545984 290098 577026 290334
rect 577582 290098 585342 290654
rect 585898 290098 592650 290654
rect -8726 290066 592650 290098
rect -8726 263334 592650 263366
rect -8726 262778 -8694 263334
rect -8138 262778 9706 263334
rect 10262 262778 45706 263334
rect 46262 262778 81706 263334
rect 82262 262778 117706 263334
rect 118262 262778 153706 263334
rect 154262 262778 189706 263334
rect 190262 262778 225706 263334
rect 226262 262778 261706 263334
rect 262262 262778 297706 263334
rect 298262 262778 333706 263334
rect 334262 262778 369706 263334
rect 370262 262778 405706 263334
rect 406262 262778 441706 263334
rect 442262 262778 477706 263334
rect 478262 262778 513706 263334
rect 514262 262778 549706 263334
rect 550262 262778 592062 263334
rect 592618 262778 592650 263334
rect -8726 262746 592650 262778
rect -8726 262094 592650 262126
rect -8726 261538 -7734 262094
rect -7178 261538 8466 262094
rect 9022 261538 44466 262094
rect 45022 261538 80466 262094
rect 81022 261538 116466 262094
rect 117022 261538 152466 262094
rect 153022 261538 188466 262094
rect 189022 261538 224466 262094
rect 225022 261538 260466 262094
rect 261022 261538 296466 262094
rect 297022 261538 332466 262094
rect 333022 261538 368466 262094
rect 369022 261538 404466 262094
rect 405022 261538 440466 262094
rect 441022 261538 476466 262094
rect 477022 261538 512466 262094
rect 513022 261538 548466 262094
rect 549022 261538 591102 262094
rect 591658 261538 592650 262094
rect -8726 261506 592650 261538
rect -8726 260854 592650 260886
rect -8726 260298 -6774 260854
rect -6218 260298 7226 260854
rect 7782 260298 43226 260854
rect 43782 260298 79226 260854
rect 79782 260298 115226 260854
rect 115782 260298 151226 260854
rect 151782 260298 187226 260854
rect 187782 260298 223226 260854
rect 223782 260298 259226 260854
rect 259782 260298 295226 260854
rect 295782 260298 331226 260854
rect 331782 260298 367226 260854
rect 367782 260298 403226 260854
rect 403782 260298 439226 260854
rect 439782 260298 475226 260854
rect 475782 260298 511226 260854
rect 511782 260298 547226 260854
rect 547782 260298 590142 260854
rect 590698 260298 592650 260854
rect -8726 260266 592650 260298
rect -8726 259614 592650 259646
rect -8726 259058 -5814 259614
rect -5258 259058 5986 259614
rect 6542 259058 41986 259614
rect 42542 259058 77986 259614
rect 78542 259058 113986 259614
rect 114542 259058 149986 259614
rect 150542 259058 185986 259614
rect 186542 259058 221986 259614
rect 222542 259058 257986 259614
rect 258542 259058 293986 259614
rect 294542 259058 329986 259614
rect 330542 259058 365986 259614
rect 366542 259058 401986 259614
rect 402542 259058 437986 259614
rect 438542 259058 473986 259614
rect 474542 259058 509986 259614
rect 510542 259058 545986 259614
rect 546542 259058 581986 259614
rect 582542 259058 589182 259614
rect 589738 259058 592650 259614
rect -8726 259026 592650 259058
rect -8726 258374 592650 258406
rect -8726 257818 -4854 258374
rect -4298 257818 4746 258374
rect 5302 257818 40746 258374
rect 41302 257818 76746 258374
rect 77302 257818 112746 258374
rect 113302 257818 148746 258374
rect 149302 257818 184746 258374
rect 185302 257818 220746 258374
rect 221302 257818 256746 258374
rect 257302 257818 292746 258374
rect 293302 257818 328746 258374
rect 329302 257818 364746 258374
rect 365302 257818 400746 258374
rect 401302 257818 436746 258374
rect 437302 257818 472746 258374
rect 473302 257818 508746 258374
rect 509302 257818 544746 258374
rect 545302 257818 580746 258374
rect 581302 257818 588222 258374
rect 588778 257818 592650 258374
rect -8726 257786 592650 257818
rect -8726 257134 592650 257166
rect -8726 256578 -3894 257134
rect -3338 256578 3506 257134
rect 4062 256578 39506 257134
rect 40062 256578 75506 257134
rect 76062 256578 111506 257134
rect 112062 256578 147506 257134
rect 148062 256578 183506 257134
rect 184062 256578 219506 257134
rect 220062 256578 255506 257134
rect 256062 256578 291506 257134
rect 292062 256578 327506 257134
rect 328062 256578 363506 257134
rect 364062 256578 399506 257134
rect 400062 256578 435506 257134
rect 436062 256578 471506 257134
rect 472062 256578 507506 257134
rect 508062 256578 543506 257134
rect 544062 256578 579506 257134
rect 580062 256578 587262 257134
rect 587818 256578 592650 257134
rect -8726 256546 592650 256578
rect -8726 255894 592650 255926
rect -8726 255338 -2934 255894
rect -2378 255338 2266 255894
rect 2822 255338 38266 255894
rect 38822 255338 74266 255894
rect 74822 255338 110266 255894
rect 110822 255338 146266 255894
rect 146822 255338 182266 255894
rect 182822 255338 218266 255894
rect 218822 255338 254266 255894
rect 254822 255338 290266 255894
rect 290822 255338 326266 255894
rect 326822 255338 362266 255894
rect 362822 255338 398266 255894
rect 398822 255338 434266 255894
rect 434822 255338 470266 255894
rect 470822 255338 506266 255894
rect 506822 255338 542266 255894
rect 542822 255338 578266 255894
rect 578822 255338 586302 255894
rect 586858 255338 592650 255894
rect -8726 255306 592650 255338
rect -8726 254654 592650 254686
rect -8726 254098 -1974 254654
rect -1418 254098 1026 254654
rect 1582 254098 37026 254654
rect 37582 254098 73026 254654
rect 73582 254098 109026 254654
rect 109582 254098 145026 254654
rect 145582 254098 181026 254654
rect 181582 254098 217026 254654
rect 217582 254098 253026 254654
rect 253582 254098 289026 254654
rect 289582 254098 325026 254654
rect 325582 254098 361026 254654
rect 361582 254098 397026 254654
rect 397582 254098 433026 254654
rect 433582 254098 469026 254654
rect 469582 254098 505026 254654
rect 505582 254098 541026 254654
rect 541582 254098 577026 254654
rect 577582 254098 585342 254654
rect 585898 254098 592650 254654
rect -8726 254066 592650 254098
rect -8726 227334 592650 227366
rect -8726 226778 -8694 227334
rect -8138 226778 9706 227334
rect 10262 226778 45706 227334
rect 46262 226778 81706 227334
rect 82262 226778 117706 227334
rect 118262 226778 153706 227334
rect 154262 226778 189706 227334
rect 190262 226778 225706 227334
rect 226262 226778 261706 227334
rect 262262 226778 297706 227334
rect 298262 226778 333706 227334
rect 334262 226778 369706 227334
rect 370262 226778 405706 227334
rect 406262 226778 441706 227334
rect 442262 226778 477706 227334
rect 478262 226778 513706 227334
rect 514262 226778 549706 227334
rect 550262 226778 592062 227334
rect 592618 226778 592650 227334
rect -8726 226746 592650 226778
rect -8726 226094 592650 226126
rect -8726 225538 -7734 226094
rect -7178 225538 8466 226094
rect 9022 225538 44466 226094
rect 45022 225538 80466 226094
rect 81022 225538 116466 226094
rect 117022 225538 152466 226094
rect 153022 225538 188466 226094
rect 189022 225538 224466 226094
rect 225022 225538 260466 226094
rect 261022 225538 296466 226094
rect 297022 225538 332466 226094
rect 333022 225538 368466 226094
rect 369022 225538 404466 226094
rect 405022 225538 440466 226094
rect 441022 225538 476466 226094
rect 477022 225538 512466 226094
rect 513022 225538 548466 226094
rect 549022 225538 591102 226094
rect 591658 225538 592650 226094
rect -8726 225506 592650 225538
rect -8726 224854 592650 224886
rect -8726 224298 -6774 224854
rect -6218 224298 7226 224854
rect 7782 224298 43226 224854
rect 43782 224298 79226 224854
rect 79782 224298 115226 224854
rect 115782 224298 151226 224854
rect 151782 224298 187226 224854
rect 187782 224298 223226 224854
rect 223782 224298 259226 224854
rect 259782 224298 295226 224854
rect 295782 224298 331226 224854
rect 331782 224298 367226 224854
rect 367782 224298 403226 224854
rect 403782 224298 439226 224854
rect 439782 224298 475226 224854
rect 475782 224298 511226 224854
rect 511782 224298 547226 224854
rect 547782 224298 590142 224854
rect 590698 224298 592650 224854
rect -8726 224266 592650 224298
rect -8726 223614 592650 223646
rect -8726 223058 -5814 223614
rect -5258 223058 5986 223614
rect 6542 223058 41986 223614
rect 42542 223058 77986 223614
rect 78542 223058 113986 223614
rect 114542 223058 149986 223614
rect 150542 223058 185986 223614
rect 186542 223058 221986 223614
rect 222542 223058 257986 223614
rect 258542 223058 293986 223614
rect 294542 223058 329986 223614
rect 330542 223058 365986 223614
rect 366542 223058 401986 223614
rect 402542 223058 437986 223614
rect 438542 223058 473986 223614
rect 474542 223058 509986 223614
rect 510542 223058 545986 223614
rect 546542 223058 581986 223614
rect 582542 223058 589182 223614
rect 589738 223058 592650 223614
rect -8726 223026 592650 223058
rect -8726 222374 592650 222406
rect -8726 221818 -4854 222374
rect -4298 221818 4746 222374
rect 5302 221818 40746 222374
rect 41302 221818 76746 222374
rect 77302 221818 112746 222374
rect 113302 221818 148746 222374
rect 149302 221818 184746 222374
rect 185302 221818 220746 222374
rect 221302 221818 256746 222374
rect 257302 221818 292746 222374
rect 293302 221818 328746 222374
rect 329302 221818 364746 222374
rect 365302 221818 400746 222374
rect 401302 221818 436746 222374
rect 437302 221818 472746 222374
rect 473302 221818 508746 222374
rect 509302 221818 544746 222374
rect 545302 221818 580746 222374
rect 581302 221818 588222 222374
rect 588778 221818 592650 222374
rect -8726 221786 592650 221818
rect -8726 221134 592650 221166
rect -8726 220578 -3894 221134
rect -3338 220578 3506 221134
rect 4062 220578 39506 221134
rect 40062 220578 75506 221134
rect 76062 220578 111506 221134
rect 112062 220578 147506 221134
rect 148062 220578 183506 221134
rect 184062 220578 219506 221134
rect 220062 220578 255506 221134
rect 256062 220578 291506 221134
rect 292062 220578 327506 221134
rect 328062 220578 363506 221134
rect 364062 220578 399506 221134
rect 400062 220578 435506 221134
rect 436062 220578 471506 221134
rect 472062 220578 507506 221134
rect 508062 220578 543506 221134
rect 544062 220578 579506 221134
rect 580062 220578 587262 221134
rect 587818 220578 592650 221134
rect -8726 220546 592650 220578
rect -8726 219894 592650 219926
rect -8726 219338 -2934 219894
rect -2378 219338 2266 219894
rect 2822 219338 38266 219894
rect 38822 219338 74266 219894
rect 74822 219338 110266 219894
rect 110822 219338 146266 219894
rect 146822 219338 182266 219894
rect 182822 219338 218266 219894
rect 218822 219338 254266 219894
rect 254822 219338 290266 219894
rect 290822 219338 326266 219894
rect 326822 219338 362266 219894
rect 362822 219338 398266 219894
rect 398822 219338 434266 219894
rect 434822 219338 470266 219894
rect 470822 219338 506266 219894
rect 506822 219338 542266 219894
rect 542822 219338 578266 219894
rect 578822 219338 586302 219894
rect 586858 219338 592650 219894
rect -8726 219306 592650 219338
rect -8726 218654 592650 218686
rect -8726 218098 -1974 218654
rect -1418 218098 1026 218654
rect 1582 218098 37026 218654
rect 37582 218098 73026 218654
rect 73582 218098 109026 218654
rect 109582 218098 145026 218654
rect 145582 218098 181026 218654
rect 181582 218098 217026 218654
rect 217582 218098 253026 218654
rect 253582 218098 289026 218654
rect 289582 218098 325026 218654
rect 325582 218098 361026 218654
rect 361582 218098 397026 218654
rect 397582 218098 433026 218654
rect 433582 218098 469026 218654
rect 469582 218098 505026 218654
rect 505582 218098 541026 218654
rect 541582 218098 577026 218654
rect 577582 218098 585342 218654
rect 585898 218098 592650 218654
rect -8726 218066 592650 218098
rect -8726 191334 592650 191366
rect -8726 190778 -8694 191334
rect -8138 190778 9706 191334
rect 10262 190778 45706 191334
rect 46262 190778 81706 191334
rect 82262 190778 117706 191334
rect 118262 190778 153706 191334
rect 154262 190778 189706 191334
rect 190262 190778 225706 191334
rect 226262 190778 261706 191334
rect 262262 190778 297706 191334
rect 298262 190778 333706 191334
rect 334262 190778 369706 191334
rect 370262 190778 405706 191334
rect 406262 190778 441706 191334
rect 442262 190778 477706 191334
rect 478262 190778 513706 191334
rect 514262 190778 549706 191334
rect 550262 190778 592062 191334
rect 592618 190778 592650 191334
rect -8726 190746 592650 190778
rect -8726 190094 592650 190126
rect -8726 189538 -7734 190094
rect -7178 189538 8466 190094
rect 9022 189538 44466 190094
rect 45022 189538 80466 190094
rect 81022 189538 116466 190094
rect 117022 189538 152466 190094
rect 153022 189538 188466 190094
rect 189022 189538 224466 190094
rect 225022 189538 260466 190094
rect 261022 189538 296466 190094
rect 297022 189538 332466 190094
rect 333022 189538 368466 190094
rect 369022 189538 404466 190094
rect 405022 189538 440466 190094
rect 441022 189538 476466 190094
rect 477022 189538 512466 190094
rect 513022 189538 548466 190094
rect 549022 189538 591102 190094
rect 591658 189538 592650 190094
rect -8726 189506 592650 189538
rect -8726 188854 592650 188886
rect -8726 188298 -6774 188854
rect -6218 188298 7226 188854
rect 7782 188298 43226 188854
rect 43782 188298 79226 188854
rect 79782 188298 115226 188854
rect 115782 188298 151226 188854
rect 151782 188298 187226 188854
rect 187782 188298 223226 188854
rect 223782 188298 259226 188854
rect 259782 188298 295226 188854
rect 295782 188298 331226 188854
rect 331782 188298 367226 188854
rect 367782 188298 403226 188854
rect 403782 188298 439226 188854
rect 439782 188298 475226 188854
rect 475782 188298 511226 188854
rect 511782 188298 547226 188854
rect 547782 188298 590142 188854
rect 590698 188298 592650 188854
rect -8726 188266 592650 188298
rect -8726 187614 592650 187646
rect -8726 187058 -5814 187614
rect -5258 187058 5986 187614
rect 6542 187058 41986 187614
rect 42542 187058 77986 187614
rect 78542 187058 113986 187614
rect 114542 187058 149986 187614
rect 150542 187058 185986 187614
rect 186542 187058 221986 187614
rect 222542 187058 257986 187614
rect 258542 187058 293986 187614
rect 294542 187058 329986 187614
rect 330542 187058 365986 187614
rect 366542 187058 401986 187614
rect 402542 187058 437986 187614
rect 438542 187058 473986 187614
rect 474542 187058 509986 187614
rect 510542 187058 545986 187614
rect 546542 187058 581986 187614
rect 582542 187058 589182 187614
rect 589738 187058 592650 187614
rect -8726 187026 592650 187058
rect -8726 186374 592650 186406
rect -8726 185818 -4854 186374
rect -4298 185818 4746 186374
rect 5302 185818 40746 186374
rect 41302 185818 76746 186374
rect 77302 185818 112746 186374
rect 113302 185818 148746 186374
rect 149302 185818 184746 186374
rect 185302 185818 220746 186374
rect 221302 185818 256746 186374
rect 257302 185818 292746 186374
rect 293302 185818 328746 186374
rect 329302 185818 364746 186374
rect 365302 185818 400746 186374
rect 401302 185818 436746 186374
rect 437302 185818 472746 186374
rect 473302 185818 508746 186374
rect 509302 185818 544746 186374
rect 545302 185818 580746 186374
rect 581302 185818 588222 186374
rect 588778 185818 592650 186374
rect -8726 185786 592650 185818
rect -8726 185134 592650 185166
rect -8726 184578 -3894 185134
rect -3338 184578 3506 185134
rect 4062 184578 39506 185134
rect 40062 184578 75506 185134
rect 76062 184578 111506 185134
rect 112062 184578 147506 185134
rect 148062 184578 183506 185134
rect 184062 184578 219506 185134
rect 220062 184578 255506 185134
rect 256062 184578 291506 185134
rect 292062 184578 327506 185134
rect 328062 184578 363506 185134
rect 364062 184578 399506 185134
rect 400062 184578 435506 185134
rect 436062 184578 471506 185134
rect 472062 184578 507506 185134
rect 508062 184578 543506 185134
rect 544062 184578 579506 185134
rect 580062 184578 587262 185134
rect 587818 184578 592650 185134
rect -8726 184546 592650 184578
rect -8726 183894 592650 183926
rect -8726 183338 -2934 183894
rect -2378 183338 2266 183894
rect 2822 183338 38266 183894
rect 38822 183338 74266 183894
rect 74822 183338 110266 183894
rect 110822 183338 146266 183894
rect 146822 183338 182266 183894
rect 182822 183338 218266 183894
rect 218822 183338 254266 183894
rect 254822 183338 290266 183894
rect 290822 183338 326266 183894
rect 326822 183338 362266 183894
rect 362822 183338 398266 183894
rect 398822 183338 434266 183894
rect 434822 183338 470266 183894
rect 470822 183338 506266 183894
rect 506822 183338 542266 183894
rect 542822 183338 578266 183894
rect 578822 183338 586302 183894
rect 586858 183338 592650 183894
rect -8726 183306 592650 183338
rect -8726 182654 592650 182686
rect -8726 182098 -1974 182654
rect -1418 182098 1026 182654
rect 1582 182098 37026 182654
rect 37582 182098 73026 182654
rect 73582 182098 109026 182654
rect 109582 182098 145026 182654
rect 145582 182098 181026 182654
rect 181582 182098 217026 182654
rect 217582 182098 253026 182654
rect 253582 182098 289026 182654
rect 289582 182098 325026 182654
rect 325582 182098 361026 182654
rect 361582 182098 397026 182654
rect 397582 182098 433026 182654
rect 433582 182098 469026 182654
rect 469582 182098 505026 182654
rect 505582 182098 541026 182654
rect 541582 182098 577026 182654
rect 577582 182098 585342 182654
rect 585898 182098 592650 182654
rect -8726 182066 592650 182098
rect -8726 155334 592650 155366
rect -8726 154778 -8694 155334
rect -8138 154778 9706 155334
rect 10262 154778 45706 155334
rect 46262 154778 81706 155334
rect 82262 154778 117706 155334
rect 118262 154778 153706 155334
rect 154262 154778 189706 155334
rect 190262 154778 225706 155334
rect 226262 154778 261706 155334
rect 262262 154778 297706 155334
rect 298262 154778 333706 155334
rect 334262 154778 369706 155334
rect 370262 154778 405706 155334
rect 406262 154778 441706 155334
rect 442262 154778 477706 155334
rect 478262 154778 513706 155334
rect 514262 154778 549706 155334
rect 550262 154778 592062 155334
rect 592618 154778 592650 155334
rect -8726 154746 592650 154778
rect -8726 154094 592650 154126
rect -8726 153538 -7734 154094
rect -7178 153538 8466 154094
rect 9022 153538 44466 154094
rect 45022 153538 80466 154094
rect 81022 153538 116466 154094
rect 117022 153538 152466 154094
rect 153022 153538 188466 154094
rect 189022 153538 224466 154094
rect 225022 153538 260466 154094
rect 261022 153538 296466 154094
rect 297022 153538 332466 154094
rect 333022 153538 368466 154094
rect 369022 153538 404466 154094
rect 405022 153538 440466 154094
rect 441022 153538 476466 154094
rect 477022 153538 512466 154094
rect 513022 153538 548466 154094
rect 549022 153538 591102 154094
rect 591658 153538 592650 154094
rect -8726 153506 592650 153538
rect -8726 152854 592650 152886
rect -8726 152298 -6774 152854
rect -6218 152298 7226 152854
rect 7782 152298 43226 152854
rect 43782 152298 79226 152854
rect 79782 152298 115226 152854
rect 115782 152298 151226 152854
rect 151782 152298 187226 152854
rect 187782 152298 223226 152854
rect 223782 152298 259226 152854
rect 259782 152298 295226 152854
rect 295782 152298 331226 152854
rect 331782 152298 367226 152854
rect 367782 152298 403226 152854
rect 403782 152298 439226 152854
rect 439782 152298 475226 152854
rect 475782 152298 511226 152854
rect 511782 152298 547226 152854
rect 547782 152298 590142 152854
rect 590698 152298 592650 152854
rect -8726 152266 592650 152298
rect -8726 151614 592650 151646
rect -8726 151058 -5814 151614
rect -5258 151058 5986 151614
rect 6542 151058 41986 151614
rect 42542 151058 77986 151614
rect 78542 151058 113986 151614
rect 114542 151058 149986 151614
rect 150542 151058 185986 151614
rect 186542 151058 221986 151614
rect 222542 151058 257986 151614
rect 258542 151058 293986 151614
rect 294542 151058 329986 151614
rect 330542 151058 365986 151614
rect 366542 151058 401986 151614
rect 402542 151058 437986 151614
rect 438542 151058 473986 151614
rect 474542 151058 509986 151614
rect 510542 151058 545986 151614
rect 546542 151058 581986 151614
rect 582542 151058 589182 151614
rect 589738 151058 592650 151614
rect -8726 151026 592650 151058
rect -8726 150374 592650 150406
rect -8726 149818 -4854 150374
rect -4298 149818 4746 150374
rect 5302 149818 40746 150374
rect 41302 149818 76746 150374
rect 77302 149818 112746 150374
rect 113302 149818 148746 150374
rect 149302 149818 184746 150374
rect 185302 149818 220746 150374
rect 221302 149818 256746 150374
rect 257302 149818 292746 150374
rect 293302 149818 328746 150374
rect 329302 149818 364746 150374
rect 365302 149818 400746 150374
rect 401302 149818 436746 150374
rect 437302 149818 472746 150374
rect 473302 149818 508746 150374
rect 509302 149818 544746 150374
rect 545302 149818 580746 150374
rect 581302 149818 588222 150374
rect 588778 149818 592650 150374
rect -8726 149786 592650 149818
rect -8726 149134 592650 149166
rect -8726 148578 -3894 149134
rect -3338 148578 3506 149134
rect 4062 148578 39506 149134
rect 40062 148578 75506 149134
rect 76062 148578 111506 149134
rect 112062 148578 147506 149134
rect 148062 148578 183506 149134
rect 184062 148578 219506 149134
rect 220062 148578 255506 149134
rect 256062 148578 291506 149134
rect 292062 148578 327506 149134
rect 328062 148578 363506 149134
rect 364062 148578 399506 149134
rect 400062 148578 435506 149134
rect 436062 148578 471506 149134
rect 472062 148578 507506 149134
rect 508062 148578 543506 149134
rect 544062 148578 579506 149134
rect 580062 148578 587262 149134
rect 587818 148578 592650 149134
rect -8726 148546 592650 148578
rect -8726 147894 592650 147926
rect -8726 147338 -2934 147894
rect -2378 147338 2266 147894
rect 2822 147338 38266 147894
rect 38822 147338 74266 147894
rect 74822 147338 110266 147894
rect 110822 147338 146266 147894
rect 146822 147338 182266 147894
rect 182822 147338 218266 147894
rect 218822 147338 254266 147894
rect 254822 147338 290266 147894
rect 290822 147338 326266 147894
rect 326822 147338 362266 147894
rect 362822 147338 398266 147894
rect 398822 147338 434266 147894
rect 434822 147338 470266 147894
rect 470822 147338 506266 147894
rect 506822 147338 542266 147894
rect 542822 147338 578266 147894
rect 578822 147338 586302 147894
rect 586858 147338 592650 147894
rect -8726 147306 592650 147338
rect -8726 146654 592650 146686
rect -8726 146098 -1974 146654
rect -1418 146098 1026 146654
rect 1582 146098 37026 146654
rect 37582 146098 73026 146654
rect 73582 146098 109026 146654
rect 109582 146098 145026 146654
rect 145582 146098 181026 146654
rect 181582 146098 217026 146654
rect 217582 146098 253026 146654
rect 253582 146098 289026 146654
rect 289582 146098 325026 146654
rect 325582 146098 361026 146654
rect 361582 146098 397026 146654
rect 397582 146098 433026 146654
rect 433582 146098 469026 146654
rect 469582 146098 505026 146654
rect 505582 146098 541026 146654
rect 541582 146098 577026 146654
rect 577582 146098 585342 146654
rect 585898 146098 592650 146654
rect -8726 146066 592650 146098
rect -8726 119334 592650 119366
rect -8726 118778 -8694 119334
rect -8138 118778 9706 119334
rect 10262 118778 45706 119334
rect 46262 118778 81706 119334
rect 82262 118778 117706 119334
rect 118262 118778 153706 119334
rect 154262 118778 189706 119334
rect 190262 118778 225706 119334
rect 226262 118778 261706 119334
rect 262262 118778 297706 119334
rect 298262 118778 333706 119334
rect 334262 118778 369706 119334
rect 370262 118778 405706 119334
rect 406262 118778 441706 119334
rect 442262 118778 477706 119334
rect 478262 118778 513706 119334
rect 514262 118778 549706 119334
rect 550262 118778 592062 119334
rect 592618 118778 592650 119334
rect -8726 118746 592650 118778
rect -8726 118094 592650 118126
rect -8726 117538 -7734 118094
rect -7178 117538 8466 118094
rect 9022 117538 44466 118094
rect 45022 117538 80466 118094
rect 81022 117538 116466 118094
rect 117022 117538 152466 118094
rect 153022 117538 188466 118094
rect 189022 117538 224466 118094
rect 225022 117538 260466 118094
rect 261022 117538 296466 118094
rect 297022 117538 332466 118094
rect 333022 117538 368466 118094
rect 369022 117538 404466 118094
rect 405022 117538 440466 118094
rect 441022 117538 476466 118094
rect 477022 117538 512466 118094
rect 513022 117538 548466 118094
rect 549022 117538 591102 118094
rect 591658 117538 592650 118094
rect -8726 117506 592650 117538
rect -8726 116854 592650 116886
rect -8726 116298 -6774 116854
rect -6218 116298 7226 116854
rect 7782 116298 43226 116854
rect 43782 116298 79226 116854
rect 79782 116298 115226 116854
rect 115782 116298 151226 116854
rect 151782 116298 187226 116854
rect 187782 116298 223226 116854
rect 223782 116298 259226 116854
rect 259782 116298 295226 116854
rect 295782 116298 331226 116854
rect 331782 116298 367226 116854
rect 367782 116298 403226 116854
rect 403782 116298 439226 116854
rect 439782 116298 475226 116854
rect 475782 116298 511226 116854
rect 511782 116298 547226 116854
rect 547782 116298 590142 116854
rect 590698 116298 592650 116854
rect -8726 116266 592650 116298
rect -8726 115614 592650 115646
rect -8726 115058 -5814 115614
rect -5258 115058 5986 115614
rect 6542 115058 41986 115614
rect 42542 115058 77986 115614
rect 78542 115058 113986 115614
rect 114542 115058 149986 115614
rect 150542 115058 185986 115614
rect 186542 115058 221986 115614
rect 222542 115058 257986 115614
rect 258542 115058 293986 115614
rect 294542 115058 329986 115614
rect 330542 115058 365986 115614
rect 366542 115058 401986 115614
rect 402542 115058 437986 115614
rect 438542 115058 473986 115614
rect 474542 115058 509986 115614
rect 510542 115058 545986 115614
rect 546542 115058 581986 115614
rect 582542 115058 589182 115614
rect 589738 115058 592650 115614
rect -8726 115026 592650 115058
rect -8726 114374 592650 114406
rect -8726 113818 -4854 114374
rect -4298 113818 4746 114374
rect 5302 113818 40746 114374
rect 41302 113818 76746 114374
rect 77302 113818 112746 114374
rect 113302 113818 148746 114374
rect 149302 113818 184746 114374
rect 185302 113818 220746 114374
rect 221302 113818 256746 114374
rect 257302 113818 292746 114374
rect 293302 113818 328746 114374
rect 329302 113818 364746 114374
rect 365302 113818 400746 114374
rect 401302 113818 436746 114374
rect 437302 113818 472746 114374
rect 473302 113818 508746 114374
rect 509302 113818 544746 114374
rect 545302 113818 580746 114374
rect 581302 113818 588222 114374
rect 588778 113818 592650 114374
rect -8726 113786 592650 113818
rect -8726 113134 592650 113166
rect -8726 112578 -3894 113134
rect -3338 112578 3506 113134
rect 4062 112578 39506 113134
rect 40062 112578 75506 113134
rect 76062 112578 111506 113134
rect 112062 112578 147506 113134
rect 148062 112578 183506 113134
rect 184062 112578 219506 113134
rect 220062 112578 255506 113134
rect 256062 112578 291506 113134
rect 292062 112578 327506 113134
rect 328062 112578 363506 113134
rect 364062 112578 399506 113134
rect 400062 112578 435506 113134
rect 436062 112578 471506 113134
rect 472062 112578 507506 113134
rect 508062 112578 543506 113134
rect 544062 112578 579506 113134
rect 580062 112578 587262 113134
rect 587818 112578 592650 113134
rect -8726 112546 592650 112578
rect -8726 111894 592650 111926
rect -8726 111338 -2934 111894
rect -2378 111338 2266 111894
rect 2822 111338 38266 111894
rect 38822 111338 74266 111894
rect 74822 111338 110266 111894
rect 110822 111338 146266 111894
rect 146822 111338 182266 111894
rect 182822 111338 218266 111894
rect 218822 111338 254266 111894
rect 254822 111338 290266 111894
rect 290822 111338 326266 111894
rect 326822 111338 362266 111894
rect 362822 111338 398266 111894
rect 398822 111338 434266 111894
rect 434822 111338 470266 111894
rect 470822 111338 506266 111894
rect 506822 111338 542266 111894
rect 542822 111338 578266 111894
rect 578822 111338 586302 111894
rect 586858 111338 592650 111894
rect -8726 111306 592650 111338
rect -8726 110654 592650 110686
rect -8726 110098 -1974 110654
rect -1418 110098 1026 110654
rect 1582 110098 37026 110654
rect 37582 110098 73026 110654
rect 73582 110098 109026 110654
rect 109582 110098 145026 110654
rect 145582 110098 181026 110654
rect 181582 110098 217026 110654
rect 217582 110098 253026 110654
rect 253582 110098 289026 110654
rect 289582 110098 325026 110654
rect 325582 110098 361026 110654
rect 361582 110098 397026 110654
rect 397582 110098 433026 110654
rect 433582 110098 469026 110654
rect 469582 110098 505026 110654
rect 505582 110098 541026 110654
rect 541582 110098 577026 110654
rect 577582 110098 585342 110654
rect 585898 110098 592650 110654
rect -8726 110066 592650 110098
rect -8726 83334 592650 83366
rect -8726 82778 -8694 83334
rect -8138 82778 9706 83334
rect 10262 82778 45706 83334
rect 46262 82778 81706 83334
rect 82262 82778 117706 83334
rect 118262 82778 153706 83334
rect 154262 82778 189706 83334
rect 190262 82778 225706 83334
rect 226262 82778 261706 83334
rect 262262 82778 297706 83334
rect 298262 82778 333706 83334
rect 334262 82778 369706 83334
rect 370262 82778 405706 83334
rect 406262 82778 441706 83334
rect 442262 82778 477706 83334
rect 478262 82778 513706 83334
rect 514262 82778 549706 83334
rect 550262 82778 592062 83334
rect 592618 82778 592650 83334
rect -8726 82746 592650 82778
rect -8726 82094 592650 82126
rect -8726 81538 -7734 82094
rect -7178 81538 8466 82094
rect 9022 81538 44466 82094
rect 45022 81538 80466 82094
rect 81022 81538 116466 82094
rect 117022 81538 152466 82094
rect 153022 81538 188466 82094
rect 189022 81538 224466 82094
rect 225022 81538 260466 82094
rect 261022 81538 296466 82094
rect 297022 81538 332466 82094
rect 333022 81538 368466 82094
rect 369022 81538 404466 82094
rect 405022 81538 440466 82094
rect 441022 81538 476466 82094
rect 477022 81538 512466 82094
rect 513022 81538 548466 82094
rect 549022 81538 591102 82094
rect 591658 81538 592650 82094
rect -8726 81506 592650 81538
rect -8726 80854 592650 80886
rect -8726 80298 -6774 80854
rect -6218 80298 7226 80854
rect 7782 80298 43226 80854
rect 43782 80298 79226 80854
rect 79782 80298 115226 80854
rect 115782 80298 151226 80854
rect 151782 80298 187226 80854
rect 187782 80298 223226 80854
rect 223782 80298 259226 80854
rect 259782 80298 295226 80854
rect 295782 80298 331226 80854
rect 331782 80298 367226 80854
rect 367782 80298 403226 80854
rect 403782 80298 439226 80854
rect 439782 80298 475226 80854
rect 475782 80298 511226 80854
rect 511782 80298 547226 80854
rect 547782 80298 590142 80854
rect 590698 80298 592650 80854
rect -8726 80266 592650 80298
rect -8726 79614 592650 79646
rect -8726 79058 -5814 79614
rect -5258 79058 5986 79614
rect 6542 79058 41986 79614
rect 42542 79058 77986 79614
rect 78542 79058 113986 79614
rect 114542 79058 149986 79614
rect 150542 79058 185986 79614
rect 186542 79058 221986 79614
rect 222542 79058 257986 79614
rect 258542 79058 293986 79614
rect 294542 79058 329986 79614
rect 330542 79058 365986 79614
rect 366542 79058 401986 79614
rect 402542 79058 437986 79614
rect 438542 79058 473986 79614
rect 474542 79058 509986 79614
rect 510542 79058 545986 79614
rect 546542 79058 581986 79614
rect 582542 79058 589182 79614
rect 589738 79058 592650 79614
rect -8726 79026 592650 79058
rect -8726 78374 592650 78406
rect -8726 77818 -4854 78374
rect -4298 77818 4746 78374
rect 5302 77818 40746 78374
rect 41302 77818 76746 78374
rect 77302 77818 112746 78374
rect 113302 77818 148746 78374
rect 149302 77818 184746 78374
rect 185302 77818 220746 78374
rect 221302 77818 256746 78374
rect 257302 77818 292746 78374
rect 293302 77818 328746 78374
rect 329302 77818 364746 78374
rect 365302 77818 400746 78374
rect 401302 77818 436746 78374
rect 437302 77818 472746 78374
rect 473302 77818 508746 78374
rect 509302 77818 544746 78374
rect 545302 77818 580746 78374
rect 581302 77818 588222 78374
rect 588778 77818 592650 78374
rect -8726 77786 592650 77818
rect -8726 77134 592650 77166
rect -8726 76578 -3894 77134
rect -3338 76578 3506 77134
rect 4062 76578 39506 77134
rect 40062 76578 75506 77134
rect 76062 76578 111506 77134
rect 112062 76578 147506 77134
rect 148062 76578 183506 77134
rect 184062 76578 219506 77134
rect 220062 76578 255506 77134
rect 256062 76578 291506 77134
rect 292062 76578 327506 77134
rect 328062 76578 363506 77134
rect 364062 76578 399506 77134
rect 400062 76578 435506 77134
rect 436062 76578 471506 77134
rect 472062 76578 507506 77134
rect 508062 76578 543506 77134
rect 544062 76578 579506 77134
rect 580062 76578 587262 77134
rect 587818 76578 592650 77134
rect -8726 76546 592650 76578
rect -8726 75894 592650 75926
rect -8726 75338 -2934 75894
rect -2378 75338 2266 75894
rect 2822 75338 38266 75894
rect 38822 75338 74266 75894
rect 74822 75338 110266 75894
rect 110822 75338 146266 75894
rect 146822 75338 182266 75894
rect 182822 75338 218266 75894
rect 218822 75338 254266 75894
rect 254822 75338 290266 75894
rect 290822 75338 326266 75894
rect 326822 75338 362266 75894
rect 362822 75338 398266 75894
rect 398822 75338 434266 75894
rect 434822 75338 470266 75894
rect 470822 75338 506266 75894
rect 506822 75338 542266 75894
rect 542822 75338 578266 75894
rect 578822 75338 586302 75894
rect 586858 75338 592650 75894
rect -8726 75306 592650 75338
rect -8726 74654 592650 74686
rect -8726 74098 -1974 74654
rect -1418 74098 1026 74654
rect 1582 74098 37026 74654
rect 37582 74098 73026 74654
rect 73582 74098 109026 74654
rect 109582 74098 145026 74654
rect 145582 74098 181026 74654
rect 181582 74098 217026 74654
rect 217582 74098 253026 74654
rect 253582 74098 289026 74654
rect 289582 74098 325026 74654
rect 325582 74098 361026 74654
rect 361582 74098 397026 74654
rect 397582 74098 433026 74654
rect 433582 74098 469026 74654
rect 469582 74098 505026 74654
rect 505582 74098 541026 74654
rect 541582 74098 577026 74654
rect 577582 74098 585342 74654
rect 585898 74098 592650 74654
rect -8726 74066 592650 74098
rect -8726 47334 592650 47366
rect -8726 46778 -8694 47334
rect -8138 46778 9706 47334
rect 10262 46778 45706 47334
rect 46262 46778 81706 47334
rect 82262 46778 117706 47334
rect 118262 46778 153706 47334
rect 154262 46778 189706 47334
rect 190262 46778 225706 47334
rect 226262 46778 261706 47334
rect 262262 46778 297706 47334
rect 298262 46778 333706 47334
rect 334262 46778 369706 47334
rect 370262 46778 405706 47334
rect 406262 46778 441706 47334
rect 442262 46778 477706 47334
rect 478262 46778 513706 47334
rect 514262 46778 549706 47334
rect 550262 46778 592062 47334
rect 592618 46778 592650 47334
rect -8726 46746 592650 46778
rect -8726 46094 592650 46126
rect -8726 45538 -7734 46094
rect -7178 45538 8466 46094
rect 9022 45538 44466 46094
rect 45022 45538 80466 46094
rect 81022 45538 116466 46094
rect 117022 45538 152466 46094
rect 153022 45538 188466 46094
rect 189022 45538 224466 46094
rect 225022 45538 260466 46094
rect 261022 45538 296466 46094
rect 297022 45538 332466 46094
rect 333022 45538 368466 46094
rect 369022 45538 404466 46094
rect 405022 45538 440466 46094
rect 441022 45538 476466 46094
rect 477022 45538 512466 46094
rect 513022 45538 548466 46094
rect 549022 45538 591102 46094
rect 591658 45538 592650 46094
rect -8726 45506 592650 45538
rect -8726 44854 592650 44886
rect -8726 44298 -6774 44854
rect -6218 44298 7226 44854
rect 7782 44298 43226 44854
rect 43782 44298 79226 44854
rect 79782 44298 115226 44854
rect 115782 44298 151226 44854
rect 151782 44298 187226 44854
rect 187782 44298 223226 44854
rect 223782 44298 259226 44854
rect 259782 44298 295226 44854
rect 295782 44298 331226 44854
rect 331782 44298 367226 44854
rect 367782 44298 403226 44854
rect 403782 44298 439226 44854
rect 439782 44298 475226 44854
rect 475782 44298 511226 44854
rect 511782 44298 547226 44854
rect 547782 44298 590142 44854
rect 590698 44298 592650 44854
rect -8726 44266 592650 44298
rect -8726 43614 592650 43646
rect -8726 43058 -5814 43614
rect -5258 43058 5986 43614
rect 6542 43058 41986 43614
rect 42542 43058 77986 43614
rect 78542 43058 113986 43614
rect 114542 43058 149986 43614
rect 150542 43058 185986 43614
rect 186542 43058 221986 43614
rect 222542 43058 257986 43614
rect 258542 43058 293986 43614
rect 294542 43058 329986 43614
rect 330542 43058 365986 43614
rect 366542 43058 401986 43614
rect 402542 43058 437986 43614
rect 438542 43058 473986 43614
rect 474542 43058 509986 43614
rect 510542 43058 545986 43614
rect 546542 43058 581986 43614
rect 582542 43058 589182 43614
rect 589738 43058 592650 43614
rect -8726 43026 592650 43058
rect -8726 42374 592650 42406
rect -8726 41818 -4854 42374
rect -4298 41818 4746 42374
rect 5302 41818 40746 42374
rect 41302 41818 76746 42374
rect 77302 41818 112746 42374
rect 113302 41818 148746 42374
rect 149302 41818 184746 42374
rect 185302 41818 220746 42374
rect 221302 41818 256746 42374
rect 257302 41818 292746 42374
rect 293302 41818 328746 42374
rect 329302 41818 364746 42374
rect 365302 41818 400746 42374
rect 401302 41818 436746 42374
rect 437302 41818 472746 42374
rect 473302 41818 508746 42374
rect 509302 41818 544746 42374
rect 545302 41818 580746 42374
rect 581302 41818 588222 42374
rect 588778 41818 592650 42374
rect -8726 41786 592650 41818
rect -8726 41134 592650 41166
rect -8726 40578 -3894 41134
rect -3338 40578 3506 41134
rect 4062 40578 39506 41134
rect 40062 40578 75506 41134
rect 76062 40578 111506 41134
rect 112062 40578 147506 41134
rect 148062 40578 183506 41134
rect 184062 40578 219506 41134
rect 220062 40578 255506 41134
rect 256062 40578 291506 41134
rect 292062 40578 327506 41134
rect 328062 40578 363506 41134
rect 364062 40578 399506 41134
rect 400062 40578 435506 41134
rect 436062 40578 471506 41134
rect 472062 40578 507506 41134
rect 508062 40578 543506 41134
rect 544062 40578 579506 41134
rect 580062 40578 587262 41134
rect 587818 40578 592650 41134
rect -8726 40546 592650 40578
rect -8726 39894 592650 39926
rect -8726 39338 -2934 39894
rect -2378 39338 2266 39894
rect 2822 39338 38266 39894
rect 38822 39338 74266 39894
rect 74822 39338 110266 39894
rect 110822 39338 146266 39894
rect 146822 39338 182266 39894
rect 182822 39338 218266 39894
rect 218822 39338 254266 39894
rect 254822 39338 290266 39894
rect 290822 39338 326266 39894
rect 326822 39338 362266 39894
rect 362822 39338 398266 39894
rect 398822 39338 434266 39894
rect 434822 39338 470266 39894
rect 470822 39338 506266 39894
rect 506822 39338 542266 39894
rect 542822 39338 578266 39894
rect 578822 39338 586302 39894
rect 586858 39338 592650 39894
rect -8726 39306 592650 39338
rect -8726 38654 592650 38686
rect -8726 38098 -1974 38654
rect -1418 38098 1026 38654
rect 1582 38098 37026 38654
rect 37582 38098 73026 38654
rect 73582 38098 109026 38654
rect 109582 38098 145026 38654
rect 145582 38098 181026 38654
rect 181582 38098 217026 38654
rect 217582 38098 253026 38654
rect 253582 38098 289026 38654
rect 289582 38098 325026 38654
rect 325582 38098 361026 38654
rect 361582 38098 397026 38654
rect 397582 38098 433026 38654
rect 433582 38098 469026 38654
rect 469582 38098 505026 38654
rect 505582 38098 541026 38654
rect 541582 38098 577026 38654
rect 577582 38098 585342 38654
rect 585898 38098 592650 38654
rect -8726 38066 592650 38098
rect -8726 11334 592650 11366
rect -8726 10778 -8694 11334
rect -8138 10778 9706 11334
rect 10262 10778 45706 11334
rect 46262 10778 81706 11334
rect 82262 10778 117706 11334
rect 118262 10778 153706 11334
rect 154262 10778 189706 11334
rect 190262 10778 225706 11334
rect 226262 10778 261706 11334
rect 262262 10778 297706 11334
rect 298262 10778 333706 11334
rect 334262 10778 369706 11334
rect 370262 10778 405706 11334
rect 406262 10778 441706 11334
rect 442262 10778 477706 11334
rect 478262 10778 513706 11334
rect 514262 10778 549706 11334
rect 550262 10778 592062 11334
rect 592618 10778 592650 11334
rect -8726 10746 592650 10778
rect -8726 10094 592650 10126
rect -8726 9538 -7734 10094
rect -7178 9538 8466 10094
rect 9022 9538 44466 10094
rect 45022 9538 80466 10094
rect 81022 9538 116466 10094
rect 117022 9538 152466 10094
rect 153022 9538 188466 10094
rect 189022 9538 224466 10094
rect 225022 9538 260466 10094
rect 261022 9538 296466 10094
rect 297022 9538 332466 10094
rect 333022 9538 368466 10094
rect 369022 9538 404466 10094
rect 405022 9538 440466 10094
rect 441022 9538 476466 10094
rect 477022 9538 512466 10094
rect 513022 9538 548466 10094
rect 549022 9538 591102 10094
rect 591658 9538 592650 10094
rect -8726 9506 592650 9538
rect -8726 8854 592650 8886
rect -8726 8298 -6774 8854
rect -6218 8298 7226 8854
rect 7782 8298 43226 8854
rect 43782 8298 79226 8854
rect 79782 8298 115226 8854
rect 115782 8298 151226 8854
rect 151782 8298 187226 8854
rect 187782 8298 223226 8854
rect 223782 8298 259226 8854
rect 259782 8298 295226 8854
rect 295782 8298 331226 8854
rect 331782 8298 367226 8854
rect 367782 8298 403226 8854
rect 403782 8298 439226 8854
rect 439782 8298 475226 8854
rect 475782 8298 511226 8854
rect 511782 8298 547226 8854
rect 547782 8298 590142 8854
rect 590698 8298 592650 8854
rect -8726 8266 592650 8298
rect -8726 7614 592650 7646
rect -8726 7058 -5814 7614
rect -5258 7058 5986 7614
rect 6542 7058 41986 7614
rect 42542 7058 77986 7614
rect 78542 7058 113986 7614
rect 114542 7058 149986 7614
rect 150542 7058 185986 7614
rect 186542 7058 221986 7614
rect 222542 7058 257986 7614
rect 258542 7058 293986 7614
rect 294542 7058 329986 7614
rect 330542 7058 365986 7614
rect 366542 7058 401986 7614
rect 402542 7058 437986 7614
rect 438542 7058 473986 7614
rect 474542 7058 509986 7614
rect 510542 7058 545986 7614
rect 546542 7058 581986 7614
rect 582542 7058 589182 7614
rect 589738 7058 592650 7614
rect -8726 7026 592650 7058
rect -8726 6374 592650 6406
rect -8726 5818 -4854 6374
rect -4298 5818 4746 6374
rect 5302 5818 40746 6374
rect 41302 5818 76746 6374
rect 77302 5818 112746 6374
rect 113302 5818 148746 6374
rect 149302 5818 184746 6374
rect 185302 5818 220746 6374
rect 221302 5818 256746 6374
rect 257302 5818 292746 6374
rect 293302 5818 328746 6374
rect 329302 5818 364746 6374
rect 365302 5818 400746 6374
rect 401302 5818 436746 6374
rect 437302 5818 472746 6374
rect 473302 5818 508746 6374
rect 509302 5818 544746 6374
rect 545302 5818 580746 6374
rect 581302 5818 588222 6374
rect 588778 5818 592650 6374
rect -8726 5786 592650 5818
rect -8726 5134 592650 5166
rect -8726 4578 -3894 5134
rect -3338 4578 3506 5134
rect 4062 4578 39506 5134
rect 40062 4578 75506 5134
rect 76062 4578 111506 5134
rect 112062 4578 147506 5134
rect 148062 4578 183506 5134
rect 184062 4578 219506 5134
rect 220062 4578 255506 5134
rect 256062 4578 291506 5134
rect 292062 4578 327506 5134
rect 328062 4578 363506 5134
rect 364062 4578 399506 5134
rect 400062 4578 435506 5134
rect 436062 4578 471506 5134
rect 472062 4578 507506 5134
rect 508062 4578 543506 5134
rect 544062 4578 579506 5134
rect 580062 4578 587262 5134
rect 587818 4578 592650 5134
rect -8726 4546 592650 4578
rect -8726 3894 592650 3926
rect -8726 3338 -2934 3894
rect -2378 3338 2266 3894
rect 2822 3338 38266 3894
rect 38822 3338 74266 3894
rect 74822 3338 110266 3894
rect 110822 3338 146266 3894
rect 146822 3338 182266 3894
rect 182822 3338 218266 3894
rect 218822 3338 254266 3894
rect 254822 3338 290266 3894
rect 290822 3338 326266 3894
rect 326822 3338 362266 3894
rect 362822 3338 398266 3894
rect 398822 3338 434266 3894
rect 434822 3338 470266 3894
rect 470822 3338 506266 3894
rect 506822 3338 542266 3894
rect 542822 3338 578266 3894
rect 578822 3338 586302 3894
rect 586858 3338 592650 3894
rect -8726 3306 592650 3338
rect -8726 2654 592650 2686
rect -8726 2098 -1974 2654
rect -1418 2098 1026 2654
rect 1582 2098 37026 2654
rect 37582 2098 73026 2654
rect 73582 2098 109026 2654
rect 109582 2098 145026 2654
rect 145582 2098 181026 2654
rect 181582 2098 217026 2654
rect 217582 2098 253026 2654
rect 253582 2098 289026 2654
rect 289582 2098 325026 2654
rect 325582 2098 361026 2654
rect 361582 2098 397026 2654
rect 397582 2098 433026 2654
rect 433582 2098 469026 2654
rect 469582 2098 505026 2654
rect 505582 2098 541026 2654
rect 541582 2098 577026 2654
rect 577582 2098 585342 2654
rect 585898 2098 592650 2654
rect -8726 2066 592650 2098
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1026 -346
rect 1582 -902 37026 -346
rect 37582 -902 73026 -346
rect 73582 -902 109026 -346
rect 109582 -902 145026 -346
rect 145582 -902 181026 -346
rect 181582 -902 217026 -346
rect 217582 -902 253026 -346
rect 253582 -902 289026 -346
rect 289582 -902 325026 -346
rect 325582 -902 361026 -346
rect 361582 -902 397026 -346
rect 397582 -902 433026 -346
rect 433582 -902 469026 -346
rect 469582 -902 505026 -346
rect 505582 -902 541026 -346
rect 541582 -902 577026 -346
rect 577582 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 2266 -1306
rect 2822 -1862 38266 -1306
rect 38822 -1862 74266 -1306
rect 74822 -1862 110266 -1306
rect 110822 -1862 146266 -1306
rect 146822 -1862 182266 -1306
rect 182822 -1862 218266 -1306
rect 218822 -1862 254266 -1306
rect 254822 -1862 290266 -1306
rect 290822 -1862 326266 -1306
rect 326822 -1862 362266 -1306
rect 362822 -1862 398266 -1306
rect 398822 -1862 434266 -1306
rect 434822 -1862 470266 -1306
rect 470822 -1862 506266 -1306
rect 506822 -1862 542266 -1306
rect 542822 -1862 578266 -1306
rect 578822 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 3506 -2266
rect 4062 -2822 39506 -2266
rect 40062 -2822 75506 -2266
rect 76062 -2822 111506 -2266
rect 112062 -2822 147506 -2266
rect 148062 -2822 183506 -2266
rect 184062 -2822 219506 -2266
rect 220062 -2822 255506 -2266
rect 256062 -2822 291506 -2266
rect 292062 -2822 327506 -2266
rect 328062 -2822 363506 -2266
rect 364062 -2822 399506 -2266
rect 400062 -2822 435506 -2266
rect 436062 -2822 471506 -2266
rect 472062 -2822 507506 -2266
rect 508062 -2822 543506 -2266
rect 544062 -2822 579506 -2266
rect 580062 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 4746 -3226
rect 5302 -3782 40746 -3226
rect 41302 -3782 76746 -3226
rect 77302 -3782 112746 -3226
rect 113302 -3782 148746 -3226
rect 149302 -3782 184746 -3226
rect 185302 -3782 220746 -3226
rect 221302 -3782 256746 -3226
rect 257302 -3782 292746 -3226
rect 293302 -3782 328746 -3226
rect 329302 -3782 364746 -3226
rect 365302 -3782 400746 -3226
rect 401302 -3782 436746 -3226
rect 437302 -3782 472746 -3226
rect 473302 -3782 508746 -3226
rect 509302 -3782 544746 -3226
rect 545302 -3782 580746 -3226
rect 581302 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 5986 -4186
rect 6542 -4742 41986 -4186
rect 42542 -4742 77986 -4186
rect 78542 -4742 113986 -4186
rect 114542 -4742 149986 -4186
rect 150542 -4742 185986 -4186
rect 186542 -4742 221986 -4186
rect 222542 -4742 257986 -4186
rect 258542 -4742 293986 -4186
rect 294542 -4742 329986 -4186
rect 330542 -4742 365986 -4186
rect 366542 -4742 401986 -4186
rect 402542 -4742 437986 -4186
rect 438542 -4742 473986 -4186
rect 474542 -4742 509986 -4186
rect 510542 -4742 545986 -4186
rect 546542 -4742 581986 -4186
rect 582542 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 7226 -5146
rect 7782 -5702 43226 -5146
rect 43782 -5702 79226 -5146
rect 79782 -5702 115226 -5146
rect 115782 -5702 151226 -5146
rect 151782 -5702 187226 -5146
rect 187782 -5702 223226 -5146
rect 223782 -5702 259226 -5146
rect 259782 -5702 295226 -5146
rect 295782 -5702 331226 -5146
rect 331782 -5702 367226 -5146
rect 367782 -5702 403226 -5146
rect 403782 -5702 439226 -5146
rect 439782 -5702 475226 -5146
rect 475782 -5702 511226 -5146
rect 511782 -5702 547226 -5146
rect 547782 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 8466 -6106
rect 9022 -6662 44466 -6106
rect 45022 -6662 80466 -6106
rect 81022 -6662 116466 -6106
rect 117022 -6662 152466 -6106
rect 153022 -6662 188466 -6106
rect 189022 -6662 224466 -6106
rect 225022 -6662 260466 -6106
rect 261022 -6662 296466 -6106
rect 297022 -6662 332466 -6106
rect 333022 -6662 368466 -6106
rect 369022 -6662 404466 -6106
rect 405022 -6662 440466 -6106
rect 441022 -6662 476466 -6106
rect 477022 -6662 512466 -6106
rect 513022 -6662 548466 -6106
rect 549022 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 9706 -7066
rect 10262 -7622 45706 -7066
rect 46262 -7622 81706 -7066
rect 82262 -7622 117706 -7066
rect 118262 -7622 153706 -7066
rect 154262 -7622 189706 -7066
rect 190262 -7622 225706 -7066
rect 226262 -7622 261706 -7066
rect 262262 -7622 297706 -7066
rect 298262 -7622 333706 -7066
rect 334262 -7622 369706 -7066
rect 370262 -7622 405706 -7066
rect 406262 -7622 441706 -7066
rect 442262 -7622 477706 -7066
rect 478262 -7622 513706 -7066
rect 514262 -7622 549706 -7066
rect 550262 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use mux16x1_project  mprj1
timestamp 1542649553
transform 1 0 538000 0 1 423800
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 1542649553
transform 1 0 538000 0 1 387800
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 1542649553
transform 1 0 538000 0 1 351800
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 1542649553
transform 1 0 538000 0 1 315800
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 1542649553
transform 1 0 538000 0 1 279800
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro1
timestamp 1542649553
transform 1 0 468600 0 1 449000
box 0 0 20145 2491
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro2
timestamp 1542649553
transform 1 0 468600 0 1 430600
box 0 0 20785 2492
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro3
timestamp 1542649553
transform 1 0 468600 0 1 409600
box 0 0 19886 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro4
timestamp 1542649553
transform 1 0 468600 0 1 388600
box 0 0 22123 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro5
timestamp 1542649553
transform 1 0 468600 0 1 356000
box 0 0 20809 2493
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro6
timestamp 1542649553
transform 1 0 468600 0 1 340000
box 0 0 20217 2494
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro7
timestamp 1542649553
transform 1 0 468600 0 1 320000
box 0 0 20783 2493
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro8
timestamp 1542649553
transform 1 0 468600 0 1 304600
box 0 0 19885 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro9
timestamp 1542649553
transform 1 0 468600 0 1 285000
box 0 0 22120 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro10
timestamp 1542649553
transform 1 0 468600 0 1 265000
box 0 0 20819 2493
use sky130_fd_sc_hd__conb_1  TIE_ZERO_zero_
timestamp 1542649553
transform 1 0 208472 0 1 69632
box -38 -48 314 592
<< labels >>
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 1200 0 0 0 analog_io[2]
port 12 nsew
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 1200 0 0 0 analog_io[3]
port 2 nsew
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 1200 0 0 0 analog_io[4]
port 3 nsew
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 1200 0 0 0 analog_io[5]
port 4 nsew
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 1200 0 0 0 analog_io[6]
port 5 nsew
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 1200 0 0 0 analog_io[7]
port 6 nsew
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 1200 0 0 0 io_in[10]
port 7 nsew
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 1200 0 0 0 io_in[11]
port 8 nsew
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 1200 0 0 0 io_in[12]
port 9 nsew
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 1200 0 0 0 io_in[13]
port 10 nsew
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 1200 0 0 0 io_in[14]
port 11 nsew
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 1200 0 0 0 io_in[9]
port 13 nsew
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 1200 0 0 0 io_oeb[10]
port 14 nsew
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 1200 0 0 0 io_oeb[11]
port 15 nsew
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 1200 0 0 0 io_oeb[12]
port 16 nsew
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 1200 0 0 0 io_oeb[13]
port 17 nsew
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 1200 0 0 0 io_oeb[14]
port 18 nsew
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 1200 0 0 0 io_oeb[8]
port 19 nsew
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 1200 0 0 0 io_oeb[9]
port 20 nsew
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 1200 0 0 0 io_out[10]
port 21 nsew
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 1200 0 0 0 io_out[11]
port 22 nsew
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 1200 0 0 0 io_out[12]
port 23 nsew
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 1200 0 0 0 io_out[13]
port 24 nsew
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 1200 0 0 0 io_out[14]
port 25 nsew
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 1200 0 0 0 io_out[8]
port 26 nsew
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 1200 0 0 0 io_out[9]
port 27 nsew
flabel metal3 s -960 436508 480 436748 0 FreeSans 1200 0 0 0 analog_io[22]
port 54 nsew
flabel metal3 s -960 384284 480 384524 0 FreeSans 1200 0 0 0 analog_io[23]
port 28 nsew
flabel metal3 s -960 697220 480 697460 0 FreeSans 1200 0 0 0 analog_io[17]
port 29 nsew
flabel metal3 s -960 644996 480 645236 0 FreeSans 1200 0 0 0 analog_io[18]
port 30 nsew
flabel metal3 s -960 592908 480 593148 0 FreeSans 1200 0 0 0 analog_io[19]
port 31 nsew
flabel metal3 s -960 658052 480 658292 0 FreeSans 1200 0 0 0 io_oeb[24]
port 33 nsew
flabel metal3 s -960 605964 480 606204 0 FreeSans 1200 0 0 0 io_oeb[25]
port 34 nsew
flabel metal3 s -960 553740 480 553980 0 FreeSans 1200 0 0 0 io_oeb[26]
port 35 nsew
flabel metal3 s -960 501652 480 501892 0 FreeSans 1200 0 0 0 io_oeb[27]
port 36 nsew
flabel metal3 s -960 449428 480 449668 0 FreeSans 1200 0 0 0 io_oeb[28]
port 37 nsew
flabel metal3 s -960 397340 480 397580 0 FreeSans 1200 0 0 0 io_oeb[29]
port 38 nsew
flabel metal3 s -960 540684 480 540924 0 FreeSans 1200 0 0 0 analog_io[20]
port 32 nsew
flabel metal3 s -960 684164 480 684404 0 FreeSans 1200 0 0 0 io_in[24]
port 39 nsew
flabel metal3 s -960 631940 480 632180 0 FreeSans 1200 0 0 0 io_in[25]
port 40 nsew
flabel metal3 s -960 579852 480 580092 0 FreeSans 1200 0 0 0 io_in[26]
port 41 nsew
flabel metal3 s -960 527764 480 528004 0 FreeSans 1200 0 0 0 io_in[27]
port 42 nsew
flabel metal3 s -960 475540 480 475780 0 FreeSans 1200 0 0 0 io_in[28]
port 43 nsew
flabel metal3 s -960 423452 480 423692 0 FreeSans 1200 0 0 0 io_in[29]
port 44 nsew
flabel metal3 s -960 671108 480 671348 0 FreeSans 1200 0 0 0 io_out[24]
port 46 nsew
flabel metal3 s -960 619020 480 619260 0 FreeSans 1200 0 0 0 io_out[25]
port 47 nsew
flabel metal3 s -960 566796 480 567036 0 FreeSans 1200 0 0 0 io_out[26]
port 48 nsew
flabel metal3 s -960 514708 480 514948 0 FreeSans 1200 0 0 0 io_out[27]
port 49 nsew
flabel metal3 s -960 462484 480 462724 0 FreeSans 1200 0 0 0 io_out[28]
port 50 nsew
flabel metal3 s -960 410396 480 410636 0 FreeSans 1200 0 0 0 io_out[29]
port 51 nsew
flabel metal3 s -960 358308 480 358548 0 FreeSans 1200 0 0 0 io_out[30]
port 52 nsew
flabel metal3 s -960 371228 480 371468 0 FreeSans 1200 0 0 0 io_in[30]
port 45 nsew
flabel metal3 s -960 488596 480 488836 0 FreeSans 1200 0 0 0 analog_io[21]
port 53 nsew
flabel metal3 s -960 136628 480 136868 0 FreeSans 1200 0 0 0 io_oeb[34]
port 55 nsew
flabel metal3 s -960 84540 480 84780 0 FreeSans 1200 0 0 0 io_oeb[35]
port 56 nsew
flabel metal3 s -960 45372 480 45612 0 FreeSans 1200 0 0 0 io_oeb[36]
port 57 nsew
flabel metal3 s -960 6340 480 6580 0 FreeSans 1200 0 0 0 io_oeb[37]
port 58 nsew
flabel metal3 s -960 175796 480 176036 0 FreeSans 1200 0 0 0 analog_io[27]
port 70 nsew
flabel metal3 s -960 123572 480 123812 0 FreeSans 1200 0 0 0 analog_io[28]
port 59 nsew
flabel metal3 s -960 332196 480 332436 0 FreeSans 1200 0 0 0 analog_io[24]
port 60 nsew
flabel metal3 s -960 279972 480 280212 0 FreeSans 1200 0 0 0 analog_io[25]
port 61 nsew
flabel metal3 s -960 227884 480 228124 0 FreeSans 1200 0 0 0 analog_io[26]
port 62 nsew
flabel metal3 s -960 319140 480 319380 0 FreeSans 1200 0 0 0 io_in[31]
port 63 nsew
flabel metal3 s -960 267052 480 267292 0 FreeSans 1200 0 0 0 io_in[32]
port 64 nsew
flabel metal3 s -960 214828 480 215068 0 FreeSans 1200 0 0 0 io_in[33]
port 65 nsew
flabel metal3 s -960 162740 480 162980 0 FreeSans 1200 0 0 0 io_in[34]
port 66 nsew
flabel metal3 s -960 110516 480 110756 0 FreeSans 1200 0 0 0 io_in[35]
port 67 nsew
flabel metal3 s -960 71484 480 71724 0 FreeSans 1200 0 0 0 io_in[36]
port 68 nsew
flabel metal3 s -960 32316 480 32556 0 FreeSans 1200 0 0 0 io_in[37]
port 69 nsew
flabel metal3 s -960 345252 480 345492 0 FreeSans 1200 0 0 0 io_oeb[30]
port 71 nsew
flabel metal3 s -960 293028 480 293268 0 FreeSans 1200 0 0 0 io_oeb[31]
port 72 nsew
flabel metal3 s -960 306084 480 306324 0 FreeSans 1200 0 0 0 io_out[31]
port 73 nsew
flabel metal3 s -960 253996 480 254236 0 FreeSans 1200 0 0 0 io_out[32]
port 74 nsew
flabel metal3 s -960 201772 480 202012 0 FreeSans 1200 0 0 0 io_out[33]
port 75 nsew
flabel metal3 s -960 149684 480 149924 0 FreeSans 1200 0 0 0 io_out[34]
port 76 nsew
flabel metal3 s -960 97460 480 97700 0 FreeSans 1200 0 0 0 io_out[35]
port 77 nsew
flabel metal3 s -960 58428 480 58668 0 FreeSans 1200 0 0 0 io_out[36]
port 78 nsew
flabel metal3 s -960 19260 480 19500 0 FreeSans 1200 0 0 0 io_out[37]
port 79 nsew
flabel metal3 s -960 240940 480 241180 0 FreeSans 1200 0 0 0 io_oeb[32]
port 80 nsew
flabel metal3 s -960 188716 480 188956 0 FreeSans 1200 0 0 0 io_oeb[33]
port 81 nsew
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 1200 0 0 0 io_in[8]
port 1 nsew
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 1200 0 0 0 analog_io[1]
port 99 nsew
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 1200 0 0 0 io_oeb[2]
port 82 nsew
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 1200 0 0 0 io_oeb[0]
port 107 nsew
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 1200 0 0 0 io_out[1]
port 85 nsew
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 1200 0 0 0 io_in[2]
port 106 nsew
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 1200 0 0 0 analog_io[0]
port 83 nsew
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 1200 0 0 0 io_in[1]
port 84 nsew
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 1200 0 0 0 io_in[0]
port 86 nsew
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 1200 0 0 0 io_in[3]
port 87 nsew
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 1200 0 0 0 io_oeb[1]
port 89 nsew
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 1200 0 0 0 io_out[2]
port 92 nsew
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 1200 0 0 0 io_in[4]
port 88 nsew
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 1200 0 0 0 io_oeb[3]
port 93 nsew
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 1200 0 0 0 io_oeb[4]
port 94 nsew
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 1200 0 0 0 io_oeb[5]
port 95 nsew
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 1200 0 0 0 io_oeb[6]
port 96 nsew
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 1200 0 0 0 io_oeb[7]
port 97 nsew
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 1200 0 0 0 io_in[5]
port 90 nsew
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 1200 0 0 0 io_in[6]
port 91 nsew
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 1200 0 0 0 io_out[3]
port 101 nsew
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 1200 0 0 0 io_out[4]
port 102 nsew
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 1200 0 0 0 io_out[5]
port 103 nsew
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 1200 0 0 0 io_out[6]
port 104 nsew
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 1200 0 0 0 io_out[7]
port 105 nsew
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 1200 0 0 0 io_out[0]
port 100 nsew
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 1200 0 0 0 io_in[7]
port 98 nsew
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 560 90 0 0 analog_io[10]
port 108 nsew
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 560 90 0 0 analog_io[11]
port 109 nsew
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 560 90 0 0 analog_io[12]
port 110 nsew
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 560 90 0 0 analog_io[8]
port 111 nsew
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 560 90 0 0 analog_io[9]
port 112 nsew
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 560 90 0 0 io_in[15]
port 113 nsew
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 560 90 0 0 io_in[16]
port 114 nsew
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 560 90 0 0 io_in[17]
port 115 nsew
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 560 90 0 0 io_in[18]
port 116 nsew
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 560 90 0 0 io_in[19]
port 117 nsew
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 560 90 0 0 io_oeb[15]
port 118 nsew
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 560 90 0 0 io_oeb[16]
port 119 nsew
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 560 90 0 0 io_oeb[17]
port 120 nsew
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 560 90 0 0 io_oeb[18]
port 121 nsew
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 560 90 0 0 io_out[15]
port 122 nsew
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 560 90 0 0 io_out[16]
port 123 nsew
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 560 90 0 0 io_out[17]
port 124 nsew
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 560 90 0 0 io_out[18]
port 125 nsew
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 560 90 0 0 analog_io[16]
port 126 nsew
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 560 90 0 0 analog_io[13]
port 127 nsew
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 560 90 0 0 analog_io[14]
port 128 nsew
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 560 90 0 0 analog_io[15]
port 129 nsew
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 560 90 0 0 io_oeb[19]
port 130 nsew
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 560 90 0 0 io_oeb[20]
port 131 nsew
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 560 90 0 0 io_oeb[21]
port 132 nsew
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 560 90 0 0 io_oeb[22]
port 133 nsew
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 560 90 0 0 io_oeb[23]
port 134 nsew
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 560 90 0 0 io_in[20]
port 135 nsew
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 560 90 0 0 io_in[21]
port 136 nsew
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 560 90 0 0 io_in[22]
port 137 nsew
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 560 90 0 0 io_in[23]
port 138 nsew
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 560 90 0 0 io_out[19]
port 139 nsew
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 560 90 0 0 io_out[20]
port 140 nsew
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 560 90 0 0 io_out[21]
port 141 nsew
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 560 90 0 0 io_out[22]
port 142 nsew
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 560 90 0 0 io_out[23]
port 143 nsew
flabel metal2 s 542 -960 654 480 0 FreeSans 560 90 0 0 wb_clk_i
port 144 nsew
flabel metal2 s 1646 -960 1758 480 0 FreeSans 560 90 0 0 wb_rst_i
port 145 nsew
flabel metal2 s 2842 -960 2954 480 0 FreeSans 560 90 0 0 wbs_ack_o
port 146 nsew
flabel metal2 s 7626 -960 7738 480 0 FreeSans 560 90 0 0 wbs_adr_i[0]
port 147 nsew
flabel metal2 s 47830 -960 47942 480 0 FreeSans 560 90 0 0 wbs_adr_i[10]
port 148 nsew
flabel metal2 s 51326 -960 51438 480 0 FreeSans 560 90 0 0 wbs_adr_i[11]
port 149 nsew
flabel metal2 s 54914 -960 55026 480 0 FreeSans 560 90 0 0 wbs_adr_i[12]
port 150 nsew
flabel metal2 s 58410 -960 58522 480 0 FreeSans 560 90 0 0 wbs_adr_i[13]
port 151 nsew
flabel metal2 s 61998 -960 62110 480 0 FreeSans 560 90 0 0 wbs_adr_i[14]
port 152 nsew
flabel metal2 s 65494 -960 65606 480 0 FreeSans 560 90 0 0 wbs_adr_i[15]
port 153 nsew
flabel metal2 s 69082 -960 69194 480 0 FreeSans 560 90 0 0 wbs_adr_i[16]
port 154 nsew
flabel metal2 s 72578 -960 72690 480 0 FreeSans 560 90 0 0 wbs_adr_i[17]
port 155 nsew
flabel metal2 s 12318 -960 12430 480 0 FreeSans 560 90 0 0 wbs_adr_i[1]
port 156 nsew
flabel metal2 s 17010 -960 17122 480 0 FreeSans 560 90 0 0 wbs_adr_i[2]
port 157 nsew
flabel metal2 s 21794 -960 21906 480 0 FreeSans 560 90 0 0 wbs_adr_i[3]
port 158 nsew
flabel metal2 s 26486 -960 26598 480 0 FreeSans 560 90 0 0 wbs_adr_i[4]
port 159 nsew
flabel metal2 s 30074 -960 30186 480 0 FreeSans 560 90 0 0 wbs_adr_i[5]
port 160 nsew
flabel metal2 s 33570 -960 33682 480 0 FreeSans 560 90 0 0 wbs_adr_i[6]
port 161 nsew
flabel metal2 s 37158 -960 37270 480 0 FreeSans 560 90 0 0 wbs_adr_i[7]
port 162 nsew
flabel metal2 s 40654 -960 40766 480 0 FreeSans 560 90 0 0 wbs_adr_i[8]
port 163 nsew
flabel metal2 s 44242 -960 44354 480 0 FreeSans 560 90 0 0 wbs_adr_i[9]
port 164 nsew
flabel metal2 s 4038 -960 4150 480 0 FreeSans 560 90 0 0 wbs_cyc_i
port 165 nsew
flabel metal2 s 8730 -960 8842 480 0 FreeSans 560 90 0 0 wbs_dat_i[0]
port 166 nsew
flabel metal2 s 48934 -960 49046 480 0 FreeSans 560 90 0 0 wbs_dat_i[10]
port 167 nsew
flabel metal2 s 52522 -960 52634 480 0 FreeSans 560 90 0 0 wbs_dat_i[11]
port 168 nsew
flabel metal2 s 56018 -960 56130 480 0 FreeSans 560 90 0 0 wbs_dat_i[12]
port 169 nsew
flabel metal2 s 59606 -960 59718 480 0 FreeSans 560 90 0 0 wbs_dat_i[13]
port 170 nsew
flabel metal2 s 63194 -960 63306 480 0 FreeSans 560 90 0 0 wbs_dat_i[14]
port 171 nsew
flabel metal2 s 66690 -960 66802 480 0 FreeSans 560 90 0 0 wbs_dat_i[15]
port 172 nsew
flabel metal2 s 70278 -960 70390 480 0 FreeSans 560 90 0 0 wbs_dat_i[16]
port 173 nsew
flabel metal2 s 13514 -960 13626 480 0 FreeSans 560 90 0 0 wbs_dat_i[1]
port 174 nsew
flabel metal2 s 18206 -960 18318 480 0 FreeSans 560 90 0 0 wbs_dat_i[2]
port 175 nsew
flabel metal2 s 22990 -960 23102 480 0 FreeSans 560 90 0 0 wbs_dat_i[3]
port 176 nsew
flabel metal2 s 27682 -960 27794 480 0 FreeSans 560 90 0 0 wbs_dat_i[4]
port 177 nsew
flabel metal2 s 31270 -960 31382 480 0 FreeSans 560 90 0 0 wbs_dat_i[5]
port 178 nsew
flabel metal2 s 34766 -960 34878 480 0 FreeSans 560 90 0 0 wbs_dat_i[6]
port 179 nsew
flabel metal2 s 38354 -960 38466 480 0 FreeSans 560 90 0 0 wbs_dat_i[7]
port 180 nsew
flabel metal2 s 41850 -960 41962 480 0 FreeSans 560 90 0 0 wbs_dat_i[8]
port 181 nsew
flabel metal2 s 45438 -960 45550 480 0 FreeSans 560 90 0 0 wbs_dat_i[9]
port 182 nsew
flabel metal2 s 9926 -960 10038 480 0 FreeSans 560 90 0 0 wbs_dat_o[0]
port 183 nsew
flabel metal2 s 50130 -960 50242 480 0 FreeSans 560 90 0 0 wbs_dat_o[10]
port 184 nsew
flabel metal2 s 53718 -960 53830 480 0 FreeSans 560 90 0 0 wbs_dat_o[11]
port 185 nsew
flabel metal2 s 57214 -960 57326 480 0 FreeSans 560 90 0 0 wbs_dat_o[12]
port 186 nsew
flabel metal2 s 60802 -960 60914 480 0 FreeSans 560 90 0 0 wbs_dat_o[13]
port 187 nsew
flabel metal2 s 64298 -960 64410 480 0 FreeSans 560 90 0 0 wbs_dat_o[14]
port 188 nsew
flabel metal2 s 67886 -960 67998 480 0 FreeSans 560 90 0 0 wbs_dat_o[15]
port 189 nsew
flabel metal2 s 71474 -960 71586 480 0 FreeSans 560 90 0 0 wbs_dat_o[16]
port 190 nsew
flabel metal2 s 14710 -960 14822 480 0 FreeSans 560 90 0 0 wbs_dat_o[1]
port 191 nsew
flabel metal2 s 19402 -960 19514 480 0 FreeSans 560 90 0 0 wbs_dat_o[2]
port 192 nsew
flabel metal2 s 24186 -960 24298 480 0 FreeSans 560 90 0 0 wbs_dat_o[3]
port 193 nsew
flabel metal2 s 28878 -960 28990 480 0 FreeSans 560 90 0 0 wbs_dat_o[4]
port 194 nsew
flabel metal2 s 32374 -960 32486 480 0 FreeSans 560 90 0 0 wbs_dat_o[5]
port 195 nsew
flabel metal2 s 35962 -960 36074 480 0 FreeSans 560 90 0 0 wbs_dat_o[6]
port 196 nsew
flabel metal2 s 39550 -960 39662 480 0 FreeSans 560 90 0 0 wbs_dat_o[7]
port 197 nsew
flabel metal2 s 43046 -960 43158 480 0 FreeSans 560 90 0 0 wbs_dat_o[8]
port 198 nsew
flabel metal2 s 46634 -960 46746 480 0 FreeSans 560 90 0 0 wbs_dat_o[9]
port 199 nsew
flabel metal2 s 11122 -960 11234 480 0 FreeSans 560 90 0 0 wbs_sel_i[0]
port 200 nsew
flabel metal2 s 15906 -960 16018 480 0 FreeSans 560 90 0 0 wbs_sel_i[1]
port 201 nsew
flabel metal2 s 20598 -960 20710 480 0 FreeSans 560 90 0 0 wbs_sel_i[2]
port 202 nsew
flabel metal2 s 25290 -960 25402 480 0 FreeSans 560 90 0 0 wbs_sel_i[3]
port 203 nsew
flabel metal2 s 5234 -960 5346 480 0 FreeSans 560 90 0 0 wbs_stb_i
port 204 nsew
flabel metal2 s 6430 -960 6542 480 0 FreeSans 560 90 0 0 wbs_we_i
port 205 nsew
flabel metal2 s 73774 -960 73886 480 0 FreeSans 560 90 0 0 wbs_dat_i[17]
port 206 nsew
flabel metal2 s 77362 -960 77474 480 0 FreeSans 560 90 0 0 wbs_dat_i[18]
port 207 nsew
flabel metal2 s 80858 -960 80970 480 0 FreeSans 560 90 0 0 wbs_dat_i[19]
port 208 nsew
flabel metal2 s 76166 -960 76278 480 0 FreeSans 560 90 0 0 wbs_adr_i[18]
port 209 nsew
flabel metal2 s 84446 -960 84558 480 0 FreeSans 560 90 0 0 wbs_dat_i[20]
port 210 nsew
flabel metal2 s 87942 -960 88054 480 0 FreeSans 560 90 0 0 wbs_dat_i[21]
port 211 nsew
flabel metal2 s 91530 -960 91642 480 0 FreeSans 560 90 0 0 wbs_dat_i[22]
port 212 nsew
flabel metal2 s 95118 -960 95230 480 0 FreeSans 560 90 0 0 wbs_dat_i[23]
port 213 nsew
flabel metal2 s 98614 -960 98726 480 0 FreeSans 560 90 0 0 wbs_dat_i[24]
port 214 nsew
flabel metal2 s 102202 -960 102314 480 0 FreeSans 560 90 0 0 wbs_dat_i[25]
port 215 nsew
flabel metal2 s 105698 -960 105810 480 0 FreeSans 560 90 0 0 wbs_dat_i[26]
port 216 nsew
flabel metal2 s 109286 -960 109398 480 0 FreeSans 560 90 0 0 wbs_dat_i[27]
port 217 nsew
flabel metal2 s 112782 -960 112894 480 0 FreeSans 560 90 0 0 wbs_dat_i[28]
port 218 nsew
flabel metal2 s 116370 -960 116482 480 0 FreeSans 560 90 0 0 wbs_dat_i[29]
port 219 nsew
flabel metal2 s 79662 -960 79774 480 0 FreeSans 560 90 0 0 wbs_adr_i[19]
port 220 nsew
flabel metal2 s 119866 -960 119978 480 0 FreeSans 560 90 0 0 wbs_dat_i[30]
port 221 nsew
flabel metal2 s 123454 -960 123566 480 0 FreeSans 560 90 0 0 wbs_dat_i[31]
port 222 nsew
flabel metal2 s 128146 -960 128258 480 0 FreeSans 560 90 0 0 la_oenb[0]
port 223 nsew
flabel metal2 s 83250 -960 83362 480 0 FreeSans 560 90 0 0 wbs_adr_i[20]
port 224 nsew
flabel metal2 s 86838 -960 86950 480 0 FreeSans 560 90 0 0 wbs_adr_i[21]
port 225 nsew
flabel metal2 s 90334 -960 90446 480 0 FreeSans 560 90 0 0 wbs_adr_i[22]
port 226 nsew
flabel metal2 s 93922 -960 94034 480 0 FreeSans 560 90 0 0 wbs_adr_i[23]
port 227 nsew
flabel metal2 s 97418 -960 97530 480 0 FreeSans 560 90 0 0 wbs_adr_i[24]
port 228 nsew
flabel metal2 s 101006 -960 101118 480 0 FreeSans 560 90 0 0 wbs_adr_i[25]
port 229 nsew
flabel metal2 s 104502 -960 104614 480 0 FreeSans 560 90 0 0 wbs_adr_i[26]
port 230 nsew
flabel metal2 s 108090 -960 108202 480 0 FreeSans 560 90 0 0 wbs_adr_i[27]
port 231 nsew
flabel metal2 s 111586 -960 111698 480 0 FreeSans 560 90 0 0 wbs_adr_i[28]
port 232 nsew
flabel metal2 s 115174 -960 115286 480 0 FreeSans 560 90 0 0 wbs_adr_i[29]
port 233 nsew
flabel metal2 s 131734 -960 131846 480 0 FreeSans 560 90 0 0 la_oenb[1]
port 234 nsew
flabel metal2 s 118762 -960 118874 480 0 FreeSans 560 90 0 0 wbs_adr_i[30]
port 235 nsew
flabel metal2 s 122258 -960 122370 480 0 FreeSans 560 90 0 0 wbs_adr_i[31]
port 236 nsew
flabel metal2 s 135230 -960 135342 480 0 FreeSans 560 90 0 0 la_oenb[2]
port 237 nsew
flabel metal2 s 74970 -960 75082 480 0 FreeSans 560 90 0 0 wbs_dat_o[17]
port 238 nsew
flabel metal2 s 78558 -960 78670 480 0 FreeSans 560 90 0 0 wbs_dat_o[18]
port 239 nsew
flabel metal2 s 82054 -960 82166 480 0 FreeSans 560 90 0 0 wbs_dat_o[19]
port 240 nsew
flabel metal2 s 138818 -960 138930 480 0 FreeSans 560 90 0 0 la_oenb[3]
port 241 nsew
flabel metal2 s 85642 -960 85754 480 0 FreeSans 560 90 0 0 wbs_dat_o[20]
port 242 nsew
flabel metal2 s 89138 -960 89250 480 0 FreeSans 560 90 0 0 wbs_dat_o[21]
port 243 nsew
flabel metal2 s 92726 -960 92838 480 0 FreeSans 560 90 0 0 wbs_dat_o[22]
port 244 nsew
flabel metal2 s 96222 -960 96334 480 0 FreeSans 560 90 0 0 wbs_dat_o[23]
port 245 nsew
flabel metal2 s 99810 -960 99922 480 0 FreeSans 560 90 0 0 wbs_dat_o[24]
port 246 nsew
flabel metal2 s 103306 -960 103418 480 0 FreeSans 560 90 0 0 wbs_dat_o[25]
port 247 nsew
flabel metal2 s 106894 -960 107006 480 0 FreeSans 560 90 0 0 wbs_dat_o[26]
port 248 nsew
flabel metal2 s 110482 -960 110594 480 0 FreeSans 560 90 0 0 wbs_dat_o[27]
port 249 nsew
flabel metal2 s 113978 -960 114090 480 0 FreeSans 560 90 0 0 wbs_dat_o[28]
port 250 nsew
flabel metal2 s 117566 -960 117678 480 0 FreeSans 560 90 0 0 wbs_dat_o[29]
port 251 nsew
flabel metal2 s 142406 -960 142518 480 0 FreeSans 560 90 0 0 la_oenb[4]
port 252 nsew
flabel metal2 s 121062 -960 121174 480 0 FreeSans 560 90 0 0 wbs_dat_o[30]
port 253 nsew
flabel metal2 s 124650 -960 124762 480 0 FreeSans 560 90 0 0 wbs_dat_o[31]
port 254 nsew
flabel metal2 s 145902 -960 146014 480 0 FreeSans 560 90 0 0 la_oenb[5]
port 255 nsew
flabel metal2 s 125846 -960 125958 480 0 FreeSans 560 90 0 0 la_data_in[0]
port 256 nsew
flabel metal2 s 129342 -960 129454 480 0 FreeSans 560 90 0 0 la_data_in[1]
port 257 nsew
flabel metal2 s 132930 -960 133042 480 0 FreeSans 560 90 0 0 la_data_in[2]
port 258 nsew
flabel metal2 s 136426 -960 136538 480 0 FreeSans 560 90 0 0 la_data_in[3]
port 259 nsew
flabel metal2 s 140014 -960 140126 480 0 FreeSans 560 90 0 0 la_data_in[4]
port 260 nsew
flabel metal2 s 143510 -960 143622 480 0 FreeSans 560 90 0 0 la_data_in[5]
port 261 nsew
flabel metal2 s 126950 -960 127062 480 0 FreeSans 560 90 0 0 la_data_out[0]
port 262 nsew
flabel metal2 s 130538 -960 130650 480 0 FreeSans 560 90 0 0 la_data_out[1]
port 263 nsew
flabel metal2 s 134126 -960 134238 480 0 FreeSans 560 90 0 0 la_data_out[2]
port 264 nsew
flabel metal2 s 137622 -960 137734 480 0 FreeSans 560 90 0 0 la_data_out[3]
port 265 nsew
flabel metal2 s 141210 -960 141322 480 0 FreeSans 560 90 0 0 la_data_out[4]
port 266 nsew
flabel metal2 s 144706 -960 144818 480 0 FreeSans 560 90 0 0 la_data_out[5]
port 267 nsew
flabel metal2 s 207358 -960 207470 480 0 FreeSans 560 90 0 0 la_data_in[23]
port 268 nsew
flabel metal2 s 210946 -960 211058 480 0 FreeSans 560 90 0 0 la_data_in[24]
port 269 nsew
flabel metal2 s 214442 -960 214554 480 0 FreeSans 560 90 0 0 la_data_in[25]
port 270 nsew
flabel metal2 s 149490 -960 149602 480 0 FreeSans 560 90 0 0 la_oenb[6]
port 271 nsew
flabel metal2 s 152986 -960 153098 480 0 FreeSans 560 90 0 0 la_oenb[7]
port 272 nsew
flabel metal2 s 156574 -960 156686 480 0 FreeSans 560 90 0 0 la_oenb[8]
port 273 nsew
flabel metal2 s 160070 -960 160182 480 0 FreeSans 560 90 0 0 la_oenb[9]
port 274 nsew
flabel metal2 s 218030 -960 218142 480 0 FreeSans 560 90 0 0 la_data_in[26]
port 275 nsew
flabel metal2 s 164854 -960 164966 480 0 FreeSans 560 90 0 0 la_data_in[11]
port 276 nsew
flabel metal2 s 168350 -960 168462 480 0 FreeSans 560 90 0 0 la_data_in[12]
port 277 nsew
flabel metal2 s 171938 -960 172050 480 0 FreeSans 560 90 0 0 la_data_in[13]
port 278 nsew
flabel metal2 s 175434 -960 175546 480 0 FreeSans 560 90 0 0 la_data_in[14]
port 279 nsew
flabel metal2 s 147098 -960 147210 480 0 FreeSans 560 90 0 0 la_data_in[6]
port 280 nsew
flabel metal2 s 150594 -960 150706 480 0 FreeSans 560 90 0 0 la_data_in[7]
port 281 nsew
flabel metal2 s 154182 -960 154294 480 0 FreeSans 560 90 0 0 la_data_in[8]
port 282 nsew
flabel metal2 s 157770 -960 157882 480 0 FreeSans 560 90 0 0 la_data_in[9]
port 283 nsew
flabel metal2 s 179022 -960 179134 480 0 FreeSans 560 90 0 0 la_data_in[15]
port 284 nsew
flabel metal2 s 162462 -960 162574 480 0 FreeSans 560 90 0 0 la_data_out[10]
port 285 nsew
flabel metal2 s 166050 -960 166162 480 0 FreeSans 560 90 0 0 la_data_out[11]
port 286 nsew
flabel metal2 s 169546 -960 169658 480 0 FreeSans 560 90 0 0 la_data_out[12]
port 287 nsew
flabel metal2 s 173134 -960 173246 480 0 FreeSans 560 90 0 0 la_data_out[13]
port 288 nsew
flabel metal2 s 176630 -960 176742 480 0 FreeSans 560 90 0 0 la_data_out[14]
port 289 nsew
flabel metal2 s 180218 -960 180330 480 0 FreeSans 560 90 0 0 la_data_out[15]
port 290 nsew
flabel metal2 s 183714 -960 183826 480 0 FreeSans 560 90 0 0 la_data_out[16]
port 291 nsew
flabel metal2 s 187302 -960 187414 480 0 FreeSans 560 90 0 0 la_data_out[17]
port 292 nsew
flabel metal2 s 190798 -960 190910 480 0 FreeSans 560 90 0 0 la_data_out[18]
port 293 nsew
flabel metal2 s 194386 -960 194498 480 0 FreeSans 560 90 0 0 la_data_out[19]
port 294 nsew
flabel metal2 s 182518 -960 182630 480 0 FreeSans 560 90 0 0 la_data_in[16]
port 295 nsew
flabel metal2 s 197882 -960 197994 480 0 FreeSans 560 90 0 0 la_data_out[20]
port 296 nsew
flabel metal2 s 201470 -960 201582 480 0 FreeSans 560 90 0 0 la_data_out[21]
port 297 nsew
flabel metal2 s 205058 -960 205170 480 0 FreeSans 560 90 0 0 la_data_out[22]
port 298 nsew
flabel metal2 s 208554 -960 208666 480 0 FreeSans 560 90 0 0 la_data_out[23]
port 299 nsew
flabel metal2 s 212142 -960 212254 480 0 FreeSans 560 90 0 0 la_data_out[24]
port 300 nsew
flabel metal2 s 215638 -960 215750 480 0 FreeSans 560 90 0 0 la_data_out[25]
port 301 nsew
flabel metal2 s 186106 -960 186218 480 0 FreeSans 560 90 0 0 la_data_in[17]
port 302 nsew
flabel metal2 s 189694 -960 189806 480 0 FreeSans 560 90 0 0 la_data_in[18]
port 303 nsew
flabel metal2 s 193190 -960 193302 480 0 FreeSans 560 90 0 0 la_data_in[19]
port 304 nsew
flabel metal2 s 161266 -960 161378 480 0 FreeSans 560 90 0 0 la_data_in[10]
port 305 nsew
flabel metal2 s 148294 -960 148406 480 0 FreeSans 560 90 0 0 la_data_out[6]
port 306 nsew
flabel metal2 s 151790 -960 151902 480 0 FreeSans 560 90 0 0 la_data_out[7]
port 307 nsew
flabel metal2 s 155378 -960 155490 480 0 FreeSans 560 90 0 0 la_data_out[8]
port 308 nsew
flabel metal2 s 158874 -960 158986 480 0 FreeSans 560 90 0 0 la_data_out[9]
port 309 nsew
flabel metal2 s 196778 -960 196890 480 0 FreeSans 560 90 0 0 la_data_in[20]
port 310 nsew
flabel metal2 s 163658 -960 163770 480 0 FreeSans 560 90 0 0 la_oenb[10]
port 311 nsew
flabel metal2 s 167154 -960 167266 480 0 FreeSans 560 90 0 0 la_oenb[11]
port 312 nsew
flabel metal2 s 170742 -960 170854 480 0 FreeSans 560 90 0 0 la_oenb[12]
port 313 nsew
flabel metal2 s 174238 -960 174350 480 0 FreeSans 560 90 0 0 la_oenb[13]
port 314 nsew
flabel metal2 s 177826 -960 177938 480 0 FreeSans 560 90 0 0 la_oenb[14]
port 315 nsew
flabel metal2 s 181414 -960 181526 480 0 FreeSans 560 90 0 0 la_oenb[15]
port 316 nsew
flabel metal2 s 184910 -960 185022 480 0 FreeSans 560 90 0 0 la_oenb[16]
port 317 nsew
flabel metal2 s 188498 -960 188610 480 0 FreeSans 560 90 0 0 la_oenb[17]
port 318 nsew
flabel metal2 s 191994 -960 192106 480 0 FreeSans 560 90 0 0 la_oenb[18]
port 319 nsew
flabel metal2 s 195582 -960 195694 480 0 FreeSans 560 90 0 0 la_oenb[19]
port 320 nsew
flabel metal2 s 200274 -960 200386 480 0 FreeSans 560 90 0 0 la_data_in[21]
port 321 nsew
flabel metal2 s 199078 -960 199190 480 0 FreeSans 560 90 0 0 la_oenb[20]
port 322 nsew
flabel metal2 s 202666 -960 202778 480 0 FreeSans 560 90 0 0 la_oenb[21]
port 323 nsew
flabel metal2 s 206162 -960 206274 480 0 FreeSans 560 90 0 0 la_oenb[22]
port 324 nsew
flabel metal2 s 209750 -960 209862 480 0 FreeSans 560 90 0 0 la_oenb[23]
port 325 nsew
flabel metal2 s 213338 -960 213450 480 0 FreeSans 560 90 0 0 la_oenb[24]
port 326 nsew
flabel metal2 s 216834 -960 216946 480 0 FreeSans 560 90 0 0 la_oenb[25]
port 327 nsew
flabel metal2 s 203862 -960 203974 480 0 FreeSans 560 90 0 0 la_data_in[22]
port 328 nsew
flabel metal2 s 264122 -960 264234 480 0 FreeSans 560 90 0 0 la_data_in[39]
port 329 nsew
flabel metal2 s 287766 -960 287878 480 0 FreeSans 560 90 0 0 la_oenb[45]
port 330 nsew
flabel metal2 s 267710 -960 267822 480 0 FreeSans 560 90 0 0 la_data_in[40]
port 331 nsew
flabel metal2 s 219226 -960 219338 480 0 FreeSans 560 90 0 0 la_data_out[26]
port 332 nsew
flabel metal2 s 222722 -960 222834 480 0 FreeSans 560 90 0 0 la_data_out[27]
port 333 nsew
flabel metal2 s 226310 -960 226422 480 0 FreeSans 560 90 0 0 la_data_out[28]
port 334 nsew
flabel metal2 s 229806 -960 229918 480 0 FreeSans 560 90 0 0 la_data_out[29]
port 335 nsew
flabel metal2 s 271206 -960 271318 480 0 FreeSans 560 90 0 0 la_data_in[41]
port 336 nsew
flabel metal2 s 233394 -960 233506 480 0 FreeSans 560 90 0 0 la_data_out[30]
port 337 nsew
flabel metal2 s 236982 -960 237094 480 0 FreeSans 560 90 0 0 la_data_out[31]
port 338 nsew
flabel metal2 s 240478 -960 240590 480 0 FreeSans 560 90 0 0 la_data_out[32]
port 339 nsew
flabel metal2 s 244066 -960 244178 480 0 FreeSans 560 90 0 0 la_data_out[33]
port 340 nsew
flabel metal2 s 247562 -960 247674 480 0 FreeSans 560 90 0 0 la_data_out[34]
port 341 nsew
flabel metal2 s 251150 -960 251262 480 0 FreeSans 560 90 0 0 la_data_out[35]
port 342 nsew
flabel metal2 s 254646 -960 254758 480 0 FreeSans 560 90 0 0 la_data_out[36]
port 343 nsew
flabel metal2 s 258234 -960 258346 480 0 FreeSans 560 90 0 0 la_data_out[37]
port 344 nsew
flabel metal2 s 261730 -960 261842 480 0 FreeSans 560 90 0 0 la_data_out[38]
port 345 nsew
flabel metal2 s 265318 -960 265430 480 0 FreeSans 560 90 0 0 la_data_out[39]
port 346 nsew
flabel metal2 s 274794 -960 274906 480 0 FreeSans 560 90 0 0 la_data_in[42]
port 347 nsew
flabel metal2 s 268814 -960 268926 480 0 FreeSans 560 90 0 0 la_data_out[40]
port 348 nsew
flabel metal2 s 272402 -960 272514 480 0 FreeSans 560 90 0 0 la_data_out[41]
port 349 nsew
flabel metal2 s 275990 -960 276102 480 0 FreeSans 560 90 0 0 la_data_out[42]
port 350 nsew
flabel metal2 s 279486 -960 279598 480 0 FreeSans 560 90 0 0 la_data_out[43]
port 351 nsew
flabel metal2 s 283074 -960 283186 480 0 FreeSans 560 90 0 0 la_data_out[44]
port 352 nsew
flabel metal2 s 286570 -960 286682 480 0 FreeSans 560 90 0 0 la_data_out[45]
port 353 nsew
flabel metal2 s 290158 -960 290270 480 0 FreeSans 560 90 0 0 la_data_out[46]
port 354 nsew
flabel metal2 s 278290 -960 278402 480 0 FreeSans 560 90 0 0 la_data_in[43]
port 355 nsew
flabel metal2 s 281878 -960 281990 480 0 FreeSans 560 90 0 0 la_data_in[44]
port 356 nsew
flabel metal2 s 285374 -960 285486 480 0 FreeSans 560 90 0 0 la_data_in[45]
port 357 nsew
flabel metal2 s 288962 -960 289074 480 0 FreeSans 560 90 0 0 la_data_in[46]
port 358 nsew
flabel metal2 s 291354 -960 291466 480 0 FreeSans 560 90 0 0 la_oenb[46]
port 359 nsew
flabel metal2 s 262926 -960 263038 480 0 FreeSans 560 90 0 0 la_oenb[38]
port 360 nsew
flabel metal2 s 266514 -960 266626 480 0 FreeSans 560 90 0 0 la_oenb[39]
port 361 nsew
flabel metal2 s 259430 -960 259542 480 0 FreeSans 560 90 0 0 la_oenb[37]
port 362 nsew
flabel metal2 s 270010 -960 270122 480 0 FreeSans 560 90 0 0 la_oenb[40]
port 363 nsew
flabel metal2 s 273598 -960 273710 480 0 FreeSans 560 90 0 0 la_oenb[41]
port 364 nsew
flabel metal2 s 277094 -960 277206 480 0 FreeSans 560 90 0 0 la_oenb[42]
port 365 nsew
flabel metal2 s 280682 -960 280794 480 0 FreeSans 560 90 0 0 la_oenb[43]
port 366 nsew
flabel metal2 s 221526 -960 221638 480 0 FreeSans 560 90 0 0 la_data_in[27]
port 367 nsew
flabel metal2 s 225114 -960 225226 480 0 FreeSans 560 90 0 0 la_data_in[28]
port 368 nsew
flabel metal2 s 228702 -960 228814 480 0 FreeSans 560 90 0 0 la_data_in[29]
port 369 nsew
flabel metal2 s 284270 -960 284382 480 0 FreeSans 560 90 0 0 la_oenb[44]
port 370 nsew
flabel metal2 s 232198 -960 232310 480 0 FreeSans 560 90 0 0 la_data_in[30]
port 371 nsew
flabel metal2 s 235786 -960 235898 480 0 FreeSans 560 90 0 0 la_data_in[31]
port 372 nsew
flabel metal2 s 239282 -960 239394 480 0 FreeSans 560 90 0 0 la_data_in[32]
port 373 nsew
flabel metal2 s 242870 -960 242982 480 0 FreeSans 560 90 0 0 la_data_in[33]
port 374 nsew
flabel metal2 s 246366 -960 246478 480 0 FreeSans 560 90 0 0 la_data_in[34]
port 375 nsew
flabel metal2 s 249954 -960 250066 480 0 FreeSans 560 90 0 0 la_data_in[35]
port 376 nsew
flabel metal2 s 253450 -960 253562 480 0 FreeSans 560 90 0 0 la_data_in[36]
port 377 nsew
flabel metal2 s 257038 -960 257150 480 0 FreeSans 560 90 0 0 la_data_in[37]
port 378 nsew
flabel metal2 s 220422 -960 220534 480 0 FreeSans 560 90 0 0 la_oenb[26]
port 379 nsew
flabel metal2 s 223918 -960 224030 480 0 FreeSans 560 90 0 0 la_oenb[27]
port 380 nsew
flabel metal2 s 227506 -960 227618 480 0 FreeSans 560 90 0 0 la_oenb[28]
port 381 nsew
flabel metal2 s 231002 -960 231114 480 0 FreeSans 560 90 0 0 la_oenb[29]
port 382 nsew
flabel metal2 s 260626 -960 260738 480 0 FreeSans 560 90 0 0 la_data_in[38]
port 383 nsew
flabel metal2 s 234590 -960 234702 480 0 FreeSans 560 90 0 0 la_oenb[30]
port 384 nsew
flabel metal2 s 238086 -960 238198 480 0 FreeSans 560 90 0 0 la_oenb[31]
port 385 nsew
flabel metal2 s 241674 -960 241786 480 0 FreeSans 560 90 0 0 la_oenb[32]
port 386 nsew
flabel metal2 s 245170 -960 245282 480 0 FreeSans 560 90 0 0 la_oenb[33]
port 387 nsew
flabel metal2 s 248758 -960 248870 480 0 FreeSans 560 90 0 0 la_oenb[34]
port 388 nsew
flabel metal2 s 252346 -960 252458 480 0 FreeSans 560 90 0 0 la_oenb[35]
port 389 nsew
flabel metal2 s 255842 -960 255954 480 0 FreeSans 560 90 0 0 la_oenb[36]
port 390 nsew
flabel metal2 s 294850 -960 294962 480 0 FreeSans 560 90 0 0 la_oenb[47]
port 391 nsew
flabel metal2 s 298438 -960 298550 480 0 FreeSans 560 90 0 0 la_oenb[48]
port 392 nsew
flabel metal2 s 301934 -960 302046 480 0 FreeSans 560 90 0 0 la_oenb[49]
port 393 nsew
flabel metal2 s 305522 -960 305634 480 0 FreeSans 560 90 0 0 la_oenb[50]
port 394 nsew
flabel metal2 s 309018 -960 309130 480 0 FreeSans 560 90 0 0 la_oenb[51]
port 395 nsew
flabel metal2 s 312606 -960 312718 480 0 FreeSans 560 90 0 0 la_oenb[52]
port 396 nsew
flabel metal2 s 316194 -960 316306 480 0 FreeSans 560 90 0 0 la_oenb[53]
port 397 nsew
flabel metal2 s 319690 -960 319802 480 0 FreeSans 560 90 0 0 la_oenb[54]
port 398 nsew
flabel metal2 s 323278 -960 323390 480 0 FreeSans 560 90 0 0 la_oenb[55]
port 399 nsew
flabel metal2 s 326774 -960 326886 480 0 FreeSans 560 90 0 0 la_oenb[56]
port 400 nsew
flabel metal2 s 330362 -960 330474 480 0 FreeSans 560 90 0 0 la_oenb[57]
port 401 nsew
flabel metal2 s 333858 -960 333970 480 0 FreeSans 560 90 0 0 la_oenb[58]
port 402 nsew
flabel metal2 s 337446 -960 337558 480 0 FreeSans 560 90 0 0 la_oenb[59]
port 403 nsew
flabel metal2 s 340942 -960 341054 480 0 FreeSans 560 90 0 0 la_oenb[60]
port 404 nsew
flabel metal2 s 344530 -960 344642 480 0 FreeSans 560 90 0 0 la_oenb[61]
port 405 nsew
flabel metal2 s 348026 -960 348138 480 0 FreeSans 560 90 0 0 la_oenb[62]
port 406 nsew
flabel metal2 s 351614 -960 351726 480 0 FreeSans 560 90 0 0 la_oenb[63]
port 407 nsew
flabel metal2 s 355202 -960 355314 480 0 FreeSans 560 90 0 0 la_oenb[64]
port 408 nsew
flabel metal2 s 358698 -960 358810 480 0 FreeSans 560 90 0 0 la_oenb[65]
port 409 nsew
flabel metal2 s 362286 -960 362398 480 0 FreeSans 560 90 0 0 la_oenb[66]
port 410 nsew
flabel metal2 s 292550 -960 292662 480 0 FreeSans 560 90 0 0 la_data_in[47]
port 411 nsew
flabel metal2 s 296046 -960 296158 480 0 FreeSans 560 90 0 0 la_data_in[48]
port 412 nsew
flabel metal2 s 299634 -960 299746 480 0 FreeSans 560 90 0 0 la_data_in[49]
port 413 nsew
flabel metal2 s 303130 -960 303242 480 0 FreeSans 560 90 0 0 la_data_in[50]
port 414 nsew
flabel metal2 s 306718 -960 306830 480 0 FreeSans 560 90 0 0 la_data_in[51]
port 415 nsew
flabel metal2 s 310214 -960 310326 480 0 FreeSans 560 90 0 0 la_data_in[52]
port 416 nsew
flabel metal2 s 313802 -960 313914 480 0 FreeSans 560 90 0 0 la_data_in[53]
port 417 nsew
flabel metal2 s 317298 -960 317410 480 0 FreeSans 560 90 0 0 la_data_in[54]
port 418 nsew
flabel metal2 s 320886 -960 320998 480 0 FreeSans 560 90 0 0 la_data_in[55]
port 419 nsew
flabel metal2 s 324382 -960 324494 480 0 FreeSans 560 90 0 0 la_data_in[56]
port 420 nsew
flabel metal2 s 327970 -960 328082 480 0 FreeSans 560 90 0 0 la_data_in[57]
port 421 nsew
flabel metal2 s 331558 -960 331670 480 0 FreeSans 560 90 0 0 la_data_in[58]
port 422 nsew
flabel metal2 s 335054 -960 335166 480 0 FreeSans 560 90 0 0 la_data_in[59]
port 423 nsew
flabel metal2 s 338642 -960 338754 480 0 FreeSans 560 90 0 0 la_data_in[60]
port 424 nsew
flabel metal2 s 342138 -960 342250 480 0 FreeSans 560 90 0 0 la_data_in[61]
port 425 nsew
flabel metal2 s 345726 -960 345838 480 0 FreeSans 560 90 0 0 la_data_in[62]
port 426 nsew
flabel metal2 s 349222 -960 349334 480 0 FreeSans 560 90 0 0 la_data_in[63]
port 427 nsew
flabel metal2 s 293654 -960 293766 480 0 FreeSans 560 90 0 0 la_data_out[47]
port 428 nsew
flabel metal2 s 297242 -960 297354 480 0 FreeSans 560 90 0 0 la_data_out[48]
port 429 nsew
flabel metal2 s 300738 -960 300850 480 0 FreeSans 560 90 0 0 la_data_out[49]
port 430 nsew
flabel metal2 s 352810 -960 352922 480 0 FreeSans 560 90 0 0 la_data_in[64]
port 431 nsew
flabel metal2 s 304326 -960 304438 480 0 FreeSans 560 90 0 0 la_data_out[50]
port 432 nsew
flabel metal2 s 307914 -960 308026 480 0 FreeSans 560 90 0 0 la_data_out[51]
port 433 nsew
flabel metal2 s 311410 -960 311522 480 0 FreeSans 560 90 0 0 la_data_out[52]
port 434 nsew
flabel metal2 s 314998 -960 315110 480 0 FreeSans 560 90 0 0 la_data_out[53]
port 435 nsew
flabel metal2 s 318494 -960 318606 480 0 FreeSans 560 90 0 0 la_data_out[54]
port 436 nsew
flabel metal2 s 322082 -960 322194 480 0 FreeSans 560 90 0 0 la_data_out[55]
port 437 nsew
flabel metal2 s 325578 -960 325690 480 0 FreeSans 560 90 0 0 la_data_out[56]
port 438 nsew
flabel metal2 s 329166 -960 329278 480 0 FreeSans 560 90 0 0 la_data_out[57]
port 439 nsew
flabel metal2 s 332662 -960 332774 480 0 FreeSans 560 90 0 0 la_data_out[58]
port 440 nsew
flabel metal2 s 336250 -960 336362 480 0 FreeSans 560 90 0 0 la_data_out[59]
port 441 nsew
flabel metal2 s 356306 -960 356418 480 0 FreeSans 560 90 0 0 la_data_in[65]
port 442 nsew
flabel metal2 s 339838 -960 339950 480 0 FreeSans 560 90 0 0 la_data_out[60]
port 443 nsew
flabel metal2 s 343334 -960 343446 480 0 FreeSans 560 90 0 0 la_data_out[61]
port 444 nsew
flabel metal2 s 346922 -960 347034 480 0 FreeSans 560 90 0 0 la_data_out[62]
port 445 nsew
flabel metal2 s 350418 -960 350530 480 0 FreeSans 560 90 0 0 la_data_out[63]
port 446 nsew
flabel metal2 s 354006 -960 354118 480 0 FreeSans 560 90 0 0 la_data_out[64]
port 447 nsew
flabel metal2 s 357502 -960 357614 480 0 FreeSans 560 90 0 0 la_data_out[65]
port 448 nsew
flabel metal2 s 361090 -960 361202 480 0 FreeSans 560 90 0 0 la_data_out[66]
port 449 nsew
flabel metal2 s 364586 -960 364698 480 0 FreeSans 560 90 0 0 la_data_out[67]
port 450 nsew
flabel metal2 s 359894 -960 360006 480 0 FreeSans 560 90 0 0 la_data_in[66]
port 451 nsew
flabel metal2 s 363482 -960 363594 480 0 FreeSans 560 90 0 0 la_data_in[67]
port 452 nsew
flabel metal2 s 381146 -960 381258 480 0 FreeSans 560 90 0 0 la_data_in[72]
port 453 nsew
flabel metal2 s 384734 -960 384846 480 0 FreeSans 560 90 0 0 la_data_in[73]
port 454 nsew
flabel metal2 s 388230 -960 388342 480 0 FreeSans 560 90 0 0 la_data_in[74]
port 455 nsew
flabel metal2 s 391818 -960 391930 480 0 FreeSans 560 90 0 0 la_data_in[75]
port 456 nsew
flabel metal2 s 395314 -960 395426 480 0 FreeSans 560 90 0 0 la_data_in[76]
port 457 nsew
flabel metal2 s 398902 -960 399014 480 0 FreeSans 560 90 0 0 la_data_in[77]
port 458 nsew
flabel metal2 s 402490 -960 402602 480 0 FreeSans 560 90 0 0 la_data_in[78]
port 459 nsew
flabel metal2 s 405986 -960 406098 480 0 FreeSans 560 90 0 0 la_data_in[79]
port 460 nsew
flabel metal2 s 409574 -960 409686 480 0 FreeSans 560 90 0 0 la_data_in[80]
port 461 nsew
flabel metal2 s 413070 -960 413182 480 0 FreeSans 560 90 0 0 la_data_in[81]
port 462 nsew
flabel metal2 s 416658 -960 416770 480 0 FreeSans 560 90 0 0 la_data_in[82]
port 463 nsew
flabel metal2 s 420154 -960 420266 480 0 FreeSans 560 90 0 0 la_data_in[83]
port 464 nsew
flabel metal2 s 423742 -960 423854 480 0 FreeSans 560 90 0 0 la_data_in[84]
port 465 nsew
flabel metal2 s 427238 -960 427350 480 0 FreeSans 560 90 0 0 la_data_in[85]
port 466 nsew
flabel metal2 s 430826 -960 430938 480 0 FreeSans 560 90 0 0 la_data_in[86]
port 467 nsew
flabel metal2 s 434414 -960 434526 480 0 FreeSans 560 90 0 0 la_data_in[87]
port 468 nsew
flabel metal2 s 370566 -960 370678 480 0 FreeSans 560 90 0 0 la_data_in[69]
port 469 nsew
flabel metal2 s 365782 -960 365894 480 0 FreeSans 560 90 0 0 la_oenb[67]
port 470 nsew
flabel metal2 s 369370 -960 369482 480 0 FreeSans 560 90 0 0 la_oenb[68]
port 471 nsew
flabel metal2 s 372866 -960 372978 480 0 FreeSans 560 90 0 0 la_oenb[69]
port 472 nsew
flabel metal2 s 376454 -960 376566 480 0 FreeSans 560 90 0 0 la_oenb[70]
port 473 nsew
flabel metal2 s 379950 -960 380062 480 0 FreeSans 560 90 0 0 la_oenb[71]
port 474 nsew
flabel metal2 s 383538 -960 383650 480 0 FreeSans 560 90 0 0 la_oenb[72]
port 475 nsew
flabel metal2 s 387126 -960 387238 480 0 FreeSans 560 90 0 0 la_oenb[73]
port 476 nsew
flabel metal2 s 390622 -960 390734 480 0 FreeSans 560 90 0 0 la_oenb[74]
port 477 nsew
flabel metal2 s 394210 -960 394322 480 0 FreeSans 560 90 0 0 la_oenb[75]
port 478 nsew
flabel metal2 s 397706 -960 397818 480 0 FreeSans 560 90 0 0 la_oenb[76]
port 479 nsew
flabel metal2 s 401294 -960 401406 480 0 FreeSans 560 90 0 0 la_oenb[77]
port 480 nsew
flabel metal2 s 404790 -960 404902 480 0 FreeSans 560 90 0 0 la_oenb[78]
port 481 nsew
flabel metal2 s 408378 -960 408490 480 0 FreeSans 560 90 0 0 la_oenb[79]
port 482 nsew
flabel metal2 s 411874 -960 411986 480 0 FreeSans 560 90 0 0 la_oenb[80]
port 483 nsew
flabel metal2 s 415462 -960 415574 480 0 FreeSans 560 90 0 0 la_oenb[81]
port 484 nsew
flabel metal2 s 418958 -960 419070 480 0 FreeSans 560 90 0 0 la_oenb[82]
port 485 nsew
flabel metal2 s 422546 -960 422658 480 0 FreeSans 560 90 0 0 la_oenb[83]
port 486 nsew
flabel metal2 s 426134 -960 426246 480 0 FreeSans 560 90 0 0 la_oenb[84]
port 487 nsew
flabel metal2 s 429630 -960 429742 480 0 FreeSans 560 90 0 0 la_oenb[85]
port 488 nsew
flabel metal2 s 433218 -960 433330 480 0 FreeSans 560 90 0 0 la_oenb[86]
port 489 nsew
flabel metal2 s 436714 -960 436826 480 0 FreeSans 560 90 0 0 la_oenb[87]
port 490 nsew
flabel metal2 s 368174 -960 368286 480 0 FreeSans 560 90 0 0 la_data_out[68]
port 491 nsew
flabel metal2 s 371670 -960 371782 480 0 FreeSans 560 90 0 0 la_data_out[69]
port 492 nsew
flabel metal2 s 374062 -960 374174 480 0 FreeSans 560 90 0 0 la_data_in[70]
port 493 nsew
flabel metal2 s 375258 -960 375370 480 0 FreeSans 560 90 0 0 la_data_out[70]
port 494 nsew
flabel metal2 s 378846 -960 378958 480 0 FreeSans 560 90 0 0 la_data_out[71]
port 495 nsew
flabel metal2 s 382342 -960 382454 480 0 FreeSans 560 90 0 0 la_data_out[72]
port 496 nsew
flabel metal2 s 385930 -960 386042 480 0 FreeSans 560 90 0 0 la_data_out[73]
port 497 nsew
flabel metal2 s 389426 -960 389538 480 0 FreeSans 560 90 0 0 la_data_out[74]
port 498 nsew
flabel metal2 s 393014 -960 393126 480 0 FreeSans 560 90 0 0 la_data_out[75]
port 499 nsew
flabel metal2 s 396510 -960 396622 480 0 FreeSans 560 90 0 0 la_data_out[76]
port 500 nsew
flabel metal2 s 400098 -960 400210 480 0 FreeSans 560 90 0 0 la_data_out[77]
port 501 nsew
flabel metal2 s 403594 -960 403706 480 0 FreeSans 560 90 0 0 la_data_out[78]
port 502 nsew
flabel metal2 s 407182 -960 407294 480 0 FreeSans 560 90 0 0 la_data_out[79]
port 503 nsew
flabel metal2 s 377650 -960 377762 480 0 FreeSans 560 90 0 0 la_data_in[71]
port 504 nsew
flabel metal2 s 410770 -960 410882 480 0 FreeSans 560 90 0 0 la_data_out[80]
port 505 nsew
flabel metal2 s 414266 -960 414378 480 0 FreeSans 560 90 0 0 la_data_out[81]
port 506 nsew
flabel metal2 s 417854 -960 417966 480 0 FreeSans 560 90 0 0 la_data_out[82]
port 507 nsew
flabel metal2 s 421350 -960 421462 480 0 FreeSans 560 90 0 0 la_data_out[83]
port 508 nsew
flabel metal2 s 424938 -960 425050 480 0 FreeSans 560 90 0 0 la_data_out[84]
port 509 nsew
flabel metal2 s 428434 -960 428546 480 0 FreeSans 560 90 0 0 la_data_out[85]
port 510 nsew
flabel metal2 s 432022 -960 432134 480 0 FreeSans 560 90 0 0 la_data_out[86]
port 511 nsew
flabel metal2 s 435518 -960 435630 480 0 FreeSans 560 90 0 0 la_data_out[87]
port 512 nsew
flabel metal2 s 366978 -960 367090 480 0 FreeSans 560 90 0 0 la_data_in[68]
port 513 nsew
flabel metal2 s 440302 -960 440414 480 0 FreeSans 560 90 0 0 la_oenb[88]
port 514 nsew
flabel metal2 s 443798 -960 443910 480 0 FreeSans 560 90 0 0 la_oenb[89]
port 515 nsew
flabel metal2 s 447386 -960 447498 480 0 FreeSans 560 90 0 0 la_oenb[90]
port 516 nsew
flabel metal2 s 450882 -960 450994 480 0 FreeSans 560 90 0 0 la_oenb[91]
port 517 nsew
flabel metal2 s 454470 -960 454582 480 0 FreeSans 560 90 0 0 la_oenb[92]
port 518 nsew
flabel metal2 s 458058 -960 458170 480 0 FreeSans 560 90 0 0 la_oenb[93]
port 519 nsew
flabel metal2 s 461554 -960 461666 480 0 FreeSans 560 90 0 0 la_oenb[94]
port 520 nsew
flabel metal2 s 465142 -960 465254 480 0 FreeSans 560 90 0 0 la_oenb[95]
port 521 nsew
flabel metal2 s 468638 -960 468750 480 0 FreeSans 560 90 0 0 la_oenb[96]
port 522 nsew
flabel metal2 s 472226 -960 472338 480 0 FreeSans 560 90 0 0 la_oenb[97]
port 523 nsew
flabel metal2 s 475722 -960 475834 480 0 FreeSans 560 90 0 0 la_oenb[98]
port 524 nsew
flabel metal2 s 479310 -960 479422 480 0 FreeSans 560 90 0 0 la_oenb[99]
port 525 nsew
flabel metal2 s 484002 -960 484114 480 0 FreeSans 560 90 0 0 la_data_in[101]
port 526 nsew
flabel metal2 s 487590 -960 487702 480 0 FreeSans 560 90 0 0 la_data_in[102]
port 527 nsew
flabel metal2 s 491086 -960 491198 480 0 FreeSans 560 90 0 0 la_data_in[103]
port 528 nsew
flabel metal2 s 494674 -960 494786 480 0 FreeSans 560 90 0 0 la_data_in[104]
port 529 nsew
flabel metal2 s 498170 -960 498282 480 0 FreeSans 560 90 0 0 la_data_in[105]
port 530 nsew
flabel metal2 s 501758 -960 501870 480 0 FreeSans 560 90 0 0 la_data_in[106]
port 531 nsew
flabel metal2 s 505346 -960 505458 480 0 FreeSans 560 90 0 0 la_data_in[107]
port 532 nsew
flabel metal2 s 508842 -960 508954 480 0 FreeSans 560 90 0 0 la_data_in[108]
port 533 nsew
flabel metal2 s 480506 -960 480618 480 0 FreeSans 560 90 0 0 la_data_in[100]
port 534 nsew
flabel metal2 s 444994 -960 445106 480 0 FreeSans 560 90 0 0 la_data_in[90]
port 535 nsew
flabel metal2 s 448582 -960 448694 480 0 FreeSans 560 90 0 0 la_data_in[91]
port 536 nsew
flabel metal2 s 452078 -960 452190 480 0 FreeSans 560 90 0 0 la_data_in[92]
port 537 nsew
flabel metal2 s 455666 -960 455778 480 0 FreeSans 560 90 0 0 la_data_in[93]
port 538 nsew
flabel metal2 s 459162 -960 459274 480 0 FreeSans 560 90 0 0 la_data_in[94]
port 539 nsew
flabel metal2 s 462750 -960 462862 480 0 FreeSans 560 90 0 0 la_data_in[95]
port 540 nsew
flabel metal2 s 466246 -960 466358 480 0 FreeSans 560 90 0 0 la_data_in[96]
port 541 nsew
flabel metal2 s 469834 -960 469946 480 0 FreeSans 560 90 0 0 la_data_in[97]
port 542 nsew
flabel metal2 s 473422 -960 473534 480 0 FreeSans 560 90 0 0 la_data_in[98]
port 543 nsew
flabel metal2 s 476918 -960 477030 480 0 FreeSans 560 90 0 0 la_data_in[99]
port 544 nsew
flabel metal2 s 481702 -960 481814 480 0 FreeSans 560 90 0 0 la_data_out[100]
port 545 nsew
flabel metal2 s 485198 -960 485310 480 0 FreeSans 560 90 0 0 la_data_out[101]
port 546 nsew
flabel metal2 s 488786 -960 488898 480 0 FreeSans 560 90 0 0 la_data_out[102]
port 547 nsew
flabel metal2 s 492282 -960 492394 480 0 FreeSans 560 90 0 0 la_data_out[103]
port 548 nsew
flabel metal2 s 495870 -960 495982 480 0 FreeSans 560 90 0 0 la_data_out[104]
port 549 nsew
flabel metal2 s 499366 -960 499478 480 0 FreeSans 560 90 0 0 la_data_out[105]
port 550 nsew
flabel metal2 s 456862 -960 456974 480 0 FreeSans 560 90 0 0 la_data_out[93]
port 551 nsew
flabel metal2 s 502954 -960 503066 480 0 FreeSans 560 90 0 0 la_data_out[106]
port 552 nsew
flabel metal2 s 460358 -960 460470 480 0 FreeSans 560 90 0 0 la_data_out[94]
port 553 nsew
flabel metal2 s 506450 -960 506562 480 0 FreeSans 560 90 0 0 la_data_out[107]
port 554 nsew
flabel metal2 s 463946 -960 464058 480 0 FreeSans 560 90 0 0 la_data_out[95]
port 555 nsew
flabel metal2 s 467442 -960 467554 480 0 FreeSans 560 90 0 0 la_data_out[96]
port 556 nsew
flabel metal2 s 510038 -960 510150 480 0 FreeSans 560 90 0 0 la_data_out[108]
port 557 nsew
flabel metal2 s 471030 -960 471142 480 0 FreeSans 560 90 0 0 la_data_out[97]
port 558 nsew
flabel metal2 s 474526 -960 474638 480 0 FreeSans 560 90 0 0 la_data_out[98]
port 559 nsew
flabel metal2 s 478114 -960 478226 480 0 FreeSans 560 90 0 0 la_data_out[99]
port 560 nsew
flabel metal2 s 453274 -960 453386 480 0 FreeSans 560 90 0 0 la_data_out[92]
port 561 nsew
flabel metal2 s 482806 -960 482918 480 0 FreeSans 560 90 0 0 la_oenb[100]
port 562 nsew
flabel metal2 s 486394 -960 486506 480 0 FreeSans 560 90 0 0 la_oenb[101]
port 563 nsew
flabel metal2 s 489890 -960 490002 480 0 FreeSans 560 90 0 0 la_oenb[102]
port 564 nsew
flabel metal2 s 493478 -960 493590 480 0 FreeSans 560 90 0 0 la_oenb[103]
port 565 nsew
flabel metal2 s 497066 -960 497178 480 0 FreeSans 560 90 0 0 la_oenb[104]
port 566 nsew
flabel metal2 s 500562 -960 500674 480 0 FreeSans 560 90 0 0 la_oenb[105]
port 567 nsew
flabel metal2 s 504150 -960 504262 480 0 FreeSans 560 90 0 0 la_oenb[106]
port 568 nsew
flabel metal2 s 507646 -960 507758 480 0 FreeSans 560 90 0 0 la_oenb[107]
port 569 nsew
flabel metal2 s 437910 -960 438022 480 0 FreeSans 560 90 0 0 la_data_in[88]
port 570 nsew
flabel metal2 s 441498 -960 441610 480 0 FreeSans 560 90 0 0 la_data_in[89]
port 571 nsew
flabel metal2 s 439106 -960 439218 480 0 FreeSans 560 90 0 0 la_data_out[88]
port 572 nsew
flabel metal2 s 442602 -960 442714 480 0 FreeSans 560 90 0 0 la_data_out[89]
port 573 nsew
flabel metal2 s 446190 -960 446302 480 0 FreeSans 560 90 0 0 la_data_out[90]
port 574 nsew
flabel metal2 s 449778 -960 449890 480 0 FreeSans 560 90 0 0 la_data_out[91]
port 575 nsew
flabel metal2 s 547850 -960 547962 480 0 FreeSans 560 90 0 0 la_data_in[119]
port 576 nsew
flabel metal2 s 552634 -960 552746 480 0 FreeSans 560 90 0 0 la_data_out[120]
port 577 nsew
flabel metal2 s 556130 -960 556242 480 0 FreeSans 560 90 0 0 la_data_out[121]
port 578 nsew
flabel metal2 s 559718 -960 559830 480 0 FreeSans 560 90 0 0 la_data_out[122]
port 579 nsew
flabel metal2 s 537178 -960 537290 480 0 FreeSans 560 90 0 0 la_data_in[116]
port 580 nsew
flabel metal2 s 540766 -960 540878 480 0 FreeSans 560 90 0 0 la_data_in[117]
port 581 nsew
flabel metal2 s 563214 -960 563326 480 0 FreeSans 560 90 0 0 la_data_out[123]
port 582 nsew
flabel metal2 s 523010 -960 523122 480 0 FreeSans 560 90 0 0 la_data_in[112]
port 583 nsew
flabel metal2 s 566802 -960 566914 480 0 FreeSans 560 90 0 0 la_data_out[124]
port 584 nsew
flabel metal2 s 570298 -960 570410 480 0 FreeSans 560 90 0 0 la_data_out[125]
port 585 nsew
flabel metal2 s 573886 -960 573998 480 0 FreeSans 560 90 0 0 la_data_out[126]
port 586 nsew
flabel metal2 s 577382 -960 577494 480 0 FreeSans 560 90 0 0 la_data_out[127]
port 587 nsew
flabel metal2 s 544354 -960 544466 480 0 FreeSans 560 90 0 0 la_data_in[118]
port 588 nsew
flabel metal2 s 514730 -960 514842 480 0 FreeSans 560 90 0 0 la_oenb[109]
port 589 nsew
flabel metal2 s 551438 -960 551550 480 0 FreeSans 560 90 0 0 la_data_in[120]
port 590 nsew
flabel metal2 s 518318 -960 518430 480 0 FreeSans 560 90 0 0 la_oenb[110]
port 591 nsew
flabel metal2 s 554934 -960 555046 480 0 FreeSans 560 90 0 0 la_data_in[121]
port 592 nsew
flabel metal2 s 521814 -960 521926 480 0 FreeSans 560 90 0 0 la_oenb[111]
port 593 nsew
flabel metal2 s 525402 -960 525514 480 0 FreeSans 560 90 0 0 la_oenb[112]
port 594 nsew
flabel metal2 s 528990 -960 529102 480 0 FreeSans 560 90 0 0 la_oenb[113]
port 595 nsew
flabel metal2 s 532486 -960 532598 480 0 FreeSans 560 90 0 0 la_oenb[114]
port 596 nsew
flabel metal2 s 536074 -960 536186 480 0 FreeSans 560 90 0 0 la_oenb[115]
port 597 nsew
flabel metal2 s 539570 -960 539682 480 0 FreeSans 560 90 0 0 la_oenb[116]
port 598 nsew
flabel metal2 s 543158 -960 543270 480 0 FreeSans 560 90 0 0 la_oenb[117]
port 599 nsew
flabel metal2 s 546654 -960 546766 480 0 FreeSans 560 90 0 0 la_oenb[118]
port 600 nsew
flabel metal2 s 550242 -960 550354 480 0 FreeSans 560 90 0 0 la_oenb[119]
port 601 nsew
flabel metal2 s 558522 -960 558634 480 0 FreeSans 560 90 0 0 la_data_in[122]
port 602 nsew
flabel metal2 s 562018 -960 562130 480 0 FreeSans 560 90 0 0 la_data_in[123]
port 603 nsew
flabel metal2 s 553738 -960 553850 480 0 FreeSans 560 90 0 0 la_oenb[120]
port 604 nsew
flabel metal2 s 557326 -960 557438 480 0 FreeSans 560 90 0 0 la_oenb[121]
port 605 nsew
flabel metal2 s 560822 -960 560934 480 0 FreeSans 560 90 0 0 la_oenb[122]
port 606 nsew
flabel metal2 s 564410 -960 564522 480 0 FreeSans 560 90 0 0 la_oenb[123]
port 607 nsew
flabel metal2 s 567998 -960 568110 480 0 FreeSans 560 90 0 0 la_oenb[124]
port 608 nsew
flabel metal2 s 571494 -960 571606 480 0 FreeSans 560 90 0 0 la_oenb[125]
port 609 nsew
flabel metal2 s 575082 -960 575194 480 0 FreeSans 560 90 0 0 la_oenb[126]
port 610 nsew
flabel metal2 s 578578 -960 578690 480 0 FreeSans 560 90 0 0 la_oenb[127]
port 611 nsew
flabel metal2 s 565606 -960 565718 480 0 FreeSans 560 90 0 0 la_data_in[124]
port 612 nsew
flabel metal2 s 569102 -960 569214 480 0 FreeSans 560 90 0 0 la_data_in[125]
port 613 nsew
flabel metal2 s 572690 -960 572802 480 0 FreeSans 560 90 0 0 la_data_in[126]
port 614 nsew
flabel metal2 s 576278 -960 576390 480 0 FreeSans 560 90 0 0 la_data_in[127]
port 615 nsew
flabel metal2 s 517122 -960 517234 480 0 FreeSans 560 90 0 0 la_data_out[110]
port 616 nsew
flabel metal2 s 579774 -960 579886 480 0 FreeSans 560 90 0 0 user_clock2
port 617 nsew
flabel metal2 s 580970 -960 581082 480 0 FreeSans 560 90 0 0 user_irq[0]
port 618 nsew
flabel metal2 s 526598 -960 526710 480 0 FreeSans 560 90 0 0 la_data_in[113]
port 619 nsew
flabel metal2 s 582166 -960 582278 480 0 FreeSans 560 90 0 0 user_irq[1]
port 620 nsew
flabel metal2 s 530094 -960 530206 480 0 FreeSans 560 90 0 0 la_data_in[114]
port 621 nsew
flabel metal2 s 583362 -960 583474 480 0 FreeSans 560 90 0 0 user_irq[2]
port 622 nsew
flabel metal2 s 520710 -960 520822 480 0 FreeSans 560 90 0 0 la_data_out[111]
port 623 nsew
flabel metal2 s 524206 -960 524318 480 0 FreeSans 560 90 0 0 la_data_out[112]
port 624 nsew
flabel metal2 s 513534 -960 513646 480 0 FreeSans 560 90 0 0 la_data_out[109]
port 625 nsew
flabel metal2 s 512430 -960 512542 480 0 FreeSans 560 90 0 0 la_data_in[109]
port 626 nsew
flabel metal2 s 527794 -960 527906 480 0 FreeSans 560 90 0 0 la_data_out[113]
port 627 nsew
flabel metal2 s 515926 -960 516038 480 0 FreeSans 560 90 0 0 la_data_in[110]
port 628 nsew
flabel metal2 s 531290 -960 531402 480 0 FreeSans 560 90 0 0 la_data_out[114]
port 629 nsew
flabel metal2 s 511234 -960 511346 480 0 FreeSans 560 90 0 0 la_oenb[108]
port 630 nsew
flabel metal2 s 534878 -960 534990 480 0 FreeSans 560 90 0 0 la_data_out[115]
port 631 nsew
flabel metal2 s 538374 -960 538486 480 0 FreeSans 560 90 0 0 la_data_out[116]
port 632 nsew
flabel metal2 s 519514 -960 519626 480 0 FreeSans 560 90 0 0 la_data_in[111]
port 633 nsew
flabel metal2 s 541962 -960 542074 480 0 FreeSans 560 90 0 0 la_data_out[117]
port 634 nsew
flabel metal2 s 533682 -960 533794 480 0 FreeSans 560 90 0 0 la_data_in[115]
port 635 nsew
flabel metal2 s 545458 -960 545570 480 0 FreeSans 560 90 0 0 la_data_out[118]
port 636 nsew
flabel metal2 s 549046 -960 549158 480 0 FreeSans 560 90 0 0 la_data_out[119]
port 637 nsew
flabel metal4 s 540994 445572 541614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 543474 445572 544094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 545954 445572 546574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 473954 359060 474574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 476434 359060 477054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 475194 359060 475814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 477674 359060 478294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 542234 445572 542854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 544714 445572 545334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 472714 359060 473334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 288994 -7654 289614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 291474 -7654 292094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 255474 -7654 256094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 219474 -7654 220094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 183474 -7654 184094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 147474 -7654 148094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 111474 -7654 112094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 75474 -7654 76094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 39474 -7654 40094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 3474 -7654 4094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 252994 -7654 253614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 216994 -7654 217614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 257954 -7654 258574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 221954 -7654 222574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 185954 -7654 186574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 149954 -7654 150574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 113954 -7654 114574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 77954 -7654 78574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 41954 -7654 42574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 5954 -7654 6574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 180994 -7654 181614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 260434 -7654 261054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 224434 -7654 225054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 188434 -7654 189054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 152434 -7654 153054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 116434 -7654 117054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 80434 -7654 81054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 44434 -7654 45054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 8434 -7654 9054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 144994 -7654 145614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 259194 -7654 259814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 223194 -7654 223814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 187194 -7654 187814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 151194 -7654 151814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 115194 -7654 115814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 79194 -7654 79814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 43194 -7654 43814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 7194 -7654 7814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 108994 -7654 109614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 261674 -7654 262294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 225674 -7654 226294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 189674 -7654 190294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 153674 -7654 154294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 117674 -7654 118294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 81674 -7654 82294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 45674 -7654 46294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 9674 -7654 10294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 72994 -7654 73614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 290234 -7654 290854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 254234 -7654 254854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 218234 -7654 218854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 182234 -7654 182854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 146234 -7654 146854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 110234 -7654 110854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 74234 -7654 74854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 38234 -7654 38854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 2234 -7654 2854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 36994 -7654 37614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 994 -7654 1614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 256714 -7654 257334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 220714 -7654 221334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 184714 -7654 185334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 148714 -7654 149334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 112714 -7654 113334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 76714 -7654 77334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 40714 -7654 41334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 4714 -7654 5334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 475194 268060 475814 354615 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 475194 -7654 475814 263615 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 439194 -7654 439814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 403194 -7654 403814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 367194 -7654 367814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 331194 -7654 331814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 295194 -7654 295814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 507474 -7654 508094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 473954 268060 474574 354615 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 473954 -7654 474574 263615 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 437954 -7654 438574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 401954 -7654 402574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 365954 -7654 366574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 329954 -7654 330574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 293954 -7654 294574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 471474 -7654 472094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 549674 -7654 550294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 513674 -7654 514294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 435474 -7654 436094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 477674 268060 478294 354615 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 477674 -7654 478294 263615 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 441674 -7654 442294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 405674 -7654 406294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 369674 -7654 370294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 333674 -7654 334294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 297674 -7654 298294 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 399474 -7654 400094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 363474 -7654 364094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 327474 -7654 328094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 468994 -7654 469614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 432994 -7654 433614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 396994 -7654 397614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 360994 -7654 361614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 4800 90 0 0 vssa2
port 643 nsew
flabel metal4 s 548434 -7654 549054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 578234 -7654 578854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 512434 -7654 513054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 542234 -7654 542854 279788 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 506234 -7654 506854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 470234 -7654 470854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 434234 -7654 434854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 398234 -7654 398854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 362234 -7654 362854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 326234 -7654 326854 711590 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 324994 -7654 325614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 476434 268060 477054 354615 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 476434 -7654 477054 263615 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 440434 -7654 441054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 404434 -7654 405054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 368434 -7654 369054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 332434 -7654 333054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 296434 -7654 297054 711590 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 576994 -7654 577614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 4800 90 0 0 vssd1
port 644 nsew
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 580714 -7654 581334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 540994 -7654 541614 279788 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 544714 -7654 545334 279788 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 508714 -7654 509334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 579474 -7654 580094 711590 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 472714 268060 473334 354615 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 472714 -7654 473334 263615 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 436714 -7654 437334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 400714 -7654 401334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 364714 -7654 365334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 328714 -7654 329334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 292714 -7654 293334 711590 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 504994 -7654 505614 711590 0 FreeSans 4800 90 0 0 vccd1
port 638 nsew
flabel metal4 s 581954 -7654 582574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 543474 -7654 544094 279788 0 FreeSans 4800 90 0 0 vccd2
port 639 nsew
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 4800 90 0 0 vdda2
port 641 nsew
flabel metal4 s 545954 -7654 546574 279788 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal4 s 547194 -7654 547814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 511194 -7654 511814 711590 0 FreeSans 4800 90 0 0 vssa1
port 642 nsew
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 4800 90 0 0 vssd2
port 645 nsew
flabel metal4 s 509954 -7654 510574 711590 0 FreeSans 4800 90 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 686066 592650 686686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 650066 592650 650686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 614066 592650 614686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 578066 592650 578686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 542066 592650 542686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 506066 592650 506686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 470066 592650 470686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 434066 592650 434686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 398066 592650 398686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 362066 592650 362686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 688546 592650 689166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 652546 592650 653166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 616546 592650 617166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 580546 592650 581166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 544546 592650 545166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 508546 592650 509166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 472546 592650 473166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 436546 592650 437166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 400546 592650 401166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 364546 592650 365166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 691026 592650 691646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 655026 592650 655646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 619026 592650 619646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 583026 592650 583646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 547026 592650 547646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 511026 592650 511646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 475026 592650 475646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 439026 592650 439646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 403026 592650 403646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 367026 592650 367646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 693506 592650 694126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 657506 592650 658126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 621506 592650 622126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 585506 592650 586126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 549506 592650 550126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 513506 592650 514126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 477506 592650 478126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 441506 592650 442126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 405506 592650 406126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 369506 592650 370126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 692266 592650 692886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 656266 592650 656886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 620266 592650 620886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 584266 592650 584886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 548266 592650 548886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 512266 592650 512886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 476266 592650 476886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 440266 592650 440886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 404266 592650 404886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 368266 592650 368886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 694746 592650 695366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 658746 592650 659366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 622746 592650 623366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 586746 592650 587366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 550746 592650 551366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 514746 592650 515366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 478746 592650 479366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 442746 592650 443366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 406746 592650 407366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 370746 592650 371366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 687306 592650 687926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 651306 592650 651926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 615306 592650 615926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 579306 592650 579926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 543306 592650 543926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 507306 592650 507926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 471306 592650 471926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 435306 592650 435926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 399306 592650 399926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 363306 592650 363926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 689786 592650 690406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 653786 592650 654406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 617786 592650 618406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 581786 592650 582406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 545786 592650 546406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 509786 592650 510406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 473786 592650 474406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 437786 592650 438406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 401786 592650 402406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 365786 592650 366406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 290066 592650 290686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 254066 592650 254686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 218066 592650 218686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 182066 592650 182686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 146066 592650 146686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 110066 592650 110686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 74066 592650 74686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 38066 592650 38686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 2066 592650 2686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 326066 592650 326686 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 332266 592650 332886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 296266 592650 296886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 260266 592650 260886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 224266 592650 224886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 188266 592650 188886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 152266 592650 152886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 116266 592650 116886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 80266 592650 80886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 44266 592650 44886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 8266 592650 8886 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 331026 592650 331646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 3200 0 0 0 vssa1
port 642 nsew
flabel metal5 s -8726 295026 592650 295646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 259026 592650 259646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 223026 592650 223646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 187026 592650 187646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 151026 592650 151646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 115026 592650 115646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 79026 592650 79646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 43026 592650 43646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 7026 592650 7646 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 328546 592650 329166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 334746 592650 335366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 298746 592650 299366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 262746 592650 263366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 226746 592650 227366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 190746 592650 191366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 154746 592650 155366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 118746 592650 119366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 82746 592650 83366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 46746 592650 47366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 10746 592650 11366 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 3200 0 0 0 vdda1
port 640 nsew
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 3200 0 0 0 vssa2
port 643 nsew
flabel metal5 s -8726 292546 592650 293166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 256546 592650 257166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 220546 592650 221166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 184546 592650 185166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 148546 592650 149166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 112546 592650 113166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 76546 592650 77166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 40546 592650 41166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 4546 592650 5166 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 3200 0 0 0 vccd1
port 638 nsew
flabel metal5 s -8726 327306 592650 327926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 291306 592650 291926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 255306 592650 255926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 219306 592650 219926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 183306 592650 183926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 147306 592650 147926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 111306 592650 111926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 75306 592650 75926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 39306 592650 39926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 3306 592650 3926 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 333506 592650 334126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 3200 0 0 0 vssd1
port 644 nsew
flabel metal5 s -8726 297506 592650 298126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 261506 592650 262126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 225506 592650 226126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 189506 592650 190126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 153506 592650 154126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 117506 592650 118126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 81506 592650 82126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 45506 592650 46126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -8726 9506 592650 10126 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 3200 0 0 0 vccd2
port 639 nsew
flabel metal5 s -8726 329786 592650 330406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 293786 592650 294406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 257786 592650 258406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 221786 592650 222406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 185786 592650 186406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 149786 592650 150406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 113786 592650 114406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 77786 592650 78406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 41786 592650 42406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -8726 5786 592650 6406 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 3200 0 0 0 vdda2
port 641 nsew
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 3200 0 0 0 vssd2
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
