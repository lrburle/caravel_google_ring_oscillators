VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r1 ;
  SIZE 81.725 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 18.055 2.21 18.225 2.38 ;
        RECT 18.05 2.205 18.22 2.375 ;
        RECT 18.05 3.685 18.22 3.855 ;
      LAYER li1 ;
        RECT 18.055 2.21 18.225 2.38 ;
        RECT 18.05 1.865 18.22 2.375 ;
        RECT 18.05 3.685 18.22 5.155 ;
      LAYER met1 ;
        RECT 17.99 3.655 18.28 3.885 ;
        RECT 17.99 2.175 18.28 2.405 ;
        RECT 18.05 2.175 18.22 3.885 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 33.835 2.21 34.005 2.38 ;
        RECT 33.83 2.205 34 2.375 ;
        RECT 33.83 3.685 34 3.855 ;
      LAYER li1 ;
        RECT 33.835 2.21 34.005 2.38 ;
        RECT 33.83 1.865 34 2.375 ;
        RECT 33.83 3.685 34 5.155 ;
      LAYER met1 ;
        RECT 33.77 3.655 34.06 3.885 ;
        RECT 33.77 2.175 34.06 2.405 ;
        RECT 33.83 2.175 34 3.885 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 49.61 2.21 49.78 2.38 ;
        RECT 49.605 2.205 49.775 2.375 ;
        RECT 49.605 3.685 49.775 3.855 ;
      LAYER li1 ;
        RECT 49.61 2.21 49.78 2.38 ;
        RECT 49.605 1.865 49.775 2.375 ;
        RECT 49.605 3.685 49.775 5.155 ;
      LAYER met1 ;
        RECT 49.545 3.655 49.835 3.885 ;
        RECT 49.545 2.175 49.835 2.405 ;
        RECT 49.605 2.175 49.775 3.885 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 65.395 2.21 65.565 2.38 ;
        RECT 65.39 2.205 65.56 2.375 ;
        RECT 65.39 3.685 65.56 3.855 ;
      LAYER li1 ;
        RECT 65.395 2.21 65.565 2.38 ;
        RECT 65.39 1.865 65.56 2.375 ;
        RECT 65.39 3.685 65.56 5.155 ;
      LAYER met1 ;
        RECT 65.33 3.655 65.62 3.885 ;
        RECT 65.33 2.175 65.62 2.405 ;
        RECT 65.39 2.175 65.56 3.885 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 81.18 2.21 81.35 2.38 ;
        RECT 81.175 2.205 81.345 2.375 ;
        RECT 81.175 3.685 81.345 3.855 ;
      LAYER li1 ;
        RECT 81.18 2.21 81.35 2.38 ;
        RECT 81.175 1.865 81.345 2.375 ;
        RECT 81.175 3.685 81.345 5.155 ;
      LAYER met1 ;
        RECT 81.115 3.655 81.405 3.885 ;
        RECT 81.115 2.175 81.405 2.405 ;
        RECT 81.175 2.175 81.345 3.885 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 13.815 8.14 14.165 8.49 ;
        RECT 13.81 4 14.16 4.35 ;
        RECT 13.885 4 14.06 8.49 ;
      LAYER li1 ;
        RECT 13.9 2.955 14.07 4.23 ;
        RECT 13.9 8.23 14.07 9.505 ;
        RECT 9.12 8.23 9.29 9.505 ;
      LAYER met1 ;
        RECT 13.81 4.06 14.3 4.23 ;
        RECT 13.81 4 14.16 4.35 ;
        RECT 9.06 8.23 14.3 8.4 ;
        RECT 13.815 8.14 14.165 8.49 ;
        RECT 9.06 8.2 9.35 8.43 ;
      LAYER via1 ;
        RECT 13.91 4.1 14.06 4.25 ;
        RECT 13.915 8.24 14.065 8.39 ;
      LAYER mcon ;
        RECT 9.12 8.23 9.29 8.4 ;
        RECT 13.9 8.23 14.07 8.4 ;
        RECT 13.9 4.06 14.07 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 29.595 8.14 29.945 8.49 ;
        RECT 29.59 4 29.94 4.35 ;
        RECT 29.665 4 29.84 8.49 ;
      LAYER li1 ;
        RECT 29.68 2.955 29.85 4.23 ;
        RECT 29.68 8.23 29.85 9.505 ;
        RECT 24.9 8.23 25.07 9.505 ;
      LAYER met1 ;
        RECT 29.59 4.06 30.08 4.23 ;
        RECT 29.59 4 29.94 4.35 ;
        RECT 24.84 8.23 30.08 8.4 ;
        RECT 29.595 8.14 29.945 8.49 ;
        RECT 24.84 8.2 25.13 8.43 ;
      LAYER via1 ;
        RECT 29.69 4.1 29.84 4.25 ;
        RECT 29.695 8.24 29.845 8.39 ;
      LAYER mcon ;
        RECT 24.9 8.23 25.07 8.4 ;
        RECT 29.68 8.23 29.85 8.4 ;
        RECT 29.68 4.06 29.85 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 45.37 8.14 45.72 8.49 ;
        RECT 45.365 4 45.715 4.35 ;
        RECT 45.44 4 45.615 8.49 ;
      LAYER li1 ;
        RECT 45.455 2.955 45.625 4.23 ;
        RECT 45.455 8.23 45.625 9.505 ;
        RECT 40.675 8.23 40.845 9.505 ;
      LAYER met1 ;
        RECT 45.365 4.06 45.855 4.23 ;
        RECT 45.365 4 45.715 4.35 ;
        RECT 40.615 8.23 45.855 8.4 ;
        RECT 45.37 8.14 45.72 8.49 ;
        RECT 40.615 8.2 40.905 8.43 ;
      LAYER via1 ;
        RECT 45.465 4.1 45.615 4.25 ;
        RECT 45.47 8.24 45.62 8.39 ;
      LAYER mcon ;
        RECT 40.675 8.23 40.845 8.4 ;
        RECT 45.455 8.23 45.625 8.4 ;
        RECT 45.455 4.06 45.625 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 61.155 8.14 61.505 8.49 ;
        RECT 61.15 4 61.5 4.35 ;
        RECT 61.225 4 61.4 8.49 ;
      LAYER li1 ;
        RECT 61.24 2.955 61.41 4.23 ;
        RECT 61.24 8.23 61.41 9.505 ;
        RECT 56.46 8.23 56.63 9.505 ;
      LAYER met1 ;
        RECT 61.15 4.06 61.64 4.23 ;
        RECT 61.15 4 61.5 4.35 ;
        RECT 56.4 8.23 61.64 8.4 ;
        RECT 61.155 8.14 61.505 8.49 ;
        RECT 56.4 8.2 56.69 8.43 ;
      LAYER via1 ;
        RECT 61.25 4.1 61.4 4.25 ;
        RECT 61.255 8.24 61.405 8.39 ;
      LAYER mcon ;
        RECT 56.46 8.23 56.63 8.4 ;
        RECT 61.24 8.23 61.41 8.4 ;
        RECT 61.24 4.06 61.41 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 76.94 8.14 77.29 8.49 ;
        RECT 76.935 4 77.285 4.35 ;
        RECT 77.01 4 77.185 8.49 ;
      LAYER li1 ;
        RECT 77.025 2.955 77.195 4.23 ;
        RECT 77.025 8.23 77.195 9.505 ;
        RECT 72.245 8.23 72.415 9.505 ;
      LAYER met1 ;
        RECT 76.935 4.06 77.425 4.23 ;
        RECT 76.935 4 77.285 4.35 ;
        RECT 72.185 8.23 77.425 8.4 ;
        RECT 76.94 8.14 77.29 8.49 ;
        RECT 72.185 8.2 72.475 8.43 ;
      LAYER via1 ;
        RECT 77.035 4.1 77.185 4.25 ;
        RECT 77.04 8.24 77.19 8.39 ;
      LAYER mcon ;
        RECT 72.245 8.23 72.415 8.4 ;
        RECT 77.025 8.23 77.195 8.4 ;
        RECT 77.025 4.06 77.195 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.23 8.23 0.4 9.505 ;
      LAYER met1 ;
        RECT 0.17 8.23 0.63 8.4 ;
        RECT 0.17 8.2 0.46 8.43 ;
      LAYER mcon ;
        RECT 0.23 8.23 0.4 8.4 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.53 81.72 7.03 ;
        RECT 2.75 5.43 81.72 7.03 ;
        RECT 65.875 5.425 81.64 7.03 ;
        RECT 79.585 5.425 81.565 7.035 ;
        RECT 80.745 4.695 80.915 7.765 ;
        RECT 79.755 4.695 79.925 7.765 ;
        RECT 77.015 4.7 77.185 7.76 ;
        RECT 75.215 4.93 75.385 7.03 ;
        RECT 74.255 4.93 74.425 7.03 ;
        RECT 72.235 5.425 72.405 7.76 ;
        RECT 71.815 4.93 71.985 7.03 ;
        RECT 70.815 4.93 70.985 7.03 ;
        RECT 69.855 4.93 70.025 7.03 ;
        RECT 67.415 4.93 67.585 7.03 ;
        RECT 50.09 5.425 65.855 7.03 ;
        RECT 63.8 5.425 65.78 7.035 ;
        RECT 64.96 4.695 65.13 7.765 ;
        RECT 63.97 4.695 64.14 7.765 ;
        RECT 61.23 4.7 61.4 7.76 ;
        RECT 59.43 4.93 59.6 7.03 ;
        RECT 58.47 4.93 58.64 7.03 ;
        RECT 56.45 5.425 56.62 7.76 ;
        RECT 56.03 4.93 56.2 7.03 ;
        RECT 55.03 4.93 55.2 7.03 ;
        RECT 54.07 4.93 54.24 7.03 ;
        RECT 51.63 4.93 51.8 7.03 ;
        RECT 34.305 5.425 50.07 7.03 ;
        RECT 48.015 5.425 49.995 7.035 ;
        RECT 49.175 4.695 49.345 7.765 ;
        RECT 48.185 4.695 48.355 7.765 ;
        RECT 45.445 4.7 45.615 7.76 ;
        RECT 43.645 4.93 43.815 7.03 ;
        RECT 42.685 4.93 42.855 7.03 ;
        RECT 40.665 5.425 40.835 7.76 ;
        RECT 40.245 4.93 40.415 7.03 ;
        RECT 39.245 4.93 39.415 7.03 ;
        RECT 38.285 4.93 38.455 7.03 ;
        RECT 35.845 4.93 36.015 7.03 ;
        RECT 18.53 5.425 34.295 7.03 ;
        RECT 32.24 5.425 34.22 7.035 ;
        RECT 33.4 4.695 33.57 7.765 ;
        RECT 32.41 4.695 32.58 7.765 ;
        RECT 29.67 4.7 29.84 7.76 ;
        RECT 27.87 4.93 28.04 7.03 ;
        RECT 26.91 4.93 27.08 7.03 ;
        RECT 24.89 5.425 25.06 7.76 ;
        RECT 24.47 4.93 24.64 7.03 ;
        RECT 23.47 4.93 23.64 7.03 ;
        RECT 22.51 4.93 22.68 7.03 ;
        RECT 20.07 4.93 20.24 7.03 ;
        RECT 2.75 5.425 18.515 7.03 ;
        RECT 16.46 5.425 18.44 7.035 ;
        RECT 17.62 4.695 17.79 7.765 ;
        RECT 16.63 4.695 16.8 7.765 ;
        RECT 13.89 4.7 14.06 7.76 ;
        RECT 12.09 4.93 12.26 7.03 ;
        RECT 11.13 4.93 11.3 7.03 ;
        RECT 9.11 5.425 9.28 7.76 ;
        RECT 8.69 4.93 8.86 7.03 ;
        RECT 7.69 4.93 7.86 7.03 ;
        RECT 6.73 4.93 6.9 7.03 ;
        RECT 4.29 4.93 4.46 7.03 ;
        RECT 0.22 5.53 0.39 7.76 ;
      LAYER met1 ;
        RECT 0 5.53 81.72 7.03 ;
        RECT 2.75 5.43 81.72 7.03 ;
        RECT 65.875 5.425 81.655 7.03 ;
        RECT 79.585 5.425 81.565 7.035 ;
        RECT 66.125 5.275 75.785 7.03 ;
        RECT 50.09 5.425 65.87 7.03 ;
        RECT 63.8 5.425 65.78 7.035 ;
        RECT 50.34 5.275 60 7.03 ;
        RECT 2.75 5.425 50.085 7.03 ;
        RECT 48.015 5.425 49.995 7.035 ;
        RECT 34.555 5.275 44.215 7.03 ;
        RECT 32.24 5.425 34.22 7.035 ;
        RECT 18.78 5.275 28.44 7.03 ;
        RECT 16.46 5.425 18.44 7.035 ;
        RECT 3 5.275 12.66 7.03 ;
      LAYER mcon ;
        RECT 2.34 6.83 2.51 7 ;
        RECT 3.145 5.43 3.315 5.6 ;
        RECT 3.605 5.43 3.775 5.6 ;
        RECT 4.065 5.43 4.235 5.6 ;
        RECT 4.525 5.43 4.695 5.6 ;
        RECT 4.985 5.43 5.155 5.6 ;
        RECT 5.445 5.43 5.615 5.6 ;
        RECT 5.905 5.43 6.075 5.6 ;
        RECT 6.365 5.43 6.535 5.6 ;
        RECT 6.825 5.43 6.995 5.6 ;
        RECT 7.285 5.43 7.455 5.6 ;
        RECT 7.745 5.43 7.915 5.6 ;
        RECT 8.205 5.43 8.375 5.6 ;
        RECT 8.665 5.43 8.835 5.6 ;
        RECT 9.125 5.43 9.295 5.6 ;
        RECT 9.585 5.43 9.755 5.6 ;
        RECT 10.045 5.43 10.215 5.6 ;
        RECT 10.505 5.43 10.675 5.6 ;
        RECT 10.965 5.43 11.135 5.6 ;
        RECT 11.23 6.83 11.4 7 ;
        RECT 11.425 5.43 11.595 5.6 ;
        RECT 11.885 5.43 12.055 5.6 ;
        RECT 12.345 5.43 12.515 5.6 ;
        RECT 16.01 6.83 16.18 7 ;
        RECT 16.01 5.46 16.18 5.63 ;
        RECT 16.71 6.835 16.88 7.005 ;
        RECT 16.71 5.455 16.88 5.625 ;
        RECT 17.7 6.835 17.87 7.005 ;
        RECT 17.7 5.455 17.87 5.625 ;
        RECT 18.925 5.43 19.095 5.6 ;
        RECT 19.385 5.43 19.555 5.6 ;
        RECT 19.845 5.43 20.015 5.6 ;
        RECT 20.305 5.43 20.475 5.6 ;
        RECT 20.765 5.43 20.935 5.6 ;
        RECT 21.225 5.43 21.395 5.6 ;
        RECT 21.685 5.43 21.855 5.6 ;
        RECT 22.145 5.43 22.315 5.6 ;
        RECT 22.605 5.43 22.775 5.6 ;
        RECT 23.065 5.43 23.235 5.6 ;
        RECT 23.525 5.43 23.695 5.6 ;
        RECT 23.985 5.43 24.155 5.6 ;
        RECT 24.445 5.43 24.615 5.6 ;
        RECT 24.905 5.43 25.075 5.6 ;
        RECT 25.365 5.43 25.535 5.6 ;
        RECT 25.825 5.43 25.995 5.6 ;
        RECT 26.285 5.43 26.455 5.6 ;
        RECT 26.745 5.43 26.915 5.6 ;
        RECT 27.01 6.83 27.18 7 ;
        RECT 27.205 5.43 27.375 5.6 ;
        RECT 27.665 5.43 27.835 5.6 ;
        RECT 28.125 5.43 28.295 5.6 ;
        RECT 31.79 6.83 31.96 7 ;
        RECT 31.79 5.46 31.96 5.63 ;
        RECT 32.49 6.835 32.66 7.005 ;
        RECT 32.49 5.455 32.66 5.625 ;
        RECT 33.48 6.835 33.65 7.005 ;
        RECT 33.48 5.455 33.65 5.625 ;
        RECT 34.7 5.43 34.87 5.6 ;
        RECT 35.16 5.43 35.33 5.6 ;
        RECT 35.62 5.43 35.79 5.6 ;
        RECT 36.08 5.43 36.25 5.6 ;
        RECT 36.54 5.43 36.71 5.6 ;
        RECT 37 5.43 37.17 5.6 ;
        RECT 37.46 5.43 37.63 5.6 ;
        RECT 37.92 5.43 38.09 5.6 ;
        RECT 38.38 5.43 38.55 5.6 ;
        RECT 38.84 5.43 39.01 5.6 ;
        RECT 39.3 5.43 39.47 5.6 ;
        RECT 39.76 5.43 39.93 5.6 ;
        RECT 40.22 5.43 40.39 5.6 ;
        RECT 40.68 5.43 40.85 5.6 ;
        RECT 41.14 5.43 41.31 5.6 ;
        RECT 41.6 5.43 41.77 5.6 ;
        RECT 42.06 5.43 42.23 5.6 ;
        RECT 42.52 5.43 42.69 5.6 ;
        RECT 42.785 6.83 42.955 7 ;
        RECT 42.98 5.43 43.15 5.6 ;
        RECT 43.44 5.43 43.61 5.6 ;
        RECT 43.9 5.43 44.07 5.6 ;
        RECT 47.565 6.83 47.735 7 ;
        RECT 47.565 5.46 47.735 5.63 ;
        RECT 48.265 6.835 48.435 7.005 ;
        RECT 48.265 5.455 48.435 5.625 ;
        RECT 49.255 6.835 49.425 7.005 ;
        RECT 49.255 5.455 49.425 5.625 ;
        RECT 50.485 5.43 50.655 5.6 ;
        RECT 50.945 5.43 51.115 5.6 ;
        RECT 51.405 5.43 51.575 5.6 ;
        RECT 51.865 5.43 52.035 5.6 ;
        RECT 52.325 5.43 52.495 5.6 ;
        RECT 52.785 5.43 52.955 5.6 ;
        RECT 53.245 5.43 53.415 5.6 ;
        RECT 53.705 5.43 53.875 5.6 ;
        RECT 54.165 5.43 54.335 5.6 ;
        RECT 54.625 5.43 54.795 5.6 ;
        RECT 55.085 5.43 55.255 5.6 ;
        RECT 55.545 5.43 55.715 5.6 ;
        RECT 56.005 5.43 56.175 5.6 ;
        RECT 56.465 5.43 56.635 5.6 ;
        RECT 56.925 5.43 57.095 5.6 ;
        RECT 57.385 5.43 57.555 5.6 ;
        RECT 57.845 5.43 58.015 5.6 ;
        RECT 58.305 5.43 58.475 5.6 ;
        RECT 58.57 6.83 58.74 7 ;
        RECT 58.765 5.43 58.935 5.6 ;
        RECT 59.225 5.43 59.395 5.6 ;
        RECT 59.685 5.43 59.855 5.6 ;
        RECT 63.35 6.83 63.52 7 ;
        RECT 63.35 5.46 63.52 5.63 ;
        RECT 64.05 6.835 64.22 7.005 ;
        RECT 64.05 5.455 64.22 5.625 ;
        RECT 65.04 6.835 65.21 7.005 ;
        RECT 65.04 5.455 65.21 5.625 ;
        RECT 66.27 5.43 66.44 5.6 ;
        RECT 66.73 5.43 66.9 5.6 ;
        RECT 67.19 5.43 67.36 5.6 ;
        RECT 67.65 5.43 67.82 5.6 ;
        RECT 68.11 5.43 68.28 5.6 ;
        RECT 68.57 5.43 68.74 5.6 ;
        RECT 69.03 5.43 69.2 5.6 ;
        RECT 69.49 5.43 69.66 5.6 ;
        RECT 69.95 5.43 70.12 5.6 ;
        RECT 70.41 5.43 70.58 5.6 ;
        RECT 70.87 5.43 71.04 5.6 ;
        RECT 71.33 5.43 71.5 5.6 ;
        RECT 71.79 5.43 71.96 5.6 ;
        RECT 72.25 5.43 72.42 5.6 ;
        RECT 72.71 5.43 72.88 5.6 ;
        RECT 73.17 5.43 73.34 5.6 ;
        RECT 73.63 5.43 73.8 5.6 ;
        RECT 74.09 5.43 74.26 5.6 ;
        RECT 74.355 6.83 74.525 7 ;
        RECT 74.55 5.43 74.72 5.6 ;
        RECT 75.01 5.43 75.18 5.6 ;
        RECT 75.47 5.43 75.64 5.6 ;
        RECT 79.135 6.83 79.305 7 ;
        RECT 79.135 5.46 79.305 5.63 ;
        RECT 79.835 6.835 80.005 7.005 ;
        RECT 79.835 5.455 80.005 5.625 ;
        RECT 80.825 6.835 80.995 7.005 ;
        RECT 80.825 5.455 80.995 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.03 10.86 81.725 12.445 ;
        RECT 0.03 10.86 81.72 12.46 ;
        RECT 80.745 10.235 80.915 12.46 ;
        RECT 79.755 10.235 79.925 12.46 ;
        RECT 77.015 10.23 77.185 12.46 ;
        RECT 72.235 10.23 72.405 12.46 ;
        RECT 64.96 10.235 65.13 12.46 ;
        RECT 63.97 10.235 64.14 12.46 ;
        RECT 61.23 10.23 61.4 12.46 ;
        RECT 56.45 10.23 56.62 12.46 ;
        RECT 49.175 10.235 49.345 12.46 ;
        RECT 48.185 10.235 48.355 12.46 ;
        RECT 45.445 10.23 45.615 12.46 ;
        RECT 40.665 10.23 40.835 12.46 ;
        RECT 33.4 10.235 33.57 12.46 ;
        RECT 32.41 10.235 32.58 12.46 ;
        RECT 29.67 10.23 29.84 12.46 ;
        RECT 24.89 10.23 25.06 12.46 ;
        RECT 17.62 10.235 17.79 12.46 ;
        RECT 16.63 10.235 16.8 12.46 ;
        RECT 13.89 10.23 14.06 12.46 ;
        RECT 9.11 10.23 9.28 12.46 ;
        RECT 0.22 10.23 0.39 12.46 ;
        RECT 73.24 8.36 73.41 10.31 ;
        RECT 73.185 10.14 73.355 10.59 ;
        RECT 73.185 7.3 73.355 8.53 ;
        RECT 57.455 8.36 57.625 10.31 ;
        RECT 57.4 10.14 57.57 10.59 ;
        RECT 57.4 7.3 57.57 8.53 ;
        RECT 41.67 8.36 41.84 10.31 ;
        RECT 41.615 10.14 41.785 10.59 ;
        RECT 41.615 7.3 41.785 8.53 ;
        RECT 25.895 8.36 26.065 10.31 ;
        RECT 25.84 10.14 26.01 10.59 ;
        RECT 25.84 7.3 26.01 8.53 ;
        RECT 10.115 8.36 10.285 10.31 ;
        RECT 10.06 10.14 10.23 10.59 ;
        RECT 10.06 7.3 10.23 8.53 ;
      LAYER met1 ;
        RECT 0.025 10.86 81.725 12.445 ;
        RECT 0.025 10.86 81.72 12.46 ;
        RECT 73.18 8.57 73.47 8.8 ;
        RECT 72.81 8.6 73.47 8.77 ;
        RECT 72.81 8.6 72.98 12.46 ;
        RECT 57.395 8.57 57.685 8.8 ;
        RECT 57.025 8.6 57.685 8.77 ;
        RECT 57.025 8.6 57.195 12.46 ;
        RECT 41.61 8.57 41.9 8.8 ;
        RECT 41.24 8.6 41.9 8.77 ;
        RECT 41.24 8.6 41.41 12.46 ;
        RECT 25.835 8.57 26.125 8.8 ;
        RECT 25.465 8.6 26.125 8.77 ;
        RECT 25.465 8.6 25.635 12.46 ;
        RECT 10.055 8.57 10.345 8.8 ;
        RECT 9.685 8.6 10.345 8.77 ;
        RECT 9.685 8.6 9.855 12.46 ;
      LAYER mcon ;
        RECT 0.3 10.89 0.47 11.06 ;
        RECT 0.98 10.89 1.15 11.06 ;
        RECT 1.66 10.89 1.83 11.06 ;
        RECT 2.34 10.89 2.51 11.06 ;
        RECT 9.19 10.89 9.36 11.06 ;
        RECT 9.87 10.89 10.04 11.06 ;
        RECT 10.115 8.6 10.285 8.77 ;
        RECT 10.55 10.89 10.72 11.06 ;
        RECT 11.23 10.89 11.4 11.06 ;
        RECT 13.97 10.89 14.14 11.06 ;
        RECT 14.65 10.89 14.82 11.06 ;
        RECT 15.33 10.89 15.5 11.06 ;
        RECT 16.01 10.89 16.18 11.06 ;
        RECT 16.71 10.895 16.88 11.065 ;
        RECT 17.7 10.895 17.87 11.065 ;
        RECT 24.97 10.89 25.14 11.06 ;
        RECT 25.65 10.89 25.82 11.06 ;
        RECT 25.895 8.6 26.065 8.77 ;
        RECT 26.33 10.89 26.5 11.06 ;
        RECT 27.01 10.89 27.18 11.06 ;
        RECT 29.75 10.89 29.92 11.06 ;
        RECT 30.43 10.89 30.6 11.06 ;
        RECT 31.11 10.89 31.28 11.06 ;
        RECT 31.79 10.89 31.96 11.06 ;
        RECT 32.49 10.895 32.66 11.065 ;
        RECT 33.48 10.895 33.65 11.065 ;
        RECT 40.745 10.89 40.915 11.06 ;
        RECT 41.425 10.89 41.595 11.06 ;
        RECT 41.67 8.6 41.84 8.77 ;
        RECT 42.105 10.89 42.275 11.06 ;
        RECT 42.785 10.89 42.955 11.06 ;
        RECT 45.525 10.89 45.695 11.06 ;
        RECT 46.205 10.89 46.375 11.06 ;
        RECT 46.885 10.89 47.055 11.06 ;
        RECT 47.565 10.89 47.735 11.06 ;
        RECT 48.265 10.895 48.435 11.065 ;
        RECT 49.255 10.895 49.425 11.065 ;
        RECT 56.53 10.89 56.7 11.06 ;
        RECT 57.21 10.89 57.38 11.06 ;
        RECT 57.455 8.6 57.625 8.77 ;
        RECT 57.89 10.89 58.06 11.06 ;
        RECT 58.57 10.89 58.74 11.06 ;
        RECT 61.31 10.89 61.48 11.06 ;
        RECT 61.99 10.89 62.16 11.06 ;
        RECT 62.67 10.89 62.84 11.06 ;
        RECT 63.35 10.89 63.52 11.06 ;
        RECT 64.05 10.895 64.22 11.065 ;
        RECT 65.04 10.895 65.21 11.065 ;
        RECT 72.315 10.89 72.485 11.06 ;
        RECT 72.995 10.89 73.165 11.06 ;
        RECT 73.24 8.6 73.41 8.77 ;
        RECT 73.675 10.89 73.845 11.06 ;
        RECT 74.355 10.89 74.525 11.06 ;
        RECT 77.095 10.89 77.265 11.06 ;
        RECT 77.775 10.89 77.945 11.06 ;
        RECT 78.455 10.89 78.625 11.06 ;
        RECT 79.135 10.89 79.305 11.06 ;
        RECT 79.835 10.895 80.005 11.065 ;
        RECT 80.825 10.895 80.995 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 73.515 9.325 73.885 9.695 ;
      RECT 73.555 9.005 73.89 9.37 ;
      RECT 73.555 9.005 73.94 9.315 ;
      RECT 73.555 9.005 76.345 9.31 ;
      RECT 76.04 4.145 76.345 9.31 ;
      RECT 76.005 4.145 76.375 4.515 ;
      RECT 75.265 2.11 75.57 5.315 ;
      RECT 75.015 4.27 75.57 5 ;
      RECT 75.225 2.11 75.595 2.48 ;
      RECT 71.375 3.145 71.705 4.04 ;
      RECT 70.495 3.31 70.825 4.04 ;
      RECT 71.37 3.145 71.74 3.945 ;
      RECT 74.535 3.145 74.865 3.875 ;
      RECT 74.495 3.03 74.675 3.68 ;
      RECT 70.505 3.145 74.865 3.515 ;
      RECT 70.995 4.83 71.325 5.16 ;
      RECT 69.79 4.845 71.325 5.145 ;
      RECT 69.79 3.725 70.09 5.145 ;
      RECT 69.535 3.71 69.865 4.04 ;
      RECT 57.73 9.325 58.1 9.695 ;
      RECT 57.77 9.005 58.105 9.37 ;
      RECT 57.77 9.005 58.155 9.315 ;
      RECT 57.77 9.005 60.56 9.31 ;
      RECT 60.255 4.145 60.56 9.31 ;
      RECT 60.22 4.145 60.59 4.515 ;
      RECT 59.48 2.11 59.785 5.315 ;
      RECT 59.23 4.27 59.785 5 ;
      RECT 59.44 2.11 59.81 2.48 ;
      RECT 55.59 3.145 55.92 4.04 ;
      RECT 54.71 3.31 55.04 4.04 ;
      RECT 55.585 3.145 55.955 3.945 ;
      RECT 58.75 3.145 59.08 3.875 ;
      RECT 58.71 3.03 58.89 3.68 ;
      RECT 54.72 3.145 59.08 3.515 ;
      RECT 55.21 4.83 55.54 5.16 ;
      RECT 54.005 4.845 55.54 5.145 ;
      RECT 54.005 3.725 54.305 5.145 ;
      RECT 53.75 3.71 54.08 4.04 ;
      RECT 41.945 9.325 42.315 9.695 ;
      RECT 41.985 9.005 42.32 9.37 ;
      RECT 41.985 9.005 42.37 9.315 ;
      RECT 41.985 9.005 44.775 9.31 ;
      RECT 44.47 4.145 44.775 9.31 ;
      RECT 44.435 4.145 44.805 4.515 ;
      RECT 43.695 2.11 44 5.315 ;
      RECT 43.445 4.27 44 5 ;
      RECT 43.655 2.11 44.025 2.48 ;
      RECT 39.805 3.145 40.135 4.04 ;
      RECT 38.925 3.31 39.255 4.04 ;
      RECT 39.8 3.145 40.17 3.945 ;
      RECT 42.965 3.145 43.295 3.875 ;
      RECT 42.925 3.03 43.105 3.68 ;
      RECT 38.935 3.145 43.295 3.515 ;
      RECT 39.425 4.83 39.755 5.16 ;
      RECT 38.22 4.845 39.755 5.145 ;
      RECT 38.22 3.725 38.52 5.145 ;
      RECT 37.965 3.71 38.295 4.04 ;
      RECT 26.17 9.325 26.54 9.695 ;
      RECT 26.21 9.005 26.545 9.37 ;
      RECT 26.21 9.005 26.595 9.315 ;
      RECT 26.21 9.005 29 9.31 ;
      RECT 28.695 4.145 29 9.31 ;
      RECT 28.66 4.145 29.03 4.515 ;
      RECT 27.92 2.11 28.225 5.315 ;
      RECT 27.67 4.27 28.225 5 ;
      RECT 27.88 2.11 28.25 2.48 ;
      RECT 24.03 3.145 24.36 4.04 ;
      RECT 23.15 3.31 23.48 4.04 ;
      RECT 24.025 3.145 24.395 3.945 ;
      RECT 27.19 3.145 27.52 3.875 ;
      RECT 27.15 3.03 27.33 3.68 ;
      RECT 23.16 3.145 27.52 3.515 ;
      RECT 23.65 4.83 23.98 5.16 ;
      RECT 22.445 4.845 23.98 5.145 ;
      RECT 22.445 3.725 22.745 5.145 ;
      RECT 22.19 3.71 22.52 4.04 ;
      RECT 10.39 9.325 10.76 9.695 ;
      RECT 10.43 9.005 10.765 9.37 ;
      RECT 10.43 9.005 10.815 9.315 ;
      RECT 10.43 9.005 13.22 9.31 ;
      RECT 12.915 4.145 13.22 9.31 ;
      RECT 12.88 4.145 13.25 4.515 ;
      RECT 12.14 2.11 12.445 5.315 ;
      RECT 11.89 4.27 12.445 5 ;
      RECT 12.1 2.11 12.47 2.48 ;
      RECT 8.25 3.145 8.58 4.04 ;
      RECT 7.37 3.31 7.7 4.04 ;
      RECT 8.245 3.145 8.615 3.945 ;
      RECT 11.41 3.145 11.74 3.875 ;
      RECT 11.37 3.03 11.55 3.68 ;
      RECT 7.38 3.145 11.74 3.515 ;
      RECT 7.87 4.83 8.2 5.16 ;
      RECT 6.665 4.845 8.2 5.145 ;
      RECT 6.665 3.725 6.965 5.145 ;
      RECT 6.41 3.71 6.74 4.04 ;
      RECT 72.935 3.87 73.265 4.6 ;
      RECT 68.815 3.71 69.145 4.44 ;
      RECT 67.815 3.15 68.145 3.88 ;
      RECT 66.375 3.87 66.705 4.6 ;
      RECT 57.15 3.87 57.48 4.6 ;
      RECT 53.03 3.71 53.36 4.44 ;
      RECT 52.03 3.15 52.36 3.88 ;
      RECT 50.59 3.87 50.92 4.6 ;
      RECT 41.365 3.87 41.695 4.6 ;
      RECT 37.245 3.71 37.575 4.44 ;
      RECT 36.245 3.15 36.575 3.88 ;
      RECT 34.805 3.87 35.135 4.6 ;
      RECT 25.59 3.87 25.92 4.6 ;
      RECT 21.47 3.71 21.8 4.44 ;
      RECT 20.47 3.15 20.8 3.88 ;
      RECT 19.03 3.87 19.36 4.6 ;
      RECT 9.81 3.87 10.14 4.6 ;
      RECT 5.69 3.71 6.02 4.44 ;
      RECT 4.69 3.15 5.02 3.88 ;
      RECT 3.25 3.87 3.58 4.6 ;
    LAYER via2 ;
      RECT 76.09 4.23 76.29 4.43 ;
      RECT 75.31 2.195 75.51 2.395 ;
      RECT 75.08 4.335 75.28 4.535 ;
      RECT 74.6 3.61 74.8 3.81 ;
      RECT 73.6 9.41 73.8 9.61 ;
      RECT 73 4.335 73.2 4.535 ;
      RECT 71.44 3.775 71.64 3.975 ;
      RECT 71.06 4.895 71.26 5.095 ;
      RECT 70.56 3.775 70.76 3.975 ;
      RECT 69.6 3.775 69.8 3.975 ;
      RECT 68.88 3.775 69.08 3.975 ;
      RECT 67.88 3.215 68.08 3.415 ;
      RECT 66.44 4.335 66.64 4.535 ;
      RECT 60.305 4.23 60.505 4.43 ;
      RECT 59.525 2.195 59.725 2.395 ;
      RECT 59.295 4.335 59.495 4.535 ;
      RECT 58.815 3.61 59.015 3.81 ;
      RECT 57.815 9.41 58.015 9.61 ;
      RECT 57.215 4.335 57.415 4.535 ;
      RECT 55.655 3.775 55.855 3.975 ;
      RECT 55.275 4.895 55.475 5.095 ;
      RECT 54.775 3.775 54.975 3.975 ;
      RECT 53.815 3.775 54.015 3.975 ;
      RECT 53.095 3.775 53.295 3.975 ;
      RECT 52.095 3.215 52.295 3.415 ;
      RECT 50.655 4.335 50.855 4.535 ;
      RECT 44.52 4.23 44.72 4.43 ;
      RECT 43.74 2.195 43.94 2.395 ;
      RECT 43.51 4.335 43.71 4.535 ;
      RECT 43.03 3.61 43.23 3.81 ;
      RECT 42.03 9.41 42.23 9.61 ;
      RECT 41.43 4.335 41.63 4.535 ;
      RECT 39.87 3.775 40.07 3.975 ;
      RECT 39.49 4.895 39.69 5.095 ;
      RECT 38.99 3.775 39.19 3.975 ;
      RECT 38.03 3.775 38.23 3.975 ;
      RECT 37.31 3.775 37.51 3.975 ;
      RECT 36.31 3.215 36.51 3.415 ;
      RECT 34.87 4.335 35.07 4.535 ;
      RECT 28.745 4.23 28.945 4.43 ;
      RECT 27.965 2.195 28.165 2.395 ;
      RECT 27.735 4.335 27.935 4.535 ;
      RECT 27.255 3.61 27.455 3.81 ;
      RECT 26.255 9.41 26.455 9.61 ;
      RECT 25.655 4.335 25.855 4.535 ;
      RECT 24.095 3.775 24.295 3.975 ;
      RECT 23.715 4.895 23.915 5.095 ;
      RECT 23.215 3.775 23.415 3.975 ;
      RECT 22.255 3.775 22.455 3.975 ;
      RECT 21.535 3.775 21.735 3.975 ;
      RECT 20.535 3.215 20.735 3.415 ;
      RECT 19.095 4.335 19.295 4.535 ;
      RECT 12.965 4.23 13.165 4.43 ;
      RECT 12.185 2.195 12.385 2.395 ;
      RECT 11.955 4.335 12.155 4.535 ;
      RECT 11.475 3.61 11.675 3.81 ;
      RECT 10.475 9.41 10.675 9.61 ;
      RECT 9.875 4.335 10.075 4.535 ;
      RECT 8.315 3.775 8.515 3.975 ;
      RECT 7.935 4.895 8.135 5.095 ;
      RECT 7.435 3.775 7.635 3.975 ;
      RECT 6.475 3.775 6.675 3.975 ;
      RECT 5.755 3.775 5.955 3.975 ;
      RECT 4.755 3.215 4.955 3.415 ;
      RECT 3.315 4.335 3.515 4.535 ;
    LAYER met2 ;
      RECT 1.23 10.685 81.35 10.855 ;
      RECT 81.18 9.56 81.35 10.855 ;
      RECT 1.23 8.54 1.4 10.855 ;
      RECT 81.15 9.56 81.5 9.91 ;
      RECT 1.165 8.54 1.455 8.89 ;
      RECT 77.99 8.505 78.31 8.83 ;
      RECT 78.02 7.98 78.19 8.83 ;
      RECT 78.02 7.98 78.195 8.33 ;
      RECT 78.02 7.98 78.995 8.155 ;
      RECT 78.82 3.26 78.995 8.155 ;
      RECT 78.765 3.26 79.115 3.61 ;
      RECT 78.79 8.94 79.115 9.265 ;
      RECT 77.675 9.03 79.115 9.2 ;
      RECT 77.675 3.69 77.835 9.2 ;
      RECT 77.99 3.66 78.31 3.98 ;
      RECT 77.675 3.69 78.31 3.86 ;
      RECT 67.76 3.215 68.02 3.475 ;
      RECT 67.815 3.175 68.12 3.455 ;
      RECT 67.815 2.715 67.99 3.475 ;
      RECT 76.33 2.635 76.68 2.985 ;
      RECT 67.815 2.715 76.68 2.89 ;
      RECT 76.005 4.145 76.375 4.515 ;
      RECT 76.09 3.53 76.26 4.515 ;
      RECT 72.11 3.75 72.345 4.01 ;
      RECT 75.255 3.53 75.42 3.79 ;
      RECT 75.16 3.52 75.175 3.79 ;
      RECT 75.255 3.53 76.26 3.71 ;
      RECT 73.76 3.09 73.8 3.23 ;
      RECT 75.175 3.525 75.255 3.79 ;
      RECT 75.12 3.52 75.16 3.756 ;
      RECT 75.106 3.52 75.12 3.756 ;
      RECT 75.02 3.525 75.106 3.758 ;
      RECT 74.975 3.532 75.02 3.76 ;
      RECT 74.945 3.532 74.975 3.762 ;
      RECT 74.92 3.527 74.945 3.764 ;
      RECT 74.89 3.523 74.92 3.773 ;
      RECT 74.88 3.52 74.89 3.785 ;
      RECT 74.875 3.52 74.88 3.793 ;
      RECT 74.87 3.52 74.875 3.798 ;
      RECT 74.86 3.519 74.87 3.808 ;
      RECT 74.855 3.518 74.86 3.818 ;
      RECT 74.84 3.517 74.855 3.823 ;
      RECT 74.812 3.514 74.84 3.85 ;
      RECT 74.726 3.506 74.812 3.85 ;
      RECT 74.64 3.495 74.726 3.85 ;
      RECT 74.6 3.48 74.64 3.85 ;
      RECT 74.56 3.454 74.6 3.85 ;
      RECT 74.555 3.436 74.56 3.662 ;
      RECT 74.545 3.432 74.555 3.652 ;
      RECT 74.53 3.422 74.545 3.639 ;
      RECT 74.51 3.406 74.53 3.624 ;
      RECT 74.495 3.391 74.51 3.609 ;
      RECT 74.485 3.38 74.495 3.599 ;
      RECT 74.46 3.364 74.485 3.588 ;
      RECT 74.455 3.351 74.46 3.578 ;
      RECT 74.45 3.347 74.455 3.573 ;
      RECT 74.395 3.333 74.45 3.551 ;
      RECT 74.356 3.314 74.395 3.515 ;
      RECT 74.27 3.288 74.356 3.468 ;
      RECT 74.266 3.27 74.27 3.434 ;
      RECT 74.18 3.251 74.266 3.412 ;
      RECT 74.175 3.233 74.18 3.39 ;
      RECT 74.17 3.231 74.175 3.388 ;
      RECT 74.16 3.23 74.17 3.383 ;
      RECT 74.1 3.217 74.16 3.369 ;
      RECT 74.055 3.195 74.1 3.348 ;
      RECT 73.995 3.172 74.055 3.327 ;
      RECT 73.931 3.147 73.995 3.302 ;
      RECT 73.845 3.117 73.931 3.271 ;
      RECT 73.83 3.097 73.845 3.25 ;
      RECT 73.8 3.092 73.83 3.241 ;
      RECT 73.747 3.09 73.76 3.23 ;
      RECT 73.661 3.09 73.747 3.232 ;
      RECT 73.575 3.09 73.661 3.234 ;
      RECT 73.555 3.09 73.575 3.238 ;
      RECT 73.51 3.092 73.555 3.249 ;
      RECT 73.47 3.102 73.51 3.265 ;
      RECT 73.466 3.111 73.47 3.273 ;
      RECT 73.38 3.131 73.466 3.289 ;
      RECT 73.37 3.15 73.38 3.307 ;
      RECT 73.365 3.152 73.37 3.31 ;
      RECT 73.355 3.156 73.365 3.313 ;
      RECT 73.335 3.161 73.355 3.323 ;
      RECT 73.305 3.171 73.335 3.343 ;
      RECT 73.3 3.178 73.305 3.357 ;
      RECT 73.29 3.182 73.3 3.364 ;
      RECT 73.275 3.19 73.29 3.375 ;
      RECT 73.265 3.2 73.275 3.386 ;
      RECT 73.255 3.207 73.265 3.394 ;
      RECT 73.23 3.22 73.255 3.409 ;
      RECT 73.166 3.256 73.23 3.448 ;
      RECT 73.08 3.319 73.166 3.512 ;
      RECT 73.045 3.37 73.08 3.565 ;
      RECT 73.04 3.387 73.045 3.582 ;
      RECT 73.025 3.396 73.04 3.589 ;
      RECT 73.005 3.411 73.025 3.603 ;
      RECT 73 3.422 73.005 3.613 ;
      RECT 72.98 3.435 73 3.623 ;
      RECT 72.975 3.445 72.98 3.633 ;
      RECT 72.96 3.45 72.975 3.642 ;
      RECT 72.95 3.46 72.96 3.653 ;
      RECT 72.92 3.477 72.95 3.67 ;
      RECT 72.91 3.495 72.92 3.688 ;
      RECT 72.895 3.506 72.91 3.699 ;
      RECT 72.855 3.53 72.895 3.715 ;
      RECT 72.82 3.564 72.855 3.732 ;
      RECT 72.79 3.587 72.82 3.744 ;
      RECT 72.775 3.597 72.79 3.753 ;
      RECT 72.735 3.607 72.775 3.764 ;
      RECT 72.715 3.618 72.735 3.776 ;
      RECT 72.71 3.622 72.715 3.783 ;
      RECT 72.695 3.626 72.71 3.788 ;
      RECT 72.685 3.631 72.695 3.793 ;
      RECT 72.68 3.634 72.685 3.796 ;
      RECT 72.65 3.64 72.68 3.803 ;
      RECT 72.615 3.65 72.65 3.817 ;
      RECT 72.555 3.665 72.615 3.837 ;
      RECT 72.5 3.685 72.555 3.861 ;
      RECT 72.471 3.7 72.5 3.879 ;
      RECT 72.385 3.72 72.471 3.904 ;
      RECT 72.38 3.735 72.385 3.924 ;
      RECT 72.37 3.738 72.38 3.925 ;
      RECT 72.345 3.745 72.37 4.01 ;
      RECT 75.04 4.238 75.32 4.575 ;
      RECT 75.04 4.248 75.325 4.533 ;
      RECT 75.04 4.257 75.33 4.43 ;
      RECT 75.04 4.272 75.335 4.298 ;
      RECT 75.04 4.1 75.3 4.575 ;
      RECT 65.34 8.94 65.69 9.29 ;
      RECT 74.165 8.895 74.515 9.245 ;
      RECT 65.34 8.97 74.515 9.17 ;
      RECT 72.76 4.98 72.77 5.17 ;
      RECT 71.02 4.855 71.3 5.135 ;
      RECT 74.065 3.795 74.07 4.28 ;
      RECT 73.96 3.795 74.02 4.055 ;
      RECT 74.285 4.765 74.29 4.84 ;
      RECT 74.275 4.632 74.285 4.875 ;
      RECT 74.265 4.467 74.275 4.896 ;
      RECT 74.26 4.337 74.265 4.912 ;
      RECT 74.25 4.227 74.26 4.928 ;
      RECT 74.245 4.126 74.25 4.945 ;
      RECT 74.24 4.108 74.245 4.955 ;
      RECT 74.235 4.09 74.24 4.965 ;
      RECT 74.225 4.065 74.235 4.98 ;
      RECT 74.22 4.045 74.225 4.995 ;
      RECT 74.2 3.795 74.22 5.02 ;
      RECT 74.185 3.795 74.2 5.053 ;
      RECT 74.155 3.795 74.185 5.075 ;
      RECT 74.135 3.795 74.155 5.089 ;
      RECT 74.115 3.795 74.135 4.605 ;
      RECT 74.13 4.672 74.135 5.094 ;
      RECT 74.125 4.702 74.13 5.096 ;
      RECT 74.12 4.715 74.125 5.099 ;
      RECT 74.115 4.725 74.12 5.103 ;
      RECT 74.11 3.795 74.115 4.523 ;
      RECT 74.11 4.735 74.115 5.105 ;
      RECT 74.105 3.795 74.11 4.5 ;
      RECT 74.095 4.757 74.11 5.105 ;
      RECT 74.09 3.795 74.105 4.445 ;
      RECT 74.085 4.782 74.095 5.105 ;
      RECT 74.085 3.795 74.09 4.39 ;
      RECT 74.075 3.795 74.085 4.338 ;
      RECT 74.08 4.795 74.085 5.106 ;
      RECT 74.075 4.807 74.08 5.107 ;
      RECT 74.07 3.795 74.075 4.298 ;
      RECT 74.07 4.82 74.075 5.108 ;
      RECT 74.055 4.835 74.07 5.109 ;
      RECT 74.06 3.795 74.065 4.26 ;
      RECT 74.055 3.795 74.06 4.225 ;
      RECT 74.05 3.795 74.055 4.2 ;
      RECT 74.045 4.862 74.055 5.111 ;
      RECT 74.04 3.795 74.05 4.158 ;
      RECT 74.04 4.88 74.045 5.112 ;
      RECT 74.035 3.795 74.04 4.118 ;
      RECT 74.035 4.887 74.04 5.113 ;
      RECT 74.03 3.795 74.035 4.09 ;
      RECT 74.025 4.905 74.035 5.114 ;
      RECT 74.02 3.795 74.03 4.07 ;
      RECT 74.015 4.925 74.025 5.116 ;
      RECT 74.005 4.942 74.015 5.117 ;
      RECT 73.97 4.965 74.005 5.12 ;
      RECT 73.915 4.983 73.97 5.126 ;
      RECT 73.829 4.991 73.915 5.135 ;
      RECT 73.743 5.002 73.829 5.146 ;
      RECT 73.657 5.012 73.743 5.157 ;
      RECT 73.571 5.022 73.657 5.169 ;
      RECT 73.485 5.032 73.571 5.18 ;
      RECT 73.465 5.038 73.485 5.186 ;
      RECT 73.385 5.04 73.465 5.19 ;
      RECT 73.38 5.039 73.385 5.195 ;
      RECT 73.372 5.038 73.38 5.195 ;
      RECT 73.286 5.034 73.372 5.193 ;
      RECT 73.2 5.026 73.286 5.19 ;
      RECT 73.114 5.017 73.2 5.186 ;
      RECT 73.028 5.009 73.114 5.183 ;
      RECT 72.942 5.001 73.028 5.179 ;
      RECT 72.856 4.992 72.942 5.176 ;
      RECT 72.77 4.984 72.856 5.172 ;
      RECT 72.715 4.977 72.76 5.17 ;
      RECT 72.63 4.97 72.715 5.168 ;
      RECT 72.556 4.962 72.63 5.164 ;
      RECT 72.47 4.954 72.556 5.161 ;
      RECT 72.467 4.95 72.47 5.159 ;
      RECT 72.381 4.946 72.467 5.158 ;
      RECT 72.295 4.938 72.381 5.155 ;
      RECT 72.21 4.933 72.295 5.152 ;
      RECT 72.124 4.93 72.21 5.149 ;
      RECT 72.038 4.928 72.124 5.146 ;
      RECT 71.952 4.925 72.038 5.143 ;
      RECT 71.866 4.922 71.952 5.14 ;
      RECT 71.78 4.919 71.866 5.137 ;
      RECT 71.704 4.917 71.78 5.134 ;
      RECT 71.618 4.914 71.704 5.131 ;
      RECT 71.532 4.911 71.618 5.129 ;
      RECT 71.446 4.909 71.532 5.126 ;
      RECT 71.36 4.906 71.446 5.123 ;
      RECT 71.3 4.897 71.36 5.121 ;
      RECT 73.81 4.515 73.885 4.775 ;
      RECT 73.79 4.495 73.795 4.775 ;
      RECT 73.11 4.28 73.215 4.575 ;
      RECT 67.555 4.255 67.625 4.515 ;
      RECT 73.45 4.13 73.455 4.501 ;
      RECT 73.44 4.185 73.445 4.501 ;
      RECT 73.745 3.355 73.805 3.615 ;
      RECT 73.8 4.51 73.81 4.775 ;
      RECT 73.795 4.5 73.8 4.775 ;
      RECT 73.715 4.447 73.79 4.775 ;
      RECT 73.74 3.355 73.745 3.635 ;
      RECT 73.73 3.355 73.74 3.655 ;
      RECT 73.715 3.355 73.73 3.685 ;
      RECT 73.7 3.355 73.715 3.728 ;
      RECT 73.695 4.39 73.715 4.775 ;
      RECT 73.685 3.355 73.7 3.765 ;
      RECT 73.68 4.37 73.695 4.775 ;
      RECT 73.68 3.355 73.685 3.788 ;
      RECT 73.67 3.355 73.68 3.813 ;
      RECT 73.64 4.337 73.68 4.775 ;
      RECT 73.645 3.355 73.67 3.863 ;
      RECT 73.64 3.355 73.645 3.918 ;
      RECT 73.635 3.355 73.64 3.96 ;
      RECT 73.625 4.3 73.64 4.775 ;
      RECT 73.63 3.355 73.635 4.003 ;
      RECT 73.625 3.355 73.63 4.068 ;
      RECT 73.62 3.355 73.625 4.09 ;
      RECT 73.62 4.288 73.625 4.64 ;
      RECT 73.615 3.355 73.62 4.158 ;
      RECT 73.615 4.28 73.62 4.623 ;
      RECT 73.61 3.355 73.615 4.203 ;
      RECT 73.605 4.262 73.615 4.6 ;
      RECT 73.605 3.355 73.61 4.24 ;
      RECT 73.595 3.355 73.605 4.58 ;
      RECT 73.59 3.355 73.595 4.563 ;
      RECT 73.585 3.355 73.59 4.548 ;
      RECT 73.58 3.355 73.585 4.533 ;
      RECT 73.56 3.355 73.58 4.523 ;
      RECT 73.555 3.355 73.56 4.513 ;
      RECT 73.545 3.355 73.555 4.509 ;
      RECT 73.54 3.632 73.545 4.508 ;
      RECT 73.535 3.655 73.54 4.507 ;
      RECT 73.53 3.685 73.535 4.506 ;
      RECT 73.525 3.712 73.53 4.505 ;
      RECT 73.52 3.74 73.525 4.505 ;
      RECT 73.515 3.767 73.52 4.505 ;
      RECT 73.51 3.787 73.515 4.505 ;
      RECT 73.505 3.815 73.51 4.505 ;
      RECT 73.495 3.857 73.505 4.505 ;
      RECT 73.485 3.902 73.495 4.504 ;
      RECT 73.48 3.955 73.485 4.503 ;
      RECT 73.475 3.987 73.48 4.502 ;
      RECT 73.47 4.007 73.475 4.501 ;
      RECT 73.465 4.045 73.47 4.501 ;
      RECT 73.46 4.067 73.465 4.501 ;
      RECT 73.455 4.092 73.46 4.501 ;
      RECT 73.445 4.157 73.45 4.501 ;
      RECT 73.43 4.217 73.44 4.501 ;
      RECT 73.415 4.227 73.43 4.501 ;
      RECT 73.395 4.237 73.415 4.501 ;
      RECT 73.365 4.242 73.395 4.498 ;
      RECT 73.305 4.252 73.365 4.495 ;
      RECT 73.285 4.261 73.305 4.5 ;
      RECT 73.26 4.267 73.285 4.513 ;
      RECT 73.24 4.272 73.26 4.528 ;
      RECT 73.215 4.277 73.24 4.575 ;
      RECT 73.086 4.279 73.11 4.575 ;
      RECT 73 4.274 73.086 4.575 ;
      RECT 72.96 4.271 73 4.575 ;
      RECT 72.91 4.273 72.96 4.555 ;
      RECT 72.88 4.277 72.91 4.555 ;
      RECT 72.801 4.287 72.88 4.555 ;
      RECT 72.715 4.302 72.801 4.556 ;
      RECT 72.665 4.312 72.715 4.557 ;
      RECT 72.657 4.315 72.665 4.557 ;
      RECT 72.571 4.317 72.657 4.558 ;
      RECT 72.485 4.321 72.571 4.558 ;
      RECT 72.399 4.325 72.485 4.559 ;
      RECT 72.313 4.328 72.399 4.56 ;
      RECT 72.227 4.332 72.313 4.56 ;
      RECT 72.141 4.336 72.227 4.561 ;
      RECT 72.055 4.339 72.141 4.562 ;
      RECT 71.969 4.343 72.055 4.562 ;
      RECT 71.883 4.347 71.969 4.563 ;
      RECT 71.797 4.351 71.883 4.564 ;
      RECT 71.711 4.354 71.797 4.564 ;
      RECT 71.625 4.358 71.711 4.565 ;
      RECT 71.595 4.36 71.625 4.565 ;
      RECT 71.509 4.363 71.595 4.566 ;
      RECT 71.423 4.367 71.509 4.567 ;
      RECT 71.337 4.371 71.423 4.568 ;
      RECT 71.251 4.374 71.337 4.568 ;
      RECT 71.165 4.378 71.251 4.569 ;
      RECT 71.13 4.383 71.165 4.57 ;
      RECT 71.075 4.393 71.13 4.577 ;
      RECT 71.05 4.405 71.075 4.587 ;
      RECT 71.015 4.418 71.05 4.595 ;
      RECT 70.975 4.435 71.015 4.618 ;
      RECT 70.955 4.448 70.975 4.645 ;
      RECT 70.925 4.46 70.955 4.673 ;
      RECT 70.92 4.468 70.925 4.693 ;
      RECT 70.915 4.471 70.92 4.703 ;
      RECT 70.865 4.483 70.915 4.737 ;
      RECT 70.855 4.498 70.865 4.77 ;
      RECT 70.845 4.504 70.855 4.783 ;
      RECT 70.835 4.511 70.845 4.795 ;
      RECT 70.81 4.524 70.835 4.813 ;
      RECT 70.795 4.539 70.81 4.835 ;
      RECT 70.785 4.547 70.795 4.851 ;
      RECT 70.77 4.556 70.785 4.866 ;
      RECT 70.76 4.566 70.77 4.88 ;
      RECT 70.741 4.579 70.76 4.897 ;
      RECT 70.655 4.624 70.741 4.962 ;
      RECT 70.64 4.669 70.655 5.02 ;
      RECT 70.635 4.678 70.64 5.033 ;
      RECT 70.625 4.685 70.635 5.038 ;
      RECT 70.62 4.69 70.625 5.042 ;
      RECT 70.6 4.7 70.62 5.049 ;
      RECT 70.575 4.72 70.6 5.063 ;
      RECT 70.54 4.745 70.575 5.083 ;
      RECT 70.525 4.768 70.54 5.098 ;
      RECT 70.515 4.778 70.525 5.103 ;
      RECT 70.505 4.786 70.515 5.11 ;
      RECT 70.495 4.795 70.505 5.116 ;
      RECT 70.475 4.807 70.495 5.118 ;
      RECT 70.465 4.82 70.475 5.12 ;
      RECT 70.44 4.835 70.465 5.123 ;
      RECT 70.42 4.852 70.44 5.127 ;
      RECT 70.38 4.88 70.42 5.133 ;
      RECT 70.315 4.927 70.38 5.142 ;
      RECT 70.3 4.96 70.315 5.15 ;
      RECT 70.295 4.967 70.3 5.152 ;
      RECT 70.245 4.992 70.295 5.157 ;
      RECT 70.23 5.016 70.245 5.164 ;
      RECT 70.18 5.021 70.23 5.165 ;
      RECT 70.094 5.025 70.18 5.165 ;
      RECT 70.008 5.025 70.094 5.165 ;
      RECT 69.922 5.025 70.008 5.166 ;
      RECT 69.836 5.025 69.922 5.166 ;
      RECT 69.75 5.025 69.836 5.166 ;
      RECT 69.684 5.025 69.75 5.166 ;
      RECT 69.598 5.025 69.684 5.167 ;
      RECT 69.512 5.025 69.598 5.167 ;
      RECT 69.426 5.026 69.512 5.168 ;
      RECT 69.34 5.026 69.426 5.168 ;
      RECT 69.254 5.026 69.34 5.168 ;
      RECT 69.168 5.026 69.254 5.169 ;
      RECT 69.082 5.026 69.168 5.169 ;
      RECT 68.996 5.027 69.082 5.17 ;
      RECT 68.91 5.027 68.996 5.17 ;
      RECT 68.89 5.027 68.91 5.17 ;
      RECT 68.804 5.027 68.89 5.17 ;
      RECT 68.718 5.027 68.804 5.17 ;
      RECT 68.632 5.028 68.718 5.17 ;
      RECT 68.546 5.028 68.632 5.17 ;
      RECT 68.46 5.028 68.546 5.17 ;
      RECT 68.374 5.029 68.46 5.17 ;
      RECT 68.288 5.029 68.374 5.17 ;
      RECT 68.202 5.029 68.288 5.17 ;
      RECT 68.116 5.029 68.202 5.17 ;
      RECT 68.03 5.03 68.116 5.17 ;
      RECT 67.98 5.027 68.03 5.17 ;
      RECT 67.97 5.025 67.98 5.169 ;
      RECT 67.966 5.025 67.97 5.168 ;
      RECT 67.88 5.02 67.966 5.163 ;
      RECT 67.858 5.013 67.88 5.157 ;
      RECT 67.772 5.004 67.858 5.151 ;
      RECT 67.686 4.991 67.772 5.142 ;
      RECT 67.6 4.977 67.686 5.132 ;
      RECT 67.555 4.967 67.6 5.125 ;
      RECT 67.535 4.255 67.555 4.533 ;
      RECT 67.535 4.96 67.555 5.121 ;
      RECT 67.505 4.255 67.535 4.555 ;
      RECT 67.495 4.927 67.535 5.118 ;
      RECT 67.49 4.255 67.505 4.575 ;
      RECT 67.49 4.892 67.495 5.116 ;
      RECT 67.485 4.255 67.49 4.7 ;
      RECT 67.485 4.852 67.49 5.116 ;
      RECT 67.475 4.255 67.485 5.116 ;
      RECT 67.4 4.255 67.475 5.11 ;
      RECT 67.37 4.255 67.4 5.1 ;
      RECT 67.365 4.255 67.37 5.092 ;
      RECT 67.36 4.297 67.365 5.085 ;
      RECT 67.35 4.366 67.36 5.076 ;
      RECT 67.345 4.436 67.35 5.028 ;
      RECT 67.34 4.5 67.345 4.925 ;
      RECT 67.335 4.535 67.34 4.88 ;
      RECT 67.333 4.572 67.335 4.772 ;
      RECT 67.33 4.58 67.333 4.765 ;
      RECT 67.325 4.645 67.33 4.708 ;
      RECT 71.4 3.735 71.68 4.015 ;
      RECT 71.39 3.735 71.68 3.878 ;
      RECT 71.345 3.6 71.605 3.86 ;
      RECT 71.345 3.715 71.66 3.86 ;
      RECT 71.345 3.685 71.655 3.86 ;
      RECT 71.345 3.672 71.645 3.86 ;
      RECT 71.345 3.662 71.64 3.86 ;
      RECT 67.32 3.645 67.58 3.905 ;
      RECT 71.09 3.195 71.35 3.455 ;
      RECT 71.08 3.22 71.35 3.415 ;
      RECT 71.075 3.22 71.08 3.414 ;
      RECT 71.005 3.215 71.075 3.406 ;
      RECT 70.92 3.202 71.005 3.389 ;
      RECT 70.916 3.194 70.92 3.379 ;
      RECT 70.83 3.187 70.916 3.369 ;
      RECT 70.821 3.179 70.83 3.359 ;
      RECT 70.735 3.172 70.821 3.347 ;
      RECT 70.715 3.163 70.735 3.333 ;
      RECT 70.66 3.158 70.715 3.325 ;
      RECT 70.65 3.152 70.66 3.319 ;
      RECT 70.63 3.15 70.65 3.315 ;
      RECT 70.622 3.149 70.63 3.311 ;
      RECT 70.536 3.141 70.622 3.3 ;
      RECT 70.45 3.127 70.536 3.28 ;
      RECT 70.39 3.115 70.45 3.265 ;
      RECT 70.38 3.11 70.39 3.26 ;
      RECT 70.33 3.11 70.38 3.262 ;
      RECT 70.283 3.112 70.33 3.266 ;
      RECT 70.197 3.119 70.283 3.271 ;
      RECT 70.111 3.127 70.197 3.277 ;
      RECT 70.025 3.136 70.111 3.283 ;
      RECT 69.966 3.142 70.025 3.288 ;
      RECT 69.88 3.147 69.966 3.294 ;
      RECT 69.805 3.152 69.88 3.3 ;
      RECT 69.766 3.154 69.805 3.305 ;
      RECT 69.68 3.151 69.766 3.31 ;
      RECT 69.595 3.149 69.68 3.317 ;
      RECT 69.563 3.148 69.595 3.32 ;
      RECT 69.477 3.147 69.563 3.321 ;
      RECT 69.391 3.146 69.477 3.322 ;
      RECT 69.305 3.145 69.391 3.322 ;
      RECT 69.219 3.144 69.305 3.323 ;
      RECT 69.133 3.143 69.219 3.324 ;
      RECT 69.047 3.142 69.133 3.325 ;
      RECT 68.961 3.141 69.047 3.325 ;
      RECT 68.875 3.14 68.961 3.326 ;
      RECT 68.825 3.14 68.875 3.327 ;
      RECT 68.811 3.141 68.825 3.327 ;
      RECT 68.725 3.148 68.811 3.328 ;
      RECT 68.651 3.159 68.725 3.329 ;
      RECT 68.565 3.168 68.651 3.33 ;
      RECT 68.53 3.175 68.565 3.345 ;
      RECT 68.505 3.178 68.53 3.375 ;
      RECT 68.48 3.187 68.505 3.404 ;
      RECT 68.47 3.198 68.48 3.424 ;
      RECT 68.46 3.206 68.47 3.438 ;
      RECT 68.455 3.212 68.46 3.448 ;
      RECT 68.43 3.229 68.455 3.465 ;
      RECT 68.415 3.251 68.43 3.493 ;
      RECT 68.385 3.277 68.415 3.523 ;
      RECT 68.365 3.306 68.385 3.553 ;
      RECT 68.36 3.321 68.365 3.57 ;
      RECT 68.34 3.336 68.36 3.585 ;
      RECT 68.33 3.354 68.34 3.603 ;
      RECT 68.32 3.365 68.33 3.618 ;
      RECT 68.27 3.397 68.32 3.644 ;
      RECT 68.265 3.427 68.27 3.664 ;
      RECT 68.255 3.44 68.265 3.67 ;
      RECT 68.246 3.45 68.255 3.678 ;
      RECT 68.235 3.461 68.246 3.686 ;
      RECT 68.23 3.471 68.235 3.692 ;
      RECT 68.215 3.492 68.23 3.699 ;
      RECT 68.2 3.522 68.215 3.707 ;
      RECT 68.165 3.552 68.2 3.713 ;
      RECT 68.14 3.57 68.165 3.72 ;
      RECT 68.09 3.578 68.14 3.729 ;
      RECT 68.065 3.583 68.09 3.738 ;
      RECT 68.01 3.589 68.065 3.748 ;
      RECT 68.005 3.594 68.01 3.756 ;
      RECT 67.991 3.597 68.005 3.758 ;
      RECT 67.905 3.609 67.991 3.77 ;
      RECT 67.895 3.621 67.905 3.783 ;
      RECT 67.81 3.634 67.895 3.795 ;
      RECT 67.766 3.651 67.81 3.809 ;
      RECT 67.68 3.668 67.766 3.825 ;
      RECT 67.65 3.682 67.68 3.839 ;
      RECT 67.64 3.687 67.65 3.844 ;
      RECT 67.58 3.69 67.64 3.853 ;
      RECT 70.47 3.96 70.73 4.22 ;
      RECT 70.47 3.96 70.75 4.073 ;
      RECT 70.47 3.96 70.775 4.04 ;
      RECT 70.47 3.96 70.78 4.02 ;
      RECT 70.52 3.735 70.8 4.015 ;
      RECT 70.075 4.47 70.335 4.73 ;
      RECT 70.065 4.327 70.26 4.668 ;
      RECT 70.06 4.435 70.275 4.66 ;
      RECT 70.055 4.485 70.335 4.65 ;
      RECT 70.045 4.562 70.335 4.635 ;
      RECT 70.065 4.41 70.275 4.668 ;
      RECT 70.075 4.285 70.26 4.73 ;
      RECT 70.075 4.18 70.24 4.73 ;
      RECT 70.085 4.167 70.24 4.73 ;
      RECT 70.085 4.125 70.23 4.73 ;
      RECT 70.09 4.05 70.23 4.73 ;
      RECT 70.12 3.7 70.23 4.73 ;
      RECT 70.125 3.43 70.25 4.053 ;
      RECT 70.095 4.005 70.25 4.053 ;
      RECT 70.11 3.807 70.23 4.73 ;
      RECT 70.1 3.917 70.25 4.053 ;
      RECT 70.125 3.43 70.265 3.91 ;
      RECT 70.125 3.43 70.285 3.785 ;
      RECT 70.09 3.43 70.35 3.69 ;
      RECT 69.56 3.735 69.84 4.015 ;
      RECT 69.545 3.735 69.84 3.995 ;
      RECT 67.6 4.6 67.86 4.86 ;
      RECT 69.385 4.455 69.645 4.715 ;
      RECT 69.365 4.475 69.645 4.69 ;
      RECT 69.322 4.475 69.365 4.689 ;
      RECT 69.236 4.476 69.322 4.686 ;
      RECT 69.15 4.477 69.236 4.682 ;
      RECT 69.075 4.479 69.15 4.679 ;
      RECT 69.052 4.48 69.075 4.677 ;
      RECT 68.966 4.481 69.052 4.675 ;
      RECT 68.88 4.482 68.966 4.672 ;
      RECT 68.856 4.483 68.88 4.67 ;
      RECT 68.77 4.485 68.856 4.667 ;
      RECT 68.685 4.487 68.77 4.668 ;
      RECT 68.628 4.488 68.685 4.674 ;
      RECT 68.542 4.49 68.628 4.684 ;
      RECT 68.456 4.493 68.542 4.697 ;
      RECT 68.37 4.495 68.456 4.709 ;
      RECT 68.356 4.496 68.37 4.716 ;
      RECT 68.27 4.497 68.356 4.724 ;
      RECT 68.23 4.499 68.27 4.733 ;
      RECT 68.221 4.5 68.23 4.736 ;
      RECT 68.135 4.508 68.221 4.742 ;
      RECT 68.115 4.517 68.135 4.75 ;
      RECT 68.03 4.532 68.115 4.758 ;
      RECT 67.97 4.555 68.03 4.769 ;
      RECT 67.96 4.567 67.97 4.774 ;
      RECT 67.92 4.577 67.96 4.778 ;
      RECT 67.865 4.594 67.92 4.786 ;
      RECT 67.86 4.604 67.865 4.79 ;
      RECT 68.926 3.735 68.985 4.132 ;
      RECT 68.84 3.735 69.045 4.123 ;
      RECT 68.835 3.765 69.045 4.118 ;
      RECT 68.801 3.765 69.045 4.116 ;
      RECT 68.715 3.765 69.045 4.11 ;
      RECT 68.67 3.765 69.065 4.088 ;
      RECT 68.67 3.765 69.085 4.043 ;
      RECT 68.63 3.765 69.085 4.033 ;
      RECT 68.84 3.735 69.12 4.015 ;
      RECT 68.575 3.735 68.835 3.995 ;
      RECT 66.4 4.295 66.68 4.575 ;
      RECT 66.37 4.257 66.625 4.56 ;
      RECT 66.365 4.258 66.625 4.558 ;
      RECT 66.36 4.259 66.625 4.552 ;
      RECT 66.355 4.262 66.625 4.545 ;
      RECT 66.35 4.295 66.68 4.538 ;
      RECT 66.32 4.265 66.625 4.525 ;
      RECT 66.32 4.292 66.645 4.525 ;
      RECT 66.32 4.282 66.64 4.525 ;
      RECT 66.32 4.267 66.635 4.525 ;
      RECT 66.4 4.254 66.615 4.575 ;
      RECT 66.486 4.252 66.615 4.575 ;
      RECT 66.572 4.25 66.6 4.575 ;
      RECT 62.205 8.505 62.525 8.83 ;
      RECT 62.235 7.98 62.405 8.83 ;
      RECT 62.235 7.98 62.41 8.33 ;
      RECT 62.235 7.98 63.21 8.155 ;
      RECT 63.035 3.26 63.21 8.155 ;
      RECT 62.98 3.26 63.33 3.61 ;
      RECT 63.005 8.94 63.33 9.265 ;
      RECT 61.89 9.03 63.33 9.2 ;
      RECT 61.89 3.69 62.05 9.2 ;
      RECT 62.205 3.66 62.525 3.98 ;
      RECT 61.89 3.69 62.525 3.86 ;
      RECT 51.975 3.215 52.235 3.475 ;
      RECT 52.03 3.175 52.335 3.455 ;
      RECT 52.03 2.715 52.205 3.475 ;
      RECT 60.545 2.635 60.895 2.985 ;
      RECT 52.03 2.715 60.895 2.89 ;
      RECT 60.22 4.145 60.59 4.515 ;
      RECT 60.305 3.53 60.475 4.515 ;
      RECT 56.325 3.75 56.56 4.01 ;
      RECT 59.47 3.53 59.635 3.79 ;
      RECT 59.375 3.52 59.39 3.79 ;
      RECT 59.47 3.53 60.475 3.71 ;
      RECT 57.975 3.09 58.015 3.23 ;
      RECT 59.39 3.525 59.47 3.79 ;
      RECT 59.335 3.52 59.375 3.756 ;
      RECT 59.321 3.52 59.335 3.756 ;
      RECT 59.235 3.525 59.321 3.758 ;
      RECT 59.19 3.532 59.235 3.76 ;
      RECT 59.16 3.532 59.19 3.762 ;
      RECT 59.135 3.527 59.16 3.764 ;
      RECT 59.105 3.523 59.135 3.773 ;
      RECT 59.095 3.52 59.105 3.785 ;
      RECT 59.09 3.52 59.095 3.793 ;
      RECT 59.085 3.52 59.09 3.798 ;
      RECT 59.075 3.519 59.085 3.808 ;
      RECT 59.07 3.518 59.075 3.818 ;
      RECT 59.055 3.517 59.07 3.823 ;
      RECT 59.027 3.514 59.055 3.85 ;
      RECT 58.941 3.506 59.027 3.85 ;
      RECT 58.855 3.495 58.941 3.85 ;
      RECT 58.815 3.48 58.855 3.85 ;
      RECT 58.775 3.454 58.815 3.85 ;
      RECT 58.77 3.436 58.775 3.662 ;
      RECT 58.76 3.432 58.77 3.652 ;
      RECT 58.745 3.422 58.76 3.639 ;
      RECT 58.725 3.406 58.745 3.624 ;
      RECT 58.71 3.391 58.725 3.609 ;
      RECT 58.7 3.38 58.71 3.599 ;
      RECT 58.675 3.364 58.7 3.588 ;
      RECT 58.67 3.351 58.675 3.578 ;
      RECT 58.665 3.347 58.67 3.573 ;
      RECT 58.61 3.333 58.665 3.551 ;
      RECT 58.571 3.314 58.61 3.515 ;
      RECT 58.485 3.288 58.571 3.468 ;
      RECT 58.481 3.27 58.485 3.434 ;
      RECT 58.395 3.251 58.481 3.412 ;
      RECT 58.39 3.233 58.395 3.39 ;
      RECT 58.385 3.231 58.39 3.388 ;
      RECT 58.375 3.23 58.385 3.383 ;
      RECT 58.315 3.217 58.375 3.369 ;
      RECT 58.27 3.195 58.315 3.348 ;
      RECT 58.21 3.172 58.27 3.327 ;
      RECT 58.146 3.147 58.21 3.302 ;
      RECT 58.06 3.117 58.146 3.271 ;
      RECT 58.045 3.097 58.06 3.25 ;
      RECT 58.015 3.092 58.045 3.241 ;
      RECT 57.962 3.09 57.975 3.23 ;
      RECT 57.876 3.09 57.962 3.232 ;
      RECT 57.79 3.09 57.876 3.234 ;
      RECT 57.77 3.09 57.79 3.238 ;
      RECT 57.725 3.092 57.77 3.249 ;
      RECT 57.685 3.102 57.725 3.265 ;
      RECT 57.681 3.111 57.685 3.273 ;
      RECT 57.595 3.131 57.681 3.289 ;
      RECT 57.585 3.15 57.595 3.307 ;
      RECT 57.58 3.152 57.585 3.31 ;
      RECT 57.57 3.156 57.58 3.313 ;
      RECT 57.55 3.161 57.57 3.323 ;
      RECT 57.52 3.171 57.55 3.343 ;
      RECT 57.515 3.178 57.52 3.357 ;
      RECT 57.505 3.182 57.515 3.364 ;
      RECT 57.49 3.19 57.505 3.375 ;
      RECT 57.48 3.2 57.49 3.386 ;
      RECT 57.47 3.207 57.48 3.394 ;
      RECT 57.445 3.22 57.47 3.409 ;
      RECT 57.381 3.256 57.445 3.448 ;
      RECT 57.295 3.319 57.381 3.512 ;
      RECT 57.26 3.37 57.295 3.565 ;
      RECT 57.255 3.387 57.26 3.582 ;
      RECT 57.24 3.396 57.255 3.589 ;
      RECT 57.22 3.411 57.24 3.603 ;
      RECT 57.215 3.422 57.22 3.613 ;
      RECT 57.195 3.435 57.215 3.623 ;
      RECT 57.19 3.445 57.195 3.633 ;
      RECT 57.175 3.45 57.19 3.642 ;
      RECT 57.165 3.46 57.175 3.653 ;
      RECT 57.135 3.477 57.165 3.67 ;
      RECT 57.125 3.495 57.135 3.688 ;
      RECT 57.11 3.506 57.125 3.699 ;
      RECT 57.07 3.53 57.11 3.715 ;
      RECT 57.035 3.564 57.07 3.732 ;
      RECT 57.005 3.587 57.035 3.744 ;
      RECT 56.99 3.597 57.005 3.753 ;
      RECT 56.95 3.607 56.99 3.764 ;
      RECT 56.93 3.618 56.95 3.776 ;
      RECT 56.925 3.622 56.93 3.783 ;
      RECT 56.91 3.626 56.925 3.788 ;
      RECT 56.9 3.631 56.91 3.793 ;
      RECT 56.895 3.634 56.9 3.796 ;
      RECT 56.865 3.64 56.895 3.803 ;
      RECT 56.83 3.65 56.865 3.817 ;
      RECT 56.77 3.665 56.83 3.837 ;
      RECT 56.715 3.685 56.77 3.861 ;
      RECT 56.686 3.7 56.715 3.879 ;
      RECT 56.6 3.72 56.686 3.904 ;
      RECT 56.595 3.735 56.6 3.924 ;
      RECT 56.585 3.738 56.595 3.925 ;
      RECT 56.56 3.745 56.585 4.01 ;
      RECT 59.255 4.238 59.535 4.575 ;
      RECT 59.255 4.248 59.54 4.533 ;
      RECT 59.255 4.257 59.545 4.43 ;
      RECT 59.255 4.272 59.55 4.298 ;
      RECT 59.255 4.1 59.515 4.575 ;
      RECT 49.555 8.94 49.905 9.29 ;
      RECT 58.38 8.895 58.73 9.245 ;
      RECT 49.555 8.97 58.73 9.17 ;
      RECT 56.975 4.98 56.985 5.17 ;
      RECT 55.235 4.855 55.515 5.135 ;
      RECT 58.28 3.795 58.285 4.28 ;
      RECT 58.175 3.795 58.235 4.055 ;
      RECT 58.5 4.765 58.505 4.84 ;
      RECT 58.49 4.632 58.5 4.875 ;
      RECT 58.48 4.467 58.49 4.896 ;
      RECT 58.475 4.337 58.48 4.912 ;
      RECT 58.465 4.227 58.475 4.928 ;
      RECT 58.46 4.126 58.465 4.945 ;
      RECT 58.455 4.108 58.46 4.955 ;
      RECT 58.45 4.09 58.455 4.965 ;
      RECT 58.44 4.065 58.45 4.98 ;
      RECT 58.435 4.045 58.44 4.995 ;
      RECT 58.415 3.795 58.435 5.02 ;
      RECT 58.4 3.795 58.415 5.053 ;
      RECT 58.37 3.795 58.4 5.075 ;
      RECT 58.35 3.795 58.37 5.089 ;
      RECT 58.33 3.795 58.35 4.605 ;
      RECT 58.345 4.672 58.35 5.094 ;
      RECT 58.34 4.702 58.345 5.096 ;
      RECT 58.335 4.715 58.34 5.099 ;
      RECT 58.33 4.725 58.335 5.103 ;
      RECT 58.325 3.795 58.33 4.523 ;
      RECT 58.325 4.735 58.33 5.105 ;
      RECT 58.32 3.795 58.325 4.5 ;
      RECT 58.31 4.757 58.325 5.105 ;
      RECT 58.305 3.795 58.32 4.445 ;
      RECT 58.3 4.782 58.31 5.105 ;
      RECT 58.3 3.795 58.305 4.39 ;
      RECT 58.29 3.795 58.3 4.338 ;
      RECT 58.295 4.795 58.3 5.106 ;
      RECT 58.29 4.807 58.295 5.107 ;
      RECT 58.285 3.795 58.29 4.298 ;
      RECT 58.285 4.82 58.29 5.108 ;
      RECT 58.27 4.835 58.285 5.109 ;
      RECT 58.275 3.795 58.28 4.26 ;
      RECT 58.27 3.795 58.275 4.225 ;
      RECT 58.265 3.795 58.27 4.2 ;
      RECT 58.26 4.862 58.27 5.111 ;
      RECT 58.255 3.795 58.265 4.158 ;
      RECT 58.255 4.88 58.26 5.112 ;
      RECT 58.25 3.795 58.255 4.118 ;
      RECT 58.25 4.887 58.255 5.113 ;
      RECT 58.245 3.795 58.25 4.09 ;
      RECT 58.24 4.905 58.25 5.114 ;
      RECT 58.235 3.795 58.245 4.07 ;
      RECT 58.23 4.925 58.24 5.116 ;
      RECT 58.22 4.942 58.23 5.117 ;
      RECT 58.185 4.965 58.22 5.12 ;
      RECT 58.13 4.983 58.185 5.126 ;
      RECT 58.044 4.991 58.13 5.135 ;
      RECT 57.958 5.002 58.044 5.146 ;
      RECT 57.872 5.012 57.958 5.157 ;
      RECT 57.786 5.022 57.872 5.169 ;
      RECT 57.7 5.032 57.786 5.18 ;
      RECT 57.68 5.038 57.7 5.186 ;
      RECT 57.6 5.04 57.68 5.19 ;
      RECT 57.595 5.039 57.6 5.195 ;
      RECT 57.587 5.038 57.595 5.195 ;
      RECT 57.501 5.034 57.587 5.193 ;
      RECT 57.415 5.026 57.501 5.19 ;
      RECT 57.329 5.017 57.415 5.186 ;
      RECT 57.243 5.009 57.329 5.183 ;
      RECT 57.157 5.001 57.243 5.179 ;
      RECT 57.071 4.992 57.157 5.176 ;
      RECT 56.985 4.984 57.071 5.172 ;
      RECT 56.93 4.977 56.975 5.17 ;
      RECT 56.845 4.97 56.93 5.168 ;
      RECT 56.771 4.962 56.845 5.164 ;
      RECT 56.685 4.954 56.771 5.161 ;
      RECT 56.682 4.95 56.685 5.159 ;
      RECT 56.596 4.946 56.682 5.158 ;
      RECT 56.51 4.938 56.596 5.155 ;
      RECT 56.425 4.933 56.51 5.152 ;
      RECT 56.339 4.93 56.425 5.149 ;
      RECT 56.253 4.928 56.339 5.146 ;
      RECT 56.167 4.925 56.253 5.143 ;
      RECT 56.081 4.922 56.167 5.14 ;
      RECT 55.995 4.919 56.081 5.137 ;
      RECT 55.919 4.917 55.995 5.134 ;
      RECT 55.833 4.914 55.919 5.131 ;
      RECT 55.747 4.911 55.833 5.129 ;
      RECT 55.661 4.909 55.747 5.126 ;
      RECT 55.575 4.906 55.661 5.123 ;
      RECT 55.515 4.897 55.575 5.121 ;
      RECT 58.025 4.515 58.1 4.775 ;
      RECT 58.005 4.495 58.01 4.775 ;
      RECT 57.325 4.28 57.43 4.575 ;
      RECT 51.77 4.255 51.84 4.515 ;
      RECT 57.665 4.13 57.67 4.501 ;
      RECT 57.655 4.185 57.66 4.501 ;
      RECT 57.96 3.355 58.02 3.615 ;
      RECT 58.015 4.51 58.025 4.775 ;
      RECT 58.01 4.5 58.015 4.775 ;
      RECT 57.93 4.447 58.005 4.775 ;
      RECT 57.955 3.355 57.96 3.635 ;
      RECT 57.945 3.355 57.955 3.655 ;
      RECT 57.93 3.355 57.945 3.685 ;
      RECT 57.915 3.355 57.93 3.728 ;
      RECT 57.91 4.39 57.93 4.775 ;
      RECT 57.9 3.355 57.915 3.765 ;
      RECT 57.895 4.37 57.91 4.775 ;
      RECT 57.895 3.355 57.9 3.788 ;
      RECT 57.885 3.355 57.895 3.813 ;
      RECT 57.855 4.337 57.895 4.775 ;
      RECT 57.86 3.355 57.885 3.863 ;
      RECT 57.855 3.355 57.86 3.918 ;
      RECT 57.85 3.355 57.855 3.96 ;
      RECT 57.84 4.3 57.855 4.775 ;
      RECT 57.845 3.355 57.85 4.003 ;
      RECT 57.84 3.355 57.845 4.068 ;
      RECT 57.835 3.355 57.84 4.09 ;
      RECT 57.835 4.288 57.84 4.64 ;
      RECT 57.83 3.355 57.835 4.158 ;
      RECT 57.83 4.28 57.835 4.623 ;
      RECT 57.825 3.355 57.83 4.203 ;
      RECT 57.82 4.262 57.83 4.6 ;
      RECT 57.82 3.355 57.825 4.24 ;
      RECT 57.81 3.355 57.82 4.58 ;
      RECT 57.805 3.355 57.81 4.563 ;
      RECT 57.8 3.355 57.805 4.548 ;
      RECT 57.795 3.355 57.8 4.533 ;
      RECT 57.775 3.355 57.795 4.523 ;
      RECT 57.77 3.355 57.775 4.513 ;
      RECT 57.76 3.355 57.77 4.509 ;
      RECT 57.755 3.632 57.76 4.508 ;
      RECT 57.75 3.655 57.755 4.507 ;
      RECT 57.745 3.685 57.75 4.506 ;
      RECT 57.74 3.712 57.745 4.505 ;
      RECT 57.735 3.74 57.74 4.505 ;
      RECT 57.73 3.767 57.735 4.505 ;
      RECT 57.725 3.787 57.73 4.505 ;
      RECT 57.72 3.815 57.725 4.505 ;
      RECT 57.71 3.857 57.72 4.505 ;
      RECT 57.7 3.902 57.71 4.504 ;
      RECT 57.695 3.955 57.7 4.503 ;
      RECT 57.69 3.987 57.695 4.502 ;
      RECT 57.685 4.007 57.69 4.501 ;
      RECT 57.68 4.045 57.685 4.501 ;
      RECT 57.675 4.067 57.68 4.501 ;
      RECT 57.67 4.092 57.675 4.501 ;
      RECT 57.66 4.157 57.665 4.501 ;
      RECT 57.645 4.217 57.655 4.501 ;
      RECT 57.63 4.227 57.645 4.501 ;
      RECT 57.61 4.237 57.63 4.501 ;
      RECT 57.58 4.242 57.61 4.498 ;
      RECT 57.52 4.252 57.58 4.495 ;
      RECT 57.5 4.261 57.52 4.5 ;
      RECT 57.475 4.267 57.5 4.513 ;
      RECT 57.455 4.272 57.475 4.528 ;
      RECT 57.43 4.277 57.455 4.575 ;
      RECT 57.301 4.279 57.325 4.575 ;
      RECT 57.215 4.274 57.301 4.575 ;
      RECT 57.175 4.271 57.215 4.575 ;
      RECT 57.125 4.273 57.175 4.555 ;
      RECT 57.095 4.277 57.125 4.555 ;
      RECT 57.016 4.287 57.095 4.555 ;
      RECT 56.93 4.302 57.016 4.556 ;
      RECT 56.88 4.312 56.93 4.557 ;
      RECT 56.872 4.315 56.88 4.557 ;
      RECT 56.786 4.317 56.872 4.558 ;
      RECT 56.7 4.321 56.786 4.558 ;
      RECT 56.614 4.325 56.7 4.559 ;
      RECT 56.528 4.328 56.614 4.56 ;
      RECT 56.442 4.332 56.528 4.56 ;
      RECT 56.356 4.336 56.442 4.561 ;
      RECT 56.27 4.339 56.356 4.562 ;
      RECT 56.184 4.343 56.27 4.562 ;
      RECT 56.098 4.347 56.184 4.563 ;
      RECT 56.012 4.351 56.098 4.564 ;
      RECT 55.926 4.354 56.012 4.564 ;
      RECT 55.84 4.358 55.926 4.565 ;
      RECT 55.81 4.36 55.84 4.565 ;
      RECT 55.724 4.363 55.81 4.566 ;
      RECT 55.638 4.367 55.724 4.567 ;
      RECT 55.552 4.371 55.638 4.568 ;
      RECT 55.466 4.374 55.552 4.568 ;
      RECT 55.38 4.378 55.466 4.569 ;
      RECT 55.345 4.383 55.38 4.57 ;
      RECT 55.29 4.393 55.345 4.577 ;
      RECT 55.265 4.405 55.29 4.587 ;
      RECT 55.23 4.418 55.265 4.595 ;
      RECT 55.19 4.435 55.23 4.618 ;
      RECT 55.17 4.448 55.19 4.645 ;
      RECT 55.14 4.46 55.17 4.673 ;
      RECT 55.135 4.468 55.14 4.693 ;
      RECT 55.13 4.471 55.135 4.703 ;
      RECT 55.08 4.483 55.13 4.737 ;
      RECT 55.07 4.498 55.08 4.77 ;
      RECT 55.06 4.504 55.07 4.783 ;
      RECT 55.05 4.511 55.06 4.795 ;
      RECT 55.025 4.524 55.05 4.813 ;
      RECT 55.01 4.539 55.025 4.835 ;
      RECT 55 4.547 55.01 4.851 ;
      RECT 54.985 4.556 55 4.866 ;
      RECT 54.975 4.566 54.985 4.88 ;
      RECT 54.956 4.579 54.975 4.897 ;
      RECT 54.87 4.624 54.956 4.962 ;
      RECT 54.855 4.669 54.87 5.02 ;
      RECT 54.85 4.678 54.855 5.033 ;
      RECT 54.84 4.685 54.85 5.038 ;
      RECT 54.835 4.69 54.84 5.042 ;
      RECT 54.815 4.7 54.835 5.049 ;
      RECT 54.79 4.72 54.815 5.063 ;
      RECT 54.755 4.745 54.79 5.083 ;
      RECT 54.74 4.768 54.755 5.098 ;
      RECT 54.73 4.778 54.74 5.103 ;
      RECT 54.72 4.786 54.73 5.11 ;
      RECT 54.71 4.795 54.72 5.116 ;
      RECT 54.69 4.807 54.71 5.118 ;
      RECT 54.68 4.82 54.69 5.12 ;
      RECT 54.655 4.835 54.68 5.123 ;
      RECT 54.635 4.852 54.655 5.127 ;
      RECT 54.595 4.88 54.635 5.133 ;
      RECT 54.53 4.927 54.595 5.142 ;
      RECT 54.515 4.96 54.53 5.15 ;
      RECT 54.51 4.967 54.515 5.152 ;
      RECT 54.46 4.992 54.51 5.157 ;
      RECT 54.445 5.016 54.46 5.164 ;
      RECT 54.395 5.021 54.445 5.165 ;
      RECT 54.309 5.025 54.395 5.165 ;
      RECT 54.223 5.025 54.309 5.165 ;
      RECT 54.137 5.025 54.223 5.166 ;
      RECT 54.051 5.025 54.137 5.166 ;
      RECT 53.965 5.025 54.051 5.166 ;
      RECT 53.899 5.025 53.965 5.166 ;
      RECT 53.813 5.025 53.899 5.167 ;
      RECT 53.727 5.025 53.813 5.167 ;
      RECT 53.641 5.026 53.727 5.168 ;
      RECT 53.555 5.026 53.641 5.168 ;
      RECT 53.469 5.026 53.555 5.168 ;
      RECT 53.383 5.026 53.469 5.169 ;
      RECT 53.297 5.026 53.383 5.169 ;
      RECT 53.211 5.027 53.297 5.17 ;
      RECT 53.125 5.027 53.211 5.17 ;
      RECT 53.105 5.027 53.125 5.17 ;
      RECT 53.019 5.027 53.105 5.17 ;
      RECT 52.933 5.027 53.019 5.17 ;
      RECT 52.847 5.028 52.933 5.17 ;
      RECT 52.761 5.028 52.847 5.17 ;
      RECT 52.675 5.028 52.761 5.17 ;
      RECT 52.589 5.029 52.675 5.17 ;
      RECT 52.503 5.029 52.589 5.17 ;
      RECT 52.417 5.029 52.503 5.17 ;
      RECT 52.331 5.029 52.417 5.17 ;
      RECT 52.245 5.03 52.331 5.17 ;
      RECT 52.195 5.027 52.245 5.17 ;
      RECT 52.185 5.025 52.195 5.169 ;
      RECT 52.181 5.025 52.185 5.168 ;
      RECT 52.095 5.02 52.181 5.163 ;
      RECT 52.073 5.013 52.095 5.157 ;
      RECT 51.987 5.004 52.073 5.151 ;
      RECT 51.901 4.991 51.987 5.142 ;
      RECT 51.815 4.977 51.901 5.132 ;
      RECT 51.77 4.967 51.815 5.125 ;
      RECT 51.75 4.255 51.77 4.533 ;
      RECT 51.75 4.96 51.77 5.121 ;
      RECT 51.72 4.255 51.75 4.555 ;
      RECT 51.71 4.927 51.75 5.118 ;
      RECT 51.705 4.255 51.72 4.575 ;
      RECT 51.705 4.892 51.71 5.116 ;
      RECT 51.7 4.255 51.705 4.7 ;
      RECT 51.7 4.852 51.705 5.116 ;
      RECT 51.69 4.255 51.7 5.116 ;
      RECT 51.615 4.255 51.69 5.11 ;
      RECT 51.585 4.255 51.615 5.1 ;
      RECT 51.58 4.255 51.585 5.092 ;
      RECT 51.575 4.297 51.58 5.085 ;
      RECT 51.565 4.366 51.575 5.076 ;
      RECT 51.56 4.436 51.565 5.028 ;
      RECT 51.555 4.5 51.56 4.925 ;
      RECT 51.55 4.535 51.555 4.88 ;
      RECT 51.548 4.572 51.55 4.772 ;
      RECT 51.545 4.58 51.548 4.765 ;
      RECT 51.54 4.645 51.545 4.708 ;
      RECT 55.615 3.735 55.895 4.015 ;
      RECT 55.605 3.735 55.895 3.878 ;
      RECT 55.56 3.6 55.82 3.86 ;
      RECT 55.56 3.715 55.875 3.86 ;
      RECT 55.56 3.685 55.87 3.86 ;
      RECT 55.56 3.672 55.86 3.86 ;
      RECT 55.56 3.662 55.855 3.86 ;
      RECT 51.535 3.645 51.795 3.905 ;
      RECT 55.305 3.195 55.565 3.455 ;
      RECT 55.295 3.22 55.565 3.415 ;
      RECT 55.29 3.22 55.295 3.414 ;
      RECT 55.22 3.215 55.29 3.406 ;
      RECT 55.135 3.202 55.22 3.389 ;
      RECT 55.131 3.194 55.135 3.379 ;
      RECT 55.045 3.187 55.131 3.369 ;
      RECT 55.036 3.179 55.045 3.359 ;
      RECT 54.95 3.172 55.036 3.347 ;
      RECT 54.93 3.163 54.95 3.333 ;
      RECT 54.875 3.158 54.93 3.325 ;
      RECT 54.865 3.152 54.875 3.319 ;
      RECT 54.845 3.15 54.865 3.315 ;
      RECT 54.837 3.149 54.845 3.311 ;
      RECT 54.751 3.141 54.837 3.3 ;
      RECT 54.665 3.127 54.751 3.28 ;
      RECT 54.605 3.115 54.665 3.265 ;
      RECT 54.595 3.11 54.605 3.26 ;
      RECT 54.545 3.11 54.595 3.262 ;
      RECT 54.498 3.112 54.545 3.266 ;
      RECT 54.412 3.119 54.498 3.271 ;
      RECT 54.326 3.127 54.412 3.277 ;
      RECT 54.24 3.136 54.326 3.283 ;
      RECT 54.181 3.142 54.24 3.288 ;
      RECT 54.095 3.147 54.181 3.294 ;
      RECT 54.02 3.152 54.095 3.3 ;
      RECT 53.981 3.154 54.02 3.305 ;
      RECT 53.895 3.151 53.981 3.31 ;
      RECT 53.81 3.149 53.895 3.317 ;
      RECT 53.778 3.148 53.81 3.32 ;
      RECT 53.692 3.147 53.778 3.321 ;
      RECT 53.606 3.146 53.692 3.322 ;
      RECT 53.52 3.145 53.606 3.322 ;
      RECT 53.434 3.144 53.52 3.323 ;
      RECT 53.348 3.143 53.434 3.324 ;
      RECT 53.262 3.142 53.348 3.325 ;
      RECT 53.176 3.141 53.262 3.325 ;
      RECT 53.09 3.14 53.176 3.326 ;
      RECT 53.04 3.14 53.09 3.327 ;
      RECT 53.026 3.141 53.04 3.327 ;
      RECT 52.94 3.148 53.026 3.328 ;
      RECT 52.866 3.159 52.94 3.329 ;
      RECT 52.78 3.168 52.866 3.33 ;
      RECT 52.745 3.175 52.78 3.345 ;
      RECT 52.72 3.178 52.745 3.375 ;
      RECT 52.695 3.187 52.72 3.404 ;
      RECT 52.685 3.198 52.695 3.424 ;
      RECT 52.675 3.206 52.685 3.438 ;
      RECT 52.67 3.212 52.675 3.448 ;
      RECT 52.645 3.229 52.67 3.465 ;
      RECT 52.63 3.251 52.645 3.493 ;
      RECT 52.6 3.277 52.63 3.523 ;
      RECT 52.58 3.306 52.6 3.553 ;
      RECT 52.575 3.321 52.58 3.57 ;
      RECT 52.555 3.336 52.575 3.585 ;
      RECT 52.545 3.354 52.555 3.603 ;
      RECT 52.535 3.365 52.545 3.618 ;
      RECT 52.485 3.397 52.535 3.644 ;
      RECT 52.48 3.427 52.485 3.664 ;
      RECT 52.47 3.44 52.48 3.67 ;
      RECT 52.461 3.45 52.47 3.678 ;
      RECT 52.45 3.461 52.461 3.686 ;
      RECT 52.445 3.471 52.45 3.692 ;
      RECT 52.43 3.492 52.445 3.699 ;
      RECT 52.415 3.522 52.43 3.707 ;
      RECT 52.38 3.552 52.415 3.713 ;
      RECT 52.355 3.57 52.38 3.72 ;
      RECT 52.305 3.578 52.355 3.729 ;
      RECT 52.28 3.583 52.305 3.738 ;
      RECT 52.225 3.589 52.28 3.748 ;
      RECT 52.22 3.594 52.225 3.756 ;
      RECT 52.206 3.597 52.22 3.758 ;
      RECT 52.12 3.609 52.206 3.77 ;
      RECT 52.11 3.621 52.12 3.783 ;
      RECT 52.025 3.634 52.11 3.795 ;
      RECT 51.981 3.651 52.025 3.809 ;
      RECT 51.895 3.668 51.981 3.825 ;
      RECT 51.865 3.682 51.895 3.839 ;
      RECT 51.855 3.687 51.865 3.844 ;
      RECT 51.795 3.69 51.855 3.853 ;
      RECT 54.685 3.96 54.945 4.22 ;
      RECT 54.685 3.96 54.965 4.073 ;
      RECT 54.685 3.96 54.99 4.04 ;
      RECT 54.685 3.96 54.995 4.02 ;
      RECT 54.735 3.735 55.015 4.015 ;
      RECT 54.29 4.47 54.55 4.73 ;
      RECT 54.28 4.327 54.475 4.668 ;
      RECT 54.275 4.435 54.49 4.66 ;
      RECT 54.27 4.485 54.55 4.65 ;
      RECT 54.26 4.562 54.55 4.635 ;
      RECT 54.28 4.41 54.49 4.668 ;
      RECT 54.29 4.285 54.475 4.73 ;
      RECT 54.29 4.18 54.455 4.73 ;
      RECT 54.3 4.167 54.455 4.73 ;
      RECT 54.3 4.125 54.445 4.73 ;
      RECT 54.305 4.05 54.445 4.73 ;
      RECT 54.335 3.7 54.445 4.73 ;
      RECT 54.34 3.43 54.465 4.053 ;
      RECT 54.31 4.005 54.465 4.053 ;
      RECT 54.325 3.807 54.445 4.73 ;
      RECT 54.315 3.917 54.465 4.053 ;
      RECT 54.34 3.43 54.48 3.91 ;
      RECT 54.34 3.43 54.5 3.785 ;
      RECT 54.305 3.43 54.565 3.69 ;
      RECT 53.775 3.735 54.055 4.015 ;
      RECT 53.76 3.735 54.055 3.995 ;
      RECT 51.815 4.6 52.075 4.86 ;
      RECT 53.6 4.455 53.86 4.715 ;
      RECT 53.58 4.475 53.86 4.69 ;
      RECT 53.537 4.475 53.58 4.689 ;
      RECT 53.451 4.476 53.537 4.686 ;
      RECT 53.365 4.477 53.451 4.682 ;
      RECT 53.29 4.479 53.365 4.679 ;
      RECT 53.267 4.48 53.29 4.677 ;
      RECT 53.181 4.481 53.267 4.675 ;
      RECT 53.095 4.482 53.181 4.672 ;
      RECT 53.071 4.483 53.095 4.67 ;
      RECT 52.985 4.485 53.071 4.667 ;
      RECT 52.9 4.487 52.985 4.668 ;
      RECT 52.843 4.488 52.9 4.674 ;
      RECT 52.757 4.49 52.843 4.684 ;
      RECT 52.671 4.493 52.757 4.697 ;
      RECT 52.585 4.495 52.671 4.709 ;
      RECT 52.571 4.496 52.585 4.716 ;
      RECT 52.485 4.497 52.571 4.724 ;
      RECT 52.445 4.499 52.485 4.733 ;
      RECT 52.436 4.5 52.445 4.736 ;
      RECT 52.35 4.508 52.436 4.742 ;
      RECT 52.33 4.517 52.35 4.75 ;
      RECT 52.245 4.532 52.33 4.758 ;
      RECT 52.185 4.555 52.245 4.769 ;
      RECT 52.175 4.567 52.185 4.774 ;
      RECT 52.135 4.577 52.175 4.778 ;
      RECT 52.08 4.594 52.135 4.786 ;
      RECT 52.075 4.604 52.08 4.79 ;
      RECT 53.141 3.735 53.2 4.132 ;
      RECT 53.055 3.735 53.26 4.123 ;
      RECT 53.05 3.765 53.26 4.118 ;
      RECT 53.016 3.765 53.26 4.116 ;
      RECT 52.93 3.765 53.26 4.11 ;
      RECT 52.885 3.765 53.28 4.088 ;
      RECT 52.885 3.765 53.3 4.043 ;
      RECT 52.845 3.765 53.3 4.033 ;
      RECT 53.055 3.735 53.335 4.015 ;
      RECT 52.79 3.735 53.05 3.995 ;
      RECT 50.615 4.295 50.895 4.575 ;
      RECT 50.585 4.257 50.84 4.56 ;
      RECT 50.58 4.258 50.84 4.558 ;
      RECT 50.575 4.259 50.84 4.552 ;
      RECT 50.57 4.262 50.84 4.545 ;
      RECT 50.565 4.295 50.895 4.538 ;
      RECT 50.535 4.265 50.84 4.525 ;
      RECT 50.535 4.292 50.86 4.525 ;
      RECT 50.535 4.282 50.855 4.525 ;
      RECT 50.535 4.267 50.85 4.525 ;
      RECT 50.615 4.254 50.83 4.575 ;
      RECT 50.701 4.252 50.83 4.575 ;
      RECT 50.787 4.25 50.815 4.575 ;
      RECT 46.42 8.505 46.74 8.83 ;
      RECT 46.45 7.98 46.62 8.83 ;
      RECT 46.45 7.98 46.625 8.33 ;
      RECT 46.45 7.98 47.425 8.155 ;
      RECT 47.25 3.26 47.425 8.155 ;
      RECT 47.195 3.26 47.545 3.61 ;
      RECT 47.22 8.94 47.545 9.265 ;
      RECT 46.105 9.03 47.545 9.2 ;
      RECT 46.105 3.69 46.265 9.2 ;
      RECT 46.42 3.66 46.74 3.98 ;
      RECT 46.105 3.69 46.74 3.86 ;
      RECT 36.19 3.215 36.45 3.475 ;
      RECT 36.245 3.175 36.55 3.455 ;
      RECT 36.245 2.715 36.42 3.475 ;
      RECT 44.76 2.635 45.11 2.985 ;
      RECT 36.245 2.715 45.11 2.89 ;
      RECT 44.435 4.145 44.805 4.515 ;
      RECT 44.52 3.53 44.69 4.515 ;
      RECT 40.54 3.75 40.775 4.01 ;
      RECT 43.685 3.53 43.85 3.79 ;
      RECT 43.59 3.52 43.605 3.79 ;
      RECT 43.685 3.53 44.69 3.71 ;
      RECT 42.19 3.09 42.23 3.23 ;
      RECT 43.605 3.525 43.685 3.79 ;
      RECT 43.55 3.52 43.59 3.756 ;
      RECT 43.536 3.52 43.55 3.756 ;
      RECT 43.45 3.525 43.536 3.758 ;
      RECT 43.405 3.532 43.45 3.76 ;
      RECT 43.375 3.532 43.405 3.762 ;
      RECT 43.35 3.527 43.375 3.764 ;
      RECT 43.32 3.523 43.35 3.773 ;
      RECT 43.31 3.52 43.32 3.785 ;
      RECT 43.305 3.52 43.31 3.793 ;
      RECT 43.3 3.52 43.305 3.798 ;
      RECT 43.29 3.519 43.3 3.808 ;
      RECT 43.285 3.518 43.29 3.818 ;
      RECT 43.27 3.517 43.285 3.823 ;
      RECT 43.242 3.514 43.27 3.85 ;
      RECT 43.156 3.506 43.242 3.85 ;
      RECT 43.07 3.495 43.156 3.85 ;
      RECT 43.03 3.48 43.07 3.85 ;
      RECT 42.99 3.454 43.03 3.85 ;
      RECT 42.985 3.436 42.99 3.662 ;
      RECT 42.975 3.432 42.985 3.652 ;
      RECT 42.96 3.422 42.975 3.639 ;
      RECT 42.94 3.406 42.96 3.624 ;
      RECT 42.925 3.391 42.94 3.609 ;
      RECT 42.915 3.38 42.925 3.599 ;
      RECT 42.89 3.364 42.915 3.588 ;
      RECT 42.885 3.351 42.89 3.578 ;
      RECT 42.88 3.347 42.885 3.573 ;
      RECT 42.825 3.333 42.88 3.551 ;
      RECT 42.786 3.314 42.825 3.515 ;
      RECT 42.7 3.288 42.786 3.468 ;
      RECT 42.696 3.27 42.7 3.434 ;
      RECT 42.61 3.251 42.696 3.412 ;
      RECT 42.605 3.233 42.61 3.39 ;
      RECT 42.6 3.231 42.605 3.388 ;
      RECT 42.59 3.23 42.6 3.383 ;
      RECT 42.53 3.217 42.59 3.369 ;
      RECT 42.485 3.195 42.53 3.348 ;
      RECT 42.425 3.172 42.485 3.327 ;
      RECT 42.361 3.147 42.425 3.302 ;
      RECT 42.275 3.117 42.361 3.271 ;
      RECT 42.26 3.097 42.275 3.25 ;
      RECT 42.23 3.092 42.26 3.241 ;
      RECT 42.177 3.09 42.19 3.23 ;
      RECT 42.091 3.09 42.177 3.232 ;
      RECT 42.005 3.09 42.091 3.234 ;
      RECT 41.985 3.09 42.005 3.238 ;
      RECT 41.94 3.092 41.985 3.249 ;
      RECT 41.9 3.102 41.94 3.265 ;
      RECT 41.896 3.111 41.9 3.273 ;
      RECT 41.81 3.131 41.896 3.289 ;
      RECT 41.8 3.15 41.81 3.307 ;
      RECT 41.795 3.152 41.8 3.31 ;
      RECT 41.785 3.156 41.795 3.313 ;
      RECT 41.765 3.161 41.785 3.323 ;
      RECT 41.735 3.171 41.765 3.343 ;
      RECT 41.73 3.178 41.735 3.357 ;
      RECT 41.72 3.182 41.73 3.364 ;
      RECT 41.705 3.19 41.72 3.375 ;
      RECT 41.695 3.2 41.705 3.386 ;
      RECT 41.685 3.207 41.695 3.394 ;
      RECT 41.66 3.22 41.685 3.409 ;
      RECT 41.596 3.256 41.66 3.448 ;
      RECT 41.51 3.319 41.596 3.512 ;
      RECT 41.475 3.37 41.51 3.565 ;
      RECT 41.47 3.387 41.475 3.582 ;
      RECT 41.455 3.396 41.47 3.589 ;
      RECT 41.435 3.411 41.455 3.603 ;
      RECT 41.43 3.422 41.435 3.613 ;
      RECT 41.41 3.435 41.43 3.623 ;
      RECT 41.405 3.445 41.41 3.633 ;
      RECT 41.39 3.45 41.405 3.642 ;
      RECT 41.38 3.46 41.39 3.653 ;
      RECT 41.35 3.477 41.38 3.67 ;
      RECT 41.34 3.495 41.35 3.688 ;
      RECT 41.325 3.506 41.34 3.699 ;
      RECT 41.285 3.53 41.325 3.715 ;
      RECT 41.25 3.564 41.285 3.732 ;
      RECT 41.22 3.587 41.25 3.744 ;
      RECT 41.205 3.597 41.22 3.753 ;
      RECT 41.165 3.607 41.205 3.764 ;
      RECT 41.145 3.618 41.165 3.776 ;
      RECT 41.14 3.622 41.145 3.783 ;
      RECT 41.125 3.626 41.14 3.788 ;
      RECT 41.115 3.631 41.125 3.793 ;
      RECT 41.11 3.634 41.115 3.796 ;
      RECT 41.08 3.64 41.11 3.803 ;
      RECT 41.045 3.65 41.08 3.817 ;
      RECT 40.985 3.665 41.045 3.837 ;
      RECT 40.93 3.685 40.985 3.861 ;
      RECT 40.901 3.7 40.93 3.879 ;
      RECT 40.815 3.72 40.901 3.904 ;
      RECT 40.81 3.735 40.815 3.924 ;
      RECT 40.8 3.738 40.81 3.925 ;
      RECT 40.775 3.745 40.8 4.01 ;
      RECT 43.47 4.238 43.75 4.575 ;
      RECT 43.47 4.248 43.755 4.533 ;
      RECT 43.47 4.257 43.76 4.43 ;
      RECT 43.47 4.272 43.765 4.298 ;
      RECT 43.47 4.1 43.73 4.575 ;
      RECT 33.825 8.945 34.175 9.295 ;
      RECT 42.65 8.9 43 9.25 ;
      RECT 33.825 8.975 43 9.175 ;
      RECT 41.19 4.98 41.2 5.17 ;
      RECT 39.45 4.855 39.73 5.135 ;
      RECT 42.495 3.795 42.5 4.28 ;
      RECT 42.39 3.795 42.45 4.055 ;
      RECT 42.715 4.765 42.72 4.84 ;
      RECT 42.705 4.632 42.715 4.875 ;
      RECT 42.695 4.467 42.705 4.896 ;
      RECT 42.69 4.337 42.695 4.912 ;
      RECT 42.68 4.227 42.69 4.928 ;
      RECT 42.675 4.126 42.68 4.945 ;
      RECT 42.67 4.108 42.675 4.955 ;
      RECT 42.665 4.09 42.67 4.965 ;
      RECT 42.655 4.065 42.665 4.98 ;
      RECT 42.65 4.045 42.655 4.995 ;
      RECT 42.63 3.795 42.65 5.02 ;
      RECT 42.615 3.795 42.63 5.053 ;
      RECT 42.585 3.795 42.615 5.075 ;
      RECT 42.565 3.795 42.585 5.089 ;
      RECT 42.545 3.795 42.565 4.605 ;
      RECT 42.56 4.672 42.565 5.094 ;
      RECT 42.555 4.702 42.56 5.096 ;
      RECT 42.55 4.715 42.555 5.099 ;
      RECT 42.545 4.725 42.55 5.103 ;
      RECT 42.54 3.795 42.545 4.523 ;
      RECT 42.54 4.735 42.545 5.105 ;
      RECT 42.535 3.795 42.54 4.5 ;
      RECT 42.525 4.757 42.54 5.105 ;
      RECT 42.52 3.795 42.535 4.445 ;
      RECT 42.515 4.782 42.525 5.105 ;
      RECT 42.515 3.795 42.52 4.39 ;
      RECT 42.505 3.795 42.515 4.338 ;
      RECT 42.51 4.795 42.515 5.106 ;
      RECT 42.505 4.807 42.51 5.107 ;
      RECT 42.5 3.795 42.505 4.298 ;
      RECT 42.5 4.82 42.505 5.108 ;
      RECT 42.485 4.835 42.5 5.109 ;
      RECT 42.49 3.795 42.495 4.26 ;
      RECT 42.485 3.795 42.49 4.225 ;
      RECT 42.48 3.795 42.485 4.2 ;
      RECT 42.475 4.862 42.485 5.111 ;
      RECT 42.47 3.795 42.48 4.158 ;
      RECT 42.47 4.88 42.475 5.112 ;
      RECT 42.465 3.795 42.47 4.118 ;
      RECT 42.465 4.887 42.47 5.113 ;
      RECT 42.46 3.795 42.465 4.09 ;
      RECT 42.455 4.905 42.465 5.114 ;
      RECT 42.45 3.795 42.46 4.07 ;
      RECT 42.445 4.925 42.455 5.116 ;
      RECT 42.435 4.942 42.445 5.117 ;
      RECT 42.4 4.965 42.435 5.12 ;
      RECT 42.345 4.983 42.4 5.126 ;
      RECT 42.259 4.991 42.345 5.135 ;
      RECT 42.173 5.002 42.259 5.146 ;
      RECT 42.087 5.012 42.173 5.157 ;
      RECT 42.001 5.022 42.087 5.169 ;
      RECT 41.915 5.032 42.001 5.18 ;
      RECT 41.895 5.038 41.915 5.186 ;
      RECT 41.815 5.04 41.895 5.19 ;
      RECT 41.81 5.039 41.815 5.195 ;
      RECT 41.802 5.038 41.81 5.195 ;
      RECT 41.716 5.034 41.802 5.193 ;
      RECT 41.63 5.026 41.716 5.19 ;
      RECT 41.544 5.017 41.63 5.186 ;
      RECT 41.458 5.009 41.544 5.183 ;
      RECT 41.372 5.001 41.458 5.179 ;
      RECT 41.286 4.992 41.372 5.176 ;
      RECT 41.2 4.984 41.286 5.172 ;
      RECT 41.145 4.977 41.19 5.17 ;
      RECT 41.06 4.97 41.145 5.168 ;
      RECT 40.986 4.962 41.06 5.164 ;
      RECT 40.9 4.954 40.986 5.161 ;
      RECT 40.897 4.95 40.9 5.159 ;
      RECT 40.811 4.946 40.897 5.158 ;
      RECT 40.725 4.938 40.811 5.155 ;
      RECT 40.64 4.933 40.725 5.152 ;
      RECT 40.554 4.93 40.64 5.149 ;
      RECT 40.468 4.928 40.554 5.146 ;
      RECT 40.382 4.925 40.468 5.143 ;
      RECT 40.296 4.922 40.382 5.14 ;
      RECT 40.21 4.919 40.296 5.137 ;
      RECT 40.134 4.917 40.21 5.134 ;
      RECT 40.048 4.914 40.134 5.131 ;
      RECT 39.962 4.911 40.048 5.129 ;
      RECT 39.876 4.909 39.962 5.126 ;
      RECT 39.79 4.906 39.876 5.123 ;
      RECT 39.73 4.897 39.79 5.121 ;
      RECT 42.24 4.515 42.315 4.775 ;
      RECT 42.22 4.495 42.225 4.775 ;
      RECT 41.54 4.28 41.645 4.575 ;
      RECT 35.985 4.255 36.055 4.515 ;
      RECT 41.88 4.13 41.885 4.501 ;
      RECT 41.87 4.185 41.875 4.501 ;
      RECT 42.175 3.355 42.235 3.615 ;
      RECT 42.23 4.51 42.24 4.775 ;
      RECT 42.225 4.5 42.23 4.775 ;
      RECT 42.145 4.447 42.22 4.775 ;
      RECT 42.17 3.355 42.175 3.635 ;
      RECT 42.16 3.355 42.17 3.655 ;
      RECT 42.145 3.355 42.16 3.685 ;
      RECT 42.13 3.355 42.145 3.728 ;
      RECT 42.125 4.39 42.145 4.775 ;
      RECT 42.115 3.355 42.13 3.765 ;
      RECT 42.11 4.37 42.125 4.775 ;
      RECT 42.11 3.355 42.115 3.788 ;
      RECT 42.1 3.355 42.11 3.813 ;
      RECT 42.07 4.337 42.11 4.775 ;
      RECT 42.075 3.355 42.1 3.863 ;
      RECT 42.07 3.355 42.075 3.918 ;
      RECT 42.065 3.355 42.07 3.96 ;
      RECT 42.055 4.3 42.07 4.775 ;
      RECT 42.06 3.355 42.065 4.003 ;
      RECT 42.055 3.355 42.06 4.068 ;
      RECT 42.05 3.355 42.055 4.09 ;
      RECT 42.05 4.288 42.055 4.64 ;
      RECT 42.045 3.355 42.05 4.158 ;
      RECT 42.045 4.28 42.05 4.623 ;
      RECT 42.04 3.355 42.045 4.203 ;
      RECT 42.035 4.262 42.045 4.6 ;
      RECT 42.035 3.355 42.04 4.24 ;
      RECT 42.025 3.355 42.035 4.58 ;
      RECT 42.02 3.355 42.025 4.563 ;
      RECT 42.015 3.355 42.02 4.548 ;
      RECT 42.01 3.355 42.015 4.533 ;
      RECT 41.99 3.355 42.01 4.523 ;
      RECT 41.985 3.355 41.99 4.513 ;
      RECT 41.975 3.355 41.985 4.509 ;
      RECT 41.97 3.632 41.975 4.508 ;
      RECT 41.965 3.655 41.97 4.507 ;
      RECT 41.96 3.685 41.965 4.506 ;
      RECT 41.955 3.712 41.96 4.505 ;
      RECT 41.95 3.74 41.955 4.505 ;
      RECT 41.945 3.767 41.95 4.505 ;
      RECT 41.94 3.787 41.945 4.505 ;
      RECT 41.935 3.815 41.94 4.505 ;
      RECT 41.925 3.857 41.935 4.505 ;
      RECT 41.915 3.902 41.925 4.504 ;
      RECT 41.91 3.955 41.915 4.503 ;
      RECT 41.905 3.987 41.91 4.502 ;
      RECT 41.9 4.007 41.905 4.501 ;
      RECT 41.895 4.045 41.9 4.501 ;
      RECT 41.89 4.067 41.895 4.501 ;
      RECT 41.885 4.092 41.89 4.501 ;
      RECT 41.875 4.157 41.88 4.501 ;
      RECT 41.86 4.217 41.87 4.501 ;
      RECT 41.845 4.227 41.86 4.501 ;
      RECT 41.825 4.237 41.845 4.501 ;
      RECT 41.795 4.242 41.825 4.498 ;
      RECT 41.735 4.252 41.795 4.495 ;
      RECT 41.715 4.261 41.735 4.5 ;
      RECT 41.69 4.267 41.715 4.513 ;
      RECT 41.67 4.272 41.69 4.528 ;
      RECT 41.645 4.277 41.67 4.575 ;
      RECT 41.516 4.279 41.54 4.575 ;
      RECT 41.43 4.274 41.516 4.575 ;
      RECT 41.39 4.271 41.43 4.575 ;
      RECT 41.34 4.273 41.39 4.555 ;
      RECT 41.31 4.277 41.34 4.555 ;
      RECT 41.231 4.287 41.31 4.555 ;
      RECT 41.145 4.302 41.231 4.556 ;
      RECT 41.095 4.312 41.145 4.557 ;
      RECT 41.087 4.315 41.095 4.557 ;
      RECT 41.001 4.317 41.087 4.558 ;
      RECT 40.915 4.321 41.001 4.558 ;
      RECT 40.829 4.325 40.915 4.559 ;
      RECT 40.743 4.328 40.829 4.56 ;
      RECT 40.657 4.332 40.743 4.56 ;
      RECT 40.571 4.336 40.657 4.561 ;
      RECT 40.485 4.339 40.571 4.562 ;
      RECT 40.399 4.343 40.485 4.562 ;
      RECT 40.313 4.347 40.399 4.563 ;
      RECT 40.227 4.351 40.313 4.564 ;
      RECT 40.141 4.354 40.227 4.564 ;
      RECT 40.055 4.358 40.141 4.565 ;
      RECT 40.025 4.36 40.055 4.565 ;
      RECT 39.939 4.363 40.025 4.566 ;
      RECT 39.853 4.367 39.939 4.567 ;
      RECT 39.767 4.371 39.853 4.568 ;
      RECT 39.681 4.374 39.767 4.568 ;
      RECT 39.595 4.378 39.681 4.569 ;
      RECT 39.56 4.383 39.595 4.57 ;
      RECT 39.505 4.393 39.56 4.577 ;
      RECT 39.48 4.405 39.505 4.587 ;
      RECT 39.445 4.418 39.48 4.595 ;
      RECT 39.405 4.435 39.445 4.618 ;
      RECT 39.385 4.448 39.405 4.645 ;
      RECT 39.355 4.46 39.385 4.673 ;
      RECT 39.35 4.468 39.355 4.693 ;
      RECT 39.345 4.471 39.35 4.703 ;
      RECT 39.295 4.483 39.345 4.737 ;
      RECT 39.285 4.498 39.295 4.77 ;
      RECT 39.275 4.504 39.285 4.783 ;
      RECT 39.265 4.511 39.275 4.795 ;
      RECT 39.24 4.524 39.265 4.813 ;
      RECT 39.225 4.539 39.24 4.835 ;
      RECT 39.215 4.547 39.225 4.851 ;
      RECT 39.2 4.556 39.215 4.866 ;
      RECT 39.19 4.566 39.2 4.88 ;
      RECT 39.171 4.579 39.19 4.897 ;
      RECT 39.085 4.624 39.171 4.962 ;
      RECT 39.07 4.669 39.085 5.02 ;
      RECT 39.065 4.678 39.07 5.033 ;
      RECT 39.055 4.685 39.065 5.038 ;
      RECT 39.05 4.69 39.055 5.042 ;
      RECT 39.03 4.7 39.05 5.049 ;
      RECT 39.005 4.72 39.03 5.063 ;
      RECT 38.97 4.745 39.005 5.083 ;
      RECT 38.955 4.768 38.97 5.098 ;
      RECT 38.945 4.778 38.955 5.103 ;
      RECT 38.935 4.786 38.945 5.11 ;
      RECT 38.925 4.795 38.935 5.116 ;
      RECT 38.905 4.807 38.925 5.118 ;
      RECT 38.895 4.82 38.905 5.12 ;
      RECT 38.87 4.835 38.895 5.123 ;
      RECT 38.85 4.852 38.87 5.127 ;
      RECT 38.81 4.88 38.85 5.133 ;
      RECT 38.745 4.927 38.81 5.142 ;
      RECT 38.73 4.96 38.745 5.15 ;
      RECT 38.725 4.967 38.73 5.152 ;
      RECT 38.675 4.992 38.725 5.157 ;
      RECT 38.66 5.016 38.675 5.164 ;
      RECT 38.61 5.021 38.66 5.165 ;
      RECT 38.524 5.025 38.61 5.165 ;
      RECT 38.438 5.025 38.524 5.165 ;
      RECT 38.352 5.025 38.438 5.166 ;
      RECT 38.266 5.025 38.352 5.166 ;
      RECT 38.18 5.025 38.266 5.166 ;
      RECT 38.114 5.025 38.18 5.166 ;
      RECT 38.028 5.025 38.114 5.167 ;
      RECT 37.942 5.025 38.028 5.167 ;
      RECT 37.856 5.026 37.942 5.168 ;
      RECT 37.77 5.026 37.856 5.168 ;
      RECT 37.684 5.026 37.77 5.168 ;
      RECT 37.598 5.026 37.684 5.169 ;
      RECT 37.512 5.026 37.598 5.169 ;
      RECT 37.426 5.027 37.512 5.17 ;
      RECT 37.34 5.027 37.426 5.17 ;
      RECT 37.32 5.027 37.34 5.17 ;
      RECT 37.234 5.027 37.32 5.17 ;
      RECT 37.148 5.027 37.234 5.17 ;
      RECT 37.062 5.028 37.148 5.17 ;
      RECT 36.976 5.028 37.062 5.17 ;
      RECT 36.89 5.028 36.976 5.17 ;
      RECT 36.804 5.029 36.89 5.17 ;
      RECT 36.718 5.029 36.804 5.17 ;
      RECT 36.632 5.029 36.718 5.17 ;
      RECT 36.546 5.029 36.632 5.17 ;
      RECT 36.46 5.03 36.546 5.17 ;
      RECT 36.41 5.027 36.46 5.17 ;
      RECT 36.4 5.025 36.41 5.169 ;
      RECT 36.396 5.025 36.4 5.168 ;
      RECT 36.31 5.02 36.396 5.163 ;
      RECT 36.288 5.013 36.31 5.157 ;
      RECT 36.202 5.004 36.288 5.151 ;
      RECT 36.116 4.991 36.202 5.142 ;
      RECT 36.03 4.977 36.116 5.132 ;
      RECT 35.985 4.967 36.03 5.125 ;
      RECT 35.965 4.255 35.985 4.533 ;
      RECT 35.965 4.96 35.985 5.121 ;
      RECT 35.935 4.255 35.965 4.555 ;
      RECT 35.925 4.927 35.965 5.118 ;
      RECT 35.92 4.255 35.935 4.575 ;
      RECT 35.92 4.892 35.925 5.116 ;
      RECT 35.915 4.255 35.92 4.7 ;
      RECT 35.915 4.852 35.92 5.116 ;
      RECT 35.905 4.255 35.915 5.116 ;
      RECT 35.83 4.255 35.905 5.11 ;
      RECT 35.8 4.255 35.83 5.1 ;
      RECT 35.795 4.255 35.8 5.092 ;
      RECT 35.79 4.297 35.795 5.085 ;
      RECT 35.78 4.366 35.79 5.076 ;
      RECT 35.775 4.436 35.78 5.028 ;
      RECT 35.77 4.5 35.775 4.925 ;
      RECT 35.765 4.535 35.77 4.88 ;
      RECT 35.763 4.572 35.765 4.772 ;
      RECT 35.76 4.58 35.763 4.765 ;
      RECT 35.755 4.645 35.76 4.708 ;
      RECT 39.83 3.735 40.11 4.015 ;
      RECT 39.82 3.735 40.11 3.878 ;
      RECT 39.775 3.6 40.035 3.86 ;
      RECT 39.775 3.715 40.09 3.86 ;
      RECT 39.775 3.685 40.085 3.86 ;
      RECT 39.775 3.672 40.075 3.86 ;
      RECT 39.775 3.662 40.07 3.86 ;
      RECT 35.75 3.645 36.01 3.905 ;
      RECT 39.52 3.195 39.78 3.455 ;
      RECT 39.51 3.22 39.78 3.415 ;
      RECT 39.505 3.22 39.51 3.414 ;
      RECT 39.435 3.215 39.505 3.406 ;
      RECT 39.35 3.202 39.435 3.389 ;
      RECT 39.346 3.194 39.35 3.379 ;
      RECT 39.26 3.187 39.346 3.369 ;
      RECT 39.251 3.179 39.26 3.359 ;
      RECT 39.165 3.172 39.251 3.347 ;
      RECT 39.145 3.163 39.165 3.333 ;
      RECT 39.09 3.158 39.145 3.325 ;
      RECT 39.08 3.152 39.09 3.319 ;
      RECT 39.06 3.15 39.08 3.315 ;
      RECT 39.052 3.149 39.06 3.311 ;
      RECT 38.966 3.141 39.052 3.3 ;
      RECT 38.88 3.127 38.966 3.28 ;
      RECT 38.82 3.115 38.88 3.265 ;
      RECT 38.81 3.11 38.82 3.26 ;
      RECT 38.76 3.11 38.81 3.262 ;
      RECT 38.713 3.112 38.76 3.266 ;
      RECT 38.627 3.119 38.713 3.271 ;
      RECT 38.541 3.127 38.627 3.277 ;
      RECT 38.455 3.136 38.541 3.283 ;
      RECT 38.396 3.142 38.455 3.288 ;
      RECT 38.31 3.147 38.396 3.294 ;
      RECT 38.235 3.152 38.31 3.3 ;
      RECT 38.196 3.154 38.235 3.305 ;
      RECT 38.11 3.151 38.196 3.31 ;
      RECT 38.025 3.149 38.11 3.317 ;
      RECT 37.993 3.148 38.025 3.32 ;
      RECT 37.907 3.147 37.993 3.321 ;
      RECT 37.821 3.146 37.907 3.322 ;
      RECT 37.735 3.145 37.821 3.322 ;
      RECT 37.649 3.144 37.735 3.323 ;
      RECT 37.563 3.143 37.649 3.324 ;
      RECT 37.477 3.142 37.563 3.325 ;
      RECT 37.391 3.141 37.477 3.325 ;
      RECT 37.305 3.14 37.391 3.326 ;
      RECT 37.255 3.14 37.305 3.327 ;
      RECT 37.241 3.141 37.255 3.327 ;
      RECT 37.155 3.148 37.241 3.328 ;
      RECT 37.081 3.159 37.155 3.329 ;
      RECT 36.995 3.168 37.081 3.33 ;
      RECT 36.96 3.175 36.995 3.345 ;
      RECT 36.935 3.178 36.96 3.375 ;
      RECT 36.91 3.187 36.935 3.404 ;
      RECT 36.9 3.198 36.91 3.424 ;
      RECT 36.89 3.206 36.9 3.438 ;
      RECT 36.885 3.212 36.89 3.448 ;
      RECT 36.86 3.229 36.885 3.465 ;
      RECT 36.845 3.251 36.86 3.493 ;
      RECT 36.815 3.277 36.845 3.523 ;
      RECT 36.795 3.306 36.815 3.553 ;
      RECT 36.79 3.321 36.795 3.57 ;
      RECT 36.77 3.336 36.79 3.585 ;
      RECT 36.76 3.354 36.77 3.603 ;
      RECT 36.75 3.365 36.76 3.618 ;
      RECT 36.7 3.397 36.75 3.644 ;
      RECT 36.695 3.427 36.7 3.664 ;
      RECT 36.685 3.44 36.695 3.67 ;
      RECT 36.676 3.45 36.685 3.678 ;
      RECT 36.665 3.461 36.676 3.686 ;
      RECT 36.66 3.471 36.665 3.692 ;
      RECT 36.645 3.492 36.66 3.699 ;
      RECT 36.63 3.522 36.645 3.707 ;
      RECT 36.595 3.552 36.63 3.713 ;
      RECT 36.57 3.57 36.595 3.72 ;
      RECT 36.52 3.578 36.57 3.729 ;
      RECT 36.495 3.583 36.52 3.738 ;
      RECT 36.44 3.589 36.495 3.748 ;
      RECT 36.435 3.594 36.44 3.756 ;
      RECT 36.421 3.597 36.435 3.758 ;
      RECT 36.335 3.609 36.421 3.77 ;
      RECT 36.325 3.621 36.335 3.783 ;
      RECT 36.24 3.634 36.325 3.795 ;
      RECT 36.196 3.651 36.24 3.809 ;
      RECT 36.11 3.668 36.196 3.825 ;
      RECT 36.08 3.682 36.11 3.839 ;
      RECT 36.07 3.687 36.08 3.844 ;
      RECT 36.01 3.69 36.07 3.853 ;
      RECT 38.9 3.96 39.16 4.22 ;
      RECT 38.9 3.96 39.18 4.073 ;
      RECT 38.9 3.96 39.205 4.04 ;
      RECT 38.9 3.96 39.21 4.02 ;
      RECT 38.95 3.735 39.23 4.015 ;
      RECT 38.505 4.47 38.765 4.73 ;
      RECT 38.495 4.327 38.69 4.668 ;
      RECT 38.49 4.435 38.705 4.66 ;
      RECT 38.485 4.485 38.765 4.65 ;
      RECT 38.475 4.562 38.765 4.635 ;
      RECT 38.495 4.41 38.705 4.668 ;
      RECT 38.505 4.285 38.69 4.73 ;
      RECT 38.505 4.18 38.67 4.73 ;
      RECT 38.515 4.167 38.67 4.73 ;
      RECT 38.515 4.125 38.66 4.73 ;
      RECT 38.52 4.05 38.66 4.73 ;
      RECT 38.55 3.7 38.66 4.73 ;
      RECT 38.555 3.43 38.68 4.053 ;
      RECT 38.525 4.005 38.68 4.053 ;
      RECT 38.54 3.807 38.66 4.73 ;
      RECT 38.53 3.917 38.68 4.053 ;
      RECT 38.555 3.43 38.695 3.91 ;
      RECT 38.555 3.43 38.715 3.785 ;
      RECT 38.52 3.43 38.78 3.69 ;
      RECT 37.99 3.735 38.27 4.015 ;
      RECT 37.975 3.735 38.27 3.995 ;
      RECT 36.03 4.6 36.29 4.86 ;
      RECT 37.815 4.455 38.075 4.715 ;
      RECT 37.795 4.475 38.075 4.69 ;
      RECT 37.752 4.475 37.795 4.689 ;
      RECT 37.666 4.476 37.752 4.686 ;
      RECT 37.58 4.477 37.666 4.682 ;
      RECT 37.505 4.479 37.58 4.679 ;
      RECT 37.482 4.48 37.505 4.677 ;
      RECT 37.396 4.481 37.482 4.675 ;
      RECT 37.31 4.482 37.396 4.672 ;
      RECT 37.286 4.483 37.31 4.67 ;
      RECT 37.2 4.485 37.286 4.667 ;
      RECT 37.115 4.487 37.2 4.668 ;
      RECT 37.058 4.488 37.115 4.674 ;
      RECT 36.972 4.49 37.058 4.684 ;
      RECT 36.886 4.493 36.972 4.697 ;
      RECT 36.8 4.495 36.886 4.709 ;
      RECT 36.786 4.496 36.8 4.716 ;
      RECT 36.7 4.497 36.786 4.724 ;
      RECT 36.66 4.499 36.7 4.733 ;
      RECT 36.651 4.5 36.66 4.736 ;
      RECT 36.565 4.508 36.651 4.742 ;
      RECT 36.545 4.517 36.565 4.75 ;
      RECT 36.46 4.532 36.545 4.758 ;
      RECT 36.4 4.555 36.46 4.769 ;
      RECT 36.39 4.567 36.4 4.774 ;
      RECT 36.35 4.577 36.39 4.778 ;
      RECT 36.295 4.594 36.35 4.786 ;
      RECT 36.29 4.604 36.295 4.79 ;
      RECT 37.356 3.735 37.415 4.132 ;
      RECT 37.27 3.735 37.475 4.123 ;
      RECT 37.265 3.765 37.475 4.118 ;
      RECT 37.231 3.765 37.475 4.116 ;
      RECT 37.145 3.765 37.475 4.11 ;
      RECT 37.1 3.765 37.495 4.088 ;
      RECT 37.1 3.765 37.515 4.043 ;
      RECT 37.06 3.765 37.515 4.033 ;
      RECT 37.27 3.735 37.55 4.015 ;
      RECT 37.005 3.735 37.265 3.995 ;
      RECT 34.83 4.295 35.11 4.575 ;
      RECT 34.8 4.257 35.055 4.56 ;
      RECT 34.795 4.258 35.055 4.558 ;
      RECT 34.79 4.259 35.055 4.552 ;
      RECT 34.785 4.262 35.055 4.545 ;
      RECT 34.78 4.295 35.11 4.538 ;
      RECT 34.75 4.265 35.055 4.525 ;
      RECT 34.75 4.292 35.075 4.525 ;
      RECT 34.75 4.282 35.07 4.525 ;
      RECT 34.75 4.267 35.065 4.525 ;
      RECT 34.83 4.254 35.045 4.575 ;
      RECT 34.916 4.252 35.045 4.575 ;
      RECT 35.002 4.25 35.03 4.575 ;
      RECT 30.645 8.505 30.965 8.83 ;
      RECT 30.675 7.98 30.845 8.83 ;
      RECT 30.675 7.98 30.85 8.33 ;
      RECT 30.675 7.98 31.65 8.155 ;
      RECT 31.475 3.26 31.65 8.155 ;
      RECT 31.42 3.26 31.77 3.61 ;
      RECT 31.445 8.94 31.77 9.265 ;
      RECT 30.33 9.03 31.77 9.2 ;
      RECT 30.33 3.69 30.49 9.2 ;
      RECT 30.645 3.66 30.965 3.98 ;
      RECT 30.33 3.69 30.965 3.86 ;
      RECT 20.415 3.215 20.675 3.475 ;
      RECT 20.47 3.175 20.775 3.455 ;
      RECT 20.47 2.715 20.645 3.475 ;
      RECT 28.985 2.635 29.335 2.985 ;
      RECT 20.47 2.715 29.335 2.89 ;
      RECT 28.66 4.145 29.03 4.515 ;
      RECT 28.745 3.53 28.915 4.515 ;
      RECT 24.765 3.75 25 4.01 ;
      RECT 27.91 3.53 28.075 3.79 ;
      RECT 27.815 3.52 27.83 3.79 ;
      RECT 27.91 3.53 28.915 3.71 ;
      RECT 26.415 3.09 26.455 3.23 ;
      RECT 27.83 3.525 27.91 3.79 ;
      RECT 27.775 3.52 27.815 3.756 ;
      RECT 27.761 3.52 27.775 3.756 ;
      RECT 27.675 3.525 27.761 3.758 ;
      RECT 27.63 3.532 27.675 3.76 ;
      RECT 27.6 3.532 27.63 3.762 ;
      RECT 27.575 3.527 27.6 3.764 ;
      RECT 27.545 3.523 27.575 3.773 ;
      RECT 27.535 3.52 27.545 3.785 ;
      RECT 27.53 3.52 27.535 3.793 ;
      RECT 27.525 3.52 27.53 3.798 ;
      RECT 27.515 3.519 27.525 3.808 ;
      RECT 27.51 3.518 27.515 3.818 ;
      RECT 27.495 3.517 27.51 3.823 ;
      RECT 27.467 3.514 27.495 3.85 ;
      RECT 27.381 3.506 27.467 3.85 ;
      RECT 27.295 3.495 27.381 3.85 ;
      RECT 27.255 3.48 27.295 3.85 ;
      RECT 27.215 3.454 27.255 3.85 ;
      RECT 27.21 3.436 27.215 3.662 ;
      RECT 27.2 3.432 27.21 3.652 ;
      RECT 27.185 3.422 27.2 3.639 ;
      RECT 27.165 3.406 27.185 3.624 ;
      RECT 27.15 3.391 27.165 3.609 ;
      RECT 27.14 3.38 27.15 3.599 ;
      RECT 27.115 3.364 27.14 3.588 ;
      RECT 27.11 3.351 27.115 3.578 ;
      RECT 27.105 3.347 27.11 3.573 ;
      RECT 27.05 3.333 27.105 3.551 ;
      RECT 27.011 3.314 27.05 3.515 ;
      RECT 26.925 3.288 27.011 3.468 ;
      RECT 26.921 3.27 26.925 3.434 ;
      RECT 26.835 3.251 26.921 3.412 ;
      RECT 26.83 3.233 26.835 3.39 ;
      RECT 26.825 3.231 26.83 3.388 ;
      RECT 26.815 3.23 26.825 3.383 ;
      RECT 26.755 3.217 26.815 3.369 ;
      RECT 26.71 3.195 26.755 3.348 ;
      RECT 26.65 3.172 26.71 3.327 ;
      RECT 26.586 3.147 26.65 3.302 ;
      RECT 26.5 3.117 26.586 3.271 ;
      RECT 26.485 3.097 26.5 3.25 ;
      RECT 26.455 3.092 26.485 3.241 ;
      RECT 26.402 3.09 26.415 3.23 ;
      RECT 26.316 3.09 26.402 3.232 ;
      RECT 26.23 3.09 26.316 3.234 ;
      RECT 26.21 3.09 26.23 3.238 ;
      RECT 26.165 3.092 26.21 3.249 ;
      RECT 26.125 3.102 26.165 3.265 ;
      RECT 26.121 3.111 26.125 3.273 ;
      RECT 26.035 3.131 26.121 3.289 ;
      RECT 26.025 3.15 26.035 3.307 ;
      RECT 26.02 3.152 26.025 3.31 ;
      RECT 26.01 3.156 26.02 3.313 ;
      RECT 25.99 3.161 26.01 3.323 ;
      RECT 25.96 3.171 25.99 3.343 ;
      RECT 25.955 3.178 25.96 3.357 ;
      RECT 25.945 3.182 25.955 3.364 ;
      RECT 25.93 3.19 25.945 3.375 ;
      RECT 25.92 3.2 25.93 3.386 ;
      RECT 25.91 3.207 25.92 3.394 ;
      RECT 25.885 3.22 25.91 3.409 ;
      RECT 25.821 3.256 25.885 3.448 ;
      RECT 25.735 3.319 25.821 3.512 ;
      RECT 25.7 3.37 25.735 3.565 ;
      RECT 25.695 3.387 25.7 3.582 ;
      RECT 25.68 3.396 25.695 3.589 ;
      RECT 25.66 3.411 25.68 3.603 ;
      RECT 25.655 3.422 25.66 3.613 ;
      RECT 25.635 3.435 25.655 3.623 ;
      RECT 25.63 3.445 25.635 3.633 ;
      RECT 25.615 3.45 25.63 3.642 ;
      RECT 25.605 3.46 25.615 3.653 ;
      RECT 25.575 3.477 25.605 3.67 ;
      RECT 25.565 3.495 25.575 3.688 ;
      RECT 25.55 3.506 25.565 3.699 ;
      RECT 25.51 3.53 25.55 3.715 ;
      RECT 25.475 3.564 25.51 3.732 ;
      RECT 25.445 3.587 25.475 3.744 ;
      RECT 25.43 3.597 25.445 3.753 ;
      RECT 25.39 3.607 25.43 3.764 ;
      RECT 25.37 3.618 25.39 3.776 ;
      RECT 25.365 3.622 25.37 3.783 ;
      RECT 25.35 3.626 25.365 3.788 ;
      RECT 25.34 3.631 25.35 3.793 ;
      RECT 25.335 3.634 25.34 3.796 ;
      RECT 25.305 3.64 25.335 3.803 ;
      RECT 25.27 3.65 25.305 3.817 ;
      RECT 25.21 3.665 25.27 3.837 ;
      RECT 25.155 3.685 25.21 3.861 ;
      RECT 25.126 3.7 25.155 3.879 ;
      RECT 25.04 3.72 25.126 3.904 ;
      RECT 25.035 3.735 25.04 3.924 ;
      RECT 25.025 3.738 25.035 3.925 ;
      RECT 25 3.745 25.025 4.01 ;
      RECT 27.695 4.238 27.975 4.575 ;
      RECT 27.695 4.248 27.98 4.533 ;
      RECT 27.695 4.257 27.985 4.43 ;
      RECT 27.695 4.272 27.99 4.298 ;
      RECT 27.695 4.1 27.955 4.575 ;
      RECT 18.045 8.94 18.395 9.29 ;
      RECT 26.87 8.895 27.22 9.245 ;
      RECT 18.045 8.97 27.22 9.17 ;
      RECT 25.415 4.98 25.425 5.17 ;
      RECT 23.675 4.855 23.955 5.135 ;
      RECT 26.72 3.795 26.725 4.28 ;
      RECT 26.615 3.795 26.675 4.055 ;
      RECT 26.94 4.765 26.945 4.84 ;
      RECT 26.93 4.632 26.94 4.875 ;
      RECT 26.92 4.467 26.93 4.896 ;
      RECT 26.915 4.337 26.92 4.912 ;
      RECT 26.905 4.227 26.915 4.928 ;
      RECT 26.9 4.126 26.905 4.945 ;
      RECT 26.895 4.108 26.9 4.955 ;
      RECT 26.89 4.09 26.895 4.965 ;
      RECT 26.88 4.065 26.89 4.98 ;
      RECT 26.875 4.045 26.88 4.995 ;
      RECT 26.855 3.795 26.875 5.02 ;
      RECT 26.84 3.795 26.855 5.053 ;
      RECT 26.81 3.795 26.84 5.075 ;
      RECT 26.79 3.795 26.81 5.089 ;
      RECT 26.77 3.795 26.79 4.605 ;
      RECT 26.785 4.672 26.79 5.094 ;
      RECT 26.78 4.702 26.785 5.096 ;
      RECT 26.775 4.715 26.78 5.099 ;
      RECT 26.77 4.725 26.775 5.103 ;
      RECT 26.765 3.795 26.77 4.523 ;
      RECT 26.765 4.735 26.77 5.105 ;
      RECT 26.76 3.795 26.765 4.5 ;
      RECT 26.75 4.757 26.765 5.105 ;
      RECT 26.745 3.795 26.76 4.445 ;
      RECT 26.74 4.782 26.75 5.105 ;
      RECT 26.74 3.795 26.745 4.39 ;
      RECT 26.73 3.795 26.74 4.338 ;
      RECT 26.735 4.795 26.74 5.106 ;
      RECT 26.73 4.807 26.735 5.107 ;
      RECT 26.725 3.795 26.73 4.298 ;
      RECT 26.725 4.82 26.73 5.108 ;
      RECT 26.71 4.835 26.725 5.109 ;
      RECT 26.715 3.795 26.72 4.26 ;
      RECT 26.71 3.795 26.715 4.225 ;
      RECT 26.705 3.795 26.71 4.2 ;
      RECT 26.7 4.862 26.71 5.111 ;
      RECT 26.695 3.795 26.705 4.158 ;
      RECT 26.695 4.88 26.7 5.112 ;
      RECT 26.69 3.795 26.695 4.118 ;
      RECT 26.69 4.887 26.695 5.113 ;
      RECT 26.685 3.795 26.69 4.09 ;
      RECT 26.68 4.905 26.69 5.114 ;
      RECT 26.675 3.795 26.685 4.07 ;
      RECT 26.67 4.925 26.68 5.116 ;
      RECT 26.66 4.942 26.67 5.117 ;
      RECT 26.625 4.965 26.66 5.12 ;
      RECT 26.57 4.983 26.625 5.126 ;
      RECT 26.484 4.991 26.57 5.135 ;
      RECT 26.398 5.002 26.484 5.146 ;
      RECT 26.312 5.012 26.398 5.157 ;
      RECT 26.226 5.022 26.312 5.169 ;
      RECT 26.14 5.032 26.226 5.18 ;
      RECT 26.12 5.038 26.14 5.186 ;
      RECT 26.04 5.04 26.12 5.19 ;
      RECT 26.035 5.039 26.04 5.195 ;
      RECT 26.027 5.038 26.035 5.195 ;
      RECT 25.941 5.034 26.027 5.193 ;
      RECT 25.855 5.026 25.941 5.19 ;
      RECT 25.769 5.017 25.855 5.186 ;
      RECT 25.683 5.009 25.769 5.183 ;
      RECT 25.597 5.001 25.683 5.179 ;
      RECT 25.511 4.992 25.597 5.176 ;
      RECT 25.425 4.984 25.511 5.172 ;
      RECT 25.37 4.977 25.415 5.17 ;
      RECT 25.285 4.97 25.37 5.168 ;
      RECT 25.211 4.962 25.285 5.164 ;
      RECT 25.125 4.954 25.211 5.161 ;
      RECT 25.122 4.95 25.125 5.159 ;
      RECT 25.036 4.946 25.122 5.158 ;
      RECT 24.95 4.938 25.036 5.155 ;
      RECT 24.865 4.933 24.95 5.152 ;
      RECT 24.779 4.93 24.865 5.149 ;
      RECT 24.693 4.928 24.779 5.146 ;
      RECT 24.607 4.925 24.693 5.143 ;
      RECT 24.521 4.922 24.607 5.14 ;
      RECT 24.435 4.919 24.521 5.137 ;
      RECT 24.359 4.917 24.435 5.134 ;
      RECT 24.273 4.914 24.359 5.131 ;
      RECT 24.187 4.911 24.273 5.129 ;
      RECT 24.101 4.909 24.187 5.126 ;
      RECT 24.015 4.906 24.101 5.123 ;
      RECT 23.955 4.897 24.015 5.121 ;
      RECT 26.465 4.515 26.54 4.775 ;
      RECT 26.445 4.495 26.45 4.775 ;
      RECT 25.765 4.28 25.87 4.575 ;
      RECT 20.21 4.255 20.28 4.515 ;
      RECT 26.105 4.13 26.11 4.501 ;
      RECT 26.095 4.185 26.1 4.501 ;
      RECT 26.4 3.355 26.46 3.615 ;
      RECT 26.455 4.51 26.465 4.775 ;
      RECT 26.45 4.5 26.455 4.775 ;
      RECT 26.37 4.447 26.445 4.775 ;
      RECT 26.395 3.355 26.4 3.635 ;
      RECT 26.385 3.355 26.395 3.655 ;
      RECT 26.37 3.355 26.385 3.685 ;
      RECT 26.355 3.355 26.37 3.728 ;
      RECT 26.35 4.39 26.37 4.775 ;
      RECT 26.34 3.355 26.355 3.765 ;
      RECT 26.335 4.37 26.35 4.775 ;
      RECT 26.335 3.355 26.34 3.788 ;
      RECT 26.325 3.355 26.335 3.813 ;
      RECT 26.295 4.337 26.335 4.775 ;
      RECT 26.3 3.355 26.325 3.863 ;
      RECT 26.295 3.355 26.3 3.918 ;
      RECT 26.29 3.355 26.295 3.96 ;
      RECT 26.28 4.3 26.295 4.775 ;
      RECT 26.285 3.355 26.29 4.003 ;
      RECT 26.28 3.355 26.285 4.068 ;
      RECT 26.275 3.355 26.28 4.09 ;
      RECT 26.275 4.288 26.28 4.64 ;
      RECT 26.27 3.355 26.275 4.158 ;
      RECT 26.27 4.28 26.275 4.623 ;
      RECT 26.265 3.355 26.27 4.203 ;
      RECT 26.26 4.262 26.27 4.6 ;
      RECT 26.26 3.355 26.265 4.24 ;
      RECT 26.25 3.355 26.26 4.58 ;
      RECT 26.245 3.355 26.25 4.563 ;
      RECT 26.24 3.355 26.245 4.548 ;
      RECT 26.235 3.355 26.24 4.533 ;
      RECT 26.215 3.355 26.235 4.523 ;
      RECT 26.21 3.355 26.215 4.513 ;
      RECT 26.2 3.355 26.21 4.509 ;
      RECT 26.195 3.632 26.2 4.508 ;
      RECT 26.19 3.655 26.195 4.507 ;
      RECT 26.185 3.685 26.19 4.506 ;
      RECT 26.18 3.712 26.185 4.505 ;
      RECT 26.175 3.74 26.18 4.505 ;
      RECT 26.17 3.767 26.175 4.505 ;
      RECT 26.165 3.787 26.17 4.505 ;
      RECT 26.16 3.815 26.165 4.505 ;
      RECT 26.15 3.857 26.16 4.505 ;
      RECT 26.14 3.902 26.15 4.504 ;
      RECT 26.135 3.955 26.14 4.503 ;
      RECT 26.13 3.987 26.135 4.502 ;
      RECT 26.125 4.007 26.13 4.501 ;
      RECT 26.12 4.045 26.125 4.501 ;
      RECT 26.115 4.067 26.12 4.501 ;
      RECT 26.11 4.092 26.115 4.501 ;
      RECT 26.1 4.157 26.105 4.501 ;
      RECT 26.085 4.217 26.095 4.501 ;
      RECT 26.07 4.227 26.085 4.501 ;
      RECT 26.05 4.237 26.07 4.501 ;
      RECT 26.02 4.242 26.05 4.498 ;
      RECT 25.96 4.252 26.02 4.495 ;
      RECT 25.94 4.261 25.96 4.5 ;
      RECT 25.915 4.267 25.94 4.513 ;
      RECT 25.895 4.272 25.915 4.528 ;
      RECT 25.87 4.277 25.895 4.575 ;
      RECT 25.741 4.279 25.765 4.575 ;
      RECT 25.655 4.274 25.741 4.575 ;
      RECT 25.615 4.271 25.655 4.575 ;
      RECT 25.565 4.273 25.615 4.555 ;
      RECT 25.535 4.277 25.565 4.555 ;
      RECT 25.456 4.287 25.535 4.555 ;
      RECT 25.37 4.302 25.456 4.556 ;
      RECT 25.32 4.312 25.37 4.557 ;
      RECT 25.312 4.315 25.32 4.557 ;
      RECT 25.226 4.317 25.312 4.558 ;
      RECT 25.14 4.321 25.226 4.558 ;
      RECT 25.054 4.325 25.14 4.559 ;
      RECT 24.968 4.328 25.054 4.56 ;
      RECT 24.882 4.332 24.968 4.56 ;
      RECT 24.796 4.336 24.882 4.561 ;
      RECT 24.71 4.339 24.796 4.562 ;
      RECT 24.624 4.343 24.71 4.562 ;
      RECT 24.538 4.347 24.624 4.563 ;
      RECT 24.452 4.351 24.538 4.564 ;
      RECT 24.366 4.354 24.452 4.564 ;
      RECT 24.28 4.358 24.366 4.565 ;
      RECT 24.25 4.36 24.28 4.565 ;
      RECT 24.164 4.363 24.25 4.566 ;
      RECT 24.078 4.367 24.164 4.567 ;
      RECT 23.992 4.371 24.078 4.568 ;
      RECT 23.906 4.374 23.992 4.568 ;
      RECT 23.82 4.378 23.906 4.569 ;
      RECT 23.785 4.383 23.82 4.57 ;
      RECT 23.73 4.393 23.785 4.577 ;
      RECT 23.705 4.405 23.73 4.587 ;
      RECT 23.67 4.418 23.705 4.595 ;
      RECT 23.63 4.435 23.67 4.618 ;
      RECT 23.61 4.448 23.63 4.645 ;
      RECT 23.58 4.46 23.61 4.673 ;
      RECT 23.575 4.468 23.58 4.693 ;
      RECT 23.57 4.471 23.575 4.703 ;
      RECT 23.52 4.483 23.57 4.737 ;
      RECT 23.51 4.498 23.52 4.77 ;
      RECT 23.5 4.504 23.51 4.783 ;
      RECT 23.49 4.511 23.5 4.795 ;
      RECT 23.465 4.524 23.49 4.813 ;
      RECT 23.45 4.539 23.465 4.835 ;
      RECT 23.44 4.547 23.45 4.851 ;
      RECT 23.425 4.556 23.44 4.866 ;
      RECT 23.415 4.566 23.425 4.88 ;
      RECT 23.396 4.579 23.415 4.897 ;
      RECT 23.31 4.624 23.396 4.962 ;
      RECT 23.295 4.669 23.31 5.02 ;
      RECT 23.29 4.678 23.295 5.033 ;
      RECT 23.28 4.685 23.29 5.038 ;
      RECT 23.275 4.69 23.28 5.042 ;
      RECT 23.255 4.7 23.275 5.049 ;
      RECT 23.23 4.72 23.255 5.063 ;
      RECT 23.195 4.745 23.23 5.083 ;
      RECT 23.18 4.768 23.195 5.098 ;
      RECT 23.17 4.778 23.18 5.103 ;
      RECT 23.16 4.786 23.17 5.11 ;
      RECT 23.15 4.795 23.16 5.116 ;
      RECT 23.13 4.807 23.15 5.118 ;
      RECT 23.12 4.82 23.13 5.12 ;
      RECT 23.095 4.835 23.12 5.123 ;
      RECT 23.075 4.852 23.095 5.127 ;
      RECT 23.035 4.88 23.075 5.133 ;
      RECT 22.97 4.927 23.035 5.142 ;
      RECT 22.955 4.96 22.97 5.15 ;
      RECT 22.95 4.967 22.955 5.152 ;
      RECT 22.9 4.992 22.95 5.157 ;
      RECT 22.885 5.016 22.9 5.164 ;
      RECT 22.835 5.021 22.885 5.165 ;
      RECT 22.749 5.025 22.835 5.165 ;
      RECT 22.663 5.025 22.749 5.165 ;
      RECT 22.577 5.025 22.663 5.166 ;
      RECT 22.491 5.025 22.577 5.166 ;
      RECT 22.405 5.025 22.491 5.166 ;
      RECT 22.339 5.025 22.405 5.166 ;
      RECT 22.253 5.025 22.339 5.167 ;
      RECT 22.167 5.025 22.253 5.167 ;
      RECT 22.081 5.026 22.167 5.168 ;
      RECT 21.995 5.026 22.081 5.168 ;
      RECT 21.909 5.026 21.995 5.168 ;
      RECT 21.823 5.026 21.909 5.169 ;
      RECT 21.737 5.026 21.823 5.169 ;
      RECT 21.651 5.027 21.737 5.17 ;
      RECT 21.565 5.027 21.651 5.17 ;
      RECT 21.545 5.027 21.565 5.17 ;
      RECT 21.459 5.027 21.545 5.17 ;
      RECT 21.373 5.027 21.459 5.17 ;
      RECT 21.287 5.028 21.373 5.17 ;
      RECT 21.201 5.028 21.287 5.17 ;
      RECT 21.115 5.028 21.201 5.17 ;
      RECT 21.029 5.029 21.115 5.17 ;
      RECT 20.943 5.029 21.029 5.17 ;
      RECT 20.857 5.029 20.943 5.17 ;
      RECT 20.771 5.029 20.857 5.17 ;
      RECT 20.685 5.03 20.771 5.17 ;
      RECT 20.635 5.027 20.685 5.17 ;
      RECT 20.625 5.025 20.635 5.169 ;
      RECT 20.621 5.025 20.625 5.168 ;
      RECT 20.535 5.02 20.621 5.163 ;
      RECT 20.513 5.013 20.535 5.157 ;
      RECT 20.427 5.004 20.513 5.151 ;
      RECT 20.341 4.991 20.427 5.142 ;
      RECT 20.255 4.977 20.341 5.132 ;
      RECT 20.21 4.967 20.255 5.125 ;
      RECT 20.19 4.255 20.21 4.533 ;
      RECT 20.19 4.96 20.21 5.121 ;
      RECT 20.16 4.255 20.19 4.555 ;
      RECT 20.15 4.927 20.19 5.118 ;
      RECT 20.145 4.255 20.16 4.575 ;
      RECT 20.145 4.892 20.15 5.116 ;
      RECT 20.14 4.255 20.145 4.7 ;
      RECT 20.14 4.852 20.145 5.116 ;
      RECT 20.13 4.255 20.14 5.116 ;
      RECT 20.055 4.255 20.13 5.11 ;
      RECT 20.025 4.255 20.055 5.1 ;
      RECT 20.02 4.255 20.025 5.092 ;
      RECT 20.015 4.297 20.02 5.085 ;
      RECT 20.005 4.366 20.015 5.076 ;
      RECT 20 4.436 20.005 5.028 ;
      RECT 19.995 4.5 20 4.925 ;
      RECT 19.99 4.535 19.995 4.88 ;
      RECT 19.988 4.572 19.99 4.772 ;
      RECT 19.985 4.58 19.988 4.765 ;
      RECT 19.98 4.645 19.985 4.708 ;
      RECT 24.055 3.735 24.335 4.015 ;
      RECT 24.045 3.735 24.335 3.878 ;
      RECT 24 3.6 24.26 3.86 ;
      RECT 24 3.715 24.315 3.86 ;
      RECT 24 3.685 24.31 3.86 ;
      RECT 24 3.672 24.3 3.86 ;
      RECT 24 3.662 24.295 3.86 ;
      RECT 19.975 3.645 20.235 3.905 ;
      RECT 23.745 3.195 24.005 3.455 ;
      RECT 23.735 3.22 24.005 3.415 ;
      RECT 23.73 3.22 23.735 3.414 ;
      RECT 23.66 3.215 23.73 3.406 ;
      RECT 23.575 3.202 23.66 3.389 ;
      RECT 23.571 3.194 23.575 3.379 ;
      RECT 23.485 3.187 23.571 3.369 ;
      RECT 23.476 3.179 23.485 3.359 ;
      RECT 23.39 3.172 23.476 3.347 ;
      RECT 23.37 3.163 23.39 3.333 ;
      RECT 23.315 3.158 23.37 3.325 ;
      RECT 23.305 3.152 23.315 3.319 ;
      RECT 23.285 3.15 23.305 3.315 ;
      RECT 23.277 3.149 23.285 3.311 ;
      RECT 23.191 3.141 23.277 3.3 ;
      RECT 23.105 3.127 23.191 3.28 ;
      RECT 23.045 3.115 23.105 3.265 ;
      RECT 23.035 3.11 23.045 3.26 ;
      RECT 22.985 3.11 23.035 3.262 ;
      RECT 22.938 3.112 22.985 3.266 ;
      RECT 22.852 3.119 22.938 3.271 ;
      RECT 22.766 3.127 22.852 3.277 ;
      RECT 22.68 3.136 22.766 3.283 ;
      RECT 22.621 3.142 22.68 3.288 ;
      RECT 22.535 3.147 22.621 3.294 ;
      RECT 22.46 3.152 22.535 3.3 ;
      RECT 22.421 3.154 22.46 3.305 ;
      RECT 22.335 3.151 22.421 3.31 ;
      RECT 22.25 3.149 22.335 3.317 ;
      RECT 22.218 3.148 22.25 3.32 ;
      RECT 22.132 3.147 22.218 3.321 ;
      RECT 22.046 3.146 22.132 3.322 ;
      RECT 21.96 3.145 22.046 3.322 ;
      RECT 21.874 3.144 21.96 3.323 ;
      RECT 21.788 3.143 21.874 3.324 ;
      RECT 21.702 3.142 21.788 3.325 ;
      RECT 21.616 3.141 21.702 3.325 ;
      RECT 21.53 3.14 21.616 3.326 ;
      RECT 21.48 3.14 21.53 3.327 ;
      RECT 21.466 3.141 21.48 3.327 ;
      RECT 21.38 3.148 21.466 3.328 ;
      RECT 21.306 3.159 21.38 3.329 ;
      RECT 21.22 3.168 21.306 3.33 ;
      RECT 21.185 3.175 21.22 3.345 ;
      RECT 21.16 3.178 21.185 3.375 ;
      RECT 21.135 3.187 21.16 3.404 ;
      RECT 21.125 3.198 21.135 3.424 ;
      RECT 21.115 3.206 21.125 3.438 ;
      RECT 21.11 3.212 21.115 3.448 ;
      RECT 21.085 3.229 21.11 3.465 ;
      RECT 21.07 3.251 21.085 3.493 ;
      RECT 21.04 3.277 21.07 3.523 ;
      RECT 21.02 3.306 21.04 3.553 ;
      RECT 21.015 3.321 21.02 3.57 ;
      RECT 20.995 3.336 21.015 3.585 ;
      RECT 20.985 3.354 20.995 3.603 ;
      RECT 20.975 3.365 20.985 3.618 ;
      RECT 20.925 3.397 20.975 3.644 ;
      RECT 20.92 3.427 20.925 3.664 ;
      RECT 20.91 3.44 20.92 3.67 ;
      RECT 20.901 3.45 20.91 3.678 ;
      RECT 20.89 3.461 20.901 3.686 ;
      RECT 20.885 3.471 20.89 3.692 ;
      RECT 20.87 3.492 20.885 3.699 ;
      RECT 20.855 3.522 20.87 3.707 ;
      RECT 20.82 3.552 20.855 3.713 ;
      RECT 20.795 3.57 20.82 3.72 ;
      RECT 20.745 3.578 20.795 3.729 ;
      RECT 20.72 3.583 20.745 3.738 ;
      RECT 20.665 3.589 20.72 3.748 ;
      RECT 20.66 3.594 20.665 3.756 ;
      RECT 20.646 3.597 20.66 3.758 ;
      RECT 20.56 3.609 20.646 3.77 ;
      RECT 20.55 3.621 20.56 3.783 ;
      RECT 20.465 3.634 20.55 3.795 ;
      RECT 20.421 3.651 20.465 3.809 ;
      RECT 20.335 3.668 20.421 3.825 ;
      RECT 20.305 3.682 20.335 3.839 ;
      RECT 20.295 3.687 20.305 3.844 ;
      RECT 20.235 3.69 20.295 3.853 ;
      RECT 23.125 3.96 23.385 4.22 ;
      RECT 23.125 3.96 23.405 4.073 ;
      RECT 23.125 3.96 23.43 4.04 ;
      RECT 23.125 3.96 23.435 4.02 ;
      RECT 23.175 3.735 23.455 4.015 ;
      RECT 22.73 4.47 22.99 4.73 ;
      RECT 22.72 4.327 22.915 4.668 ;
      RECT 22.715 4.435 22.93 4.66 ;
      RECT 22.71 4.485 22.99 4.65 ;
      RECT 22.7 4.562 22.99 4.635 ;
      RECT 22.72 4.41 22.93 4.668 ;
      RECT 22.73 4.285 22.915 4.73 ;
      RECT 22.73 4.18 22.895 4.73 ;
      RECT 22.74 4.167 22.895 4.73 ;
      RECT 22.74 4.125 22.885 4.73 ;
      RECT 22.745 4.05 22.885 4.73 ;
      RECT 22.775 3.7 22.885 4.73 ;
      RECT 22.78 3.43 22.905 4.053 ;
      RECT 22.75 4.005 22.905 4.053 ;
      RECT 22.765 3.807 22.885 4.73 ;
      RECT 22.755 3.917 22.905 4.053 ;
      RECT 22.78 3.43 22.92 3.91 ;
      RECT 22.78 3.43 22.94 3.785 ;
      RECT 22.745 3.43 23.005 3.69 ;
      RECT 22.215 3.735 22.495 4.015 ;
      RECT 22.2 3.735 22.495 3.995 ;
      RECT 20.255 4.6 20.515 4.86 ;
      RECT 22.04 4.455 22.3 4.715 ;
      RECT 22.02 4.475 22.3 4.69 ;
      RECT 21.977 4.475 22.02 4.689 ;
      RECT 21.891 4.476 21.977 4.686 ;
      RECT 21.805 4.477 21.891 4.682 ;
      RECT 21.73 4.479 21.805 4.679 ;
      RECT 21.707 4.48 21.73 4.677 ;
      RECT 21.621 4.481 21.707 4.675 ;
      RECT 21.535 4.482 21.621 4.672 ;
      RECT 21.511 4.483 21.535 4.67 ;
      RECT 21.425 4.485 21.511 4.667 ;
      RECT 21.34 4.487 21.425 4.668 ;
      RECT 21.283 4.488 21.34 4.674 ;
      RECT 21.197 4.49 21.283 4.684 ;
      RECT 21.111 4.493 21.197 4.697 ;
      RECT 21.025 4.495 21.111 4.709 ;
      RECT 21.011 4.496 21.025 4.716 ;
      RECT 20.925 4.497 21.011 4.724 ;
      RECT 20.885 4.499 20.925 4.733 ;
      RECT 20.876 4.5 20.885 4.736 ;
      RECT 20.79 4.508 20.876 4.742 ;
      RECT 20.77 4.517 20.79 4.75 ;
      RECT 20.685 4.532 20.77 4.758 ;
      RECT 20.625 4.555 20.685 4.769 ;
      RECT 20.615 4.567 20.625 4.774 ;
      RECT 20.575 4.577 20.615 4.778 ;
      RECT 20.52 4.594 20.575 4.786 ;
      RECT 20.515 4.604 20.52 4.79 ;
      RECT 21.581 3.735 21.64 4.132 ;
      RECT 21.495 3.735 21.7 4.123 ;
      RECT 21.49 3.765 21.7 4.118 ;
      RECT 21.456 3.765 21.7 4.116 ;
      RECT 21.37 3.765 21.7 4.11 ;
      RECT 21.325 3.765 21.72 4.088 ;
      RECT 21.325 3.765 21.74 4.043 ;
      RECT 21.285 3.765 21.74 4.033 ;
      RECT 21.495 3.735 21.775 4.015 ;
      RECT 21.23 3.735 21.49 3.995 ;
      RECT 19.055 4.295 19.335 4.575 ;
      RECT 19.025 4.257 19.28 4.56 ;
      RECT 19.02 4.258 19.28 4.558 ;
      RECT 19.015 4.259 19.28 4.552 ;
      RECT 19.01 4.262 19.28 4.545 ;
      RECT 19.005 4.295 19.335 4.538 ;
      RECT 18.975 4.265 19.28 4.525 ;
      RECT 18.975 4.292 19.3 4.525 ;
      RECT 18.975 4.282 19.295 4.525 ;
      RECT 18.975 4.267 19.29 4.525 ;
      RECT 19.055 4.254 19.27 4.575 ;
      RECT 19.141 4.252 19.27 4.575 ;
      RECT 19.227 4.25 19.255 4.575 ;
      RECT 14.865 8.505 15.185 8.83 ;
      RECT 14.895 7.98 15.065 8.83 ;
      RECT 14.895 7.98 15.07 8.33 ;
      RECT 14.895 7.98 15.87 8.155 ;
      RECT 15.695 3.26 15.87 8.155 ;
      RECT 15.64 3.26 15.99 3.61 ;
      RECT 15.665 8.94 15.99 9.265 ;
      RECT 14.55 9.03 15.99 9.2 ;
      RECT 14.55 3.69 14.71 9.2 ;
      RECT 14.865 3.66 15.185 3.98 ;
      RECT 14.55 3.69 15.185 3.86 ;
      RECT 4.635 3.215 4.895 3.475 ;
      RECT 4.69 3.175 4.995 3.455 ;
      RECT 4.69 2.715 4.865 3.475 ;
      RECT 13.205 2.635 13.555 2.985 ;
      RECT 4.69 2.715 13.555 2.89 ;
      RECT 12.88 4.145 13.25 4.515 ;
      RECT 12.965 3.53 13.135 4.515 ;
      RECT 8.985 3.75 9.22 4.01 ;
      RECT 12.13 3.53 12.295 3.79 ;
      RECT 12.035 3.52 12.05 3.79 ;
      RECT 12.13 3.53 13.135 3.71 ;
      RECT 10.635 3.09 10.675 3.23 ;
      RECT 12.05 3.525 12.13 3.79 ;
      RECT 11.995 3.52 12.035 3.756 ;
      RECT 11.981 3.52 11.995 3.756 ;
      RECT 11.895 3.525 11.981 3.758 ;
      RECT 11.85 3.532 11.895 3.76 ;
      RECT 11.82 3.532 11.85 3.762 ;
      RECT 11.795 3.527 11.82 3.764 ;
      RECT 11.765 3.523 11.795 3.773 ;
      RECT 11.755 3.52 11.765 3.785 ;
      RECT 11.75 3.52 11.755 3.793 ;
      RECT 11.745 3.52 11.75 3.798 ;
      RECT 11.735 3.519 11.745 3.808 ;
      RECT 11.73 3.518 11.735 3.818 ;
      RECT 11.715 3.517 11.73 3.823 ;
      RECT 11.687 3.514 11.715 3.85 ;
      RECT 11.601 3.506 11.687 3.85 ;
      RECT 11.515 3.495 11.601 3.85 ;
      RECT 11.475 3.48 11.515 3.85 ;
      RECT 11.435 3.454 11.475 3.85 ;
      RECT 11.43 3.436 11.435 3.662 ;
      RECT 11.42 3.432 11.43 3.652 ;
      RECT 11.405 3.422 11.42 3.639 ;
      RECT 11.385 3.406 11.405 3.624 ;
      RECT 11.37 3.391 11.385 3.609 ;
      RECT 11.36 3.38 11.37 3.599 ;
      RECT 11.335 3.364 11.36 3.588 ;
      RECT 11.33 3.351 11.335 3.578 ;
      RECT 11.325 3.347 11.33 3.573 ;
      RECT 11.27 3.333 11.325 3.551 ;
      RECT 11.231 3.314 11.27 3.515 ;
      RECT 11.145 3.288 11.231 3.468 ;
      RECT 11.141 3.27 11.145 3.434 ;
      RECT 11.055 3.251 11.141 3.412 ;
      RECT 11.05 3.233 11.055 3.39 ;
      RECT 11.045 3.231 11.05 3.388 ;
      RECT 11.035 3.23 11.045 3.383 ;
      RECT 10.975 3.217 11.035 3.369 ;
      RECT 10.93 3.195 10.975 3.348 ;
      RECT 10.87 3.172 10.93 3.327 ;
      RECT 10.806 3.147 10.87 3.302 ;
      RECT 10.72 3.117 10.806 3.271 ;
      RECT 10.705 3.097 10.72 3.25 ;
      RECT 10.675 3.092 10.705 3.241 ;
      RECT 10.622 3.09 10.635 3.23 ;
      RECT 10.536 3.09 10.622 3.232 ;
      RECT 10.45 3.09 10.536 3.234 ;
      RECT 10.43 3.09 10.45 3.238 ;
      RECT 10.385 3.092 10.43 3.249 ;
      RECT 10.345 3.102 10.385 3.265 ;
      RECT 10.341 3.111 10.345 3.273 ;
      RECT 10.255 3.131 10.341 3.289 ;
      RECT 10.245 3.15 10.255 3.307 ;
      RECT 10.24 3.152 10.245 3.31 ;
      RECT 10.23 3.156 10.24 3.313 ;
      RECT 10.21 3.161 10.23 3.323 ;
      RECT 10.18 3.171 10.21 3.343 ;
      RECT 10.175 3.178 10.18 3.357 ;
      RECT 10.165 3.182 10.175 3.364 ;
      RECT 10.15 3.19 10.165 3.375 ;
      RECT 10.14 3.2 10.15 3.386 ;
      RECT 10.13 3.207 10.14 3.394 ;
      RECT 10.105 3.22 10.13 3.409 ;
      RECT 10.041 3.256 10.105 3.448 ;
      RECT 9.955 3.319 10.041 3.512 ;
      RECT 9.92 3.37 9.955 3.565 ;
      RECT 9.915 3.387 9.92 3.582 ;
      RECT 9.9 3.396 9.915 3.589 ;
      RECT 9.88 3.411 9.9 3.603 ;
      RECT 9.875 3.422 9.88 3.613 ;
      RECT 9.855 3.435 9.875 3.623 ;
      RECT 9.85 3.445 9.855 3.633 ;
      RECT 9.835 3.45 9.85 3.642 ;
      RECT 9.825 3.46 9.835 3.653 ;
      RECT 9.795 3.477 9.825 3.67 ;
      RECT 9.785 3.495 9.795 3.688 ;
      RECT 9.77 3.506 9.785 3.699 ;
      RECT 9.73 3.53 9.77 3.715 ;
      RECT 9.695 3.564 9.73 3.732 ;
      RECT 9.665 3.587 9.695 3.744 ;
      RECT 9.65 3.597 9.665 3.753 ;
      RECT 9.61 3.607 9.65 3.764 ;
      RECT 9.59 3.618 9.61 3.776 ;
      RECT 9.585 3.622 9.59 3.783 ;
      RECT 9.57 3.626 9.585 3.788 ;
      RECT 9.56 3.631 9.57 3.793 ;
      RECT 9.555 3.634 9.56 3.796 ;
      RECT 9.525 3.64 9.555 3.803 ;
      RECT 9.49 3.65 9.525 3.817 ;
      RECT 9.43 3.665 9.49 3.837 ;
      RECT 9.375 3.685 9.43 3.861 ;
      RECT 9.346 3.7 9.375 3.879 ;
      RECT 9.26 3.72 9.346 3.904 ;
      RECT 9.255 3.735 9.26 3.924 ;
      RECT 9.245 3.738 9.255 3.925 ;
      RECT 9.22 3.745 9.245 4.01 ;
      RECT 11.915 4.238 12.195 4.575 ;
      RECT 11.915 4.248 12.2 4.533 ;
      RECT 11.915 4.257 12.205 4.43 ;
      RECT 11.915 4.272 12.21 4.298 ;
      RECT 11.915 4.1 12.175 4.575 ;
      RECT 1.54 9.28 1.83 9.63 ;
      RECT 1.54 9.37 2.945 9.54 ;
      RECT 2.775 8.97 2.945 9.54 ;
      RECT 11.06 8.89 11.41 9.24 ;
      RECT 2.775 8.97 11.41 9.14 ;
      RECT 9.635 4.98 9.645 5.17 ;
      RECT 7.895 4.855 8.175 5.135 ;
      RECT 10.94 3.795 10.945 4.28 ;
      RECT 10.835 3.795 10.895 4.055 ;
      RECT 11.16 4.765 11.165 4.84 ;
      RECT 11.15 4.632 11.16 4.875 ;
      RECT 11.14 4.467 11.15 4.896 ;
      RECT 11.135 4.337 11.14 4.912 ;
      RECT 11.125 4.227 11.135 4.928 ;
      RECT 11.12 4.126 11.125 4.945 ;
      RECT 11.115 4.108 11.12 4.955 ;
      RECT 11.11 4.09 11.115 4.965 ;
      RECT 11.1 4.065 11.11 4.98 ;
      RECT 11.095 4.045 11.1 4.995 ;
      RECT 11.075 3.795 11.095 5.02 ;
      RECT 11.06 3.795 11.075 5.053 ;
      RECT 11.03 3.795 11.06 5.075 ;
      RECT 11.01 3.795 11.03 5.089 ;
      RECT 10.99 3.795 11.01 4.605 ;
      RECT 11.005 4.672 11.01 5.094 ;
      RECT 11 4.702 11.005 5.096 ;
      RECT 10.995 4.715 11 5.099 ;
      RECT 10.99 4.725 10.995 5.103 ;
      RECT 10.985 3.795 10.99 4.523 ;
      RECT 10.985 4.735 10.99 5.105 ;
      RECT 10.98 3.795 10.985 4.5 ;
      RECT 10.97 4.757 10.985 5.105 ;
      RECT 10.965 3.795 10.98 4.445 ;
      RECT 10.96 4.782 10.97 5.105 ;
      RECT 10.96 3.795 10.965 4.39 ;
      RECT 10.95 3.795 10.96 4.338 ;
      RECT 10.955 4.795 10.96 5.106 ;
      RECT 10.95 4.807 10.955 5.107 ;
      RECT 10.945 3.795 10.95 4.298 ;
      RECT 10.945 4.82 10.95 5.108 ;
      RECT 10.93 4.835 10.945 5.109 ;
      RECT 10.935 3.795 10.94 4.26 ;
      RECT 10.93 3.795 10.935 4.225 ;
      RECT 10.925 3.795 10.93 4.2 ;
      RECT 10.92 4.862 10.93 5.111 ;
      RECT 10.915 3.795 10.925 4.158 ;
      RECT 10.915 4.88 10.92 5.112 ;
      RECT 10.91 3.795 10.915 4.118 ;
      RECT 10.91 4.887 10.915 5.113 ;
      RECT 10.905 3.795 10.91 4.09 ;
      RECT 10.9 4.905 10.91 5.114 ;
      RECT 10.895 3.795 10.905 4.07 ;
      RECT 10.89 4.925 10.9 5.116 ;
      RECT 10.88 4.942 10.89 5.117 ;
      RECT 10.845 4.965 10.88 5.12 ;
      RECT 10.79 4.983 10.845 5.126 ;
      RECT 10.704 4.991 10.79 5.135 ;
      RECT 10.618 5.002 10.704 5.146 ;
      RECT 10.532 5.012 10.618 5.157 ;
      RECT 10.446 5.022 10.532 5.169 ;
      RECT 10.36 5.032 10.446 5.18 ;
      RECT 10.34 5.038 10.36 5.186 ;
      RECT 10.26 5.04 10.34 5.19 ;
      RECT 10.255 5.039 10.26 5.195 ;
      RECT 10.247 5.038 10.255 5.195 ;
      RECT 10.161 5.034 10.247 5.193 ;
      RECT 10.075 5.026 10.161 5.19 ;
      RECT 9.989 5.017 10.075 5.186 ;
      RECT 9.903 5.009 9.989 5.183 ;
      RECT 9.817 5.001 9.903 5.179 ;
      RECT 9.731 4.992 9.817 5.176 ;
      RECT 9.645 4.984 9.731 5.172 ;
      RECT 9.59 4.977 9.635 5.17 ;
      RECT 9.505 4.97 9.59 5.168 ;
      RECT 9.431 4.962 9.505 5.164 ;
      RECT 9.345 4.954 9.431 5.161 ;
      RECT 9.342 4.95 9.345 5.159 ;
      RECT 9.256 4.946 9.342 5.158 ;
      RECT 9.17 4.938 9.256 5.155 ;
      RECT 9.085 4.933 9.17 5.152 ;
      RECT 8.999 4.93 9.085 5.149 ;
      RECT 8.913 4.928 8.999 5.146 ;
      RECT 8.827 4.925 8.913 5.143 ;
      RECT 8.741 4.922 8.827 5.14 ;
      RECT 8.655 4.919 8.741 5.137 ;
      RECT 8.579 4.917 8.655 5.134 ;
      RECT 8.493 4.914 8.579 5.131 ;
      RECT 8.407 4.911 8.493 5.129 ;
      RECT 8.321 4.909 8.407 5.126 ;
      RECT 8.235 4.906 8.321 5.123 ;
      RECT 8.175 4.897 8.235 5.121 ;
      RECT 10.685 4.515 10.76 4.775 ;
      RECT 10.665 4.495 10.67 4.775 ;
      RECT 9.985 4.28 10.09 4.575 ;
      RECT 4.43 4.255 4.5 4.515 ;
      RECT 10.325 4.13 10.33 4.501 ;
      RECT 10.315 4.185 10.32 4.501 ;
      RECT 10.62 3.355 10.68 3.615 ;
      RECT 10.675 4.51 10.685 4.775 ;
      RECT 10.67 4.5 10.675 4.775 ;
      RECT 10.59 4.447 10.665 4.775 ;
      RECT 10.615 3.355 10.62 3.635 ;
      RECT 10.605 3.355 10.615 3.655 ;
      RECT 10.59 3.355 10.605 3.685 ;
      RECT 10.575 3.355 10.59 3.728 ;
      RECT 10.57 4.39 10.59 4.775 ;
      RECT 10.56 3.355 10.575 3.765 ;
      RECT 10.555 4.37 10.57 4.775 ;
      RECT 10.555 3.355 10.56 3.788 ;
      RECT 10.545 3.355 10.555 3.813 ;
      RECT 10.515 4.337 10.555 4.775 ;
      RECT 10.52 3.355 10.545 3.863 ;
      RECT 10.515 3.355 10.52 3.918 ;
      RECT 10.51 3.355 10.515 3.96 ;
      RECT 10.5 4.3 10.515 4.775 ;
      RECT 10.505 3.355 10.51 4.003 ;
      RECT 10.5 3.355 10.505 4.068 ;
      RECT 10.495 3.355 10.5 4.09 ;
      RECT 10.495 4.288 10.5 4.64 ;
      RECT 10.49 3.355 10.495 4.158 ;
      RECT 10.49 4.28 10.495 4.623 ;
      RECT 10.485 3.355 10.49 4.203 ;
      RECT 10.48 4.262 10.49 4.6 ;
      RECT 10.48 3.355 10.485 4.24 ;
      RECT 10.47 3.355 10.48 4.58 ;
      RECT 10.465 3.355 10.47 4.563 ;
      RECT 10.46 3.355 10.465 4.548 ;
      RECT 10.455 3.355 10.46 4.533 ;
      RECT 10.435 3.355 10.455 4.523 ;
      RECT 10.43 3.355 10.435 4.513 ;
      RECT 10.42 3.355 10.43 4.509 ;
      RECT 10.415 3.632 10.42 4.508 ;
      RECT 10.41 3.655 10.415 4.507 ;
      RECT 10.405 3.685 10.41 4.506 ;
      RECT 10.4 3.712 10.405 4.505 ;
      RECT 10.395 3.74 10.4 4.505 ;
      RECT 10.39 3.767 10.395 4.505 ;
      RECT 10.385 3.787 10.39 4.505 ;
      RECT 10.38 3.815 10.385 4.505 ;
      RECT 10.37 3.857 10.38 4.505 ;
      RECT 10.36 3.902 10.37 4.504 ;
      RECT 10.355 3.955 10.36 4.503 ;
      RECT 10.35 3.987 10.355 4.502 ;
      RECT 10.345 4.007 10.35 4.501 ;
      RECT 10.34 4.045 10.345 4.501 ;
      RECT 10.335 4.067 10.34 4.501 ;
      RECT 10.33 4.092 10.335 4.501 ;
      RECT 10.32 4.157 10.325 4.501 ;
      RECT 10.305 4.217 10.315 4.501 ;
      RECT 10.29 4.227 10.305 4.501 ;
      RECT 10.27 4.237 10.29 4.501 ;
      RECT 10.24 4.242 10.27 4.498 ;
      RECT 10.18 4.252 10.24 4.495 ;
      RECT 10.16 4.261 10.18 4.5 ;
      RECT 10.135 4.267 10.16 4.513 ;
      RECT 10.115 4.272 10.135 4.528 ;
      RECT 10.09 4.277 10.115 4.575 ;
      RECT 9.961 4.279 9.985 4.575 ;
      RECT 9.875 4.274 9.961 4.575 ;
      RECT 9.835 4.271 9.875 4.575 ;
      RECT 9.785 4.273 9.835 4.555 ;
      RECT 9.755 4.277 9.785 4.555 ;
      RECT 9.676 4.287 9.755 4.555 ;
      RECT 9.59 4.302 9.676 4.556 ;
      RECT 9.54 4.312 9.59 4.557 ;
      RECT 9.532 4.315 9.54 4.557 ;
      RECT 9.446 4.317 9.532 4.558 ;
      RECT 9.36 4.321 9.446 4.558 ;
      RECT 9.274 4.325 9.36 4.559 ;
      RECT 9.188 4.328 9.274 4.56 ;
      RECT 9.102 4.332 9.188 4.56 ;
      RECT 9.016 4.336 9.102 4.561 ;
      RECT 8.93 4.339 9.016 4.562 ;
      RECT 8.844 4.343 8.93 4.562 ;
      RECT 8.758 4.347 8.844 4.563 ;
      RECT 8.672 4.351 8.758 4.564 ;
      RECT 8.586 4.354 8.672 4.564 ;
      RECT 8.5 4.358 8.586 4.565 ;
      RECT 8.47 4.36 8.5 4.565 ;
      RECT 8.384 4.363 8.47 4.566 ;
      RECT 8.298 4.367 8.384 4.567 ;
      RECT 8.212 4.371 8.298 4.568 ;
      RECT 8.126 4.374 8.212 4.568 ;
      RECT 8.04 4.378 8.126 4.569 ;
      RECT 8.005 4.383 8.04 4.57 ;
      RECT 7.95 4.393 8.005 4.577 ;
      RECT 7.925 4.405 7.95 4.587 ;
      RECT 7.89 4.418 7.925 4.595 ;
      RECT 7.85 4.435 7.89 4.618 ;
      RECT 7.83 4.448 7.85 4.645 ;
      RECT 7.8 4.46 7.83 4.673 ;
      RECT 7.795 4.468 7.8 4.693 ;
      RECT 7.79 4.471 7.795 4.703 ;
      RECT 7.74 4.483 7.79 4.737 ;
      RECT 7.73 4.498 7.74 4.77 ;
      RECT 7.72 4.504 7.73 4.783 ;
      RECT 7.71 4.511 7.72 4.795 ;
      RECT 7.685 4.524 7.71 4.813 ;
      RECT 7.67 4.539 7.685 4.835 ;
      RECT 7.66 4.547 7.67 4.851 ;
      RECT 7.645 4.556 7.66 4.866 ;
      RECT 7.635 4.566 7.645 4.88 ;
      RECT 7.616 4.579 7.635 4.897 ;
      RECT 7.53 4.624 7.616 4.962 ;
      RECT 7.515 4.669 7.53 5.02 ;
      RECT 7.51 4.678 7.515 5.033 ;
      RECT 7.5 4.685 7.51 5.038 ;
      RECT 7.495 4.69 7.5 5.042 ;
      RECT 7.475 4.7 7.495 5.049 ;
      RECT 7.45 4.72 7.475 5.063 ;
      RECT 7.415 4.745 7.45 5.083 ;
      RECT 7.4 4.768 7.415 5.098 ;
      RECT 7.39 4.778 7.4 5.103 ;
      RECT 7.38 4.786 7.39 5.11 ;
      RECT 7.37 4.795 7.38 5.116 ;
      RECT 7.35 4.807 7.37 5.118 ;
      RECT 7.34 4.82 7.35 5.12 ;
      RECT 7.315 4.835 7.34 5.123 ;
      RECT 7.295 4.852 7.315 5.127 ;
      RECT 7.255 4.88 7.295 5.133 ;
      RECT 7.19 4.927 7.255 5.142 ;
      RECT 7.175 4.96 7.19 5.15 ;
      RECT 7.17 4.967 7.175 5.152 ;
      RECT 7.12 4.992 7.17 5.157 ;
      RECT 7.105 5.016 7.12 5.164 ;
      RECT 7.055 5.021 7.105 5.165 ;
      RECT 6.969 5.025 7.055 5.165 ;
      RECT 6.883 5.025 6.969 5.165 ;
      RECT 6.797 5.025 6.883 5.166 ;
      RECT 6.711 5.025 6.797 5.166 ;
      RECT 6.625 5.025 6.711 5.166 ;
      RECT 6.559 5.025 6.625 5.166 ;
      RECT 6.473 5.025 6.559 5.167 ;
      RECT 6.387 5.025 6.473 5.167 ;
      RECT 6.301 5.026 6.387 5.168 ;
      RECT 6.215 5.026 6.301 5.168 ;
      RECT 6.129 5.026 6.215 5.168 ;
      RECT 6.043 5.026 6.129 5.169 ;
      RECT 5.957 5.026 6.043 5.169 ;
      RECT 5.871 5.027 5.957 5.17 ;
      RECT 5.785 5.027 5.871 5.17 ;
      RECT 5.765 5.027 5.785 5.17 ;
      RECT 5.679 5.027 5.765 5.17 ;
      RECT 5.593 5.027 5.679 5.17 ;
      RECT 5.507 5.028 5.593 5.17 ;
      RECT 5.421 5.028 5.507 5.17 ;
      RECT 5.335 5.028 5.421 5.17 ;
      RECT 5.249 5.029 5.335 5.17 ;
      RECT 5.163 5.029 5.249 5.17 ;
      RECT 5.077 5.029 5.163 5.17 ;
      RECT 4.991 5.029 5.077 5.17 ;
      RECT 4.905 5.03 4.991 5.17 ;
      RECT 4.855 5.027 4.905 5.17 ;
      RECT 4.845 5.025 4.855 5.169 ;
      RECT 4.841 5.025 4.845 5.168 ;
      RECT 4.755 5.02 4.841 5.163 ;
      RECT 4.733 5.013 4.755 5.157 ;
      RECT 4.647 5.004 4.733 5.151 ;
      RECT 4.561 4.991 4.647 5.142 ;
      RECT 4.475 4.977 4.561 5.132 ;
      RECT 4.43 4.967 4.475 5.125 ;
      RECT 4.41 4.255 4.43 4.533 ;
      RECT 4.41 4.96 4.43 5.121 ;
      RECT 4.38 4.255 4.41 4.555 ;
      RECT 4.37 4.927 4.41 5.118 ;
      RECT 4.365 4.255 4.38 4.575 ;
      RECT 4.365 4.892 4.37 5.116 ;
      RECT 4.36 4.255 4.365 4.7 ;
      RECT 4.36 4.852 4.365 5.116 ;
      RECT 4.35 4.255 4.36 5.116 ;
      RECT 4.275 4.255 4.35 5.11 ;
      RECT 4.245 4.255 4.275 5.1 ;
      RECT 4.24 4.255 4.245 5.092 ;
      RECT 4.235 4.297 4.24 5.085 ;
      RECT 4.225 4.366 4.235 5.076 ;
      RECT 4.22 4.436 4.225 5.028 ;
      RECT 4.215 4.5 4.22 4.925 ;
      RECT 4.21 4.535 4.215 4.88 ;
      RECT 4.208 4.572 4.21 4.772 ;
      RECT 4.205 4.58 4.208 4.765 ;
      RECT 4.2 4.645 4.205 4.708 ;
      RECT 8.275 3.735 8.555 4.015 ;
      RECT 8.265 3.735 8.555 3.878 ;
      RECT 8.22 3.6 8.48 3.86 ;
      RECT 8.22 3.715 8.535 3.86 ;
      RECT 8.22 3.685 8.53 3.86 ;
      RECT 8.22 3.672 8.52 3.86 ;
      RECT 8.22 3.662 8.515 3.86 ;
      RECT 4.195 3.645 4.455 3.905 ;
      RECT 7.965 3.195 8.225 3.455 ;
      RECT 7.955 3.22 8.225 3.415 ;
      RECT 7.95 3.22 7.955 3.414 ;
      RECT 7.88 3.215 7.95 3.406 ;
      RECT 7.795 3.202 7.88 3.389 ;
      RECT 7.791 3.194 7.795 3.379 ;
      RECT 7.705 3.187 7.791 3.369 ;
      RECT 7.696 3.179 7.705 3.359 ;
      RECT 7.61 3.172 7.696 3.347 ;
      RECT 7.59 3.163 7.61 3.333 ;
      RECT 7.535 3.158 7.59 3.325 ;
      RECT 7.525 3.152 7.535 3.319 ;
      RECT 7.505 3.15 7.525 3.315 ;
      RECT 7.497 3.149 7.505 3.311 ;
      RECT 7.411 3.141 7.497 3.3 ;
      RECT 7.325 3.127 7.411 3.28 ;
      RECT 7.265 3.115 7.325 3.265 ;
      RECT 7.255 3.11 7.265 3.26 ;
      RECT 7.205 3.11 7.255 3.262 ;
      RECT 7.158 3.112 7.205 3.266 ;
      RECT 7.072 3.119 7.158 3.271 ;
      RECT 6.986 3.127 7.072 3.277 ;
      RECT 6.9 3.136 6.986 3.283 ;
      RECT 6.841 3.142 6.9 3.288 ;
      RECT 6.755 3.147 6.841 3.294 ;
      RECT 6.68 3.152 6.755 3.3 ;
      RECT 6.641 3.154 6.68 3.305 ;
      RECT 6.555 3.151 6.641 3.31 ;
      RECT 6.47 3.149 6.555 3.317 ;
      RECT 6.438 3.148 6.47 3.32 ;
      RECT 6.352 3.147 6.438 3.321 ;
      RECT 6.266 3.146 6.352 3.322 ;
      RECT 6.18 3.145 6.266 3.322 ;
      RECT 6.094 3.144 6.18 3.323 ;
      RECT 6.008 3.143 6.094 3.324 ;
      RECT 5.922 3.142 6.008 3.325 ;
      RECT 5.836 3.141 5.922 3.325 ;
      RECT 5.75 3.14 5.836 3.326 ;
      RECT 5.7 3.14 5.75 3.327 ;
      RECT 5.686 3.141 5.7 3.327 ;
      RECT 5.6 3.148 5.686 3.328 ;
      RECT 5.526 3.159 5.6 3.329 ;
      RECT 5.44 3.168 5.526 3.33 ;
      RECT 5.405 3.175 5.44 3.345 ;
      RECT 5.38 3.178 5.405 3.375 ;
      RECT 5.355 3.187 5.38 3.404 ;
      RECT 5.345 3.198 5.355 3.424 ;
      RECT 5.335 3.206 5.345 3.438 ;
      RECT 5.33 3.212 5.335 3.448 ;
      RECT 5.305 3.229 5.33 3.465 ;
      RECT 5.29 3.251 5.305 3.493 ;
      RECT 5.26 3.277 5.29 3.523 ;
      RECT 5.24 3.306 5.26 3.553 ;
      RECT 5.235 3.321 5.24 3.57 ;
      RECT 5.215 3.336 5.235 3.585 ;
      RECT 5.205 3.354 5.215 3.603 ;
      RECT 5.195 3.365 5.205 3.618 ;
      RECT 5.145 3.397 5.195 3.644 ;
      RECT 5.14 3.427 5.145 3.664 ;
      RECT 5.13 3.44 5.14 3.67 ;
      RECT 5.121 3.45 5.13 3.678 ;
      RECT 5.11 3.461 5.121 3.686 ;
      RECT 5.105 3.471 5.11 3.692 ;
      RECT 5.09 3.492 5.105 3.699 ;
      RECT 5.075 3.522 5.09 3.707 ;
      RECT 5.04 3.552 5.075 3.713 ;
      RECT 5.015 3.57 5.04 3.72 ;
      RECT 4.965 3.578 5.015 3.729 ;
      RECT 4.94 3.583 4.965 3.738 ;
      RECT 4.885 3.589 4.94 3.748 ;
      RECT 4.88 3.594 4.885 3.756 ;
      RECT 4.866 3.597 4.88 3.758 ;
      RECT 4.78 3.609 4.866 3.77 ;
      RECT 4.77 3.621 4.78 3.783 ;
      RECT 4.685 3.634 4.77 3.795 ;
      RECT 4.641 3.651 4.685 3.809 ;
      RECT 4.555 3.668 4.641 3.825 ;
      RECT 4.525 3.682 4.555 3.839 ;
      RECT 4.515 3.687 4.525 3.844 ;
      RECT 4.455 3.69 4.515 3.853 ;
      RECT 7.345 3.96 7.605 4.22 ;
      RECT 7.345 3.96 7.625 4.073 ;
      RECT 7.345 3.96 7.65 4.04 ;
      RECT 7.345 3.96 7.655 4.02 ;
      RECT 7.395 3.735 7.675 4.015 ;
      RECT 6.95 4.47 7.21 4.73 ;
      RECT 6.94 4.327 7.135 4.668 ;
      RECT 6.935 4.435 7.15 4.66 ;
      RECT 6.93 4.485 7.21 4.65 ;
      RECT 6.92 4.562 7.21 4.635 ;
      RECT 6.94 4.41 7.15 4.668 ;
      RECT 6.95 4.285 7.135 4.73 ;
      RECT 6.95 4.18 7.115 4.73 ;
      RECT 6.96 4.167 7.115 4.73 ;
      RECT 6.96 4.125 7.105 4.73 ;
      RECT 6.965 4.05 7.105 4.73 ;
      RECT 6.995 3.7 7.105 4.73 ;
      RECT 7 3.43 7.125 4.053 ;
      RECT 6.97 4.005 7.125 4.053 ;
      RECT 6.985 3.807 7.105 4.73 ;
      RECT 6.975 3.917 7.125 4.053 ;
      RECT 7 3.43 7.14 3.91 ;
      RECT 7 3.43 7.16 3.785 ;
      RECT 6.965 3.43 7.225 3.69 ;
      RECT 6.435 3.735 6.715 4.015 ;
      RECT 6.42 3.735 6.715 3.995 ;
      RECT 4.475 4.6 4.735 4.86 ;
      RECT 6.26 4.455 6.52 4.715 ;
      RECT 6.24 4.475 6.52 4.69 ;
      RECT 6.197 4.475 6.24 4.689 ;
      RECT 6.111 4.476 6.197 4.686 ;
      RECT 6.025 4.477 6.111 4.682 ;
      RECT 5.95 4.479 6.025 4.679 ;
      RECT 5.927 4.48 5.95 4.677 ;
      RECT 5.841 4.481 5.927 4.675 ;
      RECT 5.755 4.482 5.841 4.672 ;
      RECT 5.731 4.483 5.755 4.67 ;
      RECT 5.645 4.485 5.731 4.667 ;
      RECT 5.56 4.487 5.645 4.668 ;
      RECT 5.503 4.488 5.56 4.674 ;
      RECT 5.417 4.49 5.503 4.684 ;
      RECT 5.331 4.493 5.417 4.697 ;
      RECT 5.245 4.495 5.331 4.709 ;
      RECT 5.231 4.496 5.245 4.716 ;
      RECT 5.145 4.497 5.231 4.724 ;
      RECT 5.105 4.499 5.145 4.733 ;
      RECT 5.096 4.5 5.105 4.736 ;
      RECT 5.01 4.508 5.096 4.742 ;
      RECT 4.99 4.517 5.01 4.75 ;
      RECT 4.905 4.532 4.99 4.758 ;
      RECT 4.845 4.555 4.905 4.769 ;
      RECT 4.835 4.567 4.845 4.774 ;
      RECT 4.795 4.577 4.835 4.778 ;
      RECT 4.74 4.594 4.795 4.786 ;
      RECT 4.735 4.604 4.74 4.79 ;
      RECT 5.801 3.735 5.86 4.132 ;
      RECT 5.715 3.735 5.92 4.123 ;
      RECT 5.71 3.765 5.92 4.118 ;
      RECT 5.676 3.765 5.92 4.116 ;
      RECT 5.59 3.765 5.92 4.11 ;
      RECT 5.545 3.765 5.94 4.088 ;
      RECT 5.545 3.765 5.96 4.043 ;
      RECT 5.505 3.765 5.96 4.033 ;
      RECT 5.715 3.735 5.995 4.015 ;
      RECT 5.45 3.735 5.71 3.995 ;
      RECT 3.275 4.295 3.555 4.575 ;
      RECT 3.245 4.257 3.5 4.56 ;
      RECT 3.24 4.258 3.5 4.558 ;
      RECT 3.235 4.259 3.5 4.552 ;
      RECT 3.23 4.262 3.5 4.545 ;
      RECT 3.225 4.295 3.555 4.538 ;
      RECT 3.195 4.265 3.5 4.525 ;
      RECT 3.195 4.292 3.52 4.525 ;
      RECT 3.195 4.282 3.515 4.525 ;
      RECT 3.195 4.267 3.51 4.525 ;
      RECT 3.275 4.254 3.49 4.575 ;
      RECT 3.361 4.252 3.49 4.575 ;
      RECT 3.447 4.25 3.475 4.575 ;
      RECT 75.225 2.11 75.595 2.48 ;
      RECT 73.515 9.325 73.885 9.695 ;
      RECT 59.44 2.11 59.81 2.48 ;
      RECT 57.73 9.325 58.1 9.695 ;
      RECT 43.655 2.11 44.025 2.48 ;
      RECT 41.945 9.325 42.315 9.695 ;
      RECT 27.88 2.11 28.25 2.48 ;
      RECT 26.17 9.325 26.54 9.695 ;
      RECT 12.1 2.11 12.47 2.48 ;
      RECT 10.39 9.325 10.76 9.695 ;
    LAYER via1 ;
      RECT 81.25 9.66 81.4 9.81 ;
      RECT 78.88 9.025 79.03 9.175 ;
      RECT 78.865 3.36 79.015 3.51 ;
      RECT 78.075 3.745 78.225 3.895 ;
      RECT 78.075 8.61 78.225 8.76 ;
      RECT 76.43 2.735 76.58 2.885 ;
      RECT 76.115 4.255 76.265 4.405 ;
      RECT 75.335 2.22 75.485 2.37 ;
      RECT 75.215 3.585 75.365 3.735 ;
      RECT 75.095 4.155 75.245 4.305 ;
      RECT 74.265 8.995 74.415 9.145 ;
      RECT 74.015 3.85 74.165 4 ;
      RECT 73.68 4.57 73.83 4.72 ;
      RECT 73.625 9.435 73.775 9.585 ;
      RECT 73.6 3.41 73.75 3.56 ;
      RECT 72.165 3.805 72.315 3.955 ;
      RECT 71.4 3.655 71.55 3.805 ;
      RECT 71.145 3.25 71.295 3.4 ;
      RECT 70.525 4.015 70.675 4.165 ;
      RECT 70.145 3.485 70.295 3.635 ;
      RECT 70.13 4.525 70.28 4.675 ;
      RECT 69.6 3.79 69.75 3.94 ;
      RECT 69.44 4.51 69.59 4.66 ;
      RECT 68.63 3.79 68.78 3.94 ;
      RECT 67.815 3.27 67.965 3.42 ;
      RECT 67.655 4.655 67.805 4.805 ;
      RECT 67.42 4.31 67.57 4.46 ;
      RECT 67.375 3.7 67.525 3.85 ;
      RECT 66.375 4.32 66.525 4.47 ;
      RECT 65.44 9.04 65.59 9.19 ;
      RECT 63.095 9.025 63.245 9.175 ;
      RECT 63.08 3.36 63.23 3.51 ;
      RECT 62.29 3.745 62.44 3.895 ;
      RECT 62.29 8.61 62.44 8.76 ;
      RECT 60.645 2.735 60.795 2.885 ;
      RECT 60.33 4.255 60.48 4.405 ;
      RECT 59.55 2.22 59.7 2.37 ;
      RECT 59.43 3.585 59.58 3.735 ;
      RECT 59.31 4.155 59.46 4.305 ;
      RECT 58.48 8.995 58.63 9.145 ;
      RECT 58.23 3.85 58.38 4 ;
      RECT 57.895 4.57 58.045 4.72 ;
      RECT 57.84 9.435 57.99 9.585 ;
      RECT 57.815 3.41 57.965 3.56 ;
      RECT 56.38 3.805 56.53 3.955 ;
      RECT 55.615 3.655 55.765 3.805 ;
      RECT 55.36 3.25 55.51 3.4 ;
      RECT 54.74 4.015 54.89 4.165 ;
      RECT 54.36 3.485 54.51 3.635 ;
      RECT 54.345 4.525 54.495 4.675 ;
      RECT 53.815 3.79 53.965 3.94 ;
      RECT 53.655 4.51 53.805 4.66 ;
      RECT 52.845 3.79 52.995 3.94 ;
      RECT 52.03 3.27 52.18 3.42 ;
      RECT 51.87 4.655 52.02 4.805 ;
      RECT 51.635 4.31 51.785 4.46 ;
      RECT 51.59 3.7 51.74 3.85 ;
      RECT 50.59 4.32 50.74 4.47 ;
      RECT 49.655 9.04 49.805 9.19 ;
      RECT 47.31 9.025 47.46 9.175 ;
      RECT 47.295 3.36 47.445 3.51 ;
      RECT 46.505 3.745 46.655 3.895 ;
      RECT 46.505 8.61 46.655 8.76 ;
      RECT 44.86 2.735 45.01 2.885 ;
      RECT 44.545 4.255 44.695 4.405 ;
      RECT 43.765 2.22 43.915 2.37 ;
      RECT 43.645 3.585 43.795 3.735 ;
      RECT 43.525 4.155 43.675 4.305 ;
      RECT 42.75 9 42.9 9.15 ;
      RECT 42.445 3.85 42.595 4 ;
      RECT 42.11 4.57 42.26 4.72 ;
      RECT 42.055 9.435 42.205 9.585 ;
      RECT 42.03 3.41 42.18 3.56 ;
      RECT 40.595 3.805 40.745 3.955 ;
      RECT 39.83 3.655 39.98 3.805 ;
      RECT 39.575 3.25 39.725 3.4 ;
      RECT 38.955 4.015 39.105 4.165 ;
      RECT 38.575 3.485 38.725 3.635 ;
      RECT 38.56 4.525 38.71 4.675 ;
      RECT 38.03 3.79 38.18 3.94 ;
      RECT 37.87 4.51 38.02 4.66 ;
      RECT 37.06 3.79 37.21 3.94 ;
      RECT 36.245 3.27 36.395 3.42 ;
      RECT 36.085 4.655 36.235 4.805 ;
      RECT 35.85 4.31 36 4.46 ;
      RECT 35.805 3.7 35.955 3.85 ;
      RECT 34.805 4.32 34.955 4.47 ;
      RECT 33.925 9.045 34.075 9.195 ;
      RECT 31.535 9.025 31.685 9.175 ;
      RECT 31.52 3.36 31.67 3.51 ;
      RECT 30.73 3.745 30.88 3.895 ;
      RECT 30.73 8.61 30.88 8.76 ;
      RECT 29.085 2.735 29.235 2.885 ;
      RECT 28.77 4.255 28.92 4.405 ;
      RECT 27.99 2.22 28.14 2.37 ;
      RECT 27.87 3.585 28.02 3.735 ;
      RECT 27.75 4.155 27.9 4.305 ;
      RECT 26.97 8.995 27.12 9.145 ;
      RECT 26.67 3.85 26.82 4 ;
      RECT 26.335 4.57 26.485 4.72 ;
      RECT 26.28 9.435 26.43 9.585 ;
      RECT 26.255 3.41 26.405 3.56 ;
      RECT 24.82 3.805 24.97 3.955 ;
      RECT 24.055 3.655 24.205 3.805 ;
      RECT 23.8 3.25 23.95 3.4 ;
      RECT 23.18 4.015 23.33 4.165 ;
      RECT 22.8 3.485 22.95 3.635 ;
      RECT 22.785 4.525 22.935 4.675 ;
      RECT 22.255 3.79 22.405 3.94 ;
      RECT 22.095 4.51 22.245 4.66 ;
      RECT 21.285 3.79 21.435 3.94 ;
      RECT 20.47 3.27 20.62 3.42 ;
      RECT 20.31 4.655 20.46 4.805 ;
      RECT 20.075 4.31 20.225 4.46 ;
      RECT 20.03 3.7 20.18 3.85 ;
      RECT 19.03 4.32 19.18 4.47 ;
      RECT 18.145 9.04 18.295 9.19 ;
      RECT 15.755 9.025 15.905 9.175 ;
      RECT 15.74 3.36 15.89 3.51 ;
      RECT 14.95 3.745 15.1 3.895 ;
      RECT 14.95 8.61 15.1 8.76 ;
      RECT 13.305 2.735 13.455 2.885 ;
      RECT 12.99 4.255 13.14 4.405 ;
      RECT 12.21 2.22 12.36 2.37 ;
      RECT 12.09 3.585 12.24 3.735 ;
      RECT 11.97 4.155 12.12 4.305 ;
      RECT 11.16 8.99 11.31 9.14 ;
      RECT 10.89 3.85 11.04 4 ;
      RECT 10.555 4.57 10.705 4.72 ;
      RECT 10.5 9.435 10.65 9.585 ;
      RECT 10.475 3.41 10.625 3.56 ;
      RECT 9.04 3.805 9.19 3.955 ;
      RECT 8.275 3.655 8.425 3.805 ;
      RECT 8.02 3.25 8.17 3.4 ;
      RECT 7.4 4.015 7.55 4.165 ;
      RECT 7.02 3.485 7.17 3.635 ;
      RECT 7.005 4.525 7.155 4.675 ;
      RECT 6.475 3.79 6.625 3.94 ;
      RECT 6.315 4.51 6.465 4.66 ;
      RECT 5.505 3.79 5.655 3.94 ;
      RECT 4.69 3.27 4.84 3.42 ;
      RECT 4.53 4.655 4.68 4.805 ;
      RECT 4.295 4.31 4.445 4.46 ;
      RECT 4.25 3.7 4.4 3.85 ;
      RECT 3.25 4.32 3.4 4.47 ;
      RECT 1.61 9.38 1.76 9.53 ;
      RECT 1.235 8.64 1.385 8.79 ;
    LAYER met1 ;
      RECT 66.125 2.555 75.785 3.035 ;
      RECT 50.34 2.555 60 3.035 ;
      RECT 34.555 2.555 44.215 3.035 ;
      RECT 18.78 2.555 28.44 3.035 ;
      RECT 3 2.555 12.66 3.035 ;
      RECT 66.125 2.555 75.84 2.885 ;
      RECT 50.34 2.555 60.055 2.885 ;
      RECT 34.555 2.555 44.27 2.885 ;
      RECT 18.78 2.555 28.495 2.885 ;
      RECT 3 2.555 12.715 2.885 ;
      RECT 66.24 0 75.955 2.88 ;
      RECT 50.455 0 60.17 2.88 ;
      RECT 34.67 0 44.385 2.88 ;
      RECT 18.895 0 28.61 2.88 ;
      RECT 3.115 0 12.83 2.88 ;
      RECT 0 0 81.72 1.6 ;
      RECT 81.115 10.055 81.405 10.285 ;
      RECT 81.175 8.575 81.345 10.285 ;
      RECT 81.15 9.56 81.5 9.91 ;
      RECT 81.115 8.575 81.405 8.805 ;
      RECT 80.71 3.69 80.815 4.26 ;
      RECT 80.71 4.025 81.035 4.255 ;
      RECT 80.71 4.055 81.205 4.225 ;
      RECT 80.71 3.69 80.9 4.255 ;
      RECT 80.125 3.655 80.415 3.885 ;
      RECT 80.125 3.69 80.9 3.86 ;
      RECT 80.185 2.175 80.355 3.885 ;
      RECT 80.125 2.175 80.415 2.405 ;
      RECT 80.125 10.055 80.415 10.285 ;
      RECT 80.185 8.575 80.355 10.285 ;
      RECT 80.125 8.575 80.415 8.805 ;
      RECT 80.125 8.61 80.98 8.77 ;
      RECT 80.81 8.205 80.98 8.77 ;
      RECT 80.125 8.605 80.52 8.77 ;
      RECT 80.745 8.205 81.035 8.435 ;
      RECT 80.745 8.235 81.205 8.405 ;
      RECT 79.755 4.025 80.045 4.255 ;
      RECT 79.755 4.055 80.215 4.225 ;
      RECT 79.82 2.95 79.985 4.255 ;
      RECT 78.335 2.92 78.625 3.15 ;
      RECT 78.335 2.95 79.985 3.12 ;
      RECT 78.395 2.18 78.565 3.15 ;
      RECT 78.335 2.18 78.625 2.41 ;
      RECT 78.335 10.05 78.625 10.28 ;
      RECT 78.395 9.31 78.565 10.28 ;
      RECT 78.395 9.405 79.985 9.575 ;
      RECT 79.815 8.205 79.985 9.575 ;
      RECT 78.335 9.31 78.625 9.54 ;
      RECT 79.755 8.205 80.045 8.435 ;
      RECT 79.755 8.235 80.215 8.405 ;
      RECT 78.765 3.26 79.115 3.61 ;
      RECT 76.43 3.32 79.115 3.49 ;
      RECT 76.43 2.635 76.6 3.49 ;
      RECT 76.33 2.635 76.68 2.985 ;
      RECT 78.79 8.94 79.115 9.265 ;
      RECT 74.165 8.895 74.515 9.245 ;
      RECT 78.765 8.94 79.115 9.17 ;
      RECT 73.985 8.94 74.515 9.17 ;
      RECT 73.815 8.97 79.115 9.14 ;
      RECT 77.99 3.66 78.31 3.98 ;
      RECT 77.96 3.66 78.31 3.89 ;
      RECT 77.79 3.69 78.31 3.86 ;
      RECT 77.99 8.54 78.31 8.83 ;
      RECT 77.96 8.57 78.31 8.8 ;
      RECT 77.79 8.6 78.31 8.77 ;
      RECT 74.625 3.76 74.81 3.97 ;
      RECT 74.615 3.765 74.825 3.963 ;
      RECT 74.615 3.765 74.911 3.94 ;
      RECT 74.615 3.765 74.97 3.915 ;
      RECT 74.615 3.765 75.025 3.895 ;
      RECT 74.615 3.765 75.035 3.883 ;
      RECT 74.615 3.765 75.23 3.822 ;
      RECT 74.615 3.765 75.26 3.805 ;
      RECT 74.615 3.765 75.28 3.795 ;
      RECT 75.16 3.53 75.42 3.79 ;
      RECT 75.145 3.62 75.16 3.837 ;
      RECT 74.68 3.752 75.42 3.79 ;
      RECT 75.131 3.631 75.145 3.843 ;
      RECT 74.72 3.745 75.42 3.79 ;
      RECT 75.045 3.671 75.131 3.862 ;
      RECT 74.97 3.732 75.42 3.79 ;
      RECT 75.04 3.707 75.045 3.879 ;
      RECT 75.025 3.717 75.42 3.79 ;
      RECT 75.035 3.712 75.04 3.881 ;
      RECT 75.33 4.217 75.335 4.309 ;
      RECT 75.325 4.195 75.33 4.326 ;
      RECT 75.32 4.185 75.325 4.338 ;
      RECT 75.31 4.176 75.32 4.348 ;
      RECT 75.305 4.171 75.31 4.356 ;
      RECT 75.3 4.03 75.305 4.359 ;
      RECT 75.266 4.03 75.3 4.37 ;
      RECT 75.18 4.03 75.266 4.405 ;
      RECT 75.1 4.03 75.18 4.453 ;
      RECT 75.071 4.03 75.1 4.477 ;
      RECT 74.985 4.03 75.071 4.483 ;
      RECT 74.98 4.214 74.985 4.488 ;
      RECT 74.945 4.225 74.98 4.491 ;
      RECT 74.92 4.24 74.945 4.495 ;
      RECT 74.906 4.249 74.92 4.497 ;
      RECT 74.82 4.276 74.906 4.503 ;
      RECT 74.755 4.317 74.82 4.512 ;
      RECT 74.74 4.337 74.755 4.517 ;
      RECT 74.71 4.347 74.74 4.52 ;
      RECT 74.705 4.357 74.71 4.523 ;
      RECT 74.675 4.362 74.705 4.525 ;
      RECT 74.655 4.367 74.675 4.529 ;
      RECT 74.57 4.37 74.655 4.536 ;
      RECT 74.555 4.367 74.57 4.542 ;
      RECT 74.545 4.364 74.555 4.544 ;
      RECT 74.525 4.361 74.545 4.546 ;
      RECT 74.505 4.357 74.525 4.547 ;
      RECT 74.49 4.353 74.505 4.549 ;
      RECT 74.48 4.35 74.49 4.55 ;
      RECT 74.44 4.344 74.48 4.548 ;
      RECT 74.43 4.339 74.44 4.546 ;
      RECT 74.415 4.336 74.43 4.542 ;
      RECT 74.39 4.331 74.415 4.535 ;
      RECT 74.34 4.322 74.39 4.523 ;
      RECT 74.27 4.308 74.34 4.505 ;
      RECT 74.212 4.293 74.27 4.487 ;
      RECT 74.126 4.276 74.212 4.467 ;
      RECT 74.04 4.255 74.126 4.442 ;
      RECT 73.99 4.24 74.04 4.423 ;
      RECT 73.986 4.234 73.99 4.415 ;
      RECT 73.9 4.224 73.986 4.402 ;
      RECT 73.865 4.209 73.9 4.385 ;
      RECT 73.85 4.202 73.865 4.378 ;
      RECT 73.79 4.19 73.85 4.366 ;
      RECT 73.77 4.177 73.79 4.354 ;
      RECT 73.73 4.168 73.77 4.346 ;
      RECT 73.725 4.16 73.73 4.339 ;
      RECT 73.645 4.15 73.725 4.325 ;
      RECT 73.63 4.137 73.645 4.31 ;
      RECT 73.625 4.135 73.63 4.308 ;
      RECT 73.546 4.123 73.625 4.295 ;
      RECT 73.46 4.098 73.546 4.27 ;
      RECT 73.445 4.067 73.46 4.255 ;
      RECT 73.43 4.042 73.445 4.251 ;
      RECT 73.415 4.035 73.43 4.247 ;
      RECT 73.24 4.04 73.245 4.243 ;
      RECT 73.235 4.045 73.24 4.238 ;
      RECT 73.245 4.035 73.415 4.245 ;
      RECT 73.96 3.795 74.065 4.055 ;
      RECT 74.775 3.32 74.78 3.545 ;
      RECT 74.905 3.32 74.96 3.53 ;
      RECT 74.96 3.325 74.97 3.523 ;
      RECT 74.866 3.32 74.905 3.533 ;
      RECT 74.78 3.32 74.866 3.54 ;
      RECT 74.76 3.325 74.775 3.546 ;
      RECT 74.75 3.365 74.76 3.548 ;
      RECT 74.72 3.375 74.75 3.55 ;
      RECT 74.715 3.38 74.72 3.552 ;
      RECT 74.69 3.385 74.715 3.554 ;
      RECT 74.675 3.39 74.69 3.556 ;
      RECT 74.66 3.392 74.675 3.558 ;
      RECT 74.655 3.397 74.66 3.56 ;
      RECT 74.605 3.405 74.655 3.563 ;
      RECT 74.58 3.414 74.605 3.568 ;
      RECT 74.57 3.421 74.58 3.573 ;
      RECT 74.565 3.424 74.57 3.577 ;
      RECT 74.545 3.427 74.565 3.586 ;
      RECT 74.515 3.435 74.545 3.606 ;
      RECT 74.486 3.448 74.515 3.628 ;
      RECT 74.4 3.482 74.486 3.672 ;
      RECT 74.395 3.508 74.4 3.71 ;
      RECT 74.39 3.512 74.395 3.719 ;
      RECT 74.355 3.525 74.39 3.752 ;
      RECT 74.345 3.539 74.355 3.79 ;
      RECT 74.34 3.543 74.345 3.803 ;
      RECT 74.335 3.547 74.34 3.808 ;
      RECT 74.325 3.555 74.335 3.82 ;
      RECT 74.32 3.562 74.325 3.835 ;
      RECT 74.295 3.575 74.32 3.86 ;
      RECT 74.255 3.604 74.295 3.915 ;
      RECT 74.24 3.629 74.255 3.97 ;
      RECT 74.23 3.64 74.24 3.993 ;
      RECT 74.225 3.647 74.23 4.005 ;
      RECT 74.22 3.651 74.225 4.013 ;
      RECT 74.165 3.679 74.22 4.055 ;
      RECT 74.145 3.715 74.165 4.055 ;
      RECT 74.13 3.73 74.145 4.055 ;
      RECT 74.075 3.762 74.13 4.055 ;
      RECT 74.065 3.792 74.075 4.055 ;
      RECT 73.675 3.407 73.86 3.645 ;
      RECT 73.66 3.409 73.87 3.64 ;
      RECT 73.545 3.355 73.805 3.615 ;
      RECT 73.54 3.392 73.805 3.569 ;
      RECT 73.535 3.402 73.805 3.566 ;
      RECT 73.53 3.442 73.87 3.56 ;
      RECT 73.525 3.475 73.87 3.55 ;
      RECT 73.535 3.417 73.885 3.488 ;
      RECT 73.832 4.515 73.845 5.045 ;
      RECT 73.746 4.515 73.845 5.044 ;
      RECT 73.746 4.515 73.85 5.043 ;
      RECT 73.66 4.515 73.85 5.041 ;
      RECT 73.655 4.515 73.85 5.038 ;
      RECT 73.655 4.515 73.86 5.036 ;
      RECT 73.65 4.807 73.86 5.033 ;
      RECT 73.65 4.817 73.865 5.03 ;
      RECT 73.65 4.885 73.87 5.026 ;
      RECT 73.64 4.89 73.87 5.025 ;
      RECT 73.64 4.982 73.875 5.022 ;
      RECT 73.625 4.515 73.885 4.775 ;
      RECT 73.555 10.05 73.845 10.28 ;
      RECT 73.615 9.31 73.785 10.28 ;
      RECT 73.53 9.34 73.87 9.685 ;
      RECT 73.555 9.31 73.845 9.685 ;
      RECT 72.855 3.505 72.9 5.04 ;
      RECT 73.055 3.505 73.085 3.72 ;
      RECT 71.43 3.245 71.55 3.455 ;
      RECT 71.09 3.195 71.35 3.455 ;
      RECT 71.09 3.24 71.385 3.445 ;
      RECT 73.095 3.521 73.1 3.575 ;
      RECT 73.09 3.514 73.095 3.708 ;
      RECT 73.085 3.508 73.09 3.715 ;
      RECT 73.04 3.505 73.055 3.728 ;
      RECT 73.035 3.505 73.04 3.75 ;
      RECT 73.03 3.505 73.035 3.798 ;
      RECT 73.025 3.505 73.03 3.818 ;
      RECT 73.015 3.505 73.025 3.925 ;
      RECT 73.01 3.505 73.015 3.988 ;
      RECT 73.005 3.505 73.01 4.045 ;
      RECT 73 3.505 73.005 4.053 ;
      RECT 72.985 3.505 73 4.16 ;
      RECT 72.975 3.505 72.985 4.295 ;
      RECT 72.965 3.505 72.975 4.405 ;
      RECT 72.955 3.505 72.965 4.462 ;
      RECT 72.95 3.505 72.955 4.502 ;
      RECT 72.945 3.505 72.95 4.538 ;
      RECT 72.935 3.505 72.945 4.578 ;
      RECT 72.93 3.505 72.935 4.62 ;
      RECT 72.91 3.505 72.93 4.685 ;
      RECT 72.915 4.83 72.92 5.01 ;
      RECT 72.91 4.812 72.915 5.018 ;
      RECT 72.905 3.505 72.91 4.748 ;
      RECT 72.905 4.792 72.91 5.025 ;
      RECT 72.9 3.505 72.905 5.035 ;
      RECT 72.845 3.505 72.855 3.805 ;
      RECT 72.85 4.052 72.855 5.04 ;
      RECT 72.845 4.117 72.85 5.04 ;
      RECT 72.84 3.506 72.845 3.795 ;
      RECT 72.835 4.182 72.845 5.04 ;
      RECT 72.83 3.507 72.84 3.785 ;
      RECT 72.82 4.295 72.835 5.04 ;
      RECT 72.825 3.508 72.83 3.775 ;
      RECT 72.805 3.509 72.825 3.753 ;
      RECT 72.81 4.392 72.82 5.04 ;
      RECT 72.805 4.467 72.81 5.04 ;
      RECT 72.795 3.508 72.805 3.73 ;
      RECT 72.8 4.51 72.805 5.04 ;
      RECT 72.795 4.537 72.8 5.04 ;
      RECT 72.785 3.506 72.795 3.718 ;
      RECT 72.79 4.58 72.795 5.04 ;
      RECT 72.785 4.607 72.79 5.04 ;
      RECT 72.775 3.505 72.785 3.705 ;
      RECT 72.78 4.622 72.785 5.04 ;
      RECT 72.74 4.68 72.78 5.04 ;
      RECT 72.77 3.504 72.775 3.69 ;
      RECT 72.765 3.502 72.77 3.683 ;
      RECT 72.755 3.499 72.765 3.673 ;
      RECT 72.75 3.496 72.755 3.658 ;
      RECT 72.735 3.492 72.75 3.651 ;
      RECT 72.73 4.735 72.74 5.04 ;
      RECT 72.73 3.489 72.735 3.646 ;
      RECT 72.715 3.485 72.73 3.64 ;
      RECT 72.725 4.752 72.73 5.04 ;
      RECT 72.715 4.815 72.725 5.04 ;
      RECT 72.635 3.47 72.715 3.62 ;
      RECT 72.71 4.822 72.715 5.035 ;
      RECT 72.705 4.83 72.71 5.025 ;
      RECT 72.625 3.456 72.635 3.604 ;
      RECT 72.61 3.452 72.625 3.602 ;
      RECT 72.6 3.447 72.61 3.598 ;
      RECT 72.575 3.44 72.6 3.59 ;
      RECT 72.57 3.435 72.575 3.585 ;
      RECT 72.56 3.435 72.57 3.583 ;
      RECT 72.55 3.433 72.56 3.581 ;
      RECT 72.52 3.425 72.55 3.575 ;
      RECT 72.505 3.417 72.52 3.568 ;
      RECT 72.485 3.412 72.505 3.561 ;
      RECT 72.48 3.408 72.485 3.556 ;
      RECT 72.45 3.401 72.48 3.55 ;
      RECT 72.425 3.392 72.45 3.54 ;
      RECT 72.395 3.385 72.425 3.532 ;
      RECT 72.37 3.375 72.395 3.523 ;
      RECT 72.355 3.367 72.37 3.517 ;
      RECT 72.33 3.362 72.355 3.512 ;
      RECT 72.32 3.358 72.33 3.507 ;
      RECT 72.3 3.353 72.32 3.502 ;
      RECT 72.265 3.348 72.3 3.495 ;
      RECT 72.205 3.343 72.265 3.488 ;
      RECT 72.192 3.339 72.205 3.486 ;
      RECT 72.106 3.334 72.192 3.483 ;
      RECT 72.02 3.324 72.106 3.479 ;
      RECT 71.979 3.317 72.02 3.476 ;
      RECT 71.893 3.31 71.979 3.473 ;
      RECT 71.807 3.3 71.893 3.469 ;
      RECT 71.721 3.29 71.807 3.464 ;
      RECT 71.635 3.28 71.721 3.46 ;
      RECT 71.625 3.265 71.635 3.458 ;
      RECT 71.615 3.25 71.625 3.458 ;
      RECT 71.55 3.245 71.615 3.457 ;
      RECT 71.385 3.242 71.43 3.45 ;
      RECT 72.63 4.147 72.635 4.338 ;
      RECT 72.625 4.142 72.63 4.345 ;
      RECT 72.611 4.14 72.625 4.351 ;
      RECT 72.525 4.14 72.611 4.353 ;
      RECT 72.521 4.14 72.525 4.356 ;
      RECT 72.435 4.14 72.521 4.374 ;
      RECT 72.425 4.145 72.435 4.393 ;
      RECT 72.415 4.2 72.425 4.397 ;
      RECT 72.39 4.215 72.415 4.404 ;
      RECT 72.35 4.235 72.39 4.417 ;
      RECT 72.345 4.247 72.35 4.427 ;
      RECT 72.33 4.253 72.345 4.432 ;
      RECT 72.325 4.258 72.33 4.436 ;
      RECT 72.305 4.265 72.325 4.441 ;
      RECT 72.235 4.29 72.305 4.458 ;
      RECT 72.195 4.318 72.235 4.478 ;
      RECT 72.19 4.328 72.195 4.486 ;
      RECT 72.17 4.335 72.19 4.488 ;
      RECT 72.165 4.342 72.17 4.491 ;
      RECT 72.135 4.35 72.165 4.494 ;
      RECT 72.13 4.355 72.135 4.498 ;
      RECT 72.056 4.359 72.13 4.506 ;
      RECT 71.97 4.368 72.056 4.522 ;
      RECT 71.966 4.373 71.97 4.531 ;
      RECT 71.88 4.378 71.966 4.541 ;
      RECT 71.84 4.386 71.88 4.553 ;
      RECT 71.79 4.392 71.84 4.56 ;
      RECT 71.705 4.401 71.79 4.575 ;
      RECT 71.63 4.412 71.705 4.593 ;
      RECT 71.595 4.419 71.63 4.603 ;
      RECT 71.52 4.427 71.595 4.608 ;
      RECT 71.465 4.436 71.52 4.608 ;
      RECT 71.44 4.441 71.465 4.606 ;
      RECT 71.43 4.444 71.44 4.604 ;
      RECT 71.395 4.446 71.43 4.602 ;
      RECT 71.365 4.448 71.395 4.598 ;
      RECT 71.32 4.447 71.365 4.594 ;
      RECT 71.3 4.442 71.32 4.591 ;
      RECT 71.25 4.427 71.3 4.588 ;
      RECT 71.24 4.412 71.25 4.583 ;
      RECT 71.19 4.397 71.24 4.573 ;
      RECT 71.14 4.372 71.19 4.553 ;
      RECT 71.13 4.357 71.14 4.535 ;
      RECT 71.125 4.355 71.13 4.529 ;
      RECT 71.105 4.35 71.125 4.524 ;
      RECT 71.1 4.342 71.105 4.518 ;
      RECT 71.085 4.336 71.1 4.511 ;
      RECT 71.08 4.331 71.085 4.503 ;
      RECT 71.06 4.326 71.08 4.495 ;
      RECT 71.045 4.319 71.06 4.488 ;
      RECT 71.03 4.313 71.045 4.479 ;
      RECT 71.025 4.307 71.03 4.472 ;
      RECT 70.98 4.282 71.025 4.458 ;
      RECT 70.965 4.252 70.98 4.44 ;
      RECT 70.95 4.235 70.965 4.431 ;
      RECT 70.925 4.215 70.95 4.419 ;
      RECT 70.885 4.185 70.925 4.399 ;
      RECT 70.875 4.155 70.885 4.384 ;
      RECT 70.86 4.145 70.875 4.377 ;
      RECT 70.805 4.11 70.86 4.356 ;
      RECT 70.79 4.073 70.805 4.335 ;
      RECT 70.78 4.06 70.79 4.327 ;
      RECT 70.73 4.03 70.78 4.309 ;
      RECT 70.715 3.96 70.73 4.29 ;
      RECT 70.67 3.96 70.715 4.273 ;
      RECT 70.645 3.96 70.67 4.255 ;
      RECT 70.635 3.96 70.645 4.248 ;
      RECT 70.556 3.96 70.635 4.241 ;
      RECT 70.47 3.96 70.556 4.233 ;
      RECT 70.455 3.992 70.47 4.228 ;
      RECT 70.38 4.002 70.455 4.224 ;
      RECT 70.36 4.012 70.38 4.219 ;
      RECT 70.335 4.012 70.36 4.216 ;
      RECT 70.325 4.002 70.335 4.215 ;
      RECT 70.315 3.975 70.325 4.214 ;
      RECT 70.275 3.97 70.315 4.212 ;
      RECT 70.23 3.97 70.275 4.208 ;
      RECT 70.205 3.97 70.23 4.203 ;
      RECT 70.155 3.97 70.205 4.19 ;
      RECT 70.115 3.975 70.125 4.175 ;
      RECT 70.125 3.97 70.155 4.18 ;
      RECT 72.11 3.75 72.37 4.01 ;
      RECT 72.105 3.772 72.37 3.968 ;
      RECT 71.345 3.6 71.565 3.965 ;
      RECT 71.327 3.687 71.565 3.964 ;
      RECT 71.31 3.692 71.565 3.961 ;
      RECT 71.31 3.692 71.585 3.96 ;
      RECT 71.28 3.702 71.585 3.958 ;
      RECT 71.275 3.717 71.585 3.954 ;
      RECT 71.275 3.717 71.59 3.953 ;
      RECT 71.27 3.775 71.59 3.951 ;
      RECT 71.27 3.775 71.6 3.948 ;
      RECT 71.265 3.84 71.6 3.943 ;
      RECT 71.345 3.6 71.605 3.86 ;
      RECT 70.09 3.43 70.35 3.69 ;
      RECT 70.09 3.473 70.436 3.664 ;
      RECT 70.09 3.473 70.48 3.663 ;
      RECT 70.09 3.473 70.5 3.661 ;
      RECT 70.09 3.473 70.6 3.66 ;
      RECT 70.09 3.473 70.62 3.658 ;
      RECT 70.09 3.473 70.63 3.653 ;
      RECT 70.5 3.44 70.69 3.65 ;
      RECT 70.5 3.442 70.695 3.648 ;
      RECT 70.49 3.447 70.7 3.64 ;
      RECT 70.436 3.471 70.7 3.64 ;
      RECT 70.48 3.465 70.49 3.662 ;
      RECT 70.49 3.445 70.695 3.648 ;
      RECT 69.445 4.505 69.65 4.735 ;
      RECT 69.385 4.455 69.44 4.715 ;
      RECT 69.445 4.455 69.645 4.735 ;
      RECT 70.415 4.77 70.42 4.797 ;
      RECT 70.405 4.68 70.415 4.802 ;
      RECT 70.4 4.602 70.405 4.808 ;
      RECT 70.39 4.592 70.4 4.815 ;
      RECT 70.385 4.582 70.39 4.821 ;
      RECT 70.375 4.577 70.385 4.823 ;
      RECT 70.36 4.569 70.375 4.831 ;
      RECT 70.345 4.56 70.36 4.843 ;
      RECT 70.335 4.552 70.345 4.853 ;
      RECT 70.3 4.47 70.335 4.871 ;
      RECT 70.265 4.47 70.3 4.89 ;
      RECT 70.25 4.47 70.265 4.898 ;
      RECT 70.195 4.47 70.25 4.898 ;
      RECT 70.161 4.47 70.195 4.889 ;
      RECT 70.075 4.47 70.161 4.865 ;
      RECT 70.065 4.53 70.075 4.847 ;
      RECT 70.025 4.532 70.065 4.838 ;
      RECT 70.02 4.534 70.025 4.828 ;
      RECT 70 4.536 70.02 4.823 ;
      RECT 69.99 4.539 70 4.818 ;
      RECT 69.98 4.54 69.99 4.813 ;
      RECT 69.956 4.541 69.98 4.805 ;
      RECT 69.87 4.546 69.956 4.783 ;
      RECT 69.815 4.545 69.87 4.756 ;
      RECT 69.8 4.538 69.815 4.743 ;
      RECT 69.765 4.533 69.8 4.739 ;
      RECT 69.71 4.525 69.765 4.738 ;
      RECT 69.65 4.512 69.71 4.736 ;
      RECT 69.44 4.455 69.445 4.723 ;
      RECT 69.515 3.825 69.7 4.035 ;
      RECT 69.505 3.83 69.715 4.028 ;
      RECT 69.545 3.735 69.805 3.995 ;
      RECT 69.5 3.892 69.805 3.918 ;
      RECT 68.845 3.685 68.85 4.485 ;
      RECT 68.79 3.735 68.82 4.485 ;
      RECT 68.78 3.735 68.785 4.045 ;
      RECT 68.765 3.735 68.77 4.04 ;
      RECT 68.31 3.78 68.325 3.995 ;
      RECT 68.24 3.78 68.325 3.99 ;
      RECT 69.505 3.36 69.575 3.57 ;
      RECT 69.575 3.367 69.585 3.565 ;
      RECT 69.471 3.36 69.505 3.577 ;
      RECT 69.385 3.36 69.471 3.601 ;
      RECT 69.375 3.365 69.385 3.62 ;
      RECT 69.37 3.377 69.375 3.623 ;
      RECT 69.355 3.392 69.37 3.627 ;
      RECT 69.35 3.41 69.355 3.631 ;
      RECT 69.31 3.42 69.35 3.64 ;
      RECT 69.295 3.427 69.31 3.652 ;
      RECT 69.28 3.432 69.295 3.657 ;
      RECT 69.265 3.435 69.28 3.662 ;
      RECT 69.255 3.437 69.265 3.666 ;
      RECT 69.22 3.444 69.255 3.674 ;
      RECT 69.185 3.452 69.22 3.688 ;
      RECT 69.175 3.458 69.185 3.697 ;
      RECT 69.17 3.46 69.175 3.699 ;
      RECT 69.15 3.463 69.17 3.705 ;
      RECT 69.12 3.47 69.15 3.716 ;
      RECT 69.11 3.476 69.12 3.723 ;
      RECT 69.085 3.479 69.11 3.73 ;
      RECT 69.075 3.483 69.085 3.738 ;
      RECT 69.07 3.484 69.075 3.76 ;
      RECT 69.065 3.485 69.07 3.775 ;
      RECT 69.06 3.486 69.065 3.79 ;
      RECT 69.055 3.487 69.06 3.805 ;
      RECT 69.05 3.488 69.055 3.835 ;
      RECT 69.04 3.49 69.05 3.868 ;
      RECT 69.025 3.494 69.04 3.915 ;
      RECT 69.015 3.497 69.025 3.96 ;
      RECT 69.01 3.5 69.015 3.988 ;
      RECT 69 3.502 69.01 4.015 ;
      RECT 68.995 3.505 69 4.05 ;
      RECT 68.965 3.51 68.995 4.108 ;
      RECT 68.96 3.515 68.965 4.193 ;
      RECT 68.955 3.517 68.96 4.228 ;
      RECT 68.95 3.519 68.955 4.31 ;
      RECT 68.945 3.521 68.95 4.398 ;
      RECT 68.935 3.523 68.945 4.48 ;
      RECT 68.92 3.537 68.935 4.485 ;
      RECT 68.885 3.582 68.92 4.485 ;
      RECT 68.875 3.622 68.885 4.485 ;
      RECT 68.86 3.65 68.875 4.485 ;
      RECT 68.855 3.667 68.86 4.485 ;
      RECT 68.85 3.675 68.855 4.485 ;
      RECT 68.84 3.69 68.845 4.485 ;
      RECT 68.835 3.697 68.84 4.485 ;
      RECT 68.825 3.717 68.835 4.485 ;
      RECT 68.82 3.73 68.825 4.485 ;
      RECT 68.785 3.735 68.79 4.07 ;
      RECT 68.77 4.125 68.79 4.485 ;
      RECT 68.77 3.735 68.78 4.043 ;
      RECT 68.765 4.165 68.77 4.485 ;
      RECT 68.715 3.735 68.765 4.038 ;
      RECT 68.76 4.202 68.765 4.485 ;
      RECT 68.75 4.225 68.76 4.485 ;
      RECT 68.745 4.27 68.75 4.485 ;
      RECT 68.735 4.28 68.745 4.478 ;
      RECT 68.661 3.735 68.715 4.032 ;
      RECT 68.575 3.735 68.661 4.025 ;
      RECT 68.526 3.782 68.575 4.018 ;
      RECT 68.44 3.79 68.526 4.011 ;
      RECT 68.425 3.787 68.44 4.006 ;
      RECT 68.411 3.78 68.425 4.005 ;
      RECT 68.325 3.78 68.411 4 ;
      RECT 68.23 3.785 68.24 3.985 ;
      RECT 67.82 3.215 67.835 3.615 ;
      RECT 68.015 3.215 68.02 3.475 ;
      RECT 67.76 3.215 67.805 3.475 ;
      RECT 68.215 4.52 68.22 4.725 ;
      RECT 68.21 4.51 68.215 4.73 ;
      RECT 68.205 4.497 68.21 4.735 ;
      RECT 68.2 4.477 68.205 4.735 ;
      RECT 68.175 4.43 68.2 4.735 ;
      RECT 68.14 4.345 68.175 4.735 ;
      RECT 68.135 4.282 68.14 4.735 ;
      RECT 68.13 4.267 68.135 4.735 ;
      RECT 68.115 4.227 68.13 4.735 ;
      RECT 68.11 4.202 68.115 4.735 ;
      RECT 68.1 4.185 68.11 4.735 ;
      RECT 68.065 4.107 68.1 4.735 ;
      RECT 68.06 4.05 68.065 4.735 ;
      RECT 68.055 4.037 68.06 4.735 ;
      RECT 68.045 4.015 68.055 4.735 ;
      RECT 68.035 3.98 68.045 4.735 ;
      RECT 68.025 3.95 68.035 4.735 ;
      RECT 68.015 3.865 68.025 4.378 ;
      RECT 68.022 4.51 68.025 4.735 ;
      RECT 68.02 4.52 68.022 4.735 ;
      RECT 68.01 4.53 68.02 4.73 ;
      RECT 68.005 3.215 68.015 3.61 ;
      RECT 68.01 3.742 68.015 4.353 ;
      RECT 68.005 3.64 68.01 4.336 ;
      RECT 67.995 3.215 68.005 4.312 ;
      RECT 67.99 3.215 67.995 4.283 ;
      RECT 67.985 3.215 67.99 4.273 ;
      RECT 67.965 3.215 67.985 4.235 ;
      RECT 67.96 3.215 67.965 4.193 ;
      RECT 67.955 3.215 67.96 4.173 ;
      RECT 67.925 3.215 67.955 4.123 ;
      RECT 67.915 3.215 67.925 4.07 ;
      RECT 67.91 3.215 67.915 4.043 ;
      RECT 67.905 3.215 67.91 4.028 ;
      RECT 67.895 3.215 67.905 4.005 ;
      RECT 67.885 3.215 67.895 3.98 ;
      RECT 67.88 3.215 67.885 3.92 ;
      RECT 67.87 3.215 67.88 3.858 ;
      RECT 67.865 3.215 67.87 3.778 ;
      RECT 67.86 3.215 67.865 3.743 ;
      RECT 67.855 3.215 67.86 3.718 ;
      RECT 67.85 3.215 67.855 3.703 ;
      RECT 67.845 3.215 67.85 3.673 ;
      RECT 67.84 3.215 67.845 3.65 ;
      RECT 67.835 3.215 67.84 3.623 ;
      RECT 67.805 3.215 67.82 3.61 ;
      RECT 66.96 4.75 67.145 4.96 ;
      RECT 66.95 4.755 67.16 4.953 ;
      RECT 66.95 4.755 67.18 4.925 ;
      RECT 66.95 4.755 67.195 4.904 ;
      RECT 66.95 4.755 67.21 4.902 ;
      RECT 66.95 4.755 67.22 4.901 ;
      RECT 66.95 4.755 67.25 4.898 ;
      RECT 67.6 4.6 67.86 4.86 ;
      RECT 67.56 4.647 67.86 4.843 ;
      RECT 67.551 4.655 67.56 4.846 ;
      RECT 67.145 4.748 67.86 4.843 ;
      RECT 67.465 4.673 67.551 4.853 ;
      RECT 67.16 4.745 67.86 4.843 ;
      RECT 67.406 4.695 67.465 4.865 ;
      RECT 67.18 4.741 67.86 4.843 ;
      RECT 67.32 4.707 67.406 4.876 ;
      RECT 67.195 4.737 67.86 4.843 ;
      RECT 67.265 4.72 67.32 4.888 ;
      RECT 67.21 4.735 67.86 4.843 ;
      RECT 67.25 4.726 67.265 4.894 ;
      RECT 67.22 4.731 67.86 4.843 ;
      RECT 67.365 4.255 67.625 4.515 ;
      RECT 67.365 4.275 67.735 4.485 ;
      RECT 67.365 4.28 67.745 4.48 ;
      RECT 67.556 3.694 67.635 3.925 ;
      RECT 67.47 3.697 67.685 3.92 ;
      RECT 67.465 3.697 67.685 3.915 ;
      RECT 67.465 3.702 67.695 3.913 ;
      RECT 67.44 3.702 67.695 3.91 ;
      RECT 67.44 3.71 67.705 3.908 ;
      RECT 67.32 3.645 67.58 3.905 ;
      RECT 67.32 3.692 67.63 3.905 ;
      RECT 66.575 4.265 66.58 4.525 ;
      RECT 66.405 4.035 66.41 4.525 ;
      RECT 66.29 4.275 66.295 4.5 ;
      RECT 67 3.37 67.005 3.58 ;
      RECT 67.005 3.375 67.02 3.575 ;
      RECT 66.94 3.37 67 3.588 ;
      RECT 66.925 3.37 66.94 3.598 ;
      RECT 66.875 3.37 66.925 3.615 ;
      RECT 66.855 3.37 66.875 3.638 ;
      RECT 66.84 3.37 66.855 3.65 ;
      RECT 66.82 3.37 66.84 3.66 ;
      RECT 66.81 3.375 66.82 3.669 ;
      RECT 66.805 3.385 66.81 3.674 ;
      RECT 66.8 3.397 66.805 3.678 ;
      RECT 66.79 3.42 66.8 3.683 ;
      RECT 66.785 3.435 66.79 3.687 ;
      RECT 66.78 3.452 66.785 3.69 ;
      RECT 66.775 3.46 66.78 3.693 ;
      RECT 66.765 3.465 66.775 3.697 ;
      RECT 66.76 3.472 66.765 3.702 ;
      RECT 66.75 3.477 66.76 3.706 ;
      RECT 66.725 3.489 66.75 3.717 ;
      RECT 66.705 3.506 66.725 3.733 ;
      RECT 66.68 3.523 66.705 3.755 ;
      RECT 66.645 3.546 66.68 3.813 ;
      RECT 66.625 3.568 66.645 3.875 ;
      RECT 66.62 3.578 66.625 3.91 ;
      RECT 66.61 3.585 66.62 3.948 ;
      RECT 66.605 3.592 66.61 3.968 ;
      RECT 66.6 3.603 66.605 4.005 ;
      RECT 66.595 3.611 66.6 4.07 ;
      RECT 66.585 3.622 66.595 4.123 ;
      RECT 66.58 3.64 66.585 4.193 ;
      RECT 66.575 3.65 66.58 4.23 ;
      RECT 66.57 3.66 66.575 4.525 ;
      RECT 66.565 3.672 66.57 4.525 ;
      RECT 66.56 3.682 66.565 4.525 ;
      RECT 66.55 3.692 66.56 4.525 ;
      RECT 66.54 3.715 66.55 4.525 ;
      RECT 66.525 3.75 66.54 4.525 ;
      RECT 66.485 3.812 66.525 4.525 ;
      RECT 66.48 3.865 66.485 4.525 ;
      RECT 66.455 3.9 66.48 4.525 ;
      RECT 66.44 3.945 66.455 4.525 ;
      RECT 66.435 3.967 66.44 4.525 ;
      RECT 66.425 3.98 66.435 4.525 ;
      RECT 66.415 4.005 66.425 4.525 ;
      RECT 66.41 4.027 66.415 4.525 ;
      RECT 66.385 4.065 66.405 4.525 ;
      RECT 66.345 4.122 66.385 4.525 ;
      RECT 66.34 4.172 66.345 4.525 ;
      RECT 66.335 4.19 66.34 4.525 ;
      RECT 66.33 4.202 66.335 4.525 ;
      RECT 66.32 4.22 66.33 4.525 ;
      RECT 66.31 4.24 66.32 4.5 ;
      RECT 66.305 4.257 66.31 4.5 ;
      RECT 66.295 4.27 66.305 4.5 ;
      RECT 66.265 4.28 66.29 4.5 ;
      RECT 66.255 4.287 66.265 4.5 ;
      RECT 66.24 4.297 66.255 4.495 ;
      RECT 65.33 10.055 65.62 10.285 ;
      RECT 65.39 8.575 65.56 10.285 ;
      RECT 65.34 8.94 65.69 9.29 ;
      RECT 65.33 8.575 65.62 8.805 ;
      RECT 64.925 3.69 65.03 4.26 ;
      RECT 64.925 4.025 65.25 4.255 ;
      RECT 64.925 4.055 65.42 4.225 ;
      RECT 64.925 3.69 65.115 4.255 ;
      RECT 64.34 3.655 64.63 3.885 ;
      RECT 64.34 3.69 65.115 3.86 ;
      RECT 64.4 2.175 64.57 3.885 ;
      RECT 64.34 2.175 64.63 2.405 ;
      RECT 64.34 10.055 64.63 10.285 ;
      RECT 64.4 8.575 64.57 10.285 ;
      RECT 64.34 8.575 64.63 8.805 ;
      RECT 64.34 8.61 65.195 8.77 ;
      RECT 65.025 8.205 65.195 8.77 ;
      RECT 64.34 8.605 64.735 8.77 ;
      RECT 64.96 8.205 65.25 8.435 ;
      RECT 64.96 8.235 65.42 8.405 ;
      RECT 63.97 4.025 64.26 4.255 ;
      RECT 63.97 4.055 64.43 4.225 ;
      RECT 64.035 2.95 64.2 4.255 ;
      RECT 62.55 2.92 62.84 3.15 ;
      RECT 62.55 2.95 64.2 3.12 ;
      RECT 62.61 2.18 62.78 3.15 ;
      RECT 62.55 2.18 62.84 2.41 ;
      RECT 62.55 10.05 62.84 10.28 ;
      RECT 62.61 9.31 62.78 10.28 ;
      RECT 62.61 9.405 64.2 9.575 ;
      RECT 64.03 8.205 64.2 9.575 ;
      RECT 62.55 9.31 62.84 9.54 ;
      RECT 63.97 8.205 64.26 8.435 ;
      RECT 63.97 8.235 64.43 8.405 ;
      RECT 62.98 3.26 63.33 3.61 ;
      RECT 60.645 3.32 63.33 3.49 ;
      RECT 60.645 2.635 60.815 3.49 ;
      RECT 60.545 2.635 60.895 2.985 ;
      RECT 63.005 8.94 63.33 9.265 ;
      RECT 58.38 8.895 58.73 9.245 ;
      RECT 62.98 8.94 63.33 9.17 ;
      RECT 58.2 8.94 58.73 9.17 ;
      RECT 58.03 8.97 63.33 9.14 ;
      RECT 62.205 3.66 62.525 3.98 ;
      RECT 62.175 3.66 62.525 3.89 ;
      RECT 62.005 3.69 62.525 3.86 ;
      RECT 62.205 8.54 62.525 8.83 ;
      RECT 62.175 8.57 62.525 8.8 ;
      RECT 62.005 8.6 62.525 8.77 ;
      RECT 58.84 3.76 59.025 3.97 ;
      RECT 58.83 3.765 59.04 3.963 ;
      RECT 58.83 3.765 59.126 3.94 ;
      RECT 58.83 3.765 59.185 3.915 ;
      RECT 58.83 3.765 59.24 3.895 ;
      RECT 58.83 3.765 59.25 3.883 ;
      RECT 58.83 3.765 59.445 3.822 ;
      RECT 58.83 3.765 59.475 3.805 ;
      RECT 58.83 3.765 59.495 3.795 ;
      RECT 59.375 3.53 59.635 3.79 ;
      RECT 59.36 3.62 59.375 3.837 ;
      RECT 58.895 3.752 59.635 3.79 ;
      RECT 59.346 3.631 59.36 3.843 ;
      RECT 58.935 3.745 59.635 3.79 ;
      RECT 59.26 3.671 59.346 3.862 ;
      RECT 59.185 3.732 59.635 3.79 ;
      RECT 59.255 3.707 59.26 3.879 ;
      RECT 59.24 3.717 59.635 3.79 ;
      RECT 59.25 3.712 59.255 3.881 ;
      RECT 59.545 4.217 59.55 4.309 ;
      RECT 59.54 4.195 59.545 4.326 ;
      RECT 59.535 4.185 59.54 4.338 ;
      RECT 59.525 4.176 59.535 4.348 ;
      RECT 59.52 4.171 59.525 4.356 ;
      RECT 59.515 4.03 59.52 4.359 ;
      RECT 59.481 4.03 59.515 4.37 ;
      RECT 59.395 4.03 59.481 4.405 ;
      RECT 59.315 4.03 59.395 4.453 ;
      RECT 59.286 4.03 59.315 4.477 ;
      RECT 59.2 4.03 59.286 4.483 ;
      RECT 59.195 4.214 59.2 4.488 ;
      RECT 59.16 4.225 59.195 4.491 ;
      RECT 59.135 4.24 59.16 4.495 ;
      RECT 59.121 4.249 59.135 4.497 ;
      RECT 59.035 4.276 59.121 4.503 ;
      RECT 58.97 4.317 59.035 4.512 ;
      RECT 58.955 4.337 58.97 4.517 ;
      RECT 58.925 4.347 58.955 4.52 ;
      RECT 58.92 4.357 58.925 4.523 ;
      RECT 58.89 4.362 58.92 4.525 ;
      RECT 58.87 4.367 58.89 4.529 ;
      RECT 58.785 4.37 58.87 4.536 ;
      RECT 58.77 4.367 58.785 4.542 ;
      RECT 58.76 4.364 58.77 4.544 ;
      RECT 58.74 4.361 58.76 4.546 ;
      RECT 58.72 4.357 58.74 4.547 ;
      RECT 58.705 4.353 58.72 4.549 ;
      RECT 58.695 4.35 58.705 4.55 ;
      RECT 58.655 4.344 58.695 4.548 ;
      RECT 58.645 4.339 58.655 4.546 ;
      RECT 58.63 4.336 58.645 4.542 ;
      RECT 58.605 4.331 58.63 4.535 ;
      RECT 58.555 4.322 58.605 4.523 ;
      RECT 58.485 4.308 58.555 4.505 ;
      RECT 58.427 4.293 58.485 4.487 ;
      RECT 58.341 4.276 58.427 4.467 ;
      RECT 58.255 4.255 58.341 4.442 ;
      RECT 58.205 4.24 58.255 4.423 ;
      RECT 58.201 4.234 58.205 4.415 ;
      RECT 58.115 4.224 58.201 4.402 ;
      RECT 58.08 4.209 58.115 4.385 ;
      RECT 58.065 4.202 58.08 4.378 ;
      RECT 58.005 4.19 58.065 4.366 ;
      RECT 57.985 4.177 58.005 4.354 ;
      RECT 57.945 4.168 57.985 4.346 ;
      RECT 57.94 4.16 57.945 4.339 ;
      RECT 57.86 4.15 57.94 4.325 ;
      RECT 57.845 4.137 57.86 4.31 ;
      RECT 57.84 4.135 57.845 4.308 ;
      RECT 57.761 4.123 57.84 4.295 ;
      RECT 57.675 4.098 57.761 4.27 ;
      RECT 57.66 4.067 57.675 4.255 ;
      RECT 57.645 4.042 57.66 4.251 ;
      RECT 57.63 4.035 57.645 4.247 ;
      RECT 57.455 4.04 57.46 4.243 ;
      RECT 57.45 4.045 57.455 4.238 ;
      RECT 57.46 4.035 57.63 4.245 ;
      RECT 58.175 3.795 58.28 4.055 ;
      RECT 58.99 3.32 58.995 3.545 ;
      RECT 59.12 3.32 59.175 3.53 ;
      RECT 59.175 3.325 59.185 3.523 ;
      RECT 59.081 3.32 59.12 3.533 ;
      RECT 58.995 3.32 59.081 3.54 ;
      RECT 58.975 3.325 58.99 3.546 ;
      RECT 58.965 3.365 58.975 3.548 ;
      RECT 58.935 3.375 58.965 3.55 ;
      RECT 58.93 3.38 58.935 3.552 ;
      RECT 58.905 3.385 58.93 3.554 ;
      RECT 58.89 3.39 58.905 3.556 ;
      RECT 58.875 3.392 58.89 3.558 ;
      RECT 58.87 3.397 58.875 3.56 ;
      RECT 58.82 3.405 58.87 3.563 ;
      RECT 58.795 3.414 58.82 3.568 ;
      RECT 58.785 3.421 58.795 3.573 ;
      RECT 58.78 3.424 58.785 3.577 ;
      RECT 58.76 3.427 58.78 3.586 ;
      RECT 58.73 3.435 58.76 3.606 ;
      RECT 58.701 3.448 58.73 3.628 ;
      RECT 58.615 3.482 58.701 3.672 ;
      RECT 58.61 3.508 58.615 3.71 ;
      RECT 58.605 3.512 58.61 3.719 ;
      RECT 58.57 3.525 58.605 3.752 ;
      RECT 58.56 3.539 58.57 3.79 ;
      RECT 58.555 3.543 58.56 3.803 ;
      RECT 58.55 3.547 58.555 3.808 ;
      RECT 58.54 3.555 58.55 3.82 ;
      RECT 58.535 3.562 58.54 3.835 ;
      RECT 58.51 3.575 58.535 3.86 ;
      RECT 58.47 3.604 58.51 3.915 ;
      RECT 58.455 3.629 58.47 3.97 ;
      RECT 58.445 3.64 58.455 3.993 ;
      RECT 58.44 3.647 58.445 4.005 ;
      RECT 58.435 3.651 58.44 4.013 ;
      RECT 58.38 3.679 58.435 4.055 ;
      RECT 58.36 3.715 58.38 4.055 ;
      RECT 58.345 3.73 58.36 4.055 ;
      RECT 58.29 3.762 58.345 4.055 ;
      RECT 58.28 3.792 58.29 4.055 ;
      RECT 57.89 3.407 58.075 3.645 ;
      RECT 57.875 3.409 58.085 3.64 ;
      RECT 57.76 3.355 58.02 3.615 ;
      RECT 57.755 3.392 58.02 3.569 ;
      RECT 57.75 3.402 58.02 3.566 ;
      RECT 57.745 3.442 58.085 3.56 ;
      RECT 57.74 3.475 58.085 3.55 ;
      RECT 57.75 3.417 58.1 3.488 ;
      RECT 58.047 4.515 58.06 5.045 ;
      RECT 57.961 4.515 58.06 5.044 ;
      RECT 57.961 4.515 58.065 5.043 ;
      RECT 57.875 4.515 58.065 5.041 ;
      RECT 57.87 4.515 58.065 5.038 ;
      RECT 57.87 4.515 58.075 5.036 ;
      RECT 57.865 4.807 58.075 5.033 ;
      RECT 57.865 4.817 58.08 5.03 ;
      RECT 57.865 4.885 58.085 5.026 ;
      RECT 57.855 4.89 58.085 5.025 ;
      RECT 57.855 4.982 58.09 5.022 ;
      RECT 57.84 4.515 58.1 4.775 ;
      RECT 57.77 10.05 58.06 10.28 ;
      RECT 57.83 9.31 58 10.28 ;
      RECT 57.745 9.34 58.085 9.685 ;
      RECT 57.77 9.31 58.06 9.685 ;
      RECT 57.07 3.505 57.115 5.04 ;
      RECT 57.27 3.505 57.3 3.72 ;
      RECT 55.645 3.245 55.765 3.455 ;
      RECT 55.305 3.195 55.565 3.455 ;
      RECT 55.305 3.24 55.6 3.445 ;
      RECT 57.31 3.521 57.315 3.575 ;
      RECT 57.305 3.514 57.31 3.708 ;
      RECT 57.3 3.508 57.305 3.715 ;
      RECT 57.255 3.505 57.27 3.728 ;
      RECT 57.25 3.505 57.255 3.75 ;
      RECT 57.245 3.505 57.25 3.798 ;
      RECT 57.24 3.505 57.245 3.818 ;
      RECT 57.23 3.505 57.24 3.925 ;
      RECT 57.225 3.505 57.23 3.988 ;
      RECT 57.22 3.505 57.225 4.045 ;
      RECT 57.215 3.505 57.22 4.053 ;
      RECT 57.2 3.505 57.215 4.16 ;
      RECT 57.19 3.505 57.2 4.295 ;
      RECT 57.18 3.505 57.19 4.405 ;
      RECT 57.17 3.505 57.18 4.462 ;
      RECT 57.165 3.505 57.17 4.502 ;
      RECT 57.16 3.505 57.165 4.538 ;
      RECT 57.15 3.505 57.16 4.578 ;
      RECT 57.145 3.505 57.15 4.62 ;
      RECT 57.125 3.505 57.145 4.685 ;
      RECT 57.13 4.83 57.135 5.01 ;
      RECT 57.125 4.812 57.13 5.018 ;
      RECT 57.12 3.505 57.125 4.748 ;
      RECT 57.12 4.792 57.125 5.025 ;
      RECT 57.115 3.505 57.12 5.035 ;
      RECT 57.06 3.505 57.07 3.805 ;
      RECT 57.065 4.052 57.07 5.04 ;
      RECT 57.06 4.117 57.065 5.04 ;
      RECT 57.055 3.506 57.06 3.795 ;
      RECT 57.05 4.182 57.06 5.04 ;
      RECT 57.045 3.507 57.055 3.785 ;
      RECT 57.035 4.295 57.05 5.04 ;
      RECT 57.04 3.508 57.045 3.775 ;
      RECT 57.02 3.509 57.04 3.753 ;
      RECT 57.025 4.392 57.035 5.04 ;
      RECT 57.02 4.467 57.025 5.04 ;
      RECT 57.01 3.508 57.02 3.73 ;
      RECT 57.015 4.51 57.02 5.04 ;
      RECT 57.01 4.537 57.015 5.04 ;
      RECT 57 3.506 57.01 3.718 ;
      RECT 57.005 4.58 57.01 5.04 ;
      RECT 57 4.607 57.005 5.04 ;
      RECT 56.99 3.505 57 3.705 ;
      RECT 56.995 4.622 57 5.04 ;
      RECT 56.955 4.68 56.995 5.04 ;
      RECT 56.985 3.504 56.99 3.69 ;
      RECT 56.98 3.502 56.985 3.683 ;
      RECT 56.97 3.499 56.98 3.673 ;
      RECT 56.965 3.496 56.97 3.658 ;
      RECT 56.95 3.492 56.965 3.651 ;
      RECT 56.945 4.735 56.955 5.04 ;
      RECT 56.945 3.489 56.95 3.646 ;
      RECT 56.93 3.485 56.945 3.64 ;
      RECT 56.94 4.752 56.945 5.04 ;
      RECT 56.93 4.815 56.94 5.04 ;
      RECT 56.85 3.47 56.93 3.62 ;
      RECT 56.925 4.822 56.93 5.035 ;
      RECT 56.92 4.83 56.925 5.025 ;
      RECT 56.84 3.456 56.85 3.604 ;
      RECT 56.825 3.452 56.84 3.602 ;
      RECT 56.815 3.447 56.825 3.598 ;
      RECT 56.79 3.44 56.815 3.59 ;
      RECT 56.785 3.435 56.79 3.585 ;
      RECT 56.775 3.435 56.785 3.583 ;
      RECT 56.765 3.433 56.775 3.581 ;
      RECT 56.735 3.425 56.765 3.575 ;
      RECT 56.72 3.417 56.735 3.568 ;
      RECT 56.7 3.412 56.72 3.561 ;
      RECT 56.695 3.408 56.7 3.556 ;
      RECT 56.665 3.401 56.695 3.55 ;
      RECT 56.64 3.392 56.665 3.54 ;
      RECT 56.61 3.385 56.64 3.532 ;
      RECT 56.585 3.375 56.61 3.523 ;
      RECT 56.57 3.367 56.585 3.517 ;
      RECT 56.545 3.362 56.57 3.512 ;
      RECT 56.535 3.358 56.545 3.507 ;
      RECT 56.515 3.353 56.535 3.502 ;
      RECT 56.48 3.348 56.515 3.495 ;
      RECT 56.42 3.343 56.48 3.488 ;
      RECT 56.407 3.339 56.42 3.486 ;
      RECT 56.321 3.334 56.407 3.483 ;
      RECT 56.235 3.324 56.321 3.479 ;
      RECT 56.194 3.317 56.235 3.476 ;
      RECT 56.108 3.31 56.194 3.473 ;
      RECT 56.022 3.3 56.108 3.469 ;
      RECT 55.936 3.29 56.022 3.464 ;
      RECT 55.85 3.28 55.936 3.46 ;
      RECT 55.84 3.265 55.85 3.458 ;
      RECT 55.83 3.25 55.84 3.458 ;
      RECT 55.765 3.245 55.83 3.457 ;
      RECT 55.6 3.242 55.645 3.45 ;
      RECT 56.845 4.147 56.85 4.338 ;
      RECT 56.84 4.142 56.845 4.345 ;
      RECT 56.826 4.14 56.84 4.351 ;
      RECT 56.74 4.14 56.826 4.353 ;
      RECT 56.736 4.14 56.74 4.356 ;
      RECT 56.65 4.14 56.736 4.374 ;
      RECT 56.64 4.145 56.65 4.393 ;
      RECT 56.63 4.2 56.64 4.397 ;
      RECT 56.605 4.215 56.63 4.404 ;
      RECT 56.565 4.235 56.605 4.417 ;
      RECT 56.56 4.247 56.565 4.427 ;
      RECT 56.545 4.253 56.56 4.432 ;
      RECT 56.54 4.258 56.545 4.436 ;
      RECT 56.52 4.265 56.54 4.441 ;
      RECT 56.45 4.29 56.52 4.458 ;
      RECT 56.41 4.318 56.45 4.478 ;
      RECT 56.405 4.328 56.41 4.486 ;
      RECT 56.385 4.335 56.405 4.488 ;
      RECT 56.38 4.342 56.385 4.491 ;
      RECT 56.35 4.35 56.38 4.494 ;
      RECT 56.345 4.355 56.35 4.498 ;
      RECT 56.271 4.359 56.345 4.506 ;
      RECT 56.185 4.368 56.271 4.522 ;
      RECT 56.181 4.373 56.185 4.531 ;
      RECT 56.095 4.378 56.181 4.541 ;
      RECT 56.055 4.386 56.095 4.553 ;
      RECT 56.005 4.392 56.055 4.56 ;
      RECT 55.92 4.401 56.005 4.575 ;
      RECT 55.845 4.412 55.92 4.593 ;
      RECT 55.81 4.419 55.845 4.603 ;
      RECT 55.735 4.427 55.81 4.608 ;
      RECT 55.68 4.436 55.735 4.608 ;
      RECT 55.655 4.441 55.68 4.606 ;
      RECT 55.645 4.444 55.655 4.604 ;
      RECT 55.61 4.446 55.645 4.602 ;
      RECT 55.58 4.448 55.61 4.598 ;
      RECT 55.535 4.447 55.58 4.594 ;
      RECT 55.515 4.442 55.535 4.591 ;
      RECT 55.465 4.427 55.515 4.588 ;
      RECT 55.455 4.412 55.465 4.583 ;
      RECT 55.405 4.397 55.455 4.573 ;
      RECT 55.355 4.372 55.405 4.553 ;
      RECT 55.345 4.357 55.355 4.535 ;
      RECT 55.34 4.355 55.345 4.529 ;
      RECT 55.32 4.35 55.34 4.524 ;
      RECT 55.315 4.342 55.32 4.518 ;
      RECT 55.3 4.336 55.315 4.511 ;
      RECT 55.295 4.331 55.3 4.503 ;
      RECT 55.275 4.326 55.295 4.495 ;
      RECT 55.26 4.319 55.275 4.488 ;
      RECT 55.245 4.313 55.26 4.479 ;
      RECT 55.24 4.307 55.245 4.472 ;
      RECT 55.195 4.282 55.24 4.458 ;
      RECT 55.18 4.252 55.195 4.44 ;
      RECT 55.165 4.235 55.18 4.431 ;
      RECT 55.14 4.215 55.165 4.419 ;
      RECT 55.1 4.185 55.14 4.399 ;
      RECT 55.09 4.155 55.1 4.384 ;
      RECT 55.075 4.145 55.09 4.377 ;
      RECT 55.02 4.11 55.075 4.356 ;
      RECT 55.005 4.073 55.02 4.335 ;
      RECT 54.995 4.06 55.005 4.327 ;
      RECT 54.945 4.03 54.995 4.309 ;
      RECT 54.93 3.96 54.945 4.29 ;
      RECT 54.885 3.96 54.93 4.273 ;
      RECT 54.86 3.96 54.885 4.255 ;
      RECT 54.85 3.96 54.86 4.248 ;
      RECT 54.771 3.96 54.85 4.241 ;
      RECT 54.685 3.96 54.771 4.233 ;
      RECT 54.67 3.992 54.685 4.228 ;
      RECT 54.595 4.002 54.67 4.224 ;
      RECT 54.575 4.012 54.595 4.219 ;
      RECT 54.55 4.012 54.575 4.216 ;
      RECT 54.54 4.002 54.55 4.215 ;
      RECT 54.53 3.975 54.54 4.214 ;
      RECT 54.49 3.97 54.53 4.212 ;
      RECT 54.445 3.97 54.49 4.208 ;
      RECT 54.42 3.97 54.445 4.203 ;
      RECT 54.37 3.97 54.42 4.19 ;
      RECT 54.33 3.975 54.34 4.175 ;
      RECT 54.34 3.97 54.37 4.18 ;
      RECT 56.325 3.75 56.585 4.01 ;
      RECT 56.32 3.772 56.585 3.968 ;
      RECT 55.56 3.6 55.78 3.965 ;
      RECT 55.542 3.687 55.78 3.964 ;
      RECT 55.525 3.692 55.78 3.961 ;
      RECT 55.525 3.692 55.8 3.96 ;
      RECT 55.495 3.702 55.8 3.958 ;
      RECT 55.49 3.717 55.8 3.954 ;
      RECT 55.49 3.717 55.805 3.953 ;
      RECT 55.485 3.775 55.805 3.951 ;
      RECT 55.485 3.775 55.815 3.948 ;
      RECT 55.48 3.84 55.815 3.943 ;
      RECT 55.56 3.6 55.82 3.86 ;
      RECT 54.305 3.43 54.565 3.69 ;
      RECT 54.305 3.473 54.651 3.664 ;
      RECT 54.305 3.473 54.695 3.663 ;
      RECT 54.305 3.473 54.715 3.661 ;
      RECT 54.305 3.473 54.815 3.66 ;
      RECT 54.305 3.473 54.835 3.658 ;
      RECT 54.305 3.473 54.845 3.653 ;
      RECT 54.715 3.44 54.905 3.65 ;
      RECT 54.715 3.442 54.91 3.648 ;
      RECT 54.705 3.447 54.915 3.64 ;
      RECT 54.651 3.471 54.915 3.64 ;
      RECT 54.695 3.465 54.705 3.662 ;
      RECT 54.705 3.445 54.91 3.648 ;
      RECT 53.66 4.505 53.865 4.735 ;
      RECT 53.6 4.455 53.655 4.715 ;
      RECT 53.66 4.455 53.86 4.735 ;
      RECT 54.63 4.77 54.635 4.797 ;
      RECT 54.62 4.68 54.63 4.802 ;
      RECT 54.615 4.602 54.62 4.808 ;
      RECT 54.605 4.592 54.615 4.815 ;
      RECT 54.6 4.582 54.605 4.821 ;
      RECT 54.59 4.577 54.6 4.823 ;
      RECT 54.575 4.569 54.59 4.831 ;
      RECT 54.56 4.56 54.575 4.843 ;
      RECT 54.55 4.552 54.56 4.853 ;
      RECT 54.515 4.47 54.55 4.871 ;
      RECT 54.48 4.47 54.515 4.89 ;
      RECT 54.465 4.47 54.48 4.898 ;
      RECT 54.41 4.47 54.465 4.898 ;
      RECT 54.376 4.47 54.41 4.889 ;
      RECT 54.29 4.47 54.376 4.865 ;
      RECT 54.28 4.53 54.29 4.847 ;
      RECT 54.24 4.532 54.28 4.838 ;
      RECT 54.235 4.534 54.24 4.828 ;
      RECT 54.215 4.536 54.235 4.823 ;
      RECT 54.205 4.539 54.215 4.818 ;
      RECT 54.195 4.54 54.205 4.813 ;
      RECT 54.171 4.541 54.195 4.805 ;
      RECT 54.085 4.546 54.171 4.783 ;
      RECT 54.03 4.545 54.085 4.756 ;
      RECT 54.015 4.538 54.03 4.743 ;
      RECT 53.98 4.533 54.015 4.739 ;
      RECT 53.925 4.525 53.98 4.738 ;
      RECT 53.865 4.512 53.925 4.736 ;
      RECT 53.655 4.455 53.66 4.723 ;
      RECT 53.73 3.825 53.915 4.035 ;
      RECT 53.72 3.83 53.93 4.028 ;
      RECT 53.76 3.735 54.02 3.995 ;
      RECT 53.715 3.892 54.02 3.918 ;
      RECT 53.06 3.685 53.065 4.485 ;
      RECT 53.005 3.735 53.035 4.485 ;
      RECT 52.995 3.735 53 4.045 ;
      RECT 52.98 3.735 52.985 4.04 ;
      RECT 52.525 3.78 52.54 3.995 ;
      RECT 52.455 3.78 52.54 3.99 ;
      RECT 53.72 3.36 53.79 3.57 ;
      RECT 53.79 3.367 53.8 3.565 ;
      RECT 53.686 3.36 53.72 3.577 ;
      RECT 53.6 3.36 53.686 3.601 ;
      RECT 53.59 3.365 53.6 3.62 ;
      RECT 53.585 3.377 53.59 3.623 ;
      RECT 53.57 3.392 53.585 3.627 ;
      RECT 53.565 3.41 53.57 3.631 ;
      RECT 53.525 3.42 53.565 3.64 ;
      RECT 53.51 3.427 53.525 3.652 ;
      RECT 53.495 3.432 53.51 3.657 ;
      RECT 53.48 3.435 53.495 3.662 ;
      RECT 53.47 3.437 53.48 3.666 ;
      RECT 53.435 3.444 53.47 3.674 ;
      RECT 53.4 3.452 53.435 3.688 ;
      RECT 53.39 3.458 53.4 3.697 ;
      RECT 53.385 3.46 53.39 3.699 ;
      RECT 53.365 3.463 53.385 3.705 ;
      RECT 53.335 3.47 53.365 3.716 ;
      RECT 53.325 3.476 53.335 3.723 ;
      RECT 53.3 3.479 53.325 3.73 ;
      RECT 53.29 3.483 53.3 3.738 ;
      RECT 53.285 3.484 53.29 3.76 ;
      RECT 53.28 3.485 53.285 3.775 ;
      RECT 53.275 3.486 53.28 3.79 ;
      RECT 53.27 3.487 53.275 3.805 ;
      RECT 53.265 3.488 53.27 3.835 ;
      RECT 53.255 3.49 53.265 3.868 ;
      RECT 53.24 3.494 53.255 3.915 ;
      RECT 53.23 3.497 53.24 3.96 ;
      RECT 53.225 3.5 53.23 3.988 ;
      RECT 53.215 3.502 53.225 4.015 ;
      RECT 53.21 3.505 53.215 4.05 ;
      RECT 53.18 3.51 53.21 4.108 ;
      RECT 53.175 3.515 53.18 4.193 ;
      RECT 53.17 3.517 53.175 4.228 ;
      RECT 53.165 3.519 53.17 4.31 ;
      RECT 53.16 3.521 53.165 4.398 ;
      RECT 53.15 3.523 53.16 4.48 ;
      RECT 53.135 3.537 53.15 4.485 ;
      RECT 53.1 3.582 53.135 4.485 ;
      RECT 53.09 3.622 53.1 4.485 ;
      RECT 53.075 3.65 53.09 4.485 ;
      RECT 53.07 3.667 53.075 4.485 ;
      RECT 53.065 3.675 53.07 4.485 ;
      RECT 53.055 3.69 53.06 4.485 ;
      RECT 53.05 3.697 53.055 4.485 ;
      RECT 53.04 3.717 53.05 4.485 ;
      RECT 53.035 3.73 53.04 4.485 ;
      RECT 53 3.735 53.005 4.07 ;
      RECT 52.985 4.125 53.005 4.485 ;
      RECT 52.985 3.735 52.995 4.043 ;
      RECT 52.98 4.165 52.985 4.485 ;
      RECT 52.93 3.735 52.98 4.038 ;
      RECT 52.975 4.202 52.98 4.485 ;
      RECT 52.965 4.225 52.975 4.485 ;
      RECT 52.96 4.27 52.965 4.485 ;
      RECT 52.95 4.28 52.96 4.478 ;
      RECT 52.876 3.735 52.93 4.032 ;
      RECT 52.79 3.735 52.876 4.025 ;
      RECT 52.741 3.782 52.79 4.018 ;
      RECT 52.655 3.79 52.741 4.011 ;
      RECT 52.64 3.787 52.655 4.006 ;
      RECT 52.626 3.78 52.64 4.005 ;
      RECT 52.54 3.78 52.626 4 ;
      RECT 52.445 3.785 52.455 3.985 ;
      RECT 52.035 3.215 52.05 3.615 ;
      RECT 52.23 3.215 52.235 3.475 ;
      RECT 51.975 3.215 52.02 3.475 ;
      RECT 52.43 4.52 52.435 4.725 ;
      RECT 52.425 4.51 52.43 4.73 ;
      RECT 52.42 4.497 52.425 4.735 ;
      RECT 52.415 4.477 52.42 4.735 ;
      RECT 52.39 4.43 52.415 4.735 ;
      RECT 52.355 4.345 52.39 4.735 ;
      RECT 52.35 4.282 52.355 4.735 ;
      RECT 52.345 4.267 52.35 4.735 ;
      RECT 52.33 4.227 52.345 4.735 ;
      RECT 52.325 4.202 52.33 4.735 ;
      RECT 52.315 4.185 52.325 4.735 ;
      RECT 52.28 4.107 52.315 4.735 ;
      RECT 52.275 4.05 52.28 4.735 ;
      RECT 52.27 4.037 52.275 4.735 ;
      RECT 52.26 4.015 52.27 4.735 ;
      RECT 52.25 3.98 52.26 4.735 ;
      RECT 52.24 3.95 52.25 4.735 ;
      RECT 52.23 3.865 52.24 4.378 ;
      RECT 52.237 4.51 52.24 4.735 ;
      RECT 52.235 4.52 52.237 4.735 ;
      RECT 52.225 4.53 52.235 4.73 ;
      RECT 52.22 3.215 52.23 3.61 ;
      RECT 52.225 3.742 52.23 4.353 ;
      RECT 52.22 3.64 52.225 4.336 ;
      RECT 52.21 3.215 52.22 4.312 ;
      RECT 52.205 3.215 52.21 4.283 ;
      RECT 52.2 3.215 52.205 4.273 ;
      RECT 52.18 3.215 52.2 4.235 ;
      RECT 52.175 3.215 52.18 4.193 ;
      RECT 52.17 3.215 52.175 4.173 ;
      RECT 52.14 3.215 52.17 4.123 ;
      RECT 52.13 3.215 52.14 4.07 ;
      RECT 52.125 3.215 52.13 4.043 ;
      RECT 52.12 3.215 52.125 4.028 ;
      RECT 52.11 3.215 52.12 4.005 ;
      RECT 52.1 3.215 52.11 3.98 ;
      RECT 52.095 3.215 52.1 3.92 ;
      RECT 52.085 3.215 52.095 3.858 ;
      RECT 52.08 3.215 52.085 3.778 ;
      RECT 52.075 3.215 52.08 3.743 ;
      RECT 52.07 3.215 52.075 3.718 ;
      RECT 52.065 3.215 52.07 3.703 ;
      RECT 52.06 3.215 52.065 3.673 ;
      RECT 52.055 3.215 52.06 3.65 ;
      RECT 52.05 3.215 52.055 3.623 ;
      RECT 52.02 3.215 52.035 3.61 ;
      RECT 51.175 4.75 51.36 4.96 ;
      RECT 51.165 4.755 51.375 4.953 ;
      RECT 51.165 4.755 51.395 4.925 ;
      RECT 51.165 4.755 51.41 4.904 ;
      RECT 51.165 4.755 51.425 4.902 ;
      RECT 51.165 4.755 51.435 4.901 ;
      RECT 51.165 4.755 51.465 4.898 ;
      RECT 51.815 4.6 52.075 4.86 ;
      RECT 51.775 4.647 52.075 4.843 ;
      RECT 51.766 4.655 51.775 4.846 ;
      RECT 51.36 4.748 52.075 4.843 ;
      RECT 51.68 4.673 51.766 4.853 ;
      RECT 51.375 4.745 52.075 4.843 ;
      RECT 51.621 4.695 51.68 4.865 ;
      RECT 51.395 4.741 52.075 4.843 ;
      RECT 51.535 4.707 51.621 4.876 ;
      RECT 51.41 4.737 52.075 4.843 ;
      RECT 51.48 4.72 51.535 4.888 ;
      RECT 51.425 4.735 52.075 4.843 ;
      RECT 51.465 4.726 51.48 4.894 ;
      RECT 51.435 4.731 52.075 4.843 ;
      RECT 51.58 4.255 51.84 4.515 ;
      RECT 51.58 4.275 51.95 4.485 ;
      RECT 51.58 4.28 51.96 4.48 ;
      RECT 51.771 3.694 51.85 3.925 ;
      RECT 51.685 3.697 51.9 3.92 ;
      RECT 51.68 3.697 51.9 3.915 ;
      RECT 51.68 3.702 51.91 3.913 ;
      RECT 51.655 3.702 51.91 3.91 ;
      RECT 51.655 3.71 51.92 3.908 ;
      RECT 51.535 3.645 51.795 3.905 ;
      RECT 51.535 3.692 51.845 3.905 ;
      RECT 50.79 4.265 50.795 4.525 ;
      RECT 50.62 4.035 50.625 4.525 ;
      RECT 50.505 4.275 50.51 4.5 ;
      RECT 51.215 3.37 51.22 3.58 ;
      RECT 51.22 3.375 51.235 3.575 ;
      RECT 51.155 3.37 51.215 3.588 ;
      RECT 51.14 3.37 51.155 3.598 ;
      RECT 51.09 3.37 51.14 3.615 ;
      RECT 51.07 3.37 51.09 3.638 ;
      RECT 51.055 3.37 51.07 3.65 ;
      RECT 51.035 3.37 51.055 3.66 ;
      RECT 51.025 3.375 51.035 3.669 ;
      RECT 51.02 3.385 51.025 3.674 ;
      RECT 51.015 3.397 51.02 3.678 ;
      RECT 51.005 3.42 51.015 3.683 ;
      RECT 51 3.435 51.005 3.687 ;
      RECT 50.995 3.452 51 3.69 ;
      RECT 50.99 3.46 50.995 3.693 ;
      RECT 50.98 3.465 50.99 3.697 ;
      RECT 50.975 3.472 50.98 3.702 ;
      RECT 50.965 3.477 50.975 3.706 ;
      RECT 50.94 3.489 50.965 3.717 ;
      RECT 50.92 3.506 50.94 3.733 ;
      RECT 50.895 3.523 50.92 3.755 ;
      RECT 50.86 3.546 50.895 3.813 ;
      RECT 50.84 3.568 50.86 3.875 ;
      RECT 50.835 3.578 50.84 3.91 ;
      RECT 50.825 3.585 50.835 3.948 ;
      RECT 50.82 3.592 50.825 3.968 ;
      RECT 50.815 3.603 50.82 4.005 ;
      RECT 50.81 3.611 50.815 4.07 ;
      RECT 50.8 3.622 50.81 4.123 ;
      RECT 50.795 3.64 50.8 4.193 ;
      RECT 50.79 3.65 50.795 4.23 ;
      RECT 50.785 3.66 50.79 4.525 ;
      RECT 50.78 3.672 50.785 4.525 ;
      RECT 50.775 3.682 50.78 4.525 ;
      RECT 50.765 3.692 50.775 4.525 ;
      RECT 50.755 3.715 50.765 4.525 ;
      RECT 50.74 3.75 50.755 4.525 ;
      RECT 50.7 3.812 50.74 4.525 ;
      RECT 50.695 3.865 50.7 4.525 ;
      RECT 50.67 3.9 50.695 4.525 ;
      RECT 50.655 3.945 50.67 4.525 ;
      RECT 50.65 3.967 50.655 4.525 ;
      RECT 50.64 3.98 50.65 4.525 ;
      RECT 50.63 4.005 50.64 4.525 ;
      RECT 50.625 4.027 50.63 4.525 ;
      RECT 50.6 4.065 50.62 4.525 ;
      RECT 50.56 4.122 50.6 4.525 ;
      RECT 50.555 4.172 50.56 4.525 ;
      RECT 50.55 4.19 50.555 4.525 ;
      RECT 50.545 4.202 50.55 4.525 ;
      RECT 50.535 4.22 50.545 4.525 ;
      RECT 50.525 4.24 50.535 4.5 ;
      RECT 50.52 4.257 50.525 4.5 ;
      RECT 50.51 4.27 50.52 4.5 ;
      RECT 50.48 4.28 50.505 4.5 ;
      RECT 50.47 4.287 50.48 4.5 ;
      RECT 50.455 4.297 50.47 4.495 ;
      RECT 49.545 10.055 49.835 10.285 ;
      RECT 49.605 8.575 49.775 10.285 ;
      RECT 49.555 8.94 49.905 9.29 ;
      RECT 49.545 8.575 49.835 8.805 ;
      RECT 49.14 3.69 49.245 4.26 ;
      RECT 49.14 4.025 49.465 4.255 ;
      RECT 49.14 4.055 49.635 4.225 ;
      RECT 49.14 3.69 49.33 4.255 ;
      RECT 48.555 3.655 48.845 3.885 ;
      RECT 48.555 3.69 49.33 3.86 ;
      RECT 48.615 2.175 48.785 3.885 ;
      RECT 48.555 2.175 48.845 2.405 ;
      RECT 48.555 10.055 48.845 10.285 ;
      RECT 48.615 8.575 48.785 10.285 ;
      RECT 48.555 8.575 48.845 8.805 ;
      RECT 48.555 8.61 49.41 8.77 ;
      RECT 49.24 8.205 49.41 8.77 ;
      RECT 48.555 8.605 48.95 8.77 ;
      RECT 49.175 8.205 49.465 8.435 ;
      RECT 49.175 8.235 49.635 8.405 ;
      RECT 48.185 4.025 48.475 4.255 ;
      RECT 48.185 4.055 48.645 4.225 ;
      RECT 48.25 2.95 48.415 4.255 ;
      RECT 46.765 2.92 47.055 3.15 ;
      RECT 46.765 2.95 48.415 3.12 ;
      RECT 46.825 2.18 46.995 3.15 ;
      RECT 46.765 2.18 47.055 2.41 ;
      RECT 46.765 10.05 47.055 10.28 ;
      RECT 46.825 9.31 46.995 10.28 ;
      RECT 46.825 9.405 48.415 9.575 ;
      RECT 48.245 8.205 48.415 9.575 ;
      RECT 46.765 9.31 47.055 9.54 ;
      RECT 48.185 8.205 48.475 8.435 ;
      RECT 48.185 8.235 48.645 8.405 ;
      RECT 47.195 3.26 47.545 3.61 ;
      RECT 44.86 3.32 47.545 3.49 ;
      RECT 44.86 2.635 45.03 3.49 ;
      RECT 44.76 2.635 45.11 2.985 ;
      RECT 47.22 8.94 47.545 9.265 ;
      RECT 42.65 8.9 43 9.25 ;
      RECT 47.195 8.94 47.545 9.17 ;
      RECT 42.415 8.94 43 9.17 ;
      RECT 42.245 8.97 47.545 9.14 ;
      RECT 46.42 3.66 46.74 3.98 ;
      RECT 46.39 3.66 46.74 3.89 ;
      RECT 46.22 3.69 46.74 3.86 ;
      RECT 46.42 8.54 46.74 8.83 ;
      RECT 46.39 8.57 46.74 8.8 ;
      RECT 46.22 8.6 46.74 8.77 ;
      RECT 43.055 3.76 43.24 3.97 ;
      RECT 43.045 3.765 43.255 3.963 ;
      RECT 43.045 3.765 43.341 3.94 ;
      RECT 43.045 3.765 43.4 3.915 ;
      RECT 43.045 3.765 43.455 3.895 ;
      RECT 43.045 3.765 43.465 3.883 ;
      RECT 43.045 3.765 43.66 3.822 ;
      RECT 43.045 3.765 43.69 3.805 ;
      RECT 43.045 3.765 43.71 3.795 ;
      RECT 43.59 3.53 43.85 3.79 ;
      RECT 43.575 3.62 43.59 3.837 ;
      RECT 43.11 3.752 43.85 3.79 ;
      RECT 43.561 3.631 43.575 3.843 ;
      RECT 43.15 3.745 43.85 3.79 ;
      RECT 43.475 3.671 43.561 3.862 ;
      RECT 43.4 3.732 43.85 3.79 ;
      RECT 43.47 3.707 43.475 3.879 ;
      RECT 43.455 3.717 43.85 3.79 ;
      RECT 43.465 3.712 43.47 3.881 ;
      RECT 43.76 4.217 43.765 4.309 ;
      RECT 43.755 4.195 43.76 4.326 ;
      RECT 43.75 4.185 43.755 4.338 ;
      RECT 43.74 4.176 43.75 4.348 ;
      RECT 43.735 4.171 43.74 4.356 ;
      RECT 43.73 4.03 43.735 4.359 ;
      RECT 43.696 4.03 43.73 4.37 ;
      RECT 43.61 4.03 43.696 4.405 ;
      RECT 43.53 4.03 43.61 4.453 ;
      RECT 43.501 4.03 43.53 4.477 ;
      RECT 43.415 4.03 43.501 4.483 ;
      RECT 43.41 4.214 43.415 4.488 ;
      RECT 43.375 4.225 43.41 4.491 ;
      RECT 43.35 4.24 43.375 4.495 ;
      RECT 43.336 4.249 43.35 4.497 ;
      RECT 43.25 4.276 43.336 4.503 ;
      RECT 43.185 4.317 43.25 4.512 ;
      RECT 43.17 4.337 43.185 4.517 ;
      RECT 43.14 4.347 43.17 4.52 ;
      RECT 43.135 4.357 43.14 4.523 ;
      RECT 43.105 4.362 43.135 4.525 ;
      RECT 43.085 4.367 43.105 4.529 ;
      RECT 43 4.37 43.085 4.536 ;
      RECT 42.985 4.367 43 4.542 ;
      RECT 42.975 4.364 42.985 4.544 ;
      RECT 42.955 4.361 42.975 4.546 ;
      RECT 42.935 4.357 42.955 4.547 ;
      RECT 42.92 4.353 42.935 4.549 ;
      RECT 42.91 4.35 42.92 4.55 ;
      RECT 42.87 4.344 42.91 4.548 ;
      RECT 42.86 4.339 42.87 4.546 ;
      RECT 42.845 4.336 42.86 4.542 ;
      RECT 42.82 4.331 42.845 4.535 ;
      RECT 42.77 4.322 42.82 4.523 ;
      RECT 42.7 4.308 42.77 4.505 ;
      RECT 42.642 4.293 42.7 4.487 ;
      RECT 42.556 4.276 42.642 4.467 ;
      RECT 42.47 4.255 42.556 4.442 ;
      RECT 42.42 4.24 42.47 4.423 ;
      RECT 42.416 4.234 42.42 4.415 ;
      RECT 42.33 4.224 42.416 4.402 ;
      RECT 42.295 4.209 42.33 4.385 ;
      RECT 42.28 4.202 42.295 4.378 ;
      RECT 42.22 4.19 42.28 4.366 ;
      RECT 42.2 4.177 42.22 4.354 ;
      RECT 42.16 4.168 42.2 4.346 ;
      RECT 42.155 4.16 42.16 4.339 ;
      RECT 42.075 4.15 42.155 4.325 ;
      RECT 42.06 4.137 42.075 4.31 ;
      RECT 42.055 4.135 42.06 4.308 ;
      RECT 41.976 4.123 42.055 4.295 ;
      RECT 41.89 4.098 41.976 4.27 ;
      RECT 41.875 4.067 41.89 4.255 ;
      RECT 41.86 4.042 41.875 4.251 ;
      RECT 41.845 4.035 41.86 4.247 ;
      RECT 41.67 4.04 41.675 4.243 ;
      RECT 41.665 4.045 41.67 4.238 ;
      RECT 41.675 4.035 41.845 4.245 ;
      RECT 42.39 3.795 42.495 4.055 ;
      RECT 43.205 3.32 43.21 3.545 ;
      RECT 43.335 3.32 43.39 3.53 ;
      RECT 43.39 3.325 43.4 3.523 ;
      RECT 43.296 3.32 43.335 3.533 ;
      RECT 43.21 3.32 43.296 3.54 ;
      RECT 43.19 3.325 43.205 3.546 ;
      RECT 43.18 3.365 43.19 3.548 ;
      RECT 43.15 3.375 43.18 3.55 ;
      RECT 43.145 3.38 43.15 3.552 ;
      RECT 43.12 3.385 43.145 3.554 ;
      RECT 43.105 3.39 43.12 3.556 ;
      RECT 43.09 3.392 43.105 3.558 ;
      RECT 43.085 3.397 43.09 3.56 ;
      RECT 43.035 3.405 43.085 3.563 ;
      RECT 43.01 3.414 43.035 3.568 ;
      RECT 43 3.421 43.01 3.573 ;
      RECT 42.995 3.424 43 3.577 ;
      RECT 42.975 3.427 42.995 3.586 ;
      RECT 42.945 3.435 42.975 3.606 ;
      RECT 42.916 3.448 42.945 3.628 ;
      RECT 42.83 3.482 42.916 3.672 ;
      RECT 42.825 3.508 42.83 3.71 ;
      RECT 42.82 3.512 42.825 3.719 ;
      RECT 42.785 3.525 42.82 3.752 ;
      RECT 42.775 3.539 42.785 3.79 ;
      RECT 42.77 3.543 42.775 3.803 ;
      RECT 42.765 3.547 42.77 3.808 ;
      RECT 42.755 3.555 42.765 3.82 ;
      RECT 42.75 3.562 42.755 3.835 ;
      RECT 42.725 3.575 42.75 3.86 ;
      RECT 42.685 3.604 42.725 3.915 ;
      RECT 42.67 3.629 42.685 3.97 ;
      RECT 42.66 3.64 42.67 3.993 ;
      RECT 42.655 3.647 42.66 4.005 ;
      RECT 42.65 3.651 42.655 4.013 ;
      RECT 42.595 3.679 42.65 4.055 ;
      RECT 42.575 3.715 42.595 4.055 ;
      RECT 42.56 3.73 42.575 4.055 ;
      RECT 42.505 3.762 42.56 4.055 ;
      RECT 42.495 3.792 42.505 4.055 ;
      RECT 42.105 3.407 42.29 3.645 ;
      RECT 42.09 3.409 42.3 3.64 ;
      RECT 41.975 3.355 42.235 3.615 ;
      RECT 41.97 3.392 42.235 3.569 ;
      RECT 41.965 3.402 42.235 3.566 ;
      RECT 41.96 3.442 42.3 3.56 ;
      RECT 41.955 3.475 42.3 3.55 ;
      RECT 41.965 3.417 42.315 3.488 ;
      RECT 42.262 4.515 42.275 5.045 ;
      RECT 42.176 4.515 42.275 5.044 ;
      RECT 42.176 4.515 42.28 5.043 ;
      RECT 42.09 4.515 42.28 5.041 ;
      RECT 42.085 4.515 42.28 5.038 ;
      RECT 42.085 4.515 42.29 5.036 ;
      RECT 42.08 4.807 42.29 5.033 ;
      RECT 42.08 4.817 42.295 5.03 ;
      RECT 42.08 4.885 42.3 5.026 ;
      RECT 42.07 4.89 42.3 5.025 ;
      RECT 42.07 4.982 42.305 5.022 ;
      RECT 42.055 4.515 42.315 4.775 ;
      RECT 41.985 10.05 42.275 10.28 ;
      RECT 42.045 9.31 42.215 10.28 ;
      RECT 41.96 9.34 42.3 9.685 ;
      RECT 41.985 9.31 42.275 9.685 ;
      RECT 41.285 3.505 41.33 5.04 ;
      RECT 41.485 3.505 41.515 3.72 ;
      RECT 39.86 3.245 39.98 3.455 ;
      RECT 39.52 3.195 39.78 3.455 ;
      RECT 39.52 3.24 39.815 3.445 ;
      RECT 41.525 3.521 41.53 3.575 ;
      RECT 41.52 3.514 41.525 3.708 ;
      RECT 41.515 3.508 41.52 3.715 ;
      RECT 41.47 3.505 41.485 3.728 ;
      RECT 41.465 3.505 41.47 3.75 ;
      RECT 41.46 3.505 41.465 3.798 ;
      RECT 41.455 3.505 41.46 3.818 ;
      RECT 41.445 3.505 41.455 3.925 ;
      RECT 41.44 3.505 41.445 3.988 ;
      RECT 41.435 3.505 41.44 4.045 ;
      RECT 41.43 3.505 41.435 4.053 ;
      RECT 41.415 3.505 41.43 4.16 ;
      RECT 41.405 3.505 41.415 4.295 ;
      RECT 41.395 3.505 41.405 4.405 ;
      RECT 41.385 3.505 41.395 4.462 ;
      RECT 41.38 3.505 41.385 4.502 ;
      RECT 41.375 3.505 41.38 4.538 ;
      RECT 41.365 3.505 41.375 4.578 ;
      RECT 41.36 3.505 41.365 4.62 ;
      RECT 41.34 3.505 41.36 4.685 ;
      RECT 41.345 4.83 41.35 5.01 ;
      RECT 41.34 4.812 41.345 5.018 ;
      RECT 41.335 3.505 41.34 4.748 ;
      RECT 41.335 4.792 41.34 5.025 ;
      RECT 41.33 3.505 41.335 5.035 ;
      RECT 41.275 3.505 41.285 3.805 ;
      RECT 41.28 4.052 41.285 5.04 ;
      RECT 41.275 4.117 41.28 5.04 ;
      RECT 41.27 3.506 41.275 3.795 ;
      RECT 41.265 4.182 41.275 5.04 ;
      RECT 41.26 3.507 41.27 3.785 ;
      RECT 41.25 4.295 41.265 5.04 ;
      RECT 41.255 3.508 41.26 3.775 ;
      RECT 41.235 3.509 41.255 3.753 ;
      RECT 41.24 4.392 41.25 5.04 ;
      RECT 41.235 4.467 41.24 5.04 ;
      RECT 41.225 3.508 41.235 3.73 ;
      RECT 41.23 4.51 41.235 5.04 ;
      RECT 41.225 4.537 41.23 5.04 ;
      RECT 41.215 3.506 41.225 3.718 ;
      RECT 41.22 4.58 41.225 5.04 ;
      RECT 41.215 4.607 41.22 5.04 ;
      RECT 41.205 3.505 41.215 3.705 ;
      RECT 41.21 4.622 41.215 5.04 ;
      RECT 41.17 4.68 41.21 5.04 ;
      RECT 41.2 3.504 41.205 3.69 ;
      RECT 41.195 3.502 41.2 3.683 ;
      RECT 41.185 3.499 41.195 3.673 ;
      RECT 41.18 3.496 41.185 3.658 ;
      RECT 41.165 3.492 41.18 3.651 ;
      RECT 41.16 4.735 41.17 5.04 ;
      RECT 41.16 3.489 41.165 3.646 ;
      RECT 41.145 3.485 41.16 3.64 ;
      RECT 41.155 4.752 41.16 5.04 ;
      RECT 41.145 4.815 41.155 5.04 ;
      RECT 41.065 3.47 41.145 3.62 ;
      RECT 41.14 4.822 41.145 5.035 ;
      RECT 41.135 4.83 41.14 5.025 ;
      RECT 41.055 3.456 41.065 3.604 ;
      RECT 41.04 3.452 41.055 3.602 ;
      RECT 41.03 3.447 41.04 3.598 ;
      RECT 41.005 3.44 41.03 3.59 ;
      RECT 41 3.435 41.005 3.585 ;
      RECT 40.99 3.435 41 3.583 ;
      RECT 40.98 3.433 40.99 3.581 ;
      RECT 40.95 3.425 40.98 3.575 ;
      RECT 40.935 3.417 40.95 3.568 ;
      RECT 40.915 3.412 40.935 3.561 ;
      RECT 40.91 3.408 40.915 3.556 ;
      RECT 40.88 3.401 40.91 3.55 ;
      RECT 40.855 3.392 40.88 3.54 ;
      RECT 40.825 3.385 40.855 3.532 ;
      RECT 40.8 3.375 40.825 3.523 ;
      RECT 40.785 3.367 40.8 3.517 ;
      RECT 40.76 3.362 40.785 3.512 ;
      RECT 40.75 3.358 40.76 3.507 ;
      RECT 40.73 3.353 40.75 3.502 ;
      RECT 40.695 3.348 40.73 3.495 ;
      RECT 40.635 3.343 40.695 3.488 ;
      RECT 40.622 3.339 40.635 3.486 ;
      RECT 40.536 3.334 40.622 3.483 ;
      RECT 40.45 3.324 40.536 3.479 ;
      RECT 40.409 3.317 40.45 3.476 ;
      RECT 40.323 3.31 40.409 3.473 ;
      RECT 40.237 3.3 40.323 3.469 ;
      RECT 40.151 3.29 40.237 3.464 ;
      RECT 40.065 3.28 40.151 3.46 ;
      RECT 40.055 3.265 40.065 3.458 ;
      RECT 40.045 3.25 40.055 3.458 ;
      RECT 39.98 3.245 40.045 3.457 ;
      RECT 39.815 3.242 39.86 3.45 ;
      RECT 41.06 4.147 41.065 4.338 ;
      RECT 41.055 4.142 41.06 4.345 ;
      RECT 41.041 4.14 41.055 4.351 ;
      RECT 40.955 4.14 41.041 4.353 ;
      RECT 40.951 4.14 40.955 4.356 ;
      RECT 40.865 4.14 40.951 4.374 ;
      RECT 40.855 4.145 40.865 4.393 ;
      RECT 40.845 4.2 40.855 4.397 ;
      RECT 40.82 4.215 40.845 4.404 ;
      RECT 40.78 4.235 40.82 4.417 ;
      RECT 40.775 4.247 40.78 4.427 ;
      RECT 40.76 4.253 40.775 4.432 ;
      RECT 40.755 4.258 40.76 4.436 ;
      RECT 40.735 4.265 40.755 4.441 ;
      RECT 40.665 4.29 40.735 4.458 ;
      RECT 40.625 4.318 40.665 4.478 ;
      RECT 40.62 4.328 40.625 4.486 ;
      RECT 40.6 4.335 40.62 4.488 ;
      RECT 40.595 4.342 40.6 4.491 ;
      RECT 40.565 4.35 40.595 4.494 ;
      RECT 40.56 4.355 40.565 4.498 ;
      RECT 40.486 4.359 40.56 4.506 ;
      RECT 40.4 4.368 40.486 4.522 ;
      RECT 40.396 4.373 40.4 4.531 ;
      RECT 40.31 4.378 40.396 4.541 ;
      RECT 40.27 4.386 40.31 4.553 ;
      RECT 40.22 4.392 40.27 4.56 ;
      RECT 40.135 4.401 40.22 4.575 ;
      RECT 40.06 4.412 40.135 4.593 ;
      RECT 40.025 4.419 40.06 4.603 ;
      RECT 39.95 4.427 40.025 4.608 ;
      RECT 39.895 4.436 39.95 4.608 ;
      RECT 39.87 4.441 39.895 4.606 ;
      RECT 39.86 4.444 39.87 4.604 ;
      RECT 39.825 4.446 39.86 4.602 ;
      RECT 39.795 4.448 39.825 4.598 ;
      RECT 39.75 4.447 39.795 4.594 ;
      RECT 39.73 4.442 39.75 4.591 ;
      RECT 39.68 4.427 39.73 4.588 ;
      RECT 39.67 4.412 39.68 4.583 ;
      RECT 39.62 4.397 39.67 4.573 ;
      RECT 39.57 4.372 39.62 4.553 ;
      RECT 39.56 4.357 39.57 4.535 ;
      RECT 39.555 4.355 39.56 4.529 ;
      RECT 39.535 4.35 39.555 4.524 ;
      RECT 39.53 4.342 39.535 4.518 ;
      RECT 39.515 4.336 39.53 4.511 ;
      RECT 39.51 4.331 39.515 4.503 ;
      RECT 39.49 4.326 39.51 4.495 ;
      RECT 39.475 4.319 39.49 4.488 ;
      RECT 39.46 4.313 39.475 4.479 ;
      RECT 39.455 4.307 39.46 4.472 ;
      RECT 39.41 4.282 39.455 4.458 ;
      RECT 39.395 4.252 39.41 4.44 ;
      RECT 39.38 4.235 39.395 4.431 ;
      RECT 39.355 4.215 39.38 4.419 ;
      RECT 39.315 4.185 39.355 4.399 ;
      RECT 39.305 4.155 39.315 4.384 ;
      RECT 39.29 4.145 39.305 4.377 ;
      RECT 39.235 4.11 39.29 4.356 ;
      RECT 39.22 4.073 39.235 4.335 ;
      RECT 39.21 4.06 39.22 4.327 ;
      RECT 39.16 4.03 39.21 4.309 ;
      RECT 39.145 3.96 39.16 4.29 ;
      RECT 39.1 3.96 39.145 4.273 ;
      RECT 39.075 3.96 39.1 4.255 ;
      RECT 39.065 3.96 39.075 4.248 ;
      RECT 38.986 3.96 39.065 4.241 ;
      RECT 38.9 3.96 38.986 4.233 ;
      RECT 38.885 3.992 38.9 4.228 ;
      RECT 38.81 4.002 38.885 4.224 ;
      RECT 38.79 4.012 38.81 4.219 ;
      RECT 38.765 4.012 38.79 4.216 ;
      RECT 38.755 4.002 38.765 4.215 ;
      RECT 38.745 3.975 38.755 4.214 ;
      RECT 38.705 3.97 38.745 4.212 ;
      RECT 38.66 3.97 38.705 4.208 ;
      RECT 38.635 3.97 38.66 4.203 ;
      RECT 38.585 3.97 38.635 4.19 ;
      RECT 38.545 3.975 38.555 4.175 ;
      RECT 38.555 3.97 38.585 4.18 ;
      RECT 40.54 3.75 40.8 4.01 ;
      RECT 40.535 3.772 40.8 3.968 ;
      RECT 39.775 3.6 39.995 3.965 ;
      RECT 39.757 3.687 39.995 3.964 ;
      RECT 39.74 3.692 39.995 3.961 ;
      RECT 39.74 3.692 40.015 3.96 ;
      RECT 39.71 3.702 40.015 3.958 ;
      RECT 39.705 3.717 40.015 3.954 ;
      RECT 39.705 3.717 40.02 3.953 ;
      RECT 39.7 3.775 40.02 3.951 ;
      RECT 39.7 3.775 40.03 3.948 ;
      RECT 39.695 3.84 40.03 3.943 ;
      RECT 39.775 3.6 40.035 3.86 ;
      RECT 38.52 3.43 38.78 3.69 ;
      RECT 38.52 3.473 38.866 3.664 ;
      RECT 38.52 3.473 38.91 3.663 ;
      RECT 38.52 3.473 38.93 3.661 ;
      RECT 38.52 3.473 39.03 3.66 ;
      RECT 38.52 3.473 39.05 3.658 ;
      RECT 38.52 3.473 39.06 3.653 ;
      RECT 38.93 3.44 39.12 3.65 ;
      RECT 38.93 3.442 39.125 3.648 ;
      RECT 38.92 3.447 39.13 3.64 ;
      RECT 38.866 3.471 39.13 3.64 ;
      RECT 38.91 3.465 38.92 3.662 ;
      RECT 38.92 3.445 39.125 3.648 ;
      RECT 37.875 4.505 38.08 4.735 ;
      RECT 37.815 4.455 37.87 4.715 ;
      RECT 37.875 4.455 38.075 4.735 ;
      RECT 38.845 4.77 38.85 4.797 ;
      RECT 38.835 4.68 38.845 4.802 ;
      RECT 38.83 4.602 38.835 4.808 ;
      RECT 38.82 4.592 38.83 4.815 ;
      RECT 38.815 4.582 38.82 4.821 ;
      RECT 38.805 4.577 38.815 4.823 ;
      RECT 38.79 4.569 38.805 4.831 ;
      RECT 38.775 4.56 38.79 4.843 ;
      RECT 38.765 4.552 38.775 4.853 ;
      RECT 38.73 4.47 38.765 4.871 ;
      RECT 38.695 4.47 38.73 4.89 ;
      RECT 38.68 4.47 38.695 4.898 ;
      RECT 38.625 4.47 38.68 4.898 ;
      RECT 38.591 4.47 38.625 4.889 ;
      RECT 38.505 4.47 38.591 4.865 ;
      RECT 38.495 4.53 38.505 4.847 ;
      RECT 38.455 4.532 38.495 4.838 ;
      RECT 38.45 4.534 38.455 4.828 ;
      RECT 38.43 4.536 38.45 4.823 ;
      RECT 38.42 4.539 38.43 4.818 ;
      RECT 38.41 4.54 38.42 4.813 ;
      RECT 38.386 4.541 38.41 4.805 ;
      RECT 38.3 4.546 38.386 4.783 ;
      RECT 38.245 4.545 38.3 4.756 ;
      RECT 38.23 4.538 38.245 4.743 ;
      RECT 38.195 4.533 38.23 4.739 ;
      RECT 38.14 4.525 38.195 4.738 ;
      RECT 38.08 4.512 38.14 4.736 ;
      RECT 37.87 4.455 37.875 4.723 ;
      RECT 37.945 3.825 38.13 4.035 ;
      RECT 37.935 3.83 38.145 4.028 ;
      RECT 37.975 3.735 38.235 3.995 ;
      RECT 37.93 3.892 38.235 3.918 ;
      RECT 37.275 3.685 37.28 4.485 ;
      RECT 37.22 3.735 37.25 4.485 ;
      RECT 37.21 3.735 37.215 4.045 ;
      RECT 37.195 3.735 37.2 4.04 ;
      RECT 36.74 3.78 36.755 3.995 ;
      RECT 36.67 3.78 36.755 3.99 ;
      RECT 37.935 3.36 38.005 3.57 ;
      RECT 38.005 3.367 38.015 3.565 ;
      RECT 37.901 3.36 37.935 3.577 ;
      RECT 37.815 3.36 37.901 3.601 ;
      RECT 37.805 3.365 37.815 3.62 ;
      RECT 37.8 3.377 37.805 3.623 ;
      RECT 37.785 3.392 37.8 3.627 ;
      RECT 37.78 3.41 37.785 3.631 ;
      RECT 37.74 3.42 37.78 3.64 ;
      RECT 37.725 3.427 37.74 3.652 ;
      RECT 37.71 3.432 37.725 3.657 ;
      RECT 37.695 3.435 37.71 3.662 ;
      RECT 37.685 3.437 37.695 3.666 ;
      RECT 37.65 3.444 37.685 3.674 ;
      RECT 37.615 3.452 37.65 3.688 ;
      RECT 37.605 3.458 37.615 3.697 ;
      RECT 37.6 3.46 37.605 3.699 ;
      RECT 37.58 3.463 37.6 3.705 ;
      RECT 37.55 3.47 37.58 3.716 ;
      RECT 37.54 3.476 37.55 3.723 ;
      RECT 37.515 3.479 37.54 3.73 ;
      RECT 37.505 3.483 37.515 3.738 ;
      RECT 37.5 3.484 37.505 3.76 ;
      RECT 37.495 3.485 37.5 3.775 ;
      RECT 37.49 3.486 37.495 3.79 ;
      RECT 37.485 3.487 37.49 3.805 ;
      RECT 37.48 3.488 37.485 3.835 ;
      RECT 37.47 3.49 37.48 3.868 ;
      RECT 37.455 3.494 37.47 3.915 ;
      RECT 37.445 3.497 37.455 3.96 ;
      RECT 37.44 3.5 37.445 3.988 ;
      RECT 37.43 3.502 37.44 4.015 ;
      RECT 37.425 3.505 37.43 4.05 ;
      RECT 37.395 3.51 37.425 4.108 ;
      RECT 37.39 3.515 37.395 4.193 ;
      RECT 37.385 3.517 37.39 4.228 ;
      RECT 37.38 3.519 37.385 4.31 ;
      RECT 37.375 3.521 37.38 4.398 ;
      RECT 37.365 3.523 37.375 4.48 ;
      RECT 37.35 3.537 37.365 4.485 ;
      RECT 37.315 3.582 37.35 4.485 ;
      RECT 37.305 3.622 37.315 4.485 ;
      RECT 37.29 3.65 37.305 4.485 ;
      RECT 37.285 3.667 37.29 4.485 ;
      RECT 37.28 3.675 37.285 4.485 ;
      RECT 37.27 3.69 37.275 4.485 ;
      RECT 37.265 3.697 37.27 4.485 ;
      RECT 37.255 3.717 37.265 4.485 ;
      RECT 37.25 3.73 37.255 4.485 ;
      RECT 37.215 3.735 37.22 4.07 ;
      RECT 37.2 4.125 37.22 4.485 ;
      RECT 37.2 3.735 37.21 4.043 ;
      RECT 37.195 4.165 37.2 4.485 ;
      RECT 37.145 3.735 37.195 4.038 ;
      RECT 37.19 4.202 37.195 4.485 ;
      RECT 37.18 4.225 37.19 4.485 ;
      RECT 37.175 4.27 37.18 4.485 ;
      RECT 37.165 4.28 37.175 4.478 ;
      RECT 37.091 3.735 37.145 4.032 ;
      RECT 37.005 3.735 37.091 4.025 ;
      RECT 36.956 3.782 37.005 4.018 ;
      RECT 36.87 3.79 36.956 4.011 ;
      RECT 36.855 3.787 36.87 4.006 ;
      RECT 36.841 3.78 36.855 4.005 ;
      RECT 36.755 3.78 36.841 4 ;
      RECT 36.66 3.785 36.67 3.985 ;
      RECT 36.25 3.215 36.265 3.615 ;
      RECT 36.445 3.215 36.45 3.475 ;
      RECT 36.19 3.215 36.235 3.475 ;
      RECT 36.645 4.52 36.65 4.725 ;
      RECT 36.64 4.51 36.645 4.73 ;
      RECT 36.635 4.497 36.64 4.735 ;
      RECT 36.63 4.477 36.635 4.735 ;
      RECT 36.605 4.43 36.63 4.735 ;
      RECT 36.57 4.345 36.605 4.735 ;
      RECT 36.565 4.282 36.57 4.735 ;
      RECT 36.56 4.267 36.565 4.735 ;
      RECT 36.545 4.227 36.56 4.735 ;
      RECT 36.54 4.202 36.545 4.735 ;
      RECT 36.53 4.185 36.54 4.735 ;
      RECT 36.495 4.107 36.53 4.735 ;
      RECT 36.49 4.05 36.495 4.735 ;
      RECT 36.485 4.037 36.49 4.735 ;
      RECT 36.475 4.015 36.485 4.735 ;
      RECT 36.465 3.98 36.475 4.735 ;
      RECT 36.455 3.95 36.465 4.735 ;
      RECT 36.445 3.865 36.455 4.378 ;
      RECT 36.452 4.51 36.455 4.735 ;
      RECT 36.45 4.52 36.452 4.735 ;
      RECT 36.44 4.53 36.45 4.73 ;
      RECT 36.435 3.215 36.445 3.61 ;
      RECT 36.44 3.742 36.445 4.353 ;
      RECT 36.435 3.64 36.44 4.336 ;
      RECT 36.425 3.215 36.435 4.312 ;
      RECT 36.42 3.215 36.425 4.283 ;
      RECT 36.415 3.215 36.42 4.273 ;
      RECT 36.395 3.215 36.415 4.235 ;
      RECT 36.39 3.215 36.395 4.193 ;
      RECT 36.385 3.215 36.39 4.173 ;
      RECT 36.355 3.215 36.385 4.123 ;
      RECT 36.345 3.215 36.355 4.07 ;
      RECT 36.34 3.215 36.345 4.043 ;
      RECT 36.335 3.215 36.34 4.028 ;
      RECT 36.325 3.215 36.335 4.005 ;
      RECT 36.315 3.215 36.325 3.98 ;
      RECT 36.31 3.215 36.315 3.92 ;
      RECT 36.3 3.215 36.31 3.858 ;
      RECT 36.295 3.215 36.3 3.778 ;
      RECT 36.29 3.215 36.295 3.743 ;
      RECT 36.285 3.215 36.29 3.718 ;
      RECT 36.28 3.215 36.285 3.703 ;
      RECT 36.275 3.215 36.28 3.673 ;
      RECT 36.27 3.215 36.275 3.65 ;
      RECT 36.265 3.215 36.27 3.623 ;
      RECT 36.235 3.215 36.25 3.61 ;
      RECT 35.39 4.75 35.575 4.96 ;
      RECT 35.38 4.755 35.59 4.953 ;
      RECT 35.38 4.755 35.61 4.925 ;
      RECT 35.38 4.755 35.625 4.904 ;
      RECT 35.38 4.755 35.64 4.902 ;
      RECT 35.38 4.755 35.65 4.901 ;
      RECT 35.38 4.755 35.68 4.898 ;
      RECT 36.03 4.6 36.29 4.86 ;
      RECT 35.99 4.647 36.29 4.843 ;
      RECT 35.981 4.655 35.99 4.846 ;
      RECT 35.575 4.748 36.29 4.843 ;
      RECT 35.895 4.673 35.981 4.853 ;
      RECT 35.59 4.745 36.29 4.843 ;
      RECT 35.836 4.695 35.895 4.865 ;
      RECT 35.61 4.741 36.29 4.843 ;
      RECT 35.75 4.707 35.836 4.876 ;
      RECT 35.625 4.737 36.29 4.843 ;
      RECT 35.695 4.72 35.75 4.888 ;
      RECT 35.64 4.735 36.29 4.843 ;
      RECT 35.68 4.726 35.695 4.894 ;
      RECT 35.65 4.731 36.29 4.843 ;
      RECT 35.795 4.255 36.055 4.515 ;
      RECT 35.795 4.275 36.165 4.485 ;
      RECT 35.795 4.28 36.175 4.48 ;
      RECT 35.986 3.694 36.065 3.925 ;
      RECT 35.9 3.697 36.115 3.92 ;
      RECT 35.895 3.697 36.115 3.915 ;
      RECT 35.895 3.702 36.125 3.913 ;
      RECT 35.87 3.702 36.125 3.91 ;
      RECT 35.87 3.71 36.135 3.908 ;
      RECT 35.75 3.645 36.01 3.905 ;
      RECT 35.75 3.692 36.06 3.905 ;
      RECT 35.005 4.265 35.01 4.525 ;
      RECT 34.835 4.035 34.84 4.525 ;
      RECT 34.72 4.275 34.725 4.5 ;
      RECT 35.43 3.37 35.435 3.58 ;
      RECT 35.435 3.375 35.45 3.575 ;
      RECT 35.37 3.37 35.43 3.588 ;
      RECT 35.355 3.37 35.37 3.598 ;
      RECT 35.305 3.37 35.355 3.615 ;
      RECT 35.285 3.37 35.305 3.638 ;
      RECT 35.27 3.37 35.285 3.65 ;
      RECT 35.25 3.37 35.27 3.66 ;
      RECT 35.24 3.375 35.25 3.669 ;
      RECT 35.235 3.385 35.24 3.674 ;
      RECT 35.23 3.397 35.235 3.678 ;
      RECT 35.22 3.42 35.23 3.683 ;
      RECT 35.215 3.435 35.22 3.687 ;
      RECT 35.21 3.452 35.215 3.69 ;
      RECT 35.205 3.46 35.21 3.693 ;
      RECT 35.195 3.465 35.205 3.697 ;
      RECT 35.19 3.472 35.195 3.702 ;
      RECT 35.18 3.477 35.19 3.706 ;
      RECT 35.155 3.489 35.18 3.717 ;
      RECT 35.135 3.506 35.155 3.733 ;
      RECT 35.11 3.523 35.135 3.755 ;
      RECT 35.075 3.546 35.11 3.813 ;
      RECT 35.055 3.568 35.075 3.875 ;
      RECT 35.05 3.578 35.055 3.91 ;
      RECT 35.04 3.585 35.05 3.948 ;
      RECT 35.035 3.592 35.04 3.968 ;
      RECT 35.03 3.603 35.035 4.005 ;
      RECT 35.025 3.611 35.03 4.07 ;
      RECT 35.015 3.622 35.025 4.123 ;
      RECT 35.01 3.64 35.015 4.193 ;
      RECT 35.005 3.65 35.01 4.23 ;
      RECT 35 3.66 35.005 4.525 ;
      RECT 34.995 3.672 35 4.525 ;
      RECT 34.99 3.682 34.995 4.525 ;
      RECT 34.98 3.692 34.99 4.525 ;
      RECT 34.97 3.715 34.98 4.525 ;
      RECT 34.955 3.75 34.97 4.525 ;
      RECT 34.915 3.812 34.955 4.525 ;
      RECT 34.91 3.865 34.915 4.525 ;
      RECT 34.885 3.9 34.91 4.525 ;
      RECT 34.87 3.945 34.885 4.525 ;
      RECT 34.865 3.967 34.87 4.525 ;
      RECT 34.855 3.98 34.865 4.525 ;
      RECT 34.845 4.005 34.855 4.525 ;
      RECT 34.84 4.027 34.845 4.525 ;
      RECT 34.815 4.065 34.835 4.525 ;
      RECT 34.775 4.122 34.815 4.525 ;
      RECT 34.77 4.172 34.775 4.525 ;
      RECT 34.765 4.19 34.77 4.525 ;
      RECT 34.76 4.202 34.765 4.525 ;
      RECT 34.75 4.22 34.76 4.525 ;
      RECT 34.74 4.24 34.75 4.5 ;
      RECT 34.735 4.257 34.74 4.5 ;
      RECT 34.725 4.27 34.735 4.5 ;
      RECT 34.695 4.28 34.72 4.5 ;
      RECT 34.685 4.287 34.695 4.5 ;
      RECT 34.67 4.297 34.685 4.495 ;
      RECT 33.77 10.055 34.06 10.285 ;
      RECT 33.83 8.575 34 10.285 ;
      RECT 33.82 8.945 34.175 9.3 ;
      RECT 33.77 8.575 34.06 8.805 ;
      RECT 33.365 3.69 33.47 4.26 ;
      RECT 33.365 4.025 33.69 4.255 ;
      RECT 33.365 4.055 33.86 4.225 ;
      RECT 33.365 3.69 33.555 4.255 ;
      RECT 32.78 3.655 33.07 3.885 ;
      RECT 32.78 3.69 33.555 3.86 ;
      RECT 32.84 2.175 33.01 3.885 ;
      RECT 32.78 2.175 33.07 2.405 ;
      RECT 32.78 10.055 33.07 10.285 ;
      RECT 32.84 8.575 33.01 10.285 ;
      RECT 32.78 8.575 33.07 8.805 ;
      RECT 32.78 8.61 33.635 8.77 ;
      RECT 33.465 8.205 33.635 8.77 ;
      RECT 32.78 8.605 33.175 8.77 ;
      RECT 33.4 8.205 33.69 8.435 ;
      RECT 33.4 8.235 33.86 8.405 ;
      RECT 32.41 4.025 32.7 4.255 ;
      RECT 32.41 4.055 32.87 4.225 ;
      RECT 32.475 2.95 32.64 4.255 ;
      RECT 30.99 2.92 31.28 3.15 ;
      RECT 30.99 2.95 32.64 3.12 ;
      RECT 31.05 2.18 31.22 3.15 ;
      RECT 30.99 2.18 31.28 2.41 ;
      RECT 30.99 10.05 31.28 10.28 ;
      RECT 31.05 9.31 31.22 10.28 ;
      RECT 31.05 9.405 32.64 9.575 ;
      RECT 32.47 8.205 32.64 9.575 ;
      RECT 30.99 9.31 31.28 9.54 ;
      RECT 32.41 8.205 32.7 8.435 ;
      RECT 32.41 8.235 32.87 8.405 ;
      RECT 31.42 3.26 31.77 3.61 ;
      RECT 29.085 3.32 31.77 3.49 ;
      RECT 29.085 2.635 29.255 3.49 ;
      RECT 28.985 2.635 29.335 2.985 ;
      RECT 31.445 8.94 31.77 9.265 ;
      RECT 26.87 8.895 27.22 9.245 ;
      RECT 31.42 8.94 31.77 9.17 ;
      RECT 26.64 8.94 27.22 9.17 ;
      RECT 26.47 8.97 31.77 9.14 ;
      RECT 30.645 3.66 30.965 3.98 ;
      RECT 30.615 3.66 30.965 3.89 ;
      RECT 30.445 3.69 30.965 3.86 ;
      RECT 30.645 8.54 30.965 8.83 ;
      RECT 30.615 8.57 30.965 8.8 ;
      RECT 30.445 8.6 30.965 8.77 ;
      RECT 27.28 3.76 27.465 3.97 ;
      RECT 27.27 3.765 27.48 3.963 ;
      RECT 27.27 3.765 27.566 3.94 ;
      RECT 27.27 3.765 27.625 3.915 ;
      RECT 27.27 3.765 27.68 3.895 ;
      RECT 27.27 3.765 27.69 3.883 ;
      RECT 27.27 3.765 27.885 3.822 ;
      RECT 27.27 3.765 27.915 3.805 ;
      RECT 27.27 3.765 27.935 3.795 ;
      RECT 27.815 3.53 28.075 3.79 ;
      RECT 27.8 3.62 27.815 3.837 ;
      RECT 27.335 3.752 28.075 3.79 ;
      RECT 27.786 3.631 27.8 3.843 ;
      RECT 27.375 3.745 28.075 3.79 ;
      RECT 27.7 3.671 27.786 3.862 ;
      RECT 27.625 3.732 28.075 3.79 ;
      RECT 27.695 3.707 27.7 3.879 ;
      RECT 27.68 3.717 28.075 3.79 ;
      RECT 27.69 3.712 27.695 3.881 ;
      RECT 27.985 4.217 27.99 4.309 ;
      RECT 27.98 4.195 27.985 4.326 ;
      RECT 27.975 4.185 27.98 4.338 ;
      RECT 27.965 4.176 27.975 4.348 ;
      RECT 27.96 4.171 27.965 4.356 ;
      RECT 27.955 4.03 27.96 4.359 ;
      RECT 27.921 4.03 27.955 4.37 ;
      RECT 27.835 4.03 27.921 4.405 ;
      RECT 27.755 4.03 27.835 4.453 ;
      RECT 27.726 4.03 27.755 4.477 ;
      RECT 27.64 4.03 27.726 4.483 ;
      RECT 27.635 4.214 27.64 4.488 ;
      RECT 27.6 4.225 27.635 4.491 ;
      RECT 27.575 4.24 27.6 4.495 ;
      RECT 27.561 4.249 27.575 4.497 ;
      RECT 27.475 4.276 27.561 4.503 ;
      RECT 27.41 4.317 27.475 4.512 ;
      RECT 27.395 4.337 27.41 4.517 ;
      RECT 27.365 4.347 27.395 4.52 ;
      RECT 27.36 4.357 27.365 4.523 ;
      RECT 27.33 4.362 27.36 4.525 ;
      RECT 27.31 4.367 27.33 4.529 ;
      RECT 27.225 4.37 27.31 4.536 ;
      RECT 27.21 4.367 27.225 4.542 ;
      RECT 27.2 4.364 27.21 4.544 ;
      RECT 27.18 4.361 27.2 4.546 ;
      RECT 27.16 4.357 27.18 4.547 ;
      RECT 27.145 4.353 27.16 4.549 ;
      RECT 27.135 4.35 27.145 4.55 ;
      RECT 27.095 4.344 27.135 4.548 ;
      RECT 27.085 4.339 27.095 4.546 ;
      RECT 27.07 4.336 27.085 4.542 ;
      RECT 27.045 4.331 27.07 4.535 ;
      RECT 26.995 4.322 27.045 4.523 ;
      RECT 26.925 4.308 26.995 4.505 ;
      RECT 26.867 4.293 26.925 4.487 ;
      RECT 26.781 4.276 26.867 4.467 ;
      RECT 26.695 4.255 26.781 4.442 ;
      RECT 26.645 4.24 26.695 4.423 ;
      RECT 26.641 4.234 26.645 4.415 ;
      RECT 26.555 4.224 26.641 4.402 ;
      RECT 26.52 4.209 26.555 4.385 ;
      RECT 26.505 4.202 26.52 4.378 ;
      RECT 26.445 4.19 26.505 4.366 ;
      RECT 26.425 4.177 26.445 4.354 ;
      RECT 26.385 4.168 26.425 4.346 ;
      RECT 26.38 4.16 26.385 4.339 ;
      RECT 26.3 4.15 26.38 4.325 ;
      RECT 26.285 4.137 26.3 4.31 ;
      RECT 26.28 4.135 26.285 4.308 ;
      RECT 26.201 4.123 26.28 4.295 ;
      RECT 26.115 4.098 26.201 4.27 ;
      RECT 26.1 4.067 26.115 4.255 ;
      RECT 26.085 4.042 26.1 4.251 ;
      RECT 26.07 4.035 26.085 4.247 ;
      RECT 25.895 4.04 25.9 4.243 ;
      RECT 25.89 4.045 25.895 4.238 ;
      RECT 25.9 4.035 26.07 4.245 ;
      RECT 26.615 3.795 26.72 4.055 ;
      RECT 27.43 3.32 27.435 3.545 ;
      RECT 27.56 3.32 27.615 3.53 ;
      RECT 27.615 3.325 27.625 3.523 ;
      RECT 27.521 3.32 27.56 3.533 ;
      RECT 27.435 3.32 27.521 3.54 ;
      RECT 27.415 3.325 27.43 3.546 ;
      RECT 27.405 3.365 27.415 3.548 ;
      RECT 27.375 3.375 27.405 3.55 ;
      RECT 27.37 3.38 27.375 3.552 ;
      RECT 27.345 3.385 27.37 3.554 ;
      RECT 27.33 3.39 27.345 3.556 ;
      RECT 27.315 3.392 27.33 3.558 ;
      RECT 27.31 3.397 27.315 3.56 ;
      RECT 27.26 3.405 27.31 3.563 ;
      RECT 27.235 3.414 27.26 3.568 ;
      RECT 27.225 3.421 27.235 3.573 ;
      RECT 27.22 3.424 27.225 3.577 ;
      RECT 27.2 3.427 27.22 3.586 ;
      RECT 27.17 3.435 27.2 3.606 ;
      RECT 27.141 3.448 27.17 3.628 ;
      RECT 27.055 3.482 27.141 3.672 ;
      RECT 27.05 3.508 27.055 3.71 ;
      RECT 27.045 3.512 27.05 3.719 ;
      RECT 27.01 3.525 27.045 3.752 ;
      RECT 27 3.539 27.01 3.79 ;
      RECT 26.995 3.543 27 3.803 ;
      RECT 26.99 3.547 26.995 3.808 ;
      RECT 26.98 3.555 26.99 3.82 ;
      RECT 26.975 3.562 26.98 3.835 ;
      RECT 26.95 3.575 26.975 3.86 ;
      RECT 26.91 3.604 26.95 3.915 ;
      RECT 26.895 3.629 26.91 3.97 ;
      RECT 26.885 3.64 26.895 3.993 ;
      RECT 26.88 3.647 26.885 4.005 ;
      RECT 26.875 3.651 26.88 4.013 ;
      RECT 26.82 3.679 26.875 4.055 ;
      RECT 26.8 3.715 26.82 4.055 ;
      RECT 26.785 3.73 26.8 4.055 ;
      RECT 26.73 3.762 26.785 4.055 ;
      RECT 26.72 3.792 26.73 4.055 ;
      RECT 26.33 3.407 26.515 3.645 ;
      RECT 26.315 3.409 26.525 3.64 ;
      RECT 26.2 3.355 26.46 3.615 ;
      RECT 26.195 3.392 26.46 3.569 ;
      RECT 26.19 3.402 26.46 3.566 ;
      RECT 26.185 3.442 26.525 3.56 ;
      RECT 26.18 3.475 26.525 3.55 ;
      RECT 26.19 3.417 26.54 3.488 ;
      RECT 26.487 4.515 26.5 5.045 ;
      RECT 26.401 4.515 26.5 5.044 ;
      RECT 26.401 4.515 26.505 5.043 ;
      RECT 26.315 4.515 26.505 5.041 ;
      RECT 26.31 4.515 26.505 5.038 ;
      RECT 26.31 4.515 26.515 5.036 ;
      RECT 26.305 4.807 26.515 5.033 ;
      RECT 26.305 4.817 26.52 5.03 ;
      RECT 26.305 4.885 26.525 5.026 ;
      RECT 26.295 4.89 26.525 5.025 ;
      RECT 26.295 4.982 26.53 5.022 ;
      RECT 26.28 4.515 26.54 4.775 ;
      RECT 26.21 10.05 26.5 10.28 ;
      RECT 26.27 9.31 26.44 10.28 ;
      RECT 26.185 9.34 26.525 9.685 ;
      RECT 26.21 9.31 26.5 9.685 ;
      RECT 25.51 3.505 25.555 5.04 ;
      RECT 25.71 3.505 25.74 3.72 ;
      RECT 24.085 3.245 24.205 3.455 ;
      RECT 23.745 3.195 24.005 3.455 ;
      RECT 23.745 3.24 24.04 3.445 ;
      RECT 25.75 3.521 25.755 3.575 ;
      RECT 25.745 3.514 25.75 3.708 ;
      RECT 25.74 3.508 25.745 3.715 ;
      RECT 25.695 3.505 25.71 3.728 ;
      RECT 25.69 3.505 25.695 3.75 ;
      RECT 25.685 3.505 25.69 3.798 ;
      RECT 25.68 3.505 25.685 3.818 ;
      RECT 25.67 3.505 25.68 3.925 ;
      RECT 25.665 3.505 25.67 3.988 ;
      RECT 25.66 3.505 25.665 4.045 ;
      RECT 25.655 3.505 25.66 4.053 ;
      RECT 25.64 3.505 25.655 4.16 ;
      RECT 25.63 3.505 25.64 4.295 ;
      RECT 25.62 3.505 25.63 4.405 ;
      RECT 25.61 3.505 25.62 4.462 ;
      RECT 25.605 3.505 25.61 4.502 ;
      RECT 25.6 3.505 25.605 4.538 ;
      RECT 25.59 3.505 25.6 4.578 ;
      RECT 25.585 3.505 25.59 4.62 ;
      RECT 25.565 3.505 25.585 4.685 ;
      RECT 25.57 4.83 25.575 5.01 ;
      RECT 25.565 4.812 25.57 5.018 ;
      RECT 25.56 3.505 25.565 4.748 ;
      RECT 25.56 4.792 25.565 5.025 ;
      RECT 25.555 3.505 25.56 5.035 ;
      RECT 25.5 3.505 25.51 3.805 ;
      RECT 25.505 4.052 25.51 5.04 ;
      RECT 25.5 4.117 25.505 5.04 ;
      RECT 25.495 3.506 25.5 3.795 ;
      RECT 25.49 4.182 25.5 5.04 ;
      RECT 25.485 3.507 25.495 3.785 ;
      RECT 25.475 4.295 25.49 5.04 ;
      RECT 25.48 3.508 25.485 3.775 ;
      RECT 25.46 3.509 25.48 3.753 ;
      RECT 25.465 4.392 25.475 5.04 ;
      RECT 25.46 4.467 25.465 5.04 ;
      RECT 25.45 3.508 25.46 3.73 ;
      RECT 25.455 4.51 25.46 5.04 ;
      RECT 25.45 4.537 25.455 5.04 ;
      RECT 25.44 3.506 25.45 3.718 ;
      RECT 25.445 4.58 25.45 5.04 ;
      RECT 25.44 4.607 25.445 5.04 ;
      RECT 25.43 3.505 25.44 3.705 ;
      RECT 25.435 4.622 25.44 5.04 ;
      RECT 25.395 4.68 25.435 5.04 ;
      RECT 25.425 3.504 25.43 3.69 ;
      RECT 25.42 3.502 25.425 3.683 ;
      RECT 25.41 3.499 25.42 3.673 ;
      RECT 25.405 3.496 25.41 3.658 ;
      RECT 25.39 3.492 25.405 3.651 ;
      RECT 25.385 4.735 25.395 5.04 ;
      RECT 25.385 3.489 25.39 3.646 ;
      RECT 25.37 3.485 25.385 3.64 ;
      RECT 25.38 4.752 25.385 5.04 ;
      RECT 25.37 4.815 25.38 5.04 ;
      RECT 25.29 3.47 25.37 3.62 ;
      RECT 25.365 4.822 25.37 5.035 ;
      RECT 25.36 4.83 25.365 5.025 ;
      RECT 25.28 3.456 25.29 3.604 ;
      RECT 25.265 3.452 25.28 3.602 ;
      RECT 25.255 3.447 25.265 3.598 ;
      RECT 25.23 3.44 25.255 3.59 ;
      RECT 25.225 3.435 25.23 3.585 ;
      RECT 25.215 3.435 25.225 3.583 ;
      RECT 25.205 3.433 25.215 3.581 ;
      RECT 25.175 3.425 25.205 3.575 ;
      RECT 25.16 3.417 25.175 3.568 ;
      RECT 25.14 3.412 25.16 3.561 ;
      RECT 25.135 3.408 25.14 3.556 ;
      RECT 25.105 3.401 25.135 3.55 ;
      RECT 25.08 3.392 25.105 3.54 ;
      RECT 25.05 3.385 25.08 3.532 ;
      RECT 25.025 3.375 25.05 3.523 ;
      RECT 25.01 3.367 25.025 3.517 ;
      RECT 24.985 3.362 25.01 3.512 ;
      RECT 24.975 3.358 24.985 3.507 ;
      RECT 24.955 3.353 24.975 3.502 ;
      RECT 24.92 3.348 24.955 3.495 ;
      RECT 24.86 3.343 24.92 3.488 ;
      RECT 24.847 3.339 24.86 3.486 ;
      RECT 24.761 3.334 24.847 3.483 ;
      RECT 24.675 3.324 24.761 3.479 ;
      RECT 24.634 3.317 24.675 3.476 ;
      RECT 24.548 3.31 24.634 3.473 ;
      RECT 24.462 3.3 24.548 3.469 ;
      RECT 24.376 3.29 24.462 3.464 ;
      RECT 24.29 3.28 24.376 3.46 ;
      RECT 24.28 3.265 24.29 3.458 ;
      RECT 24.27 3.25 24.28 3.458 ;
      RECT 24.205 3.245 24.27 3.457 ;
      RECT 24.04 3.242 24.085 3.45 ;
      RECT 25.285 4.147 25.29 4.338 ;
      RECT 25.28 4.142 25.285 4.345 ;
      RECT 25.266 4.14 25.28 4.351 ;
      RECT 25.18 4.14 25.266 4.353 ;
      RECT 25.176 4.14 25.18 4.356 ;
      RECT 25.09 4.14 25.176 4.374 ;
      RECT 25.08 4.145 25.09 4.393 ;
      RECT 25.07 4.2 25.08 4.397 ;
      RECT 25.045 4.215 25.07 4.404 ;
      RECT 25.005 4.235 25.045 4.417 ;
      RECT 25 4.247 25.005 4.427 ;
      RECT 24.985 4.253 25 4.432 ;
      RECT 24.98 4.258 24.985 4.436 ;
      RECT 24.96 4.265 24.98 4.441 ;
      RECT 24.89 4.29 24.96 4.458 ;
      RECT 24.85 4.318 24.89 4.478 ;
      RECT 24.845 4.328 24.85 4.486 ;
      RECT 24.825 4.335 24.845 4.488 ;
      RECT 24.82 4.342 24.825 4.491 ;
      RECT 24.79 4.35 24.82 4.494 ;
      RECT 24.785 4.355 24.79 4.498 ;
      RECT 24.711 4.359 24.785 4.506 ;
      RECT 24.625 4.368 24.711 4.522 ;
      RECT 24.621 4.373 24.625 4.531 ;
      RECT 24.535 4.378 24.621 4.541 ;
      RECT 24.495 4.386 24.535 4.553 ;
      RECT 24.445 4.392 24.495 4.56 ;
      RECT 24.36 4.401 24.445 4.575 ;
      RECT 24.285 4.412 24.36 4.593 ;
      RECT 24.25 4.419 24.285 4.603 ;
      RECT 24.175 4.427 24.25 4.608 ;
      RECT 24.12 4.436 24.175 4.608 ;
      RECT 24.095 4.441 24.12 4.606 ;
      RECT 24.085 4.444 24.095 4.604 ;
      RECT 24.05 4.446 24.085 4.602 ;
      RECT 24.02 4.448 24.05 4.598 ;
      RECT 23.975 4.447 24.02 4.594 ;
      RECT 23.955 4.442 23.975 4.591 ;
      RECT 23.905 4.427 23.955 4.588 ;
      RECT 23.895 4.412 23.905 4.583 ;
      RECT 23.845 4.397 23.895 4.573 ;
      RECT 23.795 4.372 23.845 4.553 ;
      RECT 23.785 4.357 23.795 4.535 ;
      RECT 23.78 4.355 23.785 4.529 ;
      RECT 23.76 4.35 23.78 4.524 ;
      RECT 23.755 4.342 23.76 4.518 ;
      RECT 23.74 4.336 23.755 4.511 ;
      RECT 23.735 4.331 23.74 4.503 ;
      RECT 23.715 4.326 23.735 4.495 ;
      RECT 23.7 4.319 23.715 4.488 ;
      RECT 23.685 4.313 23.7 4.479 ;
      RECT 23.68 4.307 23.685 4.472 ;
      RECT 23.635 4.282 23.68 4.458 ;
      RECT 23.62 4.252 23.635 4.44 ;
      RECT 23.605 4.235 23.62 4.431 ;
      RECT 23.58 4.215 23.605 4.419 ;
      RECT 23.54 4.185 23.58 4.399 ;
      RECT 23.53 4.155 23.54 4.384 ;
      RECT 23.515 4.145 23.53 4.377 ;
      RECT 23.46 4.11 23.515 4.356 ;
      RECT 23.445 4.073 23.46 4.335 ;
      RECT 23.435 4.06 23.445 4.327 ;
      RECT 23.385 4.03 23.435 4.309 ;
      RECT 23.37 3.96 23.385 4.29 ;
      RECT 23.325 3.96 23.37 4.273 ;
      RECT 23.3 3.96 23.325 4.255 ;
      RECT 23.29 3.96 23.3 4.248 ;
      RECT 23.211 3.96 23.29 4.241 ;
      RECT 23.125 3.96 23.211 4.233 ;
      RECT 23.11 3.992 23.125 4.228 ;
      RECT 23.035 4.002 23.11 4.224 ;
      RECT 23.015 4.012 23.035 4.219 ;
      RECT 22.99 4.012 23.015 4.216 ;
      RECT 22.98 4.002 22.99 4.215 ;
      RECT 22.97 3.975 22.98 4.214 ;
      RECT 22.93 3.97 22.97 4.212 ;
      RECT 22.885 3.97 22.93 4.208 ;
      RECT 22.86 3.97 22.885 4.203 ;
      RECT 22.81 3.97 22.86 4.19 ;
      RECT 22.77 3.975 22.78 4.175 ;
      RECT 22.78 3.97 22.81 4.18 ;
      RECT 24.765 3.75 25.025 4.01 ;
      RECT 24.76 3.772 25.025 3.968 ;
      RECT 24 3.6 24.22 3.965 ;
      RECT 23.982 3.687 24.22 3.964 ;
      RECT 23.965 3.692 24.22 3.961 ;
      RECT 23.965 3.692 24.24 3.96 ;
      RECT 23.935 3.702 24.24 3.958 ;
      RECT 23.93 3.717 24.24 3.954 ;
      RECT 23.93 3.717 24.245 3.953 ;
      RECT 23.925 3.775 24.245 3.951 ;
      RECT 23.925 3.775 24.255 3.948 ;
      RECT 23.92 3.84 24.255 3.943 ;
      RECT 24 3.6 24.26 3.86 ;
      RECT 22.745 3.43 23.005 3.69 ;
      RECT 22.745 3.473 23.091 3.664 ;
      RECT 22.745 3.473 23.135 3.663 ;
      RECT 22.745 3.473 23.155 3.661 ;
      RECT 22.745 3.473 23.255 3.66 ;
      RECT 22.745 3.473 23.275 3.658 ;
      RECT 22.745 3.473 23.285 3.653 ;
      RECT 23.155 3.44 23.345 3.65 ;
      RECT 23.155 3.442 23.35 3.648 ;
      RECT 23.145 3.447 23.355 3.64 ;
      RECT 23.091 3.471 23.355 3.64 ;
      RECT 23.135 3.465 23.145 3.662 ;
      RECT 23.145 3.445 23.35 3.648 ;
      RECT 22.1 4.505 22.305 4.735 ;
      RECT 22.04 4.455 22.095 4.715 ;
      RECT 22.1 4.455 22.3 4.735 ;
      RECT 23.07 4.77 23.075 4.797 ;
      RECT 23.06 4.68 23.07 4.802 ;
      RECT 23.055 4.602 23.06 4.808 ;
      RECT 23.045 4.592 23.055 4.815 ;
      RECT 23.04 4.582 23.045 4.821 ;
      RECT 23.03 4.577 23.04 4.823 ;
      RECT 23.015 4.569 23.03 4.831 ;
      RECT 23 4.56 23.015 4.843 ;
      RECT 22.99 4.552 23 4.853 ;
      RECT 22.955 4.47 22.99 4.871 ;
      RECT 22.92 4.47 22.955 4.89 ;
      RECT 22.905 4.47 22.92 4.898 ;
      RECT 22.85 4.47 22.905 4.898 ;
      RECT 22.816 4.47 22.85 4.889 ;
      RECT 22.73 4.47 22.816 4.865 ;
      RECT 22.72 4.53 22.73 4.847 ;
      RECT 22.68 4.532 22.72 4.838 ;
      RECT 22.675 4.534 22.68 4.828 ;
      RECT 22.655 4.536 22.675 4.823 ;
      RECT 22.645 4.539 22.655 4.818 ;
      RECT 22.635 4.54 22.645 4.813 ;
      RECT 22.611 4.541 22.635 4.805 ;
      RECT 22.525 4.546 22.611 4.783 ;
      RECT 22.47 4.545 22.525 4.756 ;
      RECT 22.455 4.538 22.47 4.743 ;
      RECT 22.42 4.533 22.455 4.739 ;
      RECT 22.365 4.525 22.42 4.738 ;
      RECT 22.305 4.512 22.365 4.736 ;
      RECT 22.095 4.455 22.1 4.723 ;
      RECT 22.17 3.825 22.355 4.035 ;
      RECT 22.16 3.83 22.37 4.028 ;
      RECT 22.2 3.735 22.46 3.995 ;
      RECT 22.155 3.892 22.46 3.918 ;
      RECT 21.5 3.685 21.505 4.485 ;
      RECT 21.445 3.735 21.475 4.485 ;
      RECT 21.435 3.735 21.44 4.045 ;
      RECT 21.42 3.735 21.425 4.04 ;
      RECT 20.965 3.78 20.98 3.995 ;
      RECT 20.895 3.78 20.98 3.99 ;
      RECT 22.16 3.36 22.23 3.57 ;
      RECT 22.23 3.367 22.24 3.565 ;
      RECT 22.126 3.36 22.16 3.577 ;
      RECT 22.04 3.36 22.126 3.601 ;
      RECT 22.03 3.365 22.04 3.62 ;
      RECT 22.025 3.377 22.03 3.623 ;
      RECT 22.01 3.392 22.025 3.627 ;
      RECT 22.005 3.41 22.01 3.631 ;
      RECT 21.965 3.42 22.005 3.64 ;
      RECT 21.95 3.427 21.965 3.652 ;
      RECT 21.935 3.432 21.95 3.657 ;
      RECT 21.92 3.435 21.935 3.662 ;
      RECT 21.91 3.437 21.92 3.666 ;
      RECT 21.875 3.444 21.91 3.674 ;
      RECT 21.84 3.452 21.875 3.688 ;
      RECT 21.83 3.458 21.84 3.697 ;
      RECT 21.825 3.46 21.83 3.699 ;
      RECT 21.805 3.463 21.825 3.705 ;
      RECT 21.775 3.47 21.805 3.716 ;
      RECT 21.765 3.476 21.775 3.723 ;
      RECT 21.74 3.479 21.765 3.73 ;
      RECT 21.73 3.483 21.74 3.738 ;
      RECT 21.725 3.484 21.73 3.76 ;
      RECT 21.72 3.485 21.725 3.775 ;
      RECT 21.715 3.486 21.72 3.79 ;
      RECT 21.71 3.487 21.715 3.805 ;
      RECT 21.705 3.488 21.71 3.835 ;
      RECT 21.695 3.49 21.705 3.868 ;
      RECT 21.68 3.494 21.695 3.915 ;
      RECT 21.67 3.497 21.68 3.96 ;
      RECT 21.665 3.5 21.67 3.988 ;
      RECT 21.655 3.502 21.665 4.015 ;
      RECT 21.65 3.505 21.655 4.05 ;
      RECT 21.62 3.51 21.65 4.108 ;
      RECT 21.615 3.515 21.62 4.193 ;
      RECT 21.61 3.517 21.615 4.228 ;
      RECT 21.605 3.519 21.61 4.31 ;
      RECT 21.6 3.521 21.605 4.398 ;
      RECT 21.59 3.523 21.6 4.48 ;
      RECT 21.575 3.537 21.59 4.485 ;
      RECT 21.54 3.582 21.575 4.485 ;
      RECT 21.53 3.622 21.54 4.485 ;
      RECT 21.515 3.65 21.53 4.485 ;
      RECT 21.51 3.667 21.515 4.485 ;
      RECT 21.505 3.675 21.51 4.485 ;
      RECT 21.495 3.69 21.5 4.485 ;
      RECT 21.49 3.697 21.495 4.485 ;
      RECT 21.48 3.717 21.49 4.485 ;
      RECT 21.475 3.73 21.48 4.485 ;
      RECT 21.44 3.735 21.445 4.07 ;
      RECT 21.425 4.125 21.445 4.485 ;
      RECT 21.425 3.735 21.435 4.043 ;
      RECT 21.42 4.165 21.425 4.485 ;
      RECT 21.37 3.735 21.42 4.038 ;
      RECT 21.415 4.202 21.42 4.485 ;
      RECT 21.405 4.225 21.415 4.485 ;
      RECT 21.4 4.27 21.405 4.485 ;
      RECT 21.39 4.28 21.4 4.478 ;
      RECT 21.316 3.735 21.37 4.032 ;
      RECT 21.23 3.735 21.316 4.025 ;
      RECT 21.181 3.782 21.23 4.018 ;
      RECT 21.095 3.79 21.181 4.011 ;
      RECT 21.08 3.787 21.095 4.006 ;
      RECT 21.066 3.78 21.08 4.005 ;
      RECT 20.98 3.78 21.066 4 ;
      RECT 20.885 3.785 20.895 3.985 ;
      RECT 20.475 3.215 20.49 3.615 ;
      RECT 20.67 3.215 20.675 3.475 ;
      RECT 20.415 3.215 20.46 3.475 ;
      RECT 20.87 4.52 20.875 4.725 ;
      RECT 20.865 4.51 20.87 4.73 ;
      RECT 20.86 4.497 20.865 4.735 ;
      RECT 20.855 4.477 20.86 4.735 ;
      RECT 20.83 4.43 20.855 4.735 ;
      RECT 20.795 4.345 20.83 4.735 ;
      RECT 20.79 4.282 20.795 4.735 ;
      RECT 20.785 4.267 20.79 4.735 ;
      RECT 20.77 4.227 20.785 4.735 ;
      RECT 20.765 4.202 20.77 4.735 ;
      RECT 20.755 4.185 20.765 4.735 ;
      RECT 20.72 4.107 20.755 4.735 ;
      RECT 20.715 4.05 20.72 4.735 ;
      RECT 20.71 4.037 20.715 4.735 ;
      RECT 20.7 4.015 20.71 4.735 ;
      RECT 20.69 3.98 20.7 4.735 ;
      RECT 20.68 3.95 20.69 4.735 ;
      RECT 20.67 3.865 20.68 4.378 ;
      RECT 20.677 4.51 20.68 4.735 ;
      RECT 20.675 4.52 20.677 4.735 ;
      RECT 20.665 4.53 20.675 4.73 ;
      RECT 20.66 3.215 20.67 3.61 ;
      RECT 20.665 3.742 20.67 4.353 ;
      RECT 20.66 3.64 20.665 4.336 ;
      RECT 20.65 3.215 20.66 4.312 ;
      RECT 20.645 3.215 20.65 4.283 ;
      RECT 20.64 3.215 20.645 4.273 ;
      RECT 20.62 3.215 20.64 4.235 ;
      RECT 20.615 3.215 20.62 4.193 ;
      RECT 20.61 3.215 20.615 4.173 ;
      RECT 20.58 3.215 20.61 4.123 ;
      RECT 20.57 3.215 20.58 4.07 ;
      RECT 20.565 3.215 20.57 4.043 ;
      RECT 20.56 3.215 20.565 4.028 ;
      RECT 20.55 3.215 20.56 4.005 ;
      RECT 20.54 3.215 20.55 3.98 ;
      RECT 20.535 3.215 20.54 3.92 ;
      RECT 20.525 3.215 20.535 3.858 ;
      RECT 20.52 3.215 20.525 3.778 ;
      RECT 20.515 3.215 20.52 3.743 ;
      RECT 20.51 3.215 20.515 3.718 ;
      RECT 20.505 3.215 20.51 3.703 ;
      RECT 20.5 3.215 20.505 3.673 ;
      RECT 20.495 3.215 20.5 3.65 ;
      RECT 20.49 3.215 20.495 3.623 ;
      RECT 20.46 3.215 20.475 3.61 ;
      RECT 19.615 4.75 19.8 4.96 ;
      RECT 19.605 4.755 19.815 4.953 ;
      RECT 19.605 4.755 19.835 4.925 ;
      RECT 19.605 4.755 19.85 4.904 ;
      RECT 19.605 4.755 19.865 4.902 ;
      RECT 19.605 4.755 19.875 4.901 ;
      RECT 19.605 4.755 19.905 4.898 ;
      RECT 20.255 4.6 20.515 4.86 ;
      RECT 20.215 4.647 20.515 4.843 ;
      RECT 20.206 4.655 20.215 4.846 ;
      RECT 19.8 4.748 20.515 4.843 ;
      RECT 20.12 4.673 20.206 4.853 ;
      RECT 19.815 4.745 20.515 4.843 ;
      RECT 20.061 4.695 20.12 4.865 ;
      RECT 19.835 4.741 20.515 4.843 ;
      RECT 19.975 4.707 20.061 4.876 ;
      RECT 19.85 4.737 20.515 4.843 ;
      RECT 19.92 4.72 19.975 4.888 ;
      RECT 19.865 4.735 20.515 4.843 ;
      RECT 19.905 4.726 19.92 4.894 ;
      RECT 19.875 4.731 20.515 4.843 ;
      RECT 20.02 4.255 20.28 4.515 ;
      RECT 20.02 4.275 20.39 4.485 ;
      RECT 20.02 4.28 20.4 4.48 ;
      RECT 20.211 3.694 20.29 3.925 ;
      RECT 20.125 3.697 20.34 3.92 ;
      RECT 20.12 3.697 20.34 3.915 ;
      RECT 20.12 3.702 20.35 3.913 ;
      RECT 20.095 3.702 20.35 3.91 ;
      RECT 20.095 3.71 20.36 3.908 ;
      RECT 19.975 3.645 20.235 3.905 ;
      RECT 19.975 3.692 20.285 3.905 ;
      RECT 19.23 4.265 19.235 4.525 ;
      RECT 19.06 4.035 19.065 4.525 ;
      RECT 18.945 4.275 18.95 4.5 ;
      RECT 19.655 3.37 19.66 3.58 ;
      RECT 19.66 3.375 19.675 3.575 ;
      RECT 19.595 3.37 19.655 3.588 ;
      RECT 19.58 3.37 19.595 3.598 ;
      RECT 19.53 3.37 19.58 3.615 ;
      RECT 19.51 3.37 19.53 3.638 ;
      RECT 19.495 3.37 19.51 3.65 ;
      RECT 19.475 3.37 19.495 3.66 ;
      RECT 19.465 3.375 19.475 3.669 ;
      RECT 19.46 3.385 19.465 3.674 ;
      RECT 19.455 3.397 19.46 3.678 ;
      RECT 19.445 3.42 19.455 3.683 ;
      RECT 19.44 3.435 19.445 3.687 ;
      RECT 19.435 3.452 19.44 3.69 ;
      RECT 19.43 3.46 19.435 3.693 ;
      RECT 19.42 3.465 19.43 3.697 ;
      RECT 19.415 3.472 19.42 3.702 ;
      RECT 19.405 3.477 19.415 3.706 ;
      RECT 19.38 3.489 19.405 3.717 ;
      RECT 19.36 3.506 19.38 3.733 ;
      RECT 19.335 3.523 19.36 3.755 ;
      RECT 19.3 3.546 19.335 3.813 ;
      RECT 19.28 3.568 19.3 3.875 ;
      RECT 19.275 3.578 19.28 3.91 ;
      RECT 19.265 3.585 19.275 3.948 ;
      RECT 19.26 3.592 19.265 3.968 ;
      RECT 19.255 3.603 19.26 4.005 ;
      RECT 19.25 3.611 19.255 4.07 ;
      RECT 19.24 3.622 19.25 4.123 ;
      RECT 19.235 3.64 19.24 4.193 ;
      RECT 19.23 3.65 19.235 4.23 ;
      RECT 19.225 3.66 19.23 4.525 ;
      RECT 19.22 3.672 19.225 4.525 ;
      RECT 19.215 3.682 19.22 4.525 ;
      RECT 19.205 3.692 19.215 4.525 ;
      RECT 19.195 3.715 19.205 4.525 ;
      RECT 19.18 3.75 19.195 4.525 ;
      RECT 19.14 3.812 19.18 4.525 ;
      RECT 19.135 3.865 19.14 4.525 ;
      RECT 19.11 3.9 19.135 4.525 ;
      RECT 19.095 3.945 19.11 4.525 ;
      RECT 19.09 3.967 19.095 4.525 ;
      RECT 19.08 3.98 19.09 4.525 ;
      RECT 19.07 4.005 19.08 4.525 ;
      RECT 19.065 4.027 19.07 4.525 ;
      RECT 19.04 4.065 19.06 4.525 ;
      RECT 19 4.122 19.04 4.525 ;
      RECT 18.995 4.172 19 4.525 ;
      RECT 18.99 4.19 18.995 4.525 ;
      RECT 18.985 4.202 18.99 4.525 ;
      RECT 18.975 4.22 18.985 4.525 ;
      RECT 18.965 4.24 18.975 4.5 ;
      RECT 18.96 4.257 18.965 4.5 ;
      RECT 18.95 4.27 18.96 4.5 ;
      RECT 18.92 4.28 18.945 4.5 ;
      RECT 18.91 4.287 18.92 4.5 ;
      RECT 18.895 4.297 18.91 4.495 ;
      RECT 17.99 10.055 18.28 10.285 ;
      RECT 18.05 8.575 18.22 10.285 ;
      RECT 18.045 8.94 18.395 9.29 ;
      RECT 17.99 8.575 18.28 8.805 ;
      RECT 17.585 3.69 17.69 4.26 ;
      RECT 17.585 4.025 17.91 4.255 ;
      RECT 17.585 4.055 18.08 4.225 ;
      RECT 17.585 3.69 17.775 4.255 ;
      RECT 17 3.655 17.29 3.885 ;
      RECT 17 3.69 17.775 3.86 ;
      RECT 17.06 2.175 17.23 3.885 ;
      RECT 17 2.175 17.29 2.405 ;
      RECT 17 10.055 17.29 10.285 ;
      RECT 17.06 8.575 17.23 10.285 ;
      RECT 17 8.575 17.29 8.805 ;
      RECT 17 8.61 17.855 8.77 ;
      RECT 17.685 8.205 17.855 8.77 ;
      RECT 17 8.605 17.395 8.77 ;
      RECT 17.62 8.205 17.91 8.435 ;
      RECT 17.62 8.235 18.08 8.405 ;
      RECT 16.63 4.025 16.92 4.255 ;
      RECT 16.63 4.055 17.09 4.225 ;
      RECT 16.695 2.95 16.86 4.255 ;
      RECT 15.21 2.92 15.5 3.15 ;
      RECT 15.21 2.95 16.86 3.12 ;
      RECT 15.27 2.18 15.44 3.15 ;
      RECT 15.21 2.18 15.5 2.41 ;
      RECT 15.21 10.05 15.5 10.28 ;
      RECT 15.27 9.31 15.44 10.28 ;
      RECT 15.27 9.405 16.86 9.575 ;
      RECT 16.69 8.205 16.86 9.575 ;
      RECT 15.21 9.31 15.5 9.54 ;
      RECT 16.63 8.205 16.92 8.435 ;
      RECT 16.63 8.235 17.09 8.405 ;
      RECT 15.64 3.26 15.99 3.61 ;
      RECT 13.305 3.32 15.99 3.49 ;
      RECT 13.305 2.635 13.475 3.49 ;
      RECT 13.205 2.635 13.555 2.985 ;
      RECT 15.665 8.94 15.99 9.265 ;
      RECT 11.06 8.89 11.41 9.24 ;
      RECT 15.64 8.94 15.99 9.17 ;
      RECT 10.86 8.94 11.41 9.17 ;
      RECT 10.69 8.97 15.99 9.14 ;
      RECT 14.865 3.66 15.185 3.98 ;
      RECT 14.835 3.66 15.185 3.89 ;
      RECT 14.665 3.69 15.185 3.86 ;
      RECT 14.865 8.54 15.185 8.83 ;
      RECT 14.835 8.57 15.185 8.8 ;
      RECT 14.665 8.6 15.185 8.77 ;
      RECT 11.5 3.76 11.685 3.97 ;
      RECT 11.49 3.765 11.7 3.963 ;
      RECT 11.49 3.765 11.786 3.94 ;
      RECT 11.49 3.765 11.845 3.915 ;
      RECT 11.49 3.765 11.9 3.895 ;
      RECT 11.49 3.765 11.91 3.883 ;
      RECT 11.49 3.765 12.105 3.822 ;
      RECT 11.49 3.765 12.135 3.805 ;
      RECT 11.49 3.765 12.155 3.795 ;
      RECT 12.035 3.53 12.295 3.79 ;
      RECT 12.02 3.62 12.035 3.837 ;
      RECT 11.555 3.752 12.295 3.79 ;
      RECT 12.006 3.631 12.02 3.843 ;
      RECT 11.595 3.745 12.295 3.79 ;
      RECT 11.92 3.671 12.006 3.862 ;
      RECT 11.845 3.732 12.295 3.79 ;
      RECT 11.915 3.707 11.92 3.879 ;
      RECT 11.9 3.717 12.295 3.79 ;
      RECT 11.91 3.712 11.915 3.881 ;
      RECT 12.205 4.217 12.21 4.309 ;
      RECT 12.2 4.195 12.205 4.326 ;
      RECT 12.195 4.185 12.2 4.338 ;
      RECT 12.185 4.176 12.195 4.348 ;
      RECT 12.18 4.171 12.185 4.356 ;
      RECT 12.175 4.03 12.18 4.359 ;
      RECT 12.141 4.03 12.175 4.37 ;
      RECT 12.055 4.03 12.141 4.405 ;
      RECT 11.975 4.03 12.055 4.453 ;
      RECT 11.946 4.03 11.975 4.477 ;
      RECT 11.86 4.03 11.946 4.483 ;
      RECT 11.855 4.214 11.86 4.488 ;
      RECT 11.82 4.225 11.855 4.491 ;
      RECT 11.795 4.24 11.82 4.495 ;
      RECT 11.781 4.249 11.795 4.497 ;
      RECT 11.695 4.276 11.781 4.503 ;
      RECT 11.63 4.317 11.695 4.512 ;
      RECT 11.615 4.337 11.63 4.517 ;
      RECT 11.585 4.347 11.615 4.52 ;
      RECT 11.58 4.357 11.585 4.523 ;
      RECT 11.55 4.362 11.58 4.525 ;
      RECT 11.53 4.367 11.55 4.529 ;
      RECT 11.445 4.37 11.53 4.536 ;
      RECT 11.43 4.367 11.445 4.542 ;
      RECT 11.42 4.364 11.43 4.544 ;
      RECT 11.4 4.361 11.42 4.546 ;
      RECT 11.38 4.357 11.4 4.547 ;
      RECT 11.365 4.353 11.38 4.549 ;
      RECT 11.355 4.35 11.365 4.55 ;
      RECT 11.315 4.344 11.355 4.548 ;
      RECT 11.305 4.339 11.315 4.546 ;
      RECT 11.29 4.336 11.305 4.542 ;
      RECT 11.265 4.331 11.29 4.535 ;
      RECT 11.215 4.322 11.265 4.523 ;
      RECT 11.145 4.308 11.215 4.505 ;
      RECT 11.087 4.293 11.145 4.487 ;
      RECT 11.001 4.276 11.087 4.467 ;
      RECT 10.915 4.255 11.001 4.442 ;
      RECT 10.865 4.24 10.915 4.423 ;
      RECT 10.861 4.234 10.865 4.415 ;
      RECT 10.775 4.224 10.861 4.402 ;
      RECT 10.74 4.209 10.775 4.385 ;
      RECT 10.725 4.202 10.74 4.378 ;
      RECT 10.665 4.19 10.725 4.366 ;
      RECT 10.645 4.177 10.665 4.354 ;
      RECT 10.605 4.168 10.645 4.346 ;
      RECT 10.6 4.16 10.605 4.339 ;
      RECT 10.52 4.15 10.6 4.325 ;
      RECT 10.505 4.137 10.52 4.31 ;
      RECT 10.5 4.135 10.505 4.308 ;
      RECT 10.421 4.123 10.5 4.295 ;
      RECT 10.335 4.098 10.421 4.27 ;
      RECT 10.32 4.067 10.335 4.255 ;
      RECT 10.305 4.042 10.32 4.251 ;
      RECT 10.29 4.035 10.305 4.247 ;
      RECT 10.115 4.04 10.12 4.243 ;
      RECT 10.11 4.045 10.115 4.238 ;
      RECT 10.12 4.035 10.29 4.245 ;
      RECT 10.835 3.795 10.94 4.055 ;
      RECT 11.65 3.32 11.655 3.545 ;
      RECT 11.78 3.32 11.835 3.53 ;
      RECT 11.835 3.325 11.845 3.523 ;
      RECT 11.741 3.32 11.78 3.533 ;
      RECT 11.655 3.32 11.741 3.54 ;
      RECT 11.635 3.325 11.65 3.546 ;
      RECT 11.625 3.365 11.635 3.548 ;
      RECT 11.595 3.375 11.625 3.55 ;
      RECT 11.59 3.38 11.595 3.552 ;
      RECT 11.565 3.385 11.59 3.554 ;
      RECT 11.55 3.39 11.565 3.556 ;
      RECT 11.535 3.392 11.55 3.558 ;
      RECT 11.53 3.397 11.535 3.56 ;
      RECT 11.48 3.405 11.53 3.563 ;
      RECT 11.455 3.414 11.48 3.568 ;
      RECT 11.445 3.421 11.455 3.573 ;
      RECT 11.44 3.424 11.445 3.577 ;
      RECT 11.42 3.427 11.44 3.586 ;
      RECT 11.39 3.435 11.42 3.606 ;
      RECT 11.361 3.448 11.39 3.628 ;
      RECT 11.275 3.482 11.361 3.672 ;
      RECT 11.27 3.508 11.275 3.71 ;
      RECT 11.265 3.512 11.27 3.719 ;
      RECT 11.23 3.525 11.265 3.752 ;
      RECT 11.22 3.539 11.23 3.79 ;
      RECT 11.215 3.543 11.22 3.803 ;
      RECT 11.21 3.547 11.215 3.808 ;
      RECT 11.2 3.555 11.21 3.82 ;
      RECT 11.195 3.562 11.2 3.835 ;
      RECT 11.17 3.575 11.195 3.86 ;
      RECT 11.13 3.604 11.17 3.915 ;
      RECT 11.115 3.629 11.13 3.97 ;
      RECT 11.105 3.64 11.115 3.993 ;
      RECT 11.1 3.647 11.105 4.005 ;
      RECT 11.095 3.651 11.1 4.013 ;
      RECT 11.04 3.679 11.095 4.055 ;
      RECT 11.02 3.715 11.04 4.055 ;
      RECT 11.005 3.73 11.02 4.055 ;
      RECT 10.95 3.762 11.005 4.055 ;
      RECT 10.94 3.792 10.95 4.055 ;
      RECT 10.55 3.407 10.735 3.645 ;
      RECT 10.535 3.409 10.745 3.64 ;
      RECT 10.42 3.355 10.68 3.615 ;
      RECT 10.415 3.392 10.68 3.569 ;
      RECT 10.41 3.402 10.68 3.566 ;
      RECT 10.405 3.442 10.745 3.56 ;
      RECT 10.4 3.475 10.745 3.55 ;
      RECT 10.41 3.417 10.76 3.488 ;
      RECT 10.707 4.515 10.72 5.045 ;
      RECT 10.621 4.515 10.72 5.044 ;
      RECT 10.621 4.515 10.725 5.043 ;
      RECT 10.535 4.515 10.725 5.041 ;
      RECT 10.53 4.515 10.725 5.038 ;
      RECT 10.53 4.515 10.735 5.036 ;
      RECT 10.525 4.807 10.735 5.033 ;
      RECT 10.525 4.817 10.74 5.03 ;
      RECT 10.525 4.885 10.745 5.026 ;
      RECT 10.515 4.89 10.745 5.025 ;
      RECT 10.515 4.982 10.75 5.022 ;
      RECT 10.5 4.515 10.76 4.775 ;
      RECT 10.43 10.05 10.72 10.28 ;
      RECT 10.49 9.31 10.66 10.28 ;
      RECT 10.405 9.34 10.745 9.685 ;
      RECT 10.43 9.31 10.72 9.685 ;
      RECT 9.73 3.505 9.775 5.04 ;
      RECT 9.93 3.505 9.96 3.72 ;
      RECT 8.305 3.245 8.425 3.455 ;
      RECT 7.965 3.195 8.225 3.455 ;
      RECT 7.965 3.24 8.26 3.445 ;
      RECT 9.97 3.521 9.975 3.575 ;
      RECT 9.965 3.514 9.97 3.708 ;
      RECT 9.96 3.508 9.965 3.715 ;
      RECT 9.915 3.505 9.93 3.728 ;
      RECT 9.91 3.505 9.915 3.75 ;
      RECT 9.905 3.505 9.91 3.798 ;
      RECT 9.9 3.505 9.905 3.818 ;
      RECT 9.89 3.505 9.9 3.925 ;
      RECT 9.885 3.505 9.89 3.988 ;
      RECT 9.88 3.505 9.885 4.045 ;
      RECT 9.875 3.505 9.88 4.053 ;
      RECT 9.86 3.505 9.875 4.16 ;
      RECT 9.85 3.505 9.86 4.295 ;
      RECT 9.84 3.505 9.85 4.405 ;
      RECT 9.83 3.505 9.84 4.462 ;
      RECT 9.825 3.505 9.83 4.502 ;
      RECT 9.82 3.505 9.825 4.538 ;
      RECT 9.81 3.505 9.82 4.578 ;
      RECT 9.805 3.505 9.81 4.62 ;
      RECT 9.785 3.505 9.805 4.685 ;
      RECT 9.79 4.83 9.795 5.01 ;
      RECT 9.785 4.812 9.79 5.018 ;
      RECT 9.78 3.505 9.785 4.748 ;
      RECT 9.78 4.792 9.785 5.025 ;
      RECT 9.775 3.505 9.78 5.035 ;
      RECT 9.72 3.505 9.73 3.805 ;
      RECT 9.725 4.052 9.73 5.04 ;
      RECT 9.72 4.117 9.725 5.04 ;
      RECT 9.715 3.506 9.72 3.795 ;
      RECT 9.71 4.182 9.72 5.04 ;
      RECT 9.705 3.507 9.715 3.785 ;
      RECT 9.695 4.295 9.71 5.04 ;
      RECT 9.7 3.508 9.705 3.775 ;
      RECT 9.68 3.509 9.7 3.753 ;
      RECT 9.685 4.392 9.695 5.04 ;
      RECT 9.68 4.467 9.685 5.04 ;
      RECT 9.67 3.508 9.68 3.73 ;
      RECT 9.675 4.51 9.68 5.04 ;
      RECT 9.67 4.537 9.675 5.04 ;
      RECT 9.66 3.506 9.67 3.718 ;
      RECT 9.665 4.58 9.67 5.04 ;
      RECT 9.66 4.607 9.665 5.04 ;
      RECT 9.65 3.505 9.66 3.705 ;
      RECT 9.655 4.622 9.66 5.04 ;
      RECT 9.615 4.68 9.655 5.04 ;
      RECT 9.645 3.504 9.65 3.69 ;
      RECT 9.64 3.502 9.645 3.683 ;
      RECT 9.63 3.499 9.64 3.673 ;
      RECT 9.625 3.496 9.63 3.658 ;
      RECT 9.61 3.492 9.625 3.651 ;
      RECT 9.605 4.735 9.615 5.04 ;
      RECT 9.605 3.489 9.61 3.646 ;
      RECT 9.59 3.485 9.605 3.64 ;
      RECT 9.6 4.752 9.605 5.04 ;
      RECT 9.59 4.815 9.6 5.04 ;
      RECT 9.51 3.47 9.59 3.62 ;
      RECT 9.585 4.822 9.59 5.035 ;
      RECT 9.58 4.83 9.585 5.025 ;
      RECT 9.5 3.456 9.51 3.604 ;
      RECT 9.485 3.452 9.5 3.602 ;
      RECT 9.475 3.447 9.485 3.598 ;
      RECT 9.45 3.44 9.475 3.59 ;
      RECT 9.445 3.435 9.45 3.585 ;
      RECT 9.435 3.435 9.445 3.583 ;
      RECT 9.425 3.433 9.435 3.581 ;
      RECT 9.395 3.425 9.425 3.575 ;
      RECT 9.38 3.417 9.395 3.568 ;
      RECT 9.36 3.412 9.38 3.561 ;
      RECT 9.355 3.408 9.36 3.556 ;
      RECT 9.325 3.401 9.355 3.55 ;
      RECT 9.3 3.392 9.325 3.54 ;
      RECT 9.27 3.385 9.3 3.532 ;
      RECT 9.245 3.375 9.27 3.523 ;
      RECT 9.23 3.367 9.245 3.517 ;
      RECT 9.205 3.362 9.23 3.512 ;
      RECT 9.195 3.358 9.205 3.507 ;
      RECT 9.175 3.353 9.195 3.502 ;
      RECT 9.14 3.348 9.175 3.495 ;
      RECT 9.08 3.343 9.14 3.488 ;
      RECT 9.067 3.339 9.08 3.486 ;
      RECT 8.981 3.334 9.067 3.483 ;
      RECT 8.895 3.324 8.981 3.479 ;
      RECT 8.854 3.317 8.895 3.476 ;
      RECT 8.768 3.31 8.854 3.473 ;
      RECT 8.682 3.3 8.768 3.469 ;
      RECT 8.596 3.29 8.682 3.464 ;
      RECT 8.51 3.28 8.596 3.46 ;
      RECT 8.5 3.265 8.51 3.458 ;
      RECT 8.49 3.25 8.5 3.458 ;
      RECT 8.425 3.245 8.49 3.457 ;
      RECT 8.26 3.242 8.305 3.45 ;
      RECT 9.505 4.147 9.51 4.338 ;
      RECT 9.5 4.142 9.505 4.345 ;
      RECT 9.486 4.14 9.5 4.351 ;
      RECT 9.4 4.14 9.486 4.353 ;
      RECT 9.396 4.14 9.4 4.356 ;
      RECT 9.31 4.14 9.396 4.374 ;
      RECT 9.3 4.145 9.31 4.393 ;
      RECT 9.29 4.2 9.3 4.397 ;
      RECT 9.265 4.215 9.29 4.404 ;
      RECT 9.225 4.235 9.265 4.417 ;
      RECT 9.22 4.247 9.225 4.427 ;
      RECT 9.205 4.253 9.22 4.432 ;
      RECT 9.2 4.258 9.205 4.436 ;
      RECT 9.18 4.265 9.2 4.441 ;
      RECT 9.11 4.29 9.18 4.458 ;
      RECT 9.07 4.318 9.11 4.478 ;
      RECT 9.065 4.328 9.07 4.486 ;
      RECT 9.045 4.335 9.065 4.488 ;
      RECT 9.04 4.342 9.045 4.491 ;
      RECT 9.01 4.35 9.04 4.494 ;
      RECT 9.005 4.355 9.01 4.498 ;
      RECT 8.931 4.359 9.005 4.506 ;
      RECT 8.845 4.368 8.931 4.522 ;
      RECT 8.841 4.373 8.845 4.531 ;
      RECT 8.755 4.378 8.841 4.541 ;
      RECT 8.715 4.386 8.755 4.553 ;
      RECT 8.665 4.392 8.715 4.56 ;
      RECT 8.58 4.401 8.665 4.575 ;
      RECT 8.505 4.412 8.58 4.593 ;
      RECT 8.47 4.419 8.505 4.603 ;
      RECT 8.395 4.427 8.47 4.608 ;
      RECT 8.34 4.436 8.395 4.608 ;
      RECT 8.315 4.441 8.34 4.606 ;
      RECT 8.305 4.444 8.315 4.604 ;
      RECT 8.27 4.446 8.305 4.602 ;
      RECT 8.24 4.448 8.27 4.598 ;
      RECT 8.195 4.447 8.24 4.594 ;
      RECT 8.175 4.442 8.195 4.591 ;
      RECT 8.125 4.427 8.175 4.588 ;
      RECT 8.115 4.412 8.125 4.583 ;
      RECT 8.065 4.397 8.115 4.573 ;
      RECT 8.015 4.372 8.065 4.553 ;
      RECT 8.005 4.357 8.015 4.535 ;
      RECT 8 4.355 8.005 4.529 ;
      RECT 7.98 4.35 8 4.524 ;
      RECT 7.975 4.342 7.98 4.518 ;
      RECT 7.96 4.336 7.975 4.511 ;
      RECT 7.955 4.331 7.96 4.503 ;
      RECT 7.935 4.326 7.955 4.495 ;
      RECT 7.92 4.319 7.935 4.488 ;
      RECT 7.905 4.313 7.92 4.479 ;
      RECT 7.9 4.307 7.905 4.472 ;
      RECT 7.855 4.282 7.9 4.458 ;
      RECT 7.84 4.252 7.855 4.44 ;
      RECT 7.825 4.235 7.84 4.431 ;
      RECT 7.8 4.215 7.825 4.419 ;
      RECT 7.76 4.185 7.8 4.399 ;
      RECT 7.75 4.155 7.76 4.384 ;
      RECT 7.735 4.145 7.75 4.377 ;
      RECT 7.68 4.11 7.735 4.356 ;
      RECT 7.665 4.073 7.68 4.335 ;
      RECT 7.655 4.06 7.665 4.327 ;
      RECT 7.605 4.03 7.655 4.309 ;
      RECT 7.59 3.96 7.605 4.29 ;
      RECT 7.545 3.96 7.59 4.273 ;
      RECT 7.52 3.96 7.545 4.255 ;
      RECT 7.51 3.96 7.52 4.248 ;
      RECT 7.431 3.96 7.51 4.241 ;
      RECT 7.345 3.96 7.431 4.233 ;
      RECT 7.33 3.992 7.345 4.228 ;
      RECT 7.255 4.002 7.33 4.224 ;
      RECT 7.235 4.012 7.255 4.219 ;
      RECT 7.21 4.012 7.235 4.216 ;
      RECT 7.2 4.002 7.21 4.215 ;
      RECT 7.19 3.975 7.2 4.214 ;
      RECT 7.15 3.97 7.19 4.212 ;
      RECT 7.105 3.97 7.15 4.208 ;
      RECT 7.08 3.97 7.105 4.203 ;
      RECT 7.03 3.97 7.08 4.19 ;
      RECT 6.99 3.975 7 4.175 ;
      RECT 7 3.97 7.03 4.18 ;
      RECT 8.985 3.75 9.245 4.01 ;
      RECT 8.98 3.772 9.245 3.968 ;
      RECT 8.22 3.6 8.44 3.965 ;
      RECT 8.202 3.687 8.44 3.964 ;
      RECT 8.185 3.692 8.44 3.961 ;
      RECT 8.185 3.692 8.46 3.96 ;
      RECT 8.155 3.702 8.46 3.958 ;
      RECT 8.15 3.717 8.46 3.954 ;
      RECT 8.15 3.717 8.465 3.953 ;
      RECT 8.145 3.775 8.465 3.951 ;
      RECT 8.145 3.775 8.475 3.948 ;
      RECT 8.14 3.84 8.475 3.943 ;
      RECT 8.22 3.6 8.48 3.86 ;
      RECT 6.965 3.43 7.225 3.69 ;
      RECT 6.965 3.473 7.311 3.664 ;
      RECT 6.965 3.473 7.355 3.663 ;
      RECT 6.965 3.473 7.375 3.661 ;
      RECT 6.965 3.473 7.475 3.66 ;
      RECT 6.965 3.473 7.495 3.658 ;
      RECT 6.965 3.473 7.505 3.653 ;
      RECT 7.375 3.44 7.565 3.65 ;
      RECT 7.375 3.442 7.57 3.648 ;
      RECT 7.365 3.447 7.575 3.64 ;
      RECT 7.311 3.471 7.575 3.64 ;
      RECT 7.355 3.465 7.365 3.662 ;
      RECT 7.365 3.445 7.57 3.648 ;
      RECT 6.32 4.505 6.525 4.735 ;
      RECT 6.26 4.455 6.315 4.715 ;
      RECT 6.32 4.455 6.52 4.735 ;
      RECT 7.29 4.77 7.295 4.797 ;
      RECT 7.28 4.68 7.29 4.802 ;
      RECT 7.275 4.602 7.28 4.808 ;
      RECT 7.265 4.592 7.275 4.815 ;
      RECT 7.26 4.582 7.265 4.821 ;
      RECT 7.25 4.577 7.26 4.823 ;
      RECT 7.235 4.569 7.25 4.831 ;
      RECT 7.22 4.56 7.235 4.843 ;
      RECT 7.21 4.552 7.22 4.853 ;
      RECT 7.175 4.47 7.21 4.871 ;
      RECT 7.14 4.47 7.175 4.89 ;
      RECT 7.125 4.47 7.14 4.898 ;
      RECT 7.07 4.47 7.125 4.898 ;
      RECT 7.036 4.47 7.07 4.889 ;
      RECT 6.95 4.47 7.036 4.865 ;
      RECT 6.94 4.53 6.95 4.847 ;
      RECT 6.9 4.532 6.94 4.838 ;
      RECT 6.895 4.534 6.9 4.828 ;
      RECT 6.875 4.536 6.895 4.823 ;
      RECT 6.865 4.539 6.875 4.818 ;
      RECT 6.855 4.54 6.865 4.813 ;
      RECT 6.831 4.541 6.855 4.805 ;
      RECT 6.745 4.546 6.831 4.783 ;
      RECT 6.69 4.545 6.745 4.756 ;
      RECT 6.675 4.538 6.69 4.743 ;
      RECT 6.64 4.533 6.675 4.739 ;
      RECT 6.585 4.525 6.64 4.738 ;
      RECT 6.525 4.512 6.585 4.736 ;
      RECT 6.315 4.455 6.32 4.723 ;
      RECT 6.39 3.825 6.575 4.035 ;
      RECT 6.38 3.83 6.59 4.028 ;
      RECT 6.42 3.735 6.68 3.995 ;
      RECT 6.375 3.892 6.68 3.918 ;
      RECT 5.72 3.685 5.725 4.485 ;
      RECT 5.665 3.735 5.695 4.485 ;
      RECT 5.655 3.735 5.66 4.045 ;
      RECT 5.64 3.735 5.645 4.04 ;
      RECT 5.185 3.78 5.2 3.995 ;
      RECT 5.115 3.78 5.2 3.99 ;
      RECT 6.38 3.36 6.45 3.57 ;
      RECT 6.45 3.367 6.46 3.565 ;
      RECT 6.346 3.36 6.38 3.577 ;
      RECT 6.26 3.36 6.346 3.601 ;
      RECT 6.25 3.365 6.26 3.62 ;
      RECT 6.245 3.377 6.25 3.623 ;
      RECT 6.23 3.392 6.245 3.627 ;
      RECT 6.225 3.41 6.23 3.631 ;
      RECT 6.185 3.42 6.225 3.64 ;
      RECT 6.17 3.427 6.185 3.652 ;
      RECT 6.155 3.432 6.17 3.657 ;
      RECT 6.14 3.435 6.155 3.662 ;
      RECT 6.13 3.437 6.14 3.666 ;
      RECT 6.095 3.444 6.13 3.674 ;
      RECT 6.06 3.452 6.095 3.688 ;
      RECT 6.05 3.458 6.06 3.697 ;
      RECT 6.045 3.46 6.05 3.699 ;
      RECT 6.025 3.463 6.045 3.705 ;
      RECT 5.995 3.47 6.025 3.716 ;
      RECT 5.985 3.476 5.995 3.723 ;
      RECT 5.96 3.479 5.985 3.73 ;
      RECT 5.95 3.483 5.96 3.738 ;
      RECT 5.945 3.484 5.95 3.76 ;
      RECT 5.94 3.485 5.945 3.775 ;
      RECT 5.935 3.486 5.94 3.79 ;
      RECT 5.93 3.487 5.935 3.805 ;
      RECT 5.925 3.488 5.93 3.835 ;
      RECT 5.915 3.49 5.925 3.868 ;
      RECT 5.9 3.494 5.915 3.915 ;
      RECT 5.89 3.497 5.9 3.96 ;
      RECT 5.885 3.5 5.89 3.988 ;
      RECT 5.875 3.502 5.885 4.015 ;
      RECT 5.87 3.505 5.875 4.05 ;
      RECT 5.84 3.51 5.87 4.108 ;
      RECT 5.835 3.515 5.84 4.193 ;
      RECT 5.83 3.517 5.835 4.228 ;
      RECT 5.825 3.519 5.83 4.31 ;
      RECT 5.82 3.521 5.825 4.398 ;
      RECT 5.81 3.523 5.82 4.48 ;
      RECT 5.795 3.537 5.81 4.485 ;
      RECT 5.76 3.582 5.795 4.485 ;
      RECT 5.75 3.622 5.76 4.485 ;
      RECT 5.735 3.65 5.75 4.485 ;
      RECT 5.73 3.667 5.735 4.485 ;
      RECT 5.725 3.675 5.73 4.485 ;
      RECT 5.715 3.69 5.72 4.485 ;
      RECT 5.71 3.697 5.715 4.485 ;
      RECT 5.7 3.717 5.71 4.485 ;
      RECT 5.695 3.73 5.7 4.485 ;
      RECT 5.66 3.735 5.665 4.07 ;
      RECT 5.645 4.125 5.665 4.485 ;
      RECT 5.645 3.735 5.655 4.043 ;
      RECT 5.64 4.165 5.645 4.485 ;
      RECT 5.59 3.735 5.64 4.038 ;
      RECT 5.635 4.202 5.64 4.485 ;
      RECT 5.625 4.225 5.635 4.485 ;
      RECT 5.62 4.27 5.625 4.485 ;
      RECT 5.61 4.28 5.62 4.478 ;
      RECT 5.536 3.735 5.59 4.032 ;
      RECT 5.45 3.735 5.536 4.025 ;
      RECT 5.401 3.782 5.45 4.018 ;
      RECT 5.315 3.79 5.401 4.011 ;
      RECT 5.3 3.787 5.315 4.006 ;
      RECT 5.286 3.78 5.3 4.005 ;
      RECT 5.2 3.78 5.286 4 ;
      RECT 5.105 3.785 5.115 3.985 ;
      RECT 4.695 3.215 4.71 3.615 ;
      RECT 4.89 3.215 4.895 3.475 ;
      RECT 4.635 3.215 4.68 3.475 ;
      RECT 5.09 4.52 5.095 4.725 ;
      RECT 5.085 4.51 5.09 4.73 ;
      RECT 5.08 4.497 5.085 4.735 ;
      RECT 5.075 4.477 5.08 4.735 ;
      RECT 5.05 4.43 5.075 4.735 ;
      RECT 5.015 4.345 5.05 4.735 ;
      RECT 5.01 4.282 5.015 4.735 ;
      RECT 5.005 4.267 5.01 4.735 ;
      RECT 4.99 4.227 5.005 4.735 ;
      RECT 4.985 4.202 4.99 4.735 ;
      RECT 4.975 4.185 4.985 4.735 ;
      RECT 4.94 4.107 4.975 4.735 ;
      RECT 4.935 4.05 4.94 4.735 ;
      RECT 4.93 4.037 4.935 4.735 ;
      RECT 4.92 4.015 4.93 4.735 ;
      RECT 4.91 3.98 4.92 4.735 ;
      RECT 4.9 3.95 4.91 4.735 ;
      RECT 4.89 3.865 4.9 4.378 ;
      RECT 4.897 4.51 4.9 4.735 ;
      RECT 4.895 4.52 4.897 4.735 ;
      RECT 4.885 4.53 4.895 4.73 ;
      RECT 4.88 3.215 4.89 3.61 ;
      RECT 4.885 3.742 4.89 4.353 ;
      RECT 4.88 3.64 4.885 4.336 ;
      RECT 4.87 3.215 4.88 4.312 ;
      RECT 4.865 3.215 4.87 4.283 ;
      RECT 4.86 3.215 4.865 4.273 ;
      RECT 4.84 3.215 4.86 4.235 ;
      RECT 4.835 3.215 4.84 4.193 ;
      RECT 4.83 3.215 4.835 4.173 ;
      RECT 4.8 3.215 4.83 4.123 ;
      RECT 4.79 3.215 4.8 4.07 ;
      RECT 4.785 3.215 4.79 4.043 ;
      RECT 4.78 3.215 4.785 4.028 ;
      RECT 4.77 3.215 4.78 4.005 ;
      RECT 4.76 3.215 4.77 3.98 ;
      RECT 4.755 3.215 4.76 3.92 ;
      RECT 4.745 3.215 4.755 3.858 ;
      RECT 4.74 3.215 4.745 3.778 ;
      RECT 4.735 3.215 4.74 3.743 ;
      RECT 4.73 3.215 4.735 3.718 ;
      RECT 4.725 3.215 4.73 3.703 ;
      RECT 4.72 3.215 4.725 3.673 ;
      RECT 4.715 3.215 4.72 3.65 ;
      RECT 4.71 3.215 4.715 3.623 ;
      RECT 4.68 3.215 4.695 3.61 ;
      RECT 3.835 4.75 4.02 4.96 ;
      RECT 3.825 4.755 4.035 4.953 ;
      RECT 3.825 4.755 4.055 4.925 ;
      RECT 3.825 4.755 4.07 4.904 ;
      RECT 3.825 4.755 4.085 4.902 ;
      RECT 3.825 4.755 4.095 4.901 ;
      RECT 3.825 4.755 4.125 4.898 ;
      RECT 4.475 4.6 4.735 4.86 ;
      RECT 4.435 4.647 4.735 4.843 ;
      RECT 4.426 4.655 4.435 4.846 ;
      RECT 4.02 4.748 4.735 4.843 ;
      RECT 4.34 4.673 4.426 4.853 ;
      RECT 4.035 4.745 4.735 4.843 ;
      RECT 4.281 4.695 4.34 4.865 ;
      RECT 4.055 4.741 4.735 4.843 ;
      RECT 4.195 4.707 4.281 4.876 ;
      RECT 4.07 4.737 4.735 4.843 ;
      RECT 4.14 4.72 4.195 4.888 ;
      RECT 4.085 4.735 4.735 4.843 ;
      RECT 4.125 4.726 4.14 4.894 ;
      RECT 4.095 4.731 4.735 4.843 ;
      RECT 4.24 4.255 4.5 4.515 ;
      RECT 4.24 4.275 4.61 4.485 ;
      RECT 4.24 4.28 4.62 4.48 ;
      RECT 4.431 3.694 4.51 3.925 ;
      RECT 4.345 3.697 4.56 3.92 ;
      RECT 4.34 3.697 4.56 3.915 ;
      RECT 4.34 3.702 4.57 3.913 ;
      RECT 4.315 3.702 4.57 3.91 ;
      RECT 4.315 3.71 4.58 3.908 ;
      RECT 4.195 3.645 4.455 3.905 ;
      RECT 4.195 3.692 4.505 3.905 ;
      RECT 3.45 4.265 3.455 4.525 ;
      RECT 3.28 4.035 3.285 4.525 ;
      RECT 3.165 4.275 3.17 4.5 ;
      RECT 3.875 3.37 3.88 3.58 ;
      RECT 3.88 3.375 3.895 3.575 ;
      RECT 3.815 3.37 3.875 3.588 ;
      RECT 3.8 3.37 3.815 3.598 ;
      RECT 3.75 3.37 3.8 3.615 ;
      RECT 3.73 3.37 3.75 3.638 ;
      RECT 3.715 3.37 3.73 3.65 ;
      RECT 3.695 3.37 3.715 3.66 ;
      RECT 3.685 3.375 3.695 3.669 ;
      RECT 3.68 3.385 3.685 3.674 ;
      RECT 3.675 3.397 3.68 3.678 ;
      RECT 3.665 3.42 3.675 3.683 ;
      RECT 3.66 3.435 3.665 3.687 ;
      RECT 3.655 3.452 3.66 3.69 ;
      RECT 3.65 3.46 3.655 3.693 ;
      RECT 3.64 3.465 3.65 3.697 ;
      RECT 3.635 3.472 3.64 3.702 ;
      RECT 3.625 3.477 3.635 3.706 ;
      RECT 3.6 3.489 3.625 3.717 ;
      RECT 3.58 3.506 3.6 3.733 ;
      RECT 3.555 3.523 3.58 3.755 ;
      RECT 3.52 3.546 3.555 3.813 ;
      RECT 3.5 3.568 3.52 3.875 ;
      RECT 3.495 3.578 3.5 3.91 ;
      RECT 3.485 3.585 3.495 3.948 ;
      RECT 3.48 3.592 3.485 3.968 ;
      RECT 3.475 3.603 3.48 4.005 ;
      RECT 3.47 3.611 3.475 4.07 ;
      RECT 3.46 3.622 3.47 4.123 ;
      RECT 3.455 3.64 3.46 4.193 ;
      RECT 3.45 3.65 3.455 4.23 ;
      RECT 3.445 3.66 3.45 4.525 ;
      RECT 3.44 3.672 3.445 4.525 ;
      RECT 3.435 3.682 3.44 4.525 ;
      RECT 3.425 3.692 3.435 4.525 ;
      RECT 3.415 3.715 3.425 4.525 ;
      RECT 3.4 3.75 3.415 4.525 ;
      RECT 3.36 3.812 3.4 4.525 ;
      RECT 3.355 3.865 3.36 4.525 ;
      RECT 3.33 3.9 3.355 4.525 ;
      RECT 3.315 3.945 3.33 4.525 ;
      RECT 3.31 3.967 3.315 4.525 ;
      RECT 3.3 3.98 3.31 4.525 ;
      RECT 3.29 4.005 3.3 4.525 ;
      RECT 3.285 4.027 3.29 4.525 ;
      RECT 3.26 4.065 3.28 4.525 ;
      RECT 3.22 4.122 3.26 4.525 ;
      RECT 3.215 4.172 3.22 4.525 ;
      RECT 3.21 4.19 3.215 4.525 ;
      RECT 3.205 4.202 3.21 4.525 ;
      RECT 3.195 4.22 3.205 4.525 ;
      RECT 3.185 4.24 3.195 4.5 ;
      RECT 3.18 4.257 3.185 4.5 ;
      RECT 3.17 4.27 3.18 4.5 ;
      RECT 3.14 4.28 3.165 4.5 ;
      RECT 3.13 4.287 3.14 4.5 ;
      RECT 3.115 4.297 3.13 4.495 ;
      RECT 1.97 8.94 2.26 9.17 ;
      RECT 1.8 8.97 2.26 9.14 ;
      RECT 1.54 10.05 1.83 10.28 ;
      RECT 1.6 9.31 1.77 10.28 ;
      RECT 1.51 9.31 1.86 9.6 ;
      RECT 1.135 8.57 1.485 8.86 ;
      RECT 0.995 8.6 1.485 8.77 ;
      RECT 76.005 4.145 76.375 4.515 ;
      RECT 60.22 4.145 60.59 4.515 ;
      RECT 44.435 4.145 44.805 4.515 ;
      RECT 28.66 4.145 29.03 4.515 ;
      RECT 12.88 4.145 13.25 4.515 ;
    LAYER mcon ;
      RECT 81.175 8.605 81.345 8.775 ;
      RECT 81.18 8.6 81.35 8.77 ;
      RECT 65.39 8.605 65.56 8.775 ;
      RECT 65.395 8.6 65.565 8.77 ;
      RECT 49.605 8.605 49.775 8.775 ;
      RECT 49.61 8.6 49.78 8.77 ;
      RECT 33.83 8.605 34 8.775 ;
      RECT 33.835 8.6 34.005 8.77 ;
      RECT 18.05 8.605 18.22 8.775 ;
      RECT 18.055 8.6 18.225 8.77 ;
      RECT 81.175 10.085 81.345 10.255 ;
      RECT 80.825 1.395 80.995 1.565 ;
      RECT 80.805 4.055 80.975 4.225 ;
      RECT 80.805 8.235 80.975 8.405 ;
      RECT 80.185 2.205 80.355 2.375 ;
      RECT 80.185 3.685 80.355 3.855 ;
      RECT 80.185 8.605 80.355 8.775 ;
      RECT 80.185 10.085 80.355 10.255 ;
      RECT 79.835 1.395 80.005 1.565 ;
      RECT 79.815 4.055 79.985 4.225 ;
      RECT 79.815 8.235 79.985 8.405 ;
      RECT 79.135 1.4 79.305 1.57 ;
      RECT 78.825 3.32 78.995 3.49 ;
      RECT 78.825 8.97 78.995 9.14 ;
      RECT 78.455 1.4 78.625 1.57 ;
      RECT 78.395 2.21 78.565 2.38 ;
      RECT 78.395 2.95 78.565 3.12 ;
      RECT 78.395 9.34 78.565 9.51 ;
      RECT 78.395 10.08 78.565 10.25 ;
      RECT 78.02 3.69 78.19 3.86 ;
      RECT 78.02 8.6 78.19 8.77 ;
      RECT 77.775 1.4 77.945 1.57 ;
      RECT 77.095 1.4 77.265 1.57 ;
      RECT 75.47 2.71 75.64 2.88 ;
      RECT 75.1 4.17 75.27 4.34 ;
      RECT 75.01 2.71 75.18 2.88 ;
      RECT 74.78 3.34 74.95 3.51 ;
      RECT 74.635 3.78 74.805 3.95 ;
      RECT 74.55 2.71 74.72 2.88 ;
      RECT 74.09 2.71 74.26 2.88 ;
      RECT 74.045 8.97 74.215 9.14 ;
      RECT 74.025 3.82 74.195 3.99 ;
      RECT 73.68 3.455 73.85 3.625 ;
      RECT 73.67 4.815 73.84 4.985 ;
      RECT 73.63 2.71 73.8 2.88 ;
      RECT 73.615 9.34 73.785 9.51 ;
      RECT 73.615 10.08 73.785 10.25 ;
      RECT 73.255 4.055 73.425 4.225 ;
      RECT 73.17 2.71 73.34 2.88 ;
      RECT 72.905 3.53 73.075 3.7 ;
      RECT 72.725 4.845 72.895 5.015 ;
      RECT 72.71 2.71 72.88 2.88 ;
      RECT 72.445 4.16 72.615 4.33 ;
      RECT 72.25 2.71 72.42 2.88 ;
      RECT 72.125 3.785 72.295 3.955 ;
      RECT 71.79 2.71 71.96 2.88 ;
      RECT 71.435 3.265 71.605 3.435 ;
      RECT 71.36 3.735 71.53 3.905 ;
      RECT 71.33 2.71 71.5 2.88 ;
      RECT 70.87 2.71 71.04 2.88 ;
      RECT 70.51 3.46 70.68 3.63 ;
      RECT 70.41 2.71 70.58 2.88 ;
      RECT 70.17 4.655 70.34 4.825 ;
      RECT 70.135 3.99 70.305 4.16 ;
      RECT 69.95 2.71 70.12 2.88 ;
      RECT 69.525 3.845 69.695 4.015 ;
      RECT 69.49 2.71 69.66 2.88 ;
      RECT 69.455 4.545 69.625 4.715 ;
      RECT 69.395 3.38 69.565 3.55 ;
      RECT 69.03 2.71 69.2 2.88 ;
      RECT 68.755 4.295 68.925 4.465 ;
      RECT 68.57 2.71 68.74 2.88 ;
      RECT 68.25 3.8 68.42 3.97 ;
      RECT 68.11 2.71 68.28 2.88 ;
      RECT 68.03 4.545 68.2 4.715 ;
      RECT 67.825 3.425 67.995 3.595 ;
      RECT 67.65 2.71 67.82 2.88 ;
      RECT 67.555 4.295 67.725 4.465 ;
      RECT 67.515 3.725 67.685 3.895 ;
      RECT 67.19 2.71 67.36 2.88 ;
      RECT 66.97 4.77 67.14 4.94 ;
      RECT 66.83 3.39 67 3.56 ;
      RECT 66.73 2.71 66.9 2.88 ;
      RECT 66.27 2.71 66.44 2.88 ;
      RECT 66.26 4.31 66.43 4.48 ;
      RECT 65.39 10.085 65.56 10.255 ;
      RECT 65.04 1.395 65.21 1.565 ;
      RECT 65.02 4.055 65.19 4.225 ;
      RECT 65.02 8.235 65.19 8.405 ;
      RECT 64.4 2.205 64.57 2.375 ;
      RECT 64.4 3.685 64.57 3.855 ;
      RECT 64.4 8.605 64.57 8.775 ;
      RECT 64.4 10.085 64.57 10.255 ;
      RECT 64.05 1.395 64.22 1.565 ;
      RECT 64.03 4.055 64.2 4.225 ;
      RECT 64.03 8.235 64.2 8.405 ;
      RECT 63.35 1.4 63.52 1.57 ;
      RECT 63.04 3.32 63.21 3.49 ;
      RECT 63.04 8.97 63.21 9.14 ;
      RECT 62.67 1.4 62.84 1.57 ;
      RECT 62.61 2.21 62.78 2.38 ;
      RECT 62.61 2.95 62.78 3.12 ;
      RECT 62.61 9.34 62.78 9.51 ;
      RECT 62.61 10.08 62.78 10.25 ;
      RECT 62.235 3.69 62.405 3.86 ;
      RECT 62.235 8.6 62.405 8.77 ;
      RECT 61.99 1.4 62.16 1.57 ;
      RECT 61.31 1.4 61.48 1.57 ;
      RECT 59.685 2.71 59.855 2.88 ;
      RECT 59.315 4.17 59.485 4.34 ;
      RECT 59.225 2.71 59.395 2.88 ;
      RECT 58.995 3.34 59.165 3.51 ;
      RECT 58.85 3.78 59.02 3.95 ;
      RECT 58.765 2.71 58.935 2.88 ;
      RECT 58.305 2.71 58.475 2.88 ;
      RECT 58.26 8.97 58.43 9.14 ;
      RECT 58.24 3.82 58.41 3.99 ;
      RECT 57.895 3.455 58.065 3.625 ;
      RECT 57.885 4.815 58.055 4.985 ;
      RECT 57.845 2.71 58.015 2.88 ;
      RECT 57.83 9.34 58 9.51 ;
      RECT 57.83 10.08 58 10.25 ;
      RECT 57.47 4.055 57.64 4.225 ;
      RECT 57.385 2.71 57.555 2.88 ;
      RECT 57.12 3.53 57.29 3.7 ;
      RECT 56.94 4.845 57.11 5.015 ;
      RECT 56.925 2.71 57.095 2.88 ;
      RECT 56.66 4.16 56.83 4.33 ;
      RECT 56.465 2.71 56.635 2.88 ;
      RECT 56.34 3.785 56.51 3.955 ;
      RECT 56.005 2.71 56.175 2.88 ;
      RECT 55.65 3.265 55.82 3.435 ;
      RECT 55.575 3.735 55.745 3.905 ;
      RECT 55.545 2.71 55.715 2.88 ;
      RECT 55.085 2.71 55.255 2.88 ;
      RECT 54.725 3.46 54.895 3.63 ;
      RECT 54.625 2.71 54.795 2.88 ;
      RECT 54.385 4.655 54.555 4.825 ;
      RECT 54.35 3.99 54.52 4.16 ;
      RECT 54.165 2.71 54.335 2.88 ;
      RECT 53.74 3.845 53.91 4.015 ;
      RECT 53.705 2.71 53.875 2.88 ;
      RECT 53.67 4.545 53.84 4.715 ;
      RECT 53.61 3.38 53.78 3.55 ;
      RECT 53.245 2.71 53.415 2.88 ;
      RECT 52.97 4.295 53.14 4.465 ;
      RECT 52.785 2.71 52.955 2.88 ;
      RECT 52.465 3.8 52.635 3.97 ;
      RECT 52.325 2.71 52.495 2.88 ;
      RECT 52.245 4.545 52.415 4.715 ;
      RECT 52.04 3.425 52.21 3.595 ;
      RECT 51.865 2.71 52.035 2.88 ;
      RECT 51.77 4.295 51.94 4.465 ;
      RECT 51.73 3.725 51.9 3.895 ;
      RECT 51.405 2.71 51.575 2.88 ;
      RECT 51.185 4.77 51.355 4.94 ;
      RECT 51.045 3.39 51.215 3.56 ;
      RECT 50.945 2.71 51.115 2.88 ;
      RECT 50.485 2.71 50.655 2.88 ;
      RECT 50.475 4.31 50.645 4.48 ;
      RECT 49.605 10.085 49.775 10.255 ;
      RECT 49.255 1.395 49.425 1.565 ;
      RECT 49.235 4.055 49.405 4.225 ;
      RECT 49.235 8.235 49.405 8.405 ;
      RECT 48.615 2.205 48.785 2.375 ;
      RECT 48.615 3.685 48.785 3.855 ;
      RECT 48.615 8.605 48.785 8.775 ;
      RECT 48.615 10.085 48.785 10.255 ;
      RECT 48.265 1.395 48.435 1.565 ;
      RECT 48.245 4.055 48.415 4.225 ;
      RECT 48.245 8.235 48.415 8.405 ;
      RECT 47.565 1.4 47.735 1.57 ;
      RECT 47.255 3.32 47.425 3.49 ;
      RECT 47.255 8.97 47.425 9.14 ;
      RECT 46.885 1.4 47.055 1.57 ;
      RECT 46.825 2.21 46.995 2.38 ;
      RECT 46.825 2.95 46.995 3.12 ;
      RECT 46.825 9.34 46.995 9.51 ;
      RECT 46.825 10.08 46.995 10.25 ;
      RECT 46.45 3.69 46.62 3.86 ;
      RECT 46.45 8.6 46.62 8.77 ;
      RECT 46.205 1.4 46.375 1.57 ;
      RECT 45.525 1.4 45.695 1.57 ;
      RECT 43.9 2.71 44.07 2.88 ;
      RECT 43.53 4.17 43.7 4.34 ;
      RECT 43.44 2.71 43.61 2.88 ;
      RECT 43.21 3.34 43.38 3.51 ;
      RECT 43.065 3.78 43.235 3.95 ;
      RECT 42.98 2.71 43.15 2.88 ;
      RECT 42.52 2.71 42.69 2.88 ;
      RECT 42.475 8.97 42.645 9.14 ;
      RECT 42.455 3.82 42.625 3.99 ;
      RECT 42.11 3.455 42.28 3.625 ;
      RECT 42.1 4.815 42.27 4.985 ;
      RECT 42.06 2.71 42.23 2.88 ;
      RECT 42.045 9.34 42.215 9.51 ;
      RECT 42.045 10.08 42.215 10.25 ;
      RECT 41.685 4.055 41.855 4.225 ;
      RECT 41.6 2.71 41.77 2.88 ;
      RECT 41.335 3.53 41.505 3.7 ;
      RECT 41.155 4.845 41.325 5.015 ;
      RECT 41.14 2.71 41.31 2.88 ;
      RECT 40.875 4.16 41.045 4.33 ;
      RECT 40.68 2.71 40.85 2.88 ;
      RECT 40.555 3.785 40.725 3.955 ;
      RECT 40.22 2.71 40.39 2.88 ;
      RECT 39.865 3.265 40.035 3.435 ;
      RECT 39.79 3.735 39.96 3.905 ;
      RECT 39.76 2.71 39.93 2.88 ;
      RECT 39.3 2.71 39.47 2.88 ;
      RECT 38.94 3.46 39.11 3.63 ;
      RECT 38.84 2.71 39.01 2.88 ;
      RECT 38.6 4.655 38.77 4.825 ;
      RECT 38.565 3.99 38.735 4.16 ;
      RECT 38.38 2.71 38.55 2.88 ;
      RECT 37.955 3.845 38.125 4.015 ;
      RECT 37.92 2.71 38.09 2.88 ;
      RECT 37.885 4.545 38.055 4.715 ;
      RECT 37.825 3.38 37.995 3.55 ;
      RECT 37.46 2.71 37.63 2.88 ;
      RECT 37.185 4.295 37.355 4.465 ;
      RECT 37 2.71 37.17 2.88 ;
      RECT 36.68 3.8 36.85 3.97 ;
      RECT 36.54 2.71 36.71 2.88 ;
      RECT 36.46 4.545 36.63 4.715 ;
      RECT 36.255 3.425 36.425 3.595 ;
      RECT 36.08 2.71 36.25 2.88 ;
      RECT 35.985 4.295 36.155 4.465 ;
      RECT 35.945 3.725 36.115 3.895 ;
      RECT 35.62 2.71 35.79 2.88 ;
      RECT 35.4 4.77 35.57 4.94 ;
      RECT 35.26 3.39 35.43 3.56 ;
      RECT 35.16 2.71 35.33 2.88 ;
      RECT 34.7 2.71 34.87 2.88 ;
      RECT 34.69 4.31 34.86 4.48 ;
      RECT 33.83 10.085 34 10.255 ;
      RECT 33.48 1.395 33.65 1.565 ;
      RECT 33.46 4.055 33.63 4.225 ;
      RECT 33.46 8.235 33.63 8.405 ;
      RECT 32.84 2.205 33.01 2.375 ;
      RECT 32.84 3.685 33.01 3.855 ;
      RECT 32.84 8.605 33.01 8.775 ;
      RECT 32.84 10.085 33.01 10.255 ;
      RECT 32.49 1.395 32.66 1.565 ;
      RECT 32.47 4.055 32.64 4.225 ;
      RECT 32.47 8.235 32.64 8.405 ;
      RECT 31.79 1.4 31.96 1.57 ;
      RECT 31.48 3.32 31.65 3.49 ;
      RECT 31.48 8.97 31.65 9.14 ;
      RECT 31.11 1.4 31.28 1.57 ;
      RECT 31.05 2.21 31.22 2.38 ;
      RECT 31.05 2.95 31.22 3.12 ;
      RECT 31.05 9.34 31.22 9.51 ;
      RECT 31.05 10.08 31.22 10.25 ;
      RECT 30.675 3.69 30.845 3.86 ;
      RECT 30.675 8.6 30.845 8.77 ;
      RECT 30.43 1.4 30.6 1.57 ;
      RECT 29.75 1.4 29.92 1.57 ;
      RECT 28.125 2.71 28.295 2.88 ;
      RECT 27.755 4.17 27.925 4.34 ;
      RECT 27.665 2.71 27.835 2.88 ;
      RECT 27.435 3.34 27.605 3.51 ;
      RECT 27.29 3.78 27.46 3.95 ;
      RECT 27.205 2.71 27.375 2.88 ;
      RECT 26.745 2.71 26.915 2.88 ;
      RECT 26.7 8.97 26.87 9.14 ;
      RECT 26.68 3.82 26.85 3.99 ;
      RECT 26.335 3.455 26.505 3.625 ;
      RECT 26.325 4.815 26.495 4.985 ;
      RECT 26.285 2.71 26.455 2.88 ;
      RECT 26.27 9.34 26.44 9.51 ;
      RECT 26.27 10.08 26.44 10.25 ;
      RECT 25.91 4.055 26.08 4.225 ;
      RECT 25.825 2.71 25.995 2.88 ;
      RECT 25.56 3.53 25.73 3.7 ;
      RECT 25.38 4.845 25.55 5.015 ;
      RECT 25.365 2.71 25.535 2.88 ;
      RECT 25.1 4.16 25.27 4.33 ;
      RECT 24.905 2.71 25.075 2.88 ;
      RECT 24.78 3.785 24.95 3.955 ;
      RECT 24.445 2.71 24.615 2.88 ;
      RECT 24.09 3.265 24.26 3.435 ;
      RECT 24.015 3.735 24.185 3.905 ;
      RECT 23.985 2.71 24.155 2.88 ;
      RECT 23.525 2.71 23.695 2.88 ;
      RECT 23.165 3.46 23.335 3.63 ;
      RECT 23.065 2.71 23.235 2.88 ;
      RECT 22.825 4.655 22.995 4.825 ;
      RECT 22.79 3.99 22.96 4.16 ;
      RECT 22.605 2.71 22.775 2.88 ;
      RECT 22.18 3.845 22.35 4.015 ;
      RECT 22.145 2.71 22.315 2.88 ;
      RECT 22.11 4.545 22.28 4.715 ;
      RECT 22.05 3.38 22.22 3.55 ;
      RECT 21.685 2.71 21.855 2.88 ;
      RECT 21.41 4.295 21.58 4.465 ;
      RECT 21.225 2.71 21.395 2.88 ;
      RECT 20.905 3.8 21.075 3.97 ;
      RECT 20.765 2.71 20.935 2.88 ;
      RECT 20.685 4.545 20.855 4.715 ;
      RECT 20.48 3.425 20.65 3.595 ;
      RECT 20.305 2.71 20.475 2.88 ;
      RECT 20.21 4.295 20.38 4.465 ;
      RECT 20.17 3.725 20.34 3.895 ;
      RECT 19.845 2.71 20.015 2.88 ;
      RECT 19.625 4.77 19.795 4.94 ;
      RECT 19.485 3.39 19.655 3.56 ;
      RECT 19.385 2.71 19.555 2.88 ;
      RECT 18.925 2.71 19.095 2.88 ;
      RECT 18.915 4.31 19.085 4.48 ;
      RECT 18.05 10.085 18.22 10.255 ;
      RECT 17.7 1.395 17.87 1.565 ;
      RECT 17.68 4.055 17.85 4.225 ;
      RECT 17.68 8.235 17.85 8.405 ;
      RECT 17.06 2.205 17.23 2.375 ;
      RECT 17.06 3.685 17.23 3.855 ;
      RECT 17.06 8.605 17.23 8.775 ;
      RECT 17.06 10.085 17.23 10.255 ;
      RECT 16.71 1.395 16.88 1.565 ;
      RECT 16.69 4.055 16.86 4.225 ;
      RECT 16.69 8.235 16.86 8.405 ;
      RECT 16.01 1.4 16.18 1.57 ;
      RECT 15.7 3.32 15.87 3.49 ;
      RECT 15.7 8.97 15.87 9.14 ;
      RECT 15.33 1.4 15.5 1.57 ;
      RECT 15.27 2.21 15.44 2.38 ;
      RECT 15.27 2.95 15.44 3.12 ;
      RECT 15.27 9.34 15.44 9.51 ;
      RECT 15.27 10.08 15.44 10.25 ;
      RECT 14.895 3.69 15.065 3.86 ;
      RECT 14.895 8.6 15.065 8.77 ;
      RECT 14.65 1.4 14.82 1.57 ;
      RECT 13.97 1.4 14.14 1.57 ;
      RECT 12.345 2.71 12.515 2.88 ;
      RECT 11.975 4.17 12.145 4.34 ;
      RECT 11.885 2.71 12.055 2.88 ;
      RECT 11.655 3.34 11.825 3.51 ;
      RECT 11.51 3.78 11.68 3.95 ;
      RECT 11.425 2.71 11.595 2.88 ;
      RECT 10.965 2.71 11.135 2.88 ;
      RECT 10.92 8.97 11.09 9.14 ;
      RECT 10.9 3.82 11.07 3.99 ;
      RECT 10.555 3.455 10.725 3.625 ;
      RECT 10.545 4.815 10.715 4.985 ;
      RECT 10.505 2.71 10.675 2.88 ;
      RECT 10.49 9.34 10.66 9.51 ;
      RECT 10.49 10.08 10.66 10.25 ;
      RECT 10.13 4.055 10.3 4.225 ;
      RECT 10.045 2.71 10.215 2.88 ;
      RECT 9.78 3.53 9.95 3.7 ;
      RECT 9.6 4.845 9.77 5.015 ;
      RECT 9.585 2.71 9.755 2.88 ;
      RECT 9.32 4.16 9.49 4.33 ;
      RECT 9.125 2.71 9.295 2.88 ;
      RECT 9 3.785 9.17 3.955 ;
      RECT 8.665 2.71 8.835 2.88 ;
      RECT 8.31 3.265 8.48 3.435 ;
      RECT 8.235 3.735 8.405 3.905 ;
      RECT 8.205 2.71 8.375 2.88 ;
      RECT 7.745 2.71 7.915 2.88 ;
      RECT 7.385 3.46 7.555 3.63 ;
      RECT 7.285 2.71 7.455 2.88 ;
      RECT 7.045 4.655 7.215 4.825 ;
      RECT 7.01 3.99 7.18 4.16 ;
      RECT 6.825 2.71 6.995 2.88 ;
      RECT 6.4 3.845 6.57 4.015 ;
      RECT 6.365 2.71 6.535 2.88 ;
      RECT 6.33 4.545 6.5 4.715 ;
      RECT 6.27 3.38 6.44 3.55 ;
      RECT 5.905 2.71 6.075 2.88 ;
      RECT 5.63 4.295 5.8 4.465 ;
      RECT 5.445 2.71 5.615 2.88 ;
      RECT 5.125 3.8 5.295 3.97 ;
      RECT 4.985 2.71 5.155 2.88 ;
      RECT 4.905 4.545 5.075 4.715 ;
      RECT 4.7 3.425 4.87 3.595 ;
      RECT 4.525 2.71 4.695 2.88 ;
      RECT 4.43 4.295 4.6 4.465 ;
      RECT 4.39 3.725 4.56 3.895 ;
      RECT 4.065 2.71 4.235 2.88 ;
      RECT 3.845 4.77 4.015 4.94 ;
      RECT 3.705 3.39 3.875 3.56 ;
      RECT 3.605 2.71 3.775 2.88 ;
      RECT 3.145 2.71 3.315 2.88 ;
      RECT 3.135 4.31 3.305 4.48 ;
      RECT 2.03 8.97 2.2 9.14 ;
      RECT 1.6 9.34 1.77 9.51 ;
      RECT 1.6 10.08 1.77 10.25 ;
      RECT 1.225 8.6 1.395 8.77 ;
    LAYER li1 ;
      RECT 74.255 0 74.425 3.38 ;
      RECT 72.295 0 72.465 3.38 ;
      RECT 69.855 0 70.025 3.38 ;
      RECT 68.895 0 69.065 3.38 ;
      RECT 68.375 0 68.545 3.38 ;
      RECT 67.415 0 67.585 3.38 ;
      RECT 66.455 0 66.625 3.38 ;
      RECT 58.47 0 58.64 3.38 ;
      RECT 56.51 0 56.68 3.38 ;
      RECT 54.07 0 54.24 3.38 ;
      RECT 53.11 0 53.28 3.38 ;
      RECT 52.59 0 52.76 3.38 ;
      RECT 51.63 0 51.8 3.38 ;
      RECT 50.67 0 50.84 3.38 ;
      RECT 42.685 0 42.855 3.38 ;
      RECT 40.725 0 40.895 3.38 ;
      RECT 38.285 0 38.455 3.38 ;
      RECT 37.325 0 37.495 3.38 ;
      RECT 36.805 0 36.975 3.38 ;
      RECT 35.845 0 36.015 3.38 ;
      RECT 34.885 0 35.055 3.38 ;
      RECT 26.91 0 27.08 3.38 ;
      RECT 24.95 0 25.12 3.38 ;
      RECT 22.51 0 22.68 3.38 ;
      RECT 21.55 0 21.72 3.38 ;
      RECT 21.03 0 21.2 3.38 ;
      RECT 20.07 0 20.24 3.38 ;
      RECT 19.11 0 19.28 3.38 ;
      RECT 11.13 0 11.3 3.38 ;
      RECT 9.17 0 9.34 3.38 ;
      RECT 6.73 0 6.9 3.38 ;
      RECT 5.77 0 5.94 3.38 ;
      RECT 5.25 0 5.42 3.38 ;
      RECT 4.29 0 4.46 3.38 ;
      RECT 3.33 0 3.5 3.38 ;
      RECT 66.24 0 75.84 2.885 ;
      RECT 50.455 0 60.055 2.885 ;
      RECT 34.67 0 44.27 2.885 ;
      RECT 18.895 0 28.495 2.885 ;
      RECT 3.115 0 12.715 2.885 ;
      RECT 66.125 2.71 75.955 2.88 ;
      RECT 66.24 0 75.955 2.88 ;
      RECT 50.34 2.71 60.17 2.88 ;
      RECT 50.455 0 60.17 2.88 ;
      RECT 34.555 2.71 44.385 2.88 ;
      RECT 34.67 0 44.385 2.88 ;
      RECT 18.78 2.71 28.61 2.88 ;
      RECT 18.895 0 28.61 2.88 ;
      RECT 3 2.71 12.83 2.88 ;
      RECT 3.115 0 12.83 2.88 ;
      RECT 77.015 0 77.185 2.23 ;
      RECT 61.23 0 61.4 2.23 ;
      RECT 45.445 0 45.615 2.23 ;
      RECT 29.67 0 29.84 2.23 ;
      RECT 13.89 0 14.06 2.23 ;
      RECT 80.745 0 80.915 2.225 ;
      RECT 79.755 0 79.925 2.225 ;
      RECT 64.96 0 65.13 2.225 ;
      RECT 63.97 0 64.14 2.225 ;
      RECT 49.175 0 49.345 2.225 ;
      RECT 48.185 0 48.355 2.225 ;
      RECT 33.4 0 33.57 2.225 ;
      RECT 32.41 0 32.58 2.225 ;
      RECT 17.62 0 17.79 2.225 ;
      RECT 16.63 0 16.8 2.225 ;
      RECT 0 0 81.72 1.6 ;
      RECT 81.175 7.305 81.345 8.775 ;
      RECT 81.175 8.6 81.35 8.77 ;
      RECT 80.805 3.035 80.975 4.225 ;
      RECT 80.805 3.035 81.275 3.205 ;
      RECT 80.805 9.255 81.275 9.425 ;
      RECT 80.805 8.235 80.975 9.425 ;
      RECT 79.815 3.035 79.985 4.225 ;
      RECT 79.815 3.035 80.285 3.205 ;
      RECT 79.815 9.255 80.285 9.425 ;
      RECT 79.815 8.235 79.985 9.425 ;
      RECT 77.965 3.93 78.135 5.16 ;
      RECT 78.02 2.15 78.19 4.1 ;
      RECT 77.965 1.87 78.135 2.32 ;
      RECT 77.965 10.14 78.135 10.59 ;
      RECT 78.02 8.36 78.19 10.31 ;
      RECT 77.965 7.3 78.135 8.53 ;
      RECT 77.445 1.87 77.615 5.16 ;
      RECT 77.445 3.37 77.85 3.7 ;
      RECT 77.445 2.53 77.85 2.86 ;
      RECT 77.445 7.3 77.615 10.59 ;
      RECT 77.445 9.6 77.85 9.93 ;
      RECT 77.445 8.76 77.85 9.09 ;
      RECT 74.78 3.27 75.51 3.51 ;
      RECT 75.322 3.065 75.51 3.51 ;
      RECT 75.15 3.077 75.525 3.504 ;
      RECT 75.065 3.092 75.545 3.489 ;
      RECT 75.065 3.107 75.55 3.479 ;
      RECT 75.02 3.127 75.565 3.471 ;
      RECT 74.997 3.162 75.58 3.425 ;
      RECT 74.911 3.185 75.585 3.385 ;
      RECT 74.911 3.203 75.595 3.355 ;
      RECT 74.78 3.272 75.6 3.318 ;
      RECT 74.825 3.215 75.595 3.355 ;
      RECT 74.911 3.167 75.58 3.425 ;
      RECT 74.997 3.136 75.565 3.471 ;
      RECT 75.02 3.117 75.55 3.479 ;
      RECT 75.065 3.09 75.525 3.504 ;
      RECT 75.15 3.072 75.51 3.51 ;
      RECT 75.236 3.066 75.51 3.51 ;
      RECT 75.322 3.061 75.455 3.51 ;
      RECT 75.408 3.056 75.455 3.51 ;
      RECT 75.1 3.954 75.27 4.34 ;
      RECT 75.095 3.954 75.27 4.335 ;
      RECT 75.07 3.954 75.27 4.3 ;
      RECT 75.07 3.982 75.28 4.29 ;
      RECT 75.05 3.982 75.28 4.25 ;
      RECT 75.045 3.982 75.28 4.223 ;
      RECT 75.045 4 75.285 4.215 ;
      RECT 74.99 4 75.285 4.15 ;
      RECT 74.99 4.017 75.295 4.133 ;
      RECT 74.98 4.017 75.295 4.073 ;
      RECT 74.98 4.034 75.3 4.07 ;
      RECT 74.975 3.87 75.145 4.048 ;
      RECT 74.975 3.904 75.231 4.048 ;
      RECT 74.97 4.67 74.975 4.683 ;
      RECT 74.965 4.565 74.97 4.688 ;
      RECT 74.94 4.425 74.965 4.703 ;
      RECT 74.905 4.376 74.94 4.735 ;
      RECT 74.9 4.344 74.905 4.755 ;
      RECT 74.895 4.335 74.9 4.755 ;
      RECT 74.815 4.3 74.895 4.755 ;
      RECT 74.752 4.27 74.815 4.755 ;
      RECT 74.666 4.258 74.752 4.755 ;
      RECT 74.58 4.244 74.666 4.755 ;
      RECT 74.5 4.231 74.58 4.741 ;
      RECT 74.465 4.223 74.5 4.721 ;
      RECT 74.455 4.22 74.465 4.712 ;
      RECT 74.425 4.215 74.455 4.699 ;
      RECT 74.375 4.19 74.425 4.675 ;
      RECT 74.361 4.164 74.375 4.657 ;
      RECT 74.275 4.124 74.361 4.633 ;
      RECT 74.23 4.072 74.275 4.602 ;
      RECT 74.22 4.047 74.23 4.589 ;
      RECT 74.215 3.828 74.22 3.85 ;
      RECT 74.21 4.03 74.22 4.585 ;
      RECT 74.21 3.826 74.215 3.94 ;
      RECT 74.2 3.822 74.21 4.581 ;
      RECT 74.156 3.82 74.2 4.569 ;
      RECT 74.07 3.82 74.156 4.54 ;
      RECT 74.04 3.82 74.07 4.513 ;
      RECT 74.025 3.82 74.04 4.501 ;
      RECT 73.985 3.832 74.025 4.486 ;
      RECT 73.965 3.851 73.985 4.465 ;
      RECT 73.955 3.861 73.965 4.449 ;
      RECT 73.945 3.867 73.955 4.438 ;
      RECT 73.925 3.877 73.945 4.421 ;
      RECT 73.92 3.886 73.925 4.408 ;
      RECT 73.915 3.89 73.92 4.358 ;
      RECT 73.905 3.896 73.915 4.275 ;
      RECT 73.9 3.9 73.905 4.189 ;
      RECT 73.895 3.92 73.9 4.126 ;
      RECT 73.89 3.943 73.895 4.073 ;
      RECT 73.885 3.961 73.89 4.018 ;
      RECT 74.495 3.78 74.665 4.04 ;
      RECT 74.665 3.745 74.71 4.026 ;
      RECT 74.626 3.747 74.715 4.009 ;
      RECT 74.515 3.764 74.801 3.98 ;
      RECT 74.515 3.779 74.805 3.952 ;
      RECT 74.515 3.76 74.715 4.009 ;
      RECT 74.54 3.748 74.665 4.04 ;
      RECT 74.626 3.746 74.71 4.026 ;
      RECT 73.68 3.135 73.85 3.625 ;
      RECT 73.68 3.135 73.885 3.605 ;
      RECT 73.815 3.055 73.925 3.565 ;
      RECT 73.796 3.059 73.945 3.535 ;
      RECT 73.71 3.067 73.965 3.518 ;
      RECT 73.71 3.073 73.97 3.508 ;
      RECT 73.71 3.082 73.99 3.496 ;
      RECT 73.685 3.107 74.02 3.474 ;
      RECT 73.685 3.127 74.025 3.454 ;
      RECT 73.68 3.14 74.035 3.434 ;
      RECT 73.68 3.207 74.04 3.415 ;
      RECT 73.68 3.34 74.045 3.402 ;
      RECT 73.675 3.145 74.035 3.235 ;
      RECT 73.685 3.102 73.99 3.496 ;
      RECT 73.796 3.057 73.925 3.565 ;
      RECT 73.67 4.81 73.97 5.065 ;
      RECT 73.755 4.776 73.97 5.065 ;
      RECT 73.755 4.779 73.975 4.925 ;
      RECT 73.69 4.8 73.975 4.925 ;
      RECT 73.725 4.79 73.97 5.065 ;
      RECT 73.72 4.795 73.975 4.925 ;
      RECT 73.755 4.774 73.956 5.065 ;
      RECT 73.841 4.765 73.956 5.065 ;
      RECT 73.841 4.759 73.87 5.065 ;
      RECT 73.33 4.4 73.34 4.89 ;
      RECT 72.99 4.335 73 4.635 ;
      RECT 73.505 4.507 73.51 4.726 ;
      RECT 73.495 4.487 73.505 4.743 ;
      RECT 73.485 4.467 73.495 4.773 ;
      RECT 73.48 4.457 73.485 4.788 ;
      RECT 73.475 4.453 73.48 4.793 ;
      RECT 73.46 4.445 73.475 4.8 ;
      RECT 73.42 4.425 73.46 4.825 ;
      RECT 73.395 4.407 73.42 4.858 ;
      RECT 73.39 4.405 73.395 4.871 ;
      RECT 73.37 4.402 73.39 4.875 ;
      RECT 73.34 4.4 73.37 4.885 ;
      RECT 73.27 4.402 73.33 4.886 ;
      RECT 73.25 4.402 73.27 4.88 ;
      RECT 73.225 4.4 73.25 4.877 ;
      RECT 73.19 4.395 73.225 4.873 ;
      RECT 73.17 4.389 73.19 4.86 ;
      RECT 73.16 4.386 73.17 4.848 ;
      RECT 73.14 4.383 73.16 4.833 ;
      RECT 73.12 4.379 73.14 4.815 ;
      RECT 73.115 4.376 73.12 4.805 ;
      RECT 73.11 4.375 73.115 4.803 ;
      RECT 73.1 4.372 73.11 4.795 ;
      RECT 73.09 4.366 73.1 4.778 ;
      RECT 73.08 4.36 73.09 4.76 ;
      RECT 73.07 4.354 73.08 4.748 ;
      RECT 73.06 4.348 73.07 4.728 ;
      RECT 73.055 4.344 73.06 4.713 ;
      RECT 73.05 4.342 73.055 4.705 ;
      RECT 73.045 4.34 73.05 4.698 ;
      RECT 73.04 4.338 73.045 4.688 ;
      RECT 73.035 4.336 73.04 4.682 ;
      RECT 73.025 4.335 73.035 4.672 ;
      RECT 73.015 4.335 73.025 4.663 ;
      RECT 73 4.335 73.015 4.648 ;
      RECT 72.96 4.335 72.99 4.632 ;
      RECT 72.94 4.337 72.96 4.627 ;
      RECT 72.935 4.342 72.94 4.625 ;
      RECT 72.905 4.35 72.935 4.623 ;
      RECT 72.875 4.365 72.905 4.622 ;
      RECT 72.83 4.387 72.875 4.627 ;
      RECT 72.825 4.402 72.83 4.631 ;
      RECT 72.81 4.407 72.825 4.633 ;
      RECT 72.805 4.411 72.81 4.635 ;
      RECT 72.745 4.434 72.805 4.644 ;
      RECT 72.725 4.46 72.745 4.657 ;
      RECT 72.715 4.467 72.725 4.661 ;
      RECT 72.7 4.474 72.715 4.664 ;
      RECT 72.68 4.484 72.7 4.667 ;
      RECT 72.675 4.492 72.68 4.67 ;
      RECT 72.63 4.497 72.675 4.677 ;
      RECT 72.62 4.5 72.63 4.684 ;
      RECT 72.61 4.5 72.62 4.688 ;
      RECT 72.575 4.502 72.61 4.7 ;
      RECT 72.555 4.505 72.575 4.713 ;
      RECT 72.515 4.508 72.555 4.724 ;
      RECT 72.5 4.51 72.515 4.737 ;
      RECT 72.49 4.51 72.5 4.742 ;
      RECT 72.465 4.511 72.49 4.75 ;
      RECT 72.455 4.513 72.465 4.755 ;
      RECT 72.45 4.514 72.455 4.758 ;
      RECT 72.425 4.512 72.45 4.761 ;
      RECT 72.41 4.51 72.425 4.762 ;
      RECT 72.39 4.507 72.41 4.764 ;
      RECT 72.37 4.502 72.39 4.764 ;
      RECT 72.31 4.497 72.37 4.761 ;
      RECT 72.275 4.472 72.31 4.757 ;
      RECT 72.265 4.449 72.275 4.755 ;
      RECT 72.235 4.426 72.265 4.755 ;
      RECT 72.225 4.405 72.235 4.755 ;
      RECT 72.2 4.387 72.225 4.753 ;
      RECT 72.185 4.365 72.2 4.75 ;
      RECT 72.17 4.347 72.185 4.748 ;
      RECT 72.15 4.337 72.17 4.746 ;
      RECT 72.135 4.332 72.15 4.745 ;
      RECT 72.12 4.33 72.135 4.744 ;
      RECT 72.09 4.331 72.12 4.742 ;
      RECT 72.07 4.334 72.09 4.74 ;
      RECT 72.013 4.338 72.07 4.74 ;
      RECT 71.927 4.347 72.013 4.74 ;
      RECT 71.841 4.358 71.927 4.74 ;
      RECT 71.755 4.369 71.841 4.74 ;
      RECT 71.735 4.376 71.755 4.748 ;
      RECT 71.725 4.379 71.735 4.755 ;
      RECT 71.66 4.384 71.725 4.773 ;
      RECT 71.63 4.391 71.66 4.798 ;
      RECT 71.62 4.394 71.63 4.805 ;
      RECT 71.575 4.398 71.62 4.81 ;
      RECT 71.545 4.403 71.575 4.815 ;
      RECT 71.544 4.405 71.545 4.815 ;
      RECT 71.458 4.411 71.544 4.815 ;
      RECT 71.372 4.422 71.458 4.815 ;
      RECT 71.286 4.434 71.372 4.815 ;
      RECT 71.2 4.445 71.286 4.815 ;
      RECT 71.185 4.452 71.2 4.81 ;
      RECT 71.18 4.454 71.185 4.804 ;
      RECT 71.16 4.465 71.18 4.799 ;
      RECT 71.15 4.483 71.16 4.793 ;
      RECT 71.145 4.495 71.15 4.593 ;
      RECT 73.44 3.248 73.46 3.335 ;
      RECT 73.435 3.183 73.44 3.367 ;
      RECT 73.425 3.15 73.435 3.372 ;
      RECT 73.42 3.13 73.425 3.378 ;
      RECT 73.39 3.13 73.42 3.395 ;
      RECT 73.341 3.13 73.39 3.431 ;
      RECT 73.255 3.13 73.341 3.489 ;
      RECT 73.226 3.14 73.255 3.538 ;
      RECT 73.14 3.182 73.226 3.591 ;
      RECT 73.12 3.22 73.14 3.638 ;
      RECT 73.095 3.237 73.12 3.658 ;
      RECT 73.085 3.251 73.095 3.678 ;
      RECT 73.08 3.257 73.085 3.688 ;
      RECT 73.075 3.261 73.08 3.695 ;
      RECT 73.025 3.281 73.075 3.7 ;
      RECT 72.96 3.325 73.025 3.7 ;
      RECT 72.935 3.375 72.96 3.7 ;
      RECT 72.925 3.405 72.935 3.7 ;
      RECT 72.92 3.432 72.925 3.7 ;
      RECT 72.915 3.45 72.92 3.7 ;
      RECT 72.905 3.492 72.915 3.7 ;
      RECT 73.255 4.05 73.425 4.225 ;
      RECT 73.195 3.878 73.255 4.213 ;
      RECT 73.185 3.871 73.195 4.196 ;
      RECT 73.14 4.05 73.425 4.176 ;
      RECT 73.121 4.05 73.425 4.154 ;
      RECT 73.035 4.05 73.425 4.119 ;
      RECT 73.015 3.87 73.185 4.075 ;
      RECT 73.015 4.017 73.42 4.075 ;
      RECT 73.015 3.965 73.395 4.075 ;
      RECT 73.015 3.92 73.36 4.075 ;
      RECT 73.015 3.902 73.325 4.075 ;
      RECT 73.015 3.892 73.32 4.075 ;
      RECT 72.665 7.3 72.835 10.59 ;
      RECT 72.665 9.6 73.07 9.93 ;
      RECT 72.665 8.76 73.07 9.09 ;
      RECT 72.735 4.85 72.925 5.075 ;
      RECT 72.725 4.851 72.93 5.07 ;
      RECT 72.725 4.853 72.94 5.05 ;
      RECT 72.725 4.857 72.945 5.035 ;
      RECT 72.725 4.844 72.895 5.07 ;
      RECT 72.725 4.847 72.92 5.07 ;
      RECT 72.735 4.843 72.895 5.075 ;
      RECT 72.821 4.841 72.895 5.075 ;
      RECT 72.445 4.092 72.615 4.33 ;
      RECT 72.445 4.092 72.701 4.244 ;
      RECT 72.445 4.092 72.705 4.154 ;
      RECT 72.495 3.865 72.715 4.133 ;
      RECT 72.49 3.882 72.72 4.106 ;
      RECT 72.455 4.04 72.72 4.106 ;
      RECT 72.475 3.89 72.615 4.33 ;
      RECT 72.465 3.972 72.725 4.089 ;
      RECT 72.46 4.02 72.725 4.089 ;
      RECT 72.465 3.93 72.72 4.106 ;
      RECT 72.49 3.867 72.715 4.133 ;
      RECT 72.055 3.842 72.225 4.04 ;
      RECT 72.055 3.842 72.27 4.015 ;
      RECT 72.125 3.785 72.295 3.973 ;
      RECT 72.1 3.8 72.295 3.973 ;
      RECT 71.715 3.846 71.745 4.04 ;
      RECT 71.71 3.818 71.715 4.04 ;
      RECT 71.68 3.792 71.71 4.042 ;
      RECT 71.655 3.75 71.68 4.045 ;
      RECT 71.645 3.722 71.655 4.047 ;
      RECT 71.61 3.702 71.645 4.049 ;
      RECT 71.545 3.687 71.61 4.055 ;
      RECT 71.495 3.685 71.545 4.061 ;
      RECT 71.472 3.687 71.495 4.066 ;
      RECT 71.386 3.698 71.472 4.072 ;
      RECT 71.3 3.716 71.386 4.082 ;
      RECT 71.285 3.727 71.3 4.088 ;
      RECT 71.215 3.75 71.285 4.094 ;
      RECT 71.16 3.782 71.215 4.102 ;
      RECT 71.12 3.805 71.16 4.108 ;
      RECT 71.106 3.818 71.12 4.111 ;
      RECT 71.02 3.84 71.106 4.117 ;
      RECT 71.005 3.865 71.02 4.123 ;
      RECT 70.965 3.88 71.005 4.127 ;
      RECT 70.915 3.895 70.965 4.132 ;
      RECT 70.89 3.902 70.915 4.136 ;
      RECT 70.83 3.897 70.89 4.14 ;
      RECT 70.815 3.888 70.83 4.144 ;
      RECT 70.745 3.878 70.815 4.14 ;
      RECT 70.72 3.87 70.74 4.13 ;
      RECT 70.661 3.87 70.72 4.108 ;
      RECT 70.575 3.87 70.661 4.065 ;
      RECT 70.74 3.87 70.745 4.135 ;
      RECT 71.435 3.101 71.605 3.435 ;
      RECT 71.405 3.101 71.605 3.43 ;
      RECT 71.345 3.068 71.405 3.418 ;
      RECT 71.345 3.124 71.615 3.413 ;
      RECT 71.32 3.124 71.615 3.407 ;
      RECT 71.315 3.065 71.345 3.404 ;
      RECT 71.3 3.071 71.435 3.402 ;
      RECT 71.295 3.079 71.52 3.39 ;
      RECT 71.295 3.131 71.63 3.343 ;
      RECT 71.28 3.087 71.52 3.338 ;
      RECT 71.28 3.157 71.64 3.279 ;
      RECT 71.25 3.107 71.605 3.24 ;
      RECT 71.25 3.197 71.65 3.236 ;
      RECT 71.3 3.076 71.52 3.402 ;
      RECT 70.64 3.406 70.695 3.67 ;
      RECT 70.64 3.406 70.76 3.669 ;
      RECT 70.64 3.406 70.785 3.668 ;
      RECT 70.64 3.406 70.85 3.667 ;
      RECT 70.785 3.372 70.865 3.666 ;
      RECT 70.6 3.416 71.01 3.665 ;
      RECT 70.64 3.413 71.01 3.665 ;
      RECT 70.6 3.421 71.015 3.658 ;
      RECT 70.585 3.423 71.015 3.657 ;
      RECT 70.585 3.43 71.02 3.653 ;
      RECT 70.565 3.429 71.015 3.649 ;
      RECT 70.565 3.437 71.025 3.648 ;
      RECT 70.56 3.434 71.02 3.644 ;
      RECT 70.56 3.447 71.035 3.643 ;
      RECT 70.545 3.437 71.025 3.642 ;
      RECT 70.51 3.45 71.035 3.635 ;
      RECT 70.695 3.405 71.005 3.665 ;
      RECT 70.695 3.39 70.955 3.665 ;
      RECT 70.76 3.377 70.89 3.665 ;
      RECT 70.305 4.466 70.32 4.859 ;
      RECT 70.27 4.471 70.32 4.858 ;
      RECT 70.305 4.47 70.365 4.857 ;
      RECT 70.25 4.481 70.365 4.856 ;
      RECT 70.265 4.477 70.365 4.856 ;
      RECT 70.23 4.487 70.44 4.853 ;
      RECT 70.23 4.506 70.485 4.851 ;
      RECT 70.23 4.513 70.49 4.848 ;
      RECT 70.215 4.49 70.44 4.845 ;
      RECT 70.195 4.495 70.44 4.838 ;
      RECT 70.19 4.499 70.44 4.834 ;
      RECT 70.19 4.516 70.5 4.833 ;
      RECT 70.17 4.51 70.485 4.829 ;
      RECT 70.17 4.519 70.505 4.823 ;
      RECT 70.165 4.525 70.505 4.595 ;
      RECT 70.23 4.485 70.365 4.853 ;
      RECT 70.105 3.848 70.305 4.16 ;
      RECT 70.18 3.826 70.305 4.16 ;
      RECT 70.12 3.845 70.31 4.145 ;
      RECT 70.09 3.856 70.31 4.143 ;
      RECT 70.105 3.851 70.315 4.109 ;
      RECT 70.09 3.955 70.32 4.076 ;
      RECT 70.12 3.827 70.305 4.16 ;
      RECT 70.18 3.805 70.28 4.16 ;
      RECT 70.205 3.802 70.28 4.16 ;
      RECT 70.205 3.797 70.225 4.16 ;
      RECT 69.61 3.865 69.785 4.04 ;
      RECT 69.605 3.865 69.785 4.038 ;
      RECT 69.58 3.865 69.785 4.033 ;
      RECT 69.525 3.845 69.695 4.023 ;
      RECT 69.525 3.852 69.76 4.023 ;
      RECT 69.61 4.532 69.625 4.715 ;
      RECT 69.6 4.51 69.61 4.715 ;
      RECT 69.585 4.49 69.6 4.715 ;
      RECT 69.575 4.465 69.585 4.715 ;
      RECT 69.545 4.43 69.575 4.715 ;
      RECT 69.51 4.37 69.545 4.715 ;
      RECT 69.505 4.332 69.51 4.715 ;
      RECT 69.455 4.283 69.505 4.715 ;
      RECT 69.445 4.233 69.455 4.703 ;
      RECT 69.43 4.212 69.445 4.663 ;
      RECT 69.41 4.18 69.43 4.613 ;
      RECT 69.385 4.136 69.41 4.553 ;
      RECT 69.38 4.108 69.385 4.508 ;
      RECT 69.375 4.099 69.38 4.494 ;
      RECT 69.37 4.092 69.375 4.481 ;
      RECT 69.365 4.087 69.37 4.47 ;
      RECT 69.36 4.072 69.365 4.46 ;
      RECT 69.355 4.05 69.36 4.447 ;
      RECT 69.345 4.01 69.355 4.422 ;
      RECT 69.32 3.94 69.345 4.378 ;
      RECT 69.315 3.88 69.32 4.343 ;
      RECT 69.3 3.86 69.315 4.31 ;
      RECT 69.295 3.86 69.3 4.285 ;
      RECT 69.265 3.86 69.295 4.24 ;
      RECT 69.22 3.86 69.265 4.18 ;
      RECT 69.145 3.86 69.22 4.128 ;
      RECT 69.14 3.86 69.145 4.093 ;
      RECT 69.135 3.86 69.14 4.083 ;
      RECT 69.13 3.86 69.135 4.063 ;
      RECT 69.395 3.08 69.565 3.55 ;
      RECT 69.34 3.073 69.535 3.534 ;
      RECT 69.34 3.087 69.57 3.533 ;
      RECT 69.325 3.088 69.57 3.514 ;
      RECT 69.32 3.106 69.57 3.5 ;
      RECT 69.325 3.089 69.575 3.498 ;
      RECT 69.31 3.12 69.575 3.483 ;
      RECT 69.325 3.095 69.58 3.468 ;
      RECT 69.305 3.135 69.58 3.465 ;
      RECT 69.32 3.107 69.585 3.45 ;
      RECT 69.32 3.119 69.59 3.43 ;
      RECT 69.305 3.135 69.595 3.413 ;
      RECT 69.305 3.145 69.6 3.268 ;
      RECT 69.3 3.145 69.6 3.225 ;
      RECT 69.3 3.16 69.605 3.203 ;
      RECT 69.395 3.07 69.535 3.55 ;
      RECT 69.395 3.068 69.505 3.55 ;
      RECT 69.481 3.065 69.505 3.55 ;
      RECT 69.14 4.732 69.145 4.778 ;
      RECT 69.13 4.58 69.14 4.802 ;
      RECT 69.125 4.425 69.13 4.827 ;
      RECT 69.11 4.387 69.125 4.838 ;
      RECT 69.105 4.37 69.11 4.845 ;
      RECT 69.095 4.358 69.105 4.852 ;
      RECT 69.09 4.349 69.095 4.854 ;
      RECT 69.085 4.347 69.09 4.858 ;
      RECT 69.04 4.338 69.085 4.873 ;
      RECT 69.035 4.33 69.04 4.887 ;
      RECT 69.03 4.327 69.035 4.891 ;
      RECT 69.015 4.322 69.03 4.899 ;
      RECT 68.96 4.312 69.015 4.91 ;
      RECT 68.925 4.3 68.96 4.911 ;
      RECT 68.916 4.295 68.925 4.905 ;
      RECT 68.83 4.295 68.916 4.895 ;
      RECT 68.8 4.295 68.83 4.873 ;
      RECT 68.79 4.295 68.795 4.853 ;
      RECT 68.785 4.295 68.79 4.815 ;
      RECT 68.78 4.295 68.785 4.773 ;
      RECT 68.775 4.295 68.78 4.733 ;
      RECT 68.77 4.295 68.775 4.663 ;
      RECT 68.76 4.295 68.77 4.585 ;
      RECT 68.755 4.295 68.76 4.485 ;
      RECT 68.795 4.295 68.8 4.855 ;
      RECT 68.29 4.377 68.38 4.855 ;
      RECT 68.275 4.38 68.395 4.853 ;
      RECT 68.29 4.379 68.395 4.853 ;
      RECT 68.255 4.386 68.42 4.843 ;
      RECT 68.275 4.38 68.42 4.843 ;
      RECT 68.24 4.392 68.42 4.831 ;
      RECT 68.275 4.383 68.47 4.824 ;
      RECT 68.226 4.4 68.47 4.822 ;
      RECT 68.255 4.39 68.48 4.81 ;
      RECT 68.226 4.411 68.51 4.801 ;
      RECT 68.14 4.435 68.51 4.795 ;
      RECT 68.14 4.448 68.55 4.778 ;
      RECT 68.135 4.47 68.55 4.771 ;
      RECT 68.105 4.485 68.55 4.761 ;
      RECT 68.1 4.496 68.55 4.751 ;
      RECT 68.07 4.509 68.55 4.742 ;
      RECT 68.055 4.527 68.55 4.731 ;
      RECT 68.03 4.54 68.55 4.721 ;
      RECT 68.29 4.376 68.3 4.855 ;
      RECT 68.336 3.8 68.375 4.045 ;
      RECT 68.25 3.8 68.385 4.043 ;
      RECT 68.135 3.825 68.385 4.04 ;
      RECT 68.135 3.825 68.39 4.038 ;
      RECT 68.135 3.825 68.405 4.033 ;
      RECT 68.241 3.8 68.42 4.013 ;
      RECT 68.155 3.808 68.42 4.013 ;
      RECT 67.825 3.16 67.995 3.595 ;
      RECT 67.815 3.194 67.995 3.578 ;
      RECT 67.895 3.13 68.065 3.565 ;
      RECT 67.8 3.205 68.065 3.543 ;
      RECT 67.895 3.14 68.07 3.533 ;
      RECT 67.825 3.192 68.1 3.518 ;
      RECT 67.785 3.218 68.1 3.503 ;
      RECT 67.785 3.26 68.11 3.483 ;
      RECT 67.78 3.285 68.115 3.465 ;
      RECT 67.78 3.295 68.12 3.45 ;
      RECT 67.775 3.232 68.1 3.448 ;
      RECT 67.775 3.305 68.125 3.433 ;
      RECT 67.77 3.242 68.1 3.43 ;
      RECT 67.765 3.326 68.13 3.413 ;
      RECT 67.765 3.358 68.135 3.393 ;
      RECT 67.76 3.272 68.11 3.385 ;
      RECT 67.765 3.257 68.1 3.413 ;
      RECT 67.78 3.227 68.1 3.465 ;
      RECT 67.625 3.814 67.85 4.07 ;
      RECT 67.625 3.847 67.87 4.06 ;
      RECT 67.59 3.847 67.87 4.058 ;
      RECT 67.59 3.86 67.875 4.048 ;
      RECT 67.59 3.88 67.885 4.04 ;
      RECT 67.59 3.977 67.89 4.033 ;
      RECT 67.57 3.725 67.7 4.023 ;
      RECT 67.525 3.88 67.885 3.965 ;
      RECT 67.515 3.725 67.7 3.91 ;
      RECT 67.515 3.757 67.786 3.91 ;
      RECT 67.48 4.287 67.5 4.465 ;
      RECT 67.445 4.24 67.48 4.465 ;
      RECT 67.43 4.18 67.445 4.465 ;
      RECT 67.405 4.127 67.43 4.465 ;
      RECT 67.39 4.08 67.405 4.465 ;
      RECT 67.37 4.057 67.39 4.465 ;
      RECT 67.345 4.022 67.37 4.465 ;
      RECT 67.335 3.868 67.345 4.465 ;
      RECT 67.305 3.863 67.335 4.456 ;
      RECT 67.3 3.86 67.305 4.446 ;
      RECT 67.285 3.86 67.3 4.42 ;
      RECT 67.28 3.86 67.285 4.383 ;
      RECT 67.255 3.86 67.28 4.335 ;
      RECT 67.235 3.86 67.255 4.26 ;
      RECT 67.225 3.86 67.235 4.22 ;
      RECT 67.22 3.86 67.225 4.195 ;
      RECT 67.215 3.86 67.22 4.178 ;
      RECT 67.21 3.86 67.215 4.16 ;
      RECT 67.205 3.861 67.21 4.15 ;
      RECT 67.195 3.863 67.205 4.118 ;
      RECT 67.185 3.865 67.195 4.085 ;
      RECT 67.175 3.868 67.185 4.058 ;
      RECT 67.5 4.295 67.725 4.465 ;
      RECT 66.83 3.107 67 3.56 ;
      RECT 66.83 3.107 67.09 3.526 ;
      RECT 66.83 3.107 67.12 3.51 ;
      RECT 66.83 3.107 67.15 3.483 ;
      RECT 67.086 3.085 67.165 3.465 ;
      RECT 66.865 3.092 67.17 3.45 ;
      RECT 66.865 3.1 67.18 3.413 ;
      RECT 66.825 3.127 67.18 3.385 ;
      RECT 66.81 3.14 67.18 3.35 ;
      RECT 66.83 3.115 67.2 3.34 ;
      RECT 66.805 3.18 67.2 3.31 ;
      RECT 66.805 3.21 67.205 3.293 ;
      RECT 66.8 3.24 67.205 3.28 ;
      RECT 66.865 3.089 67.165 3.465 ;
      RECT 67 3.086 67.086 3.544 ;
      RECT 66.951 3.087 67.165 3.465 ;
      RECT 67.095 4.747 67.14 4.94 ;
      RECT 67.085 4.717 67.095 4.94 ;
      RECT 67.08 4.702 67.085 4.94 ;
      RECT 67.04 4.612 67.08 4.94 ;
      RECT 67.035 4.525 67.04 4.94 ;
      RECT 67.025 4.495 67.035 4.94 ;
      RECT 67.02 4.455 67.025 4.94 ;
      RECT 67.01 4.417 67.02 4.94 ;
      RECT 67.005 4.382 67.01 4.94 ;
      RECT 66.985 4.335 67.005 4.94 ;
      RECT 66.97 4.26 66.985 4.94 ;
      RECT 66.965 4.215 66.97 4.935 ;
      RECT 66.96 4.195 66.965 4.908 ;
      RECT 66.955 4.175 66.96 4.893 ;
      RECT 66.95 4.15 66.955 4.873 ;
      RECT 66.945 4.128 66.95 4.858 ;
      RECT 66.94 4.106 66.945 4.84 ;
      RECT 66.935 4.085 66.94 4.83 ;
      RECT 66.925 4.057 66.935 4.8 ;
      RECT 66.915 4.02 66.925 4.768 ;
      RECT 66.905 3.98 66.915 4.735 ;
      RECT 66.895 3.958 66.905 4.705 ;
      RECT 66.865 3.91 66.895 4.637 ;
      RECT 66.85 3.87 66.865 4.564 ;
      RECT 66.84 3.87 66.85 4.53 ;
      RECT 66.835 3.87 66.84 4.505 ;
      RECT 66.83 3.87 66.835 4.49 ;
      RECT 66.825 3.87 66.83 4.468 ;
      RECT 66.82 3.87 66.825 4.455 ;
      RECT 66.805 3.87 66.82 4.42 ;
      RECT 66.785 3.87 66.805 4.36 ;
      RECT 66.775 3.87 66.785 4.31 ;
      RECT 66.755 3.87 66.775 4.258 ;
      RECT 66.735 3.87 66.755 4.215 ;
      RECT 66.725 3.87 66.735 4.203 ;
      RECT 66.695 3.87 66.725 4.19 ;
      RECT 66.665 3.891 66.695 4.17 ;
      RECT 66.655 3.919 66.665 4.15 ;
      RECT 66.64 3.936 66.655 4.118 ;
      RECT 66.635 3.95 66.64 4.085 ;
      RECT 66.63 3.958 66.635 4.058 ;
      RECT 66.625 3.966 66.63 4.02 ;
      RECT 66.63 4.49 66.635 4.825 ;
      RECT 66.595 4.477 66.63 4.824 ;
      RECT 66.525 4.417 66.595 4.823 ;
      RECT 66.445 4.36 66.525 4.822 ;
      RECT 66.31 4.32 66.445 4.821 ;
      RECT 66.31 4.507 66.645 4.81 ;
      RECT 66.27 4.507 66.645 4.8 ;
      RECT 66.27 4.525 66.65 4.795 ;
      RECT 66.27 4.615 66.655 4.785 ;
      RECT 66.265 4.31 66.43 4.765 ;
      RECT 66.26 4.31 66.43 4.508 ;
      RECT 66.26 4.467 66.625 4.508 ;
      RECT 66.26 4.455 66.62 4.508 ;
      RECT 65.39 7.305 65.56 8.775 ;
      RECT 65.39 8.6 65.565 8.77 ;
      RECT 65.02 3.035 65.19 4.225 ;
      RECT 65.02 3.035 65.49 3.205 ;
      RECT 65.02 9.255 65.49 9.425 ;
      RECT 65.02 8.235 65.19 9.425 ;
      RECT 64.03 3.035 64.2 4.225 ;
      RECT 64.03 3.035 64.5 3.205 ;
      RECT 64.03 9.255 64.5 9.425 ;
      RECT 64.03 8.235 64.2 9.425 ;
      RECT 62.18 3.93 62.35 5.16 ;
      RECT 62.235 2.15 62.405 4.1 ;
      RECT 62.18 1.87 62.35 2.32 ;
      RECT 62.18 10.14 62.35 10.59 ;
      RECT 62.235 8.36 62.405 10.31 ;
      RECT 62.18 7.3 62.35 8.53 ;
      RECT 61.66 1.87 61.83 5.16 ;
      RECT 61.66 3.37 62.065 3.7 ;
      RECT 61.66 2.53 62.065 2.86 ;
      RECT 61.66 7.3 61.83 10.59 ;
      RECT 61.66 9.6 62.065 9.93 ;
      RECT 61.66 8.76 62.065 9.09 ;
      RECT 58.995 3.27 59.725 3.51 ;
      RECT 59.537 3.065 59.725 3.51 ;
      RECT 59.365 3.077 59.74 3.504 ;
      RECT 59.28 3.092 59.76 3.489 ;
      RECT 59.28 3.107 59.765 3.479 ;
      RECT 59.235 3.127 59.78 3.471 ;
      RECT 59.212 3.162 59.795 3.425 ;
      RECT 59.126 3.185 59.8 3.385 ;
      RECT 59.126 3.203 59.81 3.355 ;
      RECT 58.995 3.272 59.815 3.318 ;
      RECT 59.04 3.215 59.81 3.355 ;
      RECT 59.126 3.167 59.795 3.425 ;
      RECT 59.212 3.136 59.78 3.471 ;
      RECT 59.235 3.117 59.765 3.479 ;
      RECT 59.28 3.09 59.74 3.504 ;
      RECT 59.365 3.072 59.725 3.51 ;
      RECT 59.451 3.066 59.725 3.51 ;
      RECT 59.537 3.061 59.67 3.51 ;
      RECT 59.623 3.056 59.67 3.51 ;
      RECT 59.315 3.954 59.485 4.34 ;
      RECT 59.31 3.954 59.485 4.335 ;
      RECT 59.285 3.954 59.485 4.3 ;
      RECT 59.285 3.982 59.495 4.29 ;
      RECT 59.265 3.982 59.495 4.25 ;
      RECT 59.26 3.982 59.495 4.223 ;
      RECT 59.26 4 59.5 4.215 ;
      RECT 59.205 4 59.5 4.15 ;
      RECT 59.205 4.017 59.51 4.133 ;
      RECT 59.195 4.017 59.51 4.073 ;
      RECT 59.195 4.034 59.515 4.07 ;
      RECT 59.19 3.87 59.36 4.048 ;
      RECT 59.19 3.904 59.446 4.048 ;
      RECT 59.185 4.67 59.19 4.683 ;
      RECT 59.18 4.565 59.185 4.688 ;
      RECT 59.155 4.425 59.18 4.703 ;
      RECT 59.12 4.376 59.155 4.735 ;
      RECT 59.115 4.344 59.12 4.755 ;
      RECT 59.11 4.335 59.115 4.755 ;
      RECT 59.03 4.3 59.11 4.755 ;
      RECT 58.967 4.27 59.03 4.755 ;
      RECT 58.881 4.258 58.967 4.755 ;
      RECT 58.795 4.244 58.881 4.755 ;
      RECT 58.715 4.231 58.795 4.741 ;
      RECT 58.68 4.223 58.715 4.721 ;
      RECT 58.67 4.22 58.68 4.712 ;
      RECT 58.64 4.215 58.67 4.699 ;
      RECT 58.59 4.19 58.64 4.675 ;
      RECT 58.576 4.164 58.59 4.657 ;
      RECT 58.49 4.124 58.576 4.633 ;
      RECT 58.445 4.072 58.49 4.602 ;
      RECT 58.435 4.047 58.445 4.589 ;
      RECT 58.43 3.828 58.435 3.85 ;
      RECT 58.425 4.03 58.435 4.585 ;
      RECT 58.425 3.826 58.43 3.94 ;
      RECT 58.415 3.822 58.425 4.581 ;
      RECT 58.371 3.82 58.415 4.569 ;
      RECT 58.285 3.82 58.371 4.54 ;
      RECT 58.255 3.82 58.285 4.513 ;
      RECT 58.24 3.82 58.255 4.501 ;
      RECT 58.2 3.832 58.24 4.486 ;
      RECT 58.18 3.851 58.2 4.465 ;
      RECT 58.17 3.861 58.18 4.449 ;
      RECT 58.16 3.867 58.17 4.438 ;
      RECT 58.14 3.877 58.16 4.421 ;
      RECT 58.135 3.886 58.14 4.408 ;
      RECT 58.13 3.89 58.135 4.358 ;
      RECT 58.12 3.896 58.13 4.275 ;
      RECT 58.115 3.9 58.12 4.189 ;
      RECT 58.11 3.92 58.115 4.126 ;
      RECT 58.105 3.943 58.11 4.073 ;
      RECT 58.1 3.961 58.105 4.018 ;
      RECT 58.71 3.78 58.88 4.04 ;
      RECT 58.88 3.745 58.925 4.026 ;
      RECT 58.841 3.747 58.93 4.009 ;
      RECT 58.73 3.764 59.016 3.98 ;
      RECT 58.73 3.779 59.02 3.952 ;
      RECT 58.73 3.76 58.93 4.009 ;
      RECT 58.755 3.748 58.88 4.04 ;
      RECT 58.841 3.746 58.925 4.026 ;
      RECT 57.895 3.135 58.065 3.625 ;
      RECT 57.895 3.135 58.1 3.605 ;
      RECT 58.03 3.055 58.14 3.565 ;
      RECT 58.011 3.059 58.16 3.535 ;
      RECT 57.925 3.067 58.18 3.518 ;
      RECT 57.925 3.073 58.185 3.508 ;
      RECT 57.925 3.082 58.205 3.496 ;
      RECT 57.9 3.107 58.235 3.474 ;
      RECT 57.9 3.127 58.24 3.454 ;
      RECT 57.895 3.14 58.25 3.434 ;
      RECT 57.895 3.207 58.255 3.415 ;
      RECT 57.895 3.34 58.26 3.402 ;
      RECT 57.89 3.145 58.25 3.235 ;
      RECT 57.9 3.102 58.205 3.496 ;
      RECT 58.011 3.057 58.14 3.565 ;
      RECT 57.885 4.81 58.185 5.065 ;
      RECT 57.97 4.776 58.185 5.065 ;
      RECT 57.97 4.779 58.19 4.925 ;
      RECT 57.905 4.8 58.19 4.925 ;
      RECT 57.94 4.79 58.185 5.065 ;
      RECT 57.935 4.795 58.19 4.925 ;
      RECT 57.97 4.774 58.171 5.065 ;
      RECT 58.056 4.765 58.171 5.065 ;
      RECT 58.056 4.759 58.085 5.065 ;
      RECT 57.545 4.4 57.555 4.89 ;
      RECT 57.205 4.335 57.215 4.635 ;
      RECT 57.72 4.507 57.725 4.726 ;
      RECT 57.71 4.487 57.72 4.743 ;
      RECT 57.7 4.467 57.71 4.773 ;
      RECT 57.695 4.457 57.7 4.788 ;
      RECT 57.69 4.453 57.695 4.793 ;
      RECT 57.675 4.445 57.69 4.8 ;
      RECT 57.635 4.425 57.675 4.825 ;
      RECT 57.61 4.407 57.635 4.858 ;
      RECT 57.605 4.405 57.61 4.871 ;
      RECT 57.585 4.402 57.605 4.875 ;
      RECT 57.555 4.4 57.585 4.885 ;
      RECT 57.485 4.402 57.545 4.886 ;
      RECT 57.465 4.402 57.485 4.88 ;
      RECT 57.44 4.4 57.465 4.877 ;
      RECT 57.405 4.395 57.44 4.873 ;
      RECT 57.385 4.389 57.405 4.86 ;
      RECT 57.375 4.386 57.385 4.848 ;
      RECT 57.355 4.383 57.375 4.833 ;
      RECT 57.335 4.379 57.355 4.815 ;
      RECT 57.33 4.376 57.335 4.805 ;
      RECT 57.325 4.375 57.33 4.803 ;
      RECT 57.315 4.372 57.325 4.795 ;
      RECT 57.305 4.366 57.315 4.778 ;
      RECT 57.295 4.36 57.305 4.76 ;
      RECT 57.285 4.354 57.295 4.748 ;
      RECT 57.275 4.348 57.285 4.728 ;
      RECT 57.27 4.344 57.275 4.713 ;
      RECT 57.265 4.342 57.27 4.705 ;
      RECT 57.26 4.34 57.265 4.698 ;
      RECT 57.255 4.338 57.26 4.688 ;
      RECT 57.25 4.336 57.255 4.682 ;
      RECT 57.24 4.335 57.25 4.672 ;
      RECT 57.23 4.335 57.24 4.663 ;
      RECT 57.215 4.335 57.23 4.648 ;
      RECT 57.175 4.335 57.205 4.632 ;
      RECT 57.155 4.337 57.175 4.627 ;
      RECT 57.15 4.342 57.155 4.625 ;
      RECT 57.12 4.35 57.15 4.623 ;
      RECT 57.09 4.365 57.12 4.622 ;
      RECT 57.045 4.387 57.09 4.627 ;
      RECT 57.04 4.402 57.045 4.631 ;
      RECT 57.025 4.407 57.04 4.633 ;
      RECT 57.02 4.411 57.025 4.635 ;
      RECT 56.96 4.434 57.02 4.644 ;
      RECT 56.94 4.46 56.96 4.657 ;
      RECT 56.93 4.467 56.94 4.661 ;
      RECT 56.915 4.474 56.93 4.664 ;
      RECT 56.895 4.484 56.915 4.667 ;
      RECT 56.89 4.492 56.895 4.67 ;
      RECT 56.845 4.497 56.89 4.677 ;
      RECT 56.835 4.5 56.845 4.684 ;
      RECT 56.825 4.5 56.835 4.688 ;
      RECT 56.79 4.502 56.825 4.7 ;
      RECT 56.77 4.505 56.79 4.713 ;
      RECT 56.73 4.508 56.77 4.724 ;
      RECT 56.715 4.51 56.73 4.737 ;
      RECT 56.705 4.51 56.715 4.742 ;
      RECT 56.68 4.511 56.705 4.75 ;
      RECT 56.67 4.513 56.68 4.755 ;
      RECT 56.665 4.514 56.67 4.758 ;
      RECT 56.64 4.512 56.665 4.761 ;
      RECT 56.625 4.51 56.64 4.762 ;
      RECT 56.605 4.507 56.625 4.764 ;
      RECT 56.585 4.502 56.605 4.764 ;
      RECT 56.525 4.497 56.585 4.761 ;
      RECT 56.49 4.472 56.525 4.757 ;
      RECT 56.48 4.449 56.49 4.755 ;
      RECT 56.45 4.426 56.48 4.755 ;
      RECT 56.44 4.405 56.45 4.755 ;
      RECT 56.415 4.387 56.44 4.753 ;
      RECT 56.4 4.365 56.415 4.75 ;
      RECT 56.385 4.347 56.4 4.748 ;
      RECT 56.365 4.337 56.385 4.746 ;
      RECT 56.35 4.332 56.365 4.745 ;
      RECT 56.335 4.33 56.35 4.744 ;
      RECT 56.305 4.331 56.335 4.742 ;
      RECT 56.285 4.334 56.305 4.74 ;
      RECT 56.228 4.338 56.285 4.74 ;
      RECT 56.142 4.347 56.228 4.74 ;
      RECT 56.056 4.358 56.142 4.74 ;
      RECT 55.97 4.369 56.056 4.74 ;
      RECT 55.95 4.376 55.97 4.748 ;
      RECT 55.94 4.379 55.95 4.755 ;
      RECT 55.875 4.384 55.94 4.773 ;
      RECT 55.845 4.391 55.875 4.798 ;
      RECT 55.835 4.394 55.845 4.805 ;
      RECT 55.79 4.398 55.835 4.81 ;
      RECT 55.76 4.403 55.79 4.815 ;
      RECT 55.759 4.405 55.76 4.815 ;
      RECT 55.673 4.411 55.759 4.815 ;
      RECT 55.587 4.422 55.673 4.815 ;
      RECT 55.501 4.434 55.587 4.815 ;
      RECT 55.415 4.445 55.501 4.815 ;
      RECT 55.4 4.452 55.415 4.81 ;
      RECT 55.395 4.454 55.4 4.804 ;
      RECT 55.375 4.465 55.395 4.799 ;
      RECT 55.365 4.483 55.375 4.793 ;
      RECT 55.36 4.495 55.365 4.593 ;
      RECT 57.655 3.248 57.675 3.335 ;
      RECT 57.65 3.183 57.655 3.367 ;
      RECT 57.64 3.15 57.65 3.372 ;
      RECT 57.635 3.13 57.64 3.378 ;
      RECT 57.605 3.13 57.635 3.395 ;
      RECT 57.556 3.13 57.605 3.431 ;
      RECT 57.47 3.13 57.556 3.489 ;
      RECT 57.441 3.14 57.47 3.538 ;
      RECT 57.355 3.182 57.441 3.591 ;
      RECT 57.335 3.22 57.355 3.638 ;
      RECT 57.31 3.237 57.335 3.658 ;
      RECT 57.3 3.251 57.31 3.678 ;
      RECT 57.295 3.257 57.3 3.688 ;
      RECT 57.29 3.261 57.295 3.695 ;
      RECT 57.24 3.281 57.29 3.7 ;
      RECT 57.175 3.325 57.24 3.7 ;
      RECT 57.15 3.375 57.175 3.7 ;
      RECT 57.14 3.405 57.15 3.7 ;
      RECT 57.135 3.432 57.14 3.7 ;
      RECT 57.13 3.45 57.135 3.7 ;
      RECT 57.12 3.492 57.13 3.7 ;
      RECT 57.47 4.05 57.64 4.225 ;
      RECT 57.41 3.878 57.47 4.213 ;
      RECT 57.4 3.871 57.41 4.196 ;
      RECT 57.355 4.05 57.64 4.176 ;
      RECT 57.336 4.05 57.64 4.154 ;
      RECT 57.25 4.05 57.64 4.119 ;
      RECT 57.23 3.87 57.4 4.075 ;
      RECT 57.23 4.017 57.635 4.075 ;
      RECT 57.23 3.965 57.61 4.075 ;
      RECT 57.23 3.92 57.575 4.075 ;
      RECT 57.23 3.902 57.54 4.075 ;
      RECT 57.23 3.892 57.535 4.075 ;
      RECT 56.88 7.3 57.05 10.59 ;
      RECT 56.88 9.6 57.285 9.93 ;
      RECT 56.88 8.76 57.285 9.09 ;
      RECT 56.95 4.85 57.14 5.075 ;
      RECT 56.94 4.851 57.145 5.07 ;
      RECT 56.94 4.853 57.155 5.05 ;
      RECT 56.94 4.857 57.16 5.035 ;
      RECT 56.94 4.844 57.11 5.07 ;
      RECT 56.94 4.847 57.135 5.07 ;
      RECT 56.95 4.843 57.11 5.075 ;
      RECT 57.036 4.841 57.11 5.075 ;
      RECT 56.66 4.092 56.83 4.33 ;
      RECT 56.66 4.092 56.916 4.244 ;
      RECT 56.66 4.092 56.92 4.154 ;
      RECT 56.71 3.865 56.93 4.133 ;
      RECT 56.705 3.882 56.935 4.106 ;
      RECT 56.67 4.04 56.935 4.106 ;
      RECT 56.69 3.89 56.83 4.33 ;
      RECT 56.68 3.972 56.94 4.089 ;
      RECT 56.675 4.02 56.94 4.089 ;
      RECT 56.68 3.93 56.935 4.106 ;
      RECT 56.705 3.867 56.93 4.133 ;
      RECT 56.27 3.842 56.44 4.04 ;
      RECT 56.27 3.842 56.485 4.015 ;
      RECT 56.34 3.785 56.51 3.973 ;
      RECT 56.315 3.8 56.51 3.973 ;
      RECT 55.93 3.846 55.96 4.04 ;
      RECT 55.925 3.818 55.93 4.04 ;
      RECT 55.895 3.792 55.925 4.042 ;
      RECT 55.87 3.75 55.895 4.045 ;
      RECT 55.86 3.722 55.87 4.047 ;
      RECT 55.825 3.702 55.86 4.049 ;
      RECT 55.76 3.687 55.825 4.055 ;
      RECT 55.71 3.685 55.76 4.061 ;
      RECT 55.687 3.687 55.71 4.066 ;
      RECT 55.601 3.698 55.687 4.072 ;
      RECT 55.515 3.716 55.601 4.082 ;
      RECT 55.5 3.727 55.515 4.088 ;
      RECT 55.43 3.75 55.5 4.094 ;
      RECT 55.375 3.782 55.43 4.102 ;
      RECT 55.335 3.805 55.375 4.108 ;
      RECT 55.321 3.818 55.335 4.111 ;
      RECT 55.235 3.84 55.321 4.117 ;
      RECT 55.22 3.865 55.235 4.123 ;
      RECT 55.18 3.88 55.22 4.127 ;
      RECT 55.13 3.895 55.18 4.132 ;
      RECT 55.105 3.902 55.13 4.136 ;
      RECT 55.045 3.897 55.105 4.14 ;
      RECT 55.03 3.888 55.045 4.144 ;
      RECT 54.96 3.878 55.03 4.14 ;
      RECT 54.935 3.87 54.955 4.13 ;
      RECT 54.876 3.87 54.935 4.108 ;
      RECT 54.79 3.87 54.876 4.065 ;
      RECT 54.955 3.87 54.96 4.135 ;
      RECT 55.65 3.101 55.82 3.435 ;
      RECT 55.62 3.101 55.82 3.43 ;
      RECT 55.56 3.068 55.62 3.418 ;
      RECT 55.56 3.124 55.83 3.413 ;
      RECT 55.535 3.124 55.83 3.407 ;
      RECT 55.53 3.065 55.56 3.404 ;
      RECT 55.515 3.071 55.65 3.402 ;
      RECT 55.51 3.079 55.735 3.39 ;
      RECT 55.51 3.131 55.845 3.343 ;
      RECT 55.495 3.087 55.735 3.338 ;
      RECT 55.495 3.157 55.855 3.279 ;
      RECT 55.465 3.107 55.82 3.24 ;
      RECT 55.465 3.197 55.865 3.236 ;
      RECT 55.515 3.076 55.735 3.402 ;
      RECT 54.855 3.406 54.91 3.67 ;
      RECT 54.855 3.406 54.975 3.669 ;
      RECT 54.855 3.406 55 3.668 ;
      RECT 54.855 3.406 55.065 3.667 ;
      RECT 55 3.372 55.08 3.666 ;
      RECT 54.815 3.416 55.225 3.665 ;
      RECT 54.855 3.413 55.225 3.665 ;
      RECT 54.815 3.421 55.23 3.658 ;
      RECT 54.8 3.423 55.23 3.657 ;
      RECT 54.8 3.43 55.235 3.653 ;
      RECT 54.78 3.429 55.23 3.649 ;
      RECT 54.78 3.437 55.24 3.648 ;
      RECT 54.775 3.434 55.235 3.644 ;
      RECT 54.775 3.447 55.25 3.643 ;
      RECT 54.76 3.437 55.24 3.642 ;
      RECT 54.725 3.45 55.25 3.635 ;
      RECT 54.91 3.405 55.22 3.665 ;
      RECT 54.91 3.39 55.17 3.665 ;
      RECT 54.975 3.377 55.105 3.665 ;
      RECT 54.52 4.466 54.535 4.859 ;
      RECT 54.485 4.471 54.535 4.858 ;
      RECT 54.52 4.47 54.58 4.857 ;
      RECT 54.465 4.481 54.58 4.856 ;
      RECT 54.48 4.477 54.58 4.856 ;
      RECT 54.445 4.487 54.655 4.853 ;
      RECT 54.445 4.506 54.7 4.851 ;
      RECT 54.445 4.513 54.705 4.848 ;
      RECT 54.43 4.49 54.655 4.845 ;
      RECT 54.41 4.495 54.655 4.838 ;
      RECT 54.405 4.499 54.655 4.834 ;
      RECT 54.405 4.516 54.715 4.833 ;
      RECT 54.385 4.51 54.7 4.829 ;
      RECT 54.385 4.519 54.72 4.823 ;
      RECT 54.38 4.525 54.72 4.595 ;
      RECT 54.445 4.485 54.58 4.853 ;
      RECT 54.32 3.848 54.52 4.16 ;
      RECT 54.395 3.826 54.52 4.16 ;
      RECT 54.335 3.845 54.525 4.145 ;
      RECT 54.305 3.856 54.525 4.143 ;
      RECT 54.32 3.851 54.53 4.109 ;
      RECT 54.305 3.955 54.535 4.076 ;
      RECT 54.335 3.827 54.52 4.16 ;
      RECT 54.395 3.805 54.495 4.16 ;
      RECT 54.42 3.802 54.495 4.16 ;
      RECT 54.42 3.797 54.44 4.16 ;
      RECT 53.825 3.865 54 4.04 ;
      RECT 53.82 3.865 54 4.038 ;
      RECT 53.795 3.865 54 4.033 ;
      RECT 53.74 3.845 53.91 4.023 ;
      RECT 53.74 3.852 53.975 4.023 ;
      RECT 53.825 4.532 53.84 4.715 ;
      RECT 53.815 4.51 53.825 4.715 ;
      RECT 53.8 4.49 53.815 4.715 ;
      RECT 53.79 4.465 53.8 4.715 ;
      RECT 53.76 4.43 53.79 4.715 ;
      RECT 53.725 4.37 53.76 4.715 ;
      RECT 53.72 4.332 53.725 4.715 ;
      RECT 53.67 4.283 53.72 4.715 ;
      RECT 53.66 4.233 53.67 4.703 ;
      RECT 53.645 4.212 53.66 4.663 ;
      RECT 53.625 4.18 53.645 4.613 ;
      RECT 53.6 4.136 53.625 4.553 ;
      RECT 53.595 4.108 53.6 4.508 ;
      RECT 53.59 4.099 53.595 4.494 ;
      RECT 53.585 4.092 53.59 4.481 ;
      RECT 53.58 4.087 53.585 4.47 ;
      RECT 53.575 4.072 53.58 4.46 ;
      RECT 53.57 4.05 53.575 4.447 ;
      RECT 53.56 4.01 53.57 4.422 ;
      RECT 53.535 3.94 53.56 4.378 ;
      RECT 53.53 3.88 53.535 4.343 ;
      RECT 53.515 3.86 53.53 4.31 ;
      RECT 53.51 3.86 53.515 4.285 ;
      RECT 53.48 3.86 53.51 4.24 ;
      RECT 53.435 3.86 53.48 4.18 ;
      RECT 53.36 3.86 53.435 4.128 ;
      RECT 53.355 3.86 53.36 4.093 ;
      RECT 53.35 3.86 53.355 4.083 ;
      RECT 53.345 3.86 53.35 4.063 ;
      RECT 53.61 3.08 53.78 3.55 ;
      RECT 53.555 3.073 53.75 3.534 ;
      RECT 53.555 3.087 53.785 3.533 ;
      RECT 53.54 3.088 53.785 3.514 ;
      RECT 53.535 3.106 53.785 3.5 ;
      RECT 53.54 3.089 53.79 3.498 ;
      RECT 53.525 3.12 53.79 3.483 ;
      RECT 53.54 3.095 53.795 3.468 ;
      RECT 53.52 3.135 53.795 3.465 ;
      RECT 53.535 3.107 53.8 3.45 ;
      RECT 53.535 3.119 53.805 3.43 ;
      RECT 53.52 3.135 53.81 3.413 ;
      RECT 53.52 3.145 53.815 3.268 ;
      RECT 53.515 3.145 53.815 3.225 ;
      RECT 53.515 3.16 53.82 3.203 ;
      RECT 53.61 3.07 53.75 3.55 ;
      RECT 53.61 3.068 53.72 3.55 ;
      RECT 53.696 3.065 53.72 3.55 ;
      RECT 53.355 4.732 53.36 4.778 ;
      RECT 53.345 4.58 53.355 4.802 ;
      RECT 53.34 4.425 53.345 4.827 ;
      RECT 53.325 4.387 53.34 4.838 ;
      RECT 53.32 4.37 53.325 4.845 ;
      RECT 53.31 4.358 53.32 4.852 ;
      RECT 53.305 4.349 53.31 4.854 ;
      RECT 53.3 4.347 53.305 4.858 ;
      RECT 53.255 4.338 53.3 4.873 ;
      RECT 53.25 4.33 53.255 4.887 ;
      RECT 53.245 4.327 53.25 4.891 ;
      RECT 53.23 4.322 53.245 4.899 ;
      RECT 53.175 4.312 53.23 4.91 ;
      RECT 53.14 4.3 53.175 4.911 ;
      RECT 53.131 4.295 53.14 4.905 ;
      RECT 53.045 4.295 53.131 4.895 ;
      RECT 53.015 4.295 53.045 4.873 ;
      RECT 53.005 4.295 53.01 4.853 ;
      RECT 53 4.295 53.005 4.815 ;
      RECT 52.995 4.295 53 4.773 ;
      RECT 52.99 4.295 52.995 4.733 ;
      RECT 52.985 4.295 52.99 4.663 ;
      RECT 52.975 4.295 52.985 4.585 ;
      RECT 52.97 4.295 52.975 4.485 ;
      RECT 53.01 4.295 53.015 4.855 ;
      RECT 52.505 4.377 52.595 4.855 ;
      RECT 52.49 4.38 52.61 4.853 ;
      RECT 52.505 4.379 52.61 4.853 ;
      RECT 52.47 4.386 52.635 4.843 ;
      RECT 52.49 4.38 52.635 4.843 ;
      RECT 52.455 4.392 52.635 4.831 ;
      RECT 52.49 4.383 52.685 4.824 ;
      RECT 52.441 4.4 52.685 4.822 ;
      RECT 52.47 4.39 52.695 4.81 ;
      RECT 52.441 4.411 52.725 4.801 ;
      RECT 52.355 4.435 52.725 4.795 ;
      RECT 52.355 4.448 52.765 4.778 ;
      RECT 52.35 4.47 52.765 4.771 ;
      RECT 52.32 4.485 52.765 4.761 ;
      RECT 52.315 4.496 52.765 4.751 ;
      RECT 52.285 4.509 52.765 4.742 ;
      RECT 52.27 4.527 52.765 4.731 ;
      RECT 52.245 4.54 52.765 4.721 ;
      RECT 52.505 4.376 52.515 4.855 ;
      RECT 52.551 3.8 52.59 4.045 ;
      RECT 52.465 3.8 52.6 4.043 ;
      RECT 52.35 3.825 52.6 4.04 ;
      RECT 52.35 3.825 52.605 4.038 ;
      RECT 52.35 3.825 52.62 4.033 ;
      RECT 52.456 3.8 52.635 4.013 ;
      RECT 52.37 3.808 52.635 4.013 ;
      RECT 52.04 3.16 52.21 3.595 ;
      RECT 52.03 3.194 52.21 3.578 ;
      RECT 52.11 3.13 52.28 3.565 ;
      RECT 52.015 3.205 52.28 3.543 ;
      RECT 52.11 3.14 52.285 3.533 ;
      RECT 52.04 3.192 52.315 3.518 ;
      RECT 52 3.218 52.315 3.503 ;
      RECT 52 3.26 52.325 3.483 ;
      RECT 51.995 3.285 52.33 3.465 ;
      RECT 51.995 3.295 52.335 3.45 ;
      RECT 51.99 3.232 52.315 3.448 ;
      RECT 51.99 3.305 52.34 3.433 ;
      RECT 51.985 3.242 52.315 3.43 ;
      RECT 51.98 3.326 52.345 3.413 ;
      RECT 51.98 3.358 52.35 3.393 ;
      RECT 51.975 3.272 52.325 3.385 ;
      RECT 51.98 3.257 52.315 3.413 ;
      RECT 51.995 3.227 52.315 3.465 ;
      RECT 51.84 3.814 52.065 4.07 ;
      RECT 51.84 3.847 52.085 4.06 ;
      RECT 51.805 3.847 52.085 4.058 ;
      RECT 51.805 3.86 52.09 4.048 ;
      RECT 51.805 3.88 52.1 4.04 ;
      RECT 51.805 3.977 52.105 4.033 ;
      RECT 51.785 3.725 51.915 4.023 ;
      RECT 51.74 3.88 52.1 3.965 ;
      RECT 51.73 3.725 51.915 3.91 ;
      RECT 51.73 3.757 52.001 3.91 ;
      RECT 51.695 4.287 51.715 4.465 ;
      RECT 51.66 4.24 51.695 4.465 ;
      RECT 51.645 4.18 51.66 4.465 ;
      RECT 51.62 4.127 51.645 4.465 ;
      RECT 51.605 4.08 51.62 4.465 ;
      RECT 51.585 4.057 51.605 4.465 ;
      RECT 51.56 4.022 51.585 4.465 ;
      RECT 51.55 3.868 51.56 4.465 ;
      RECT 51.52 3.863 51.55 4.456 ;
      RECT 51.515 3.86 51.52 4.446 ;
      RECT 51.5 3.86 51.515 4.42 ;
      RECT 51.495 3.86 51.5 4.383 ;
      RECT 51.47 3.86 51.495 4.335 ;
      RECT 51.45 3.86 51.47 4.26 ;
      RECT 51.44 3.86 51.45 4.22 ;
      RECT 51.435 3.86 51.44 4.195 ;
      RECT 51.43 3.86 51.435 4.178 ;
      RECT 51.425 3.86 51.43 4.16 ;
      RECT 51.42 3.861 51.425 4.15 ;
      RECT 51.41 3.863 51.42 4.118 ;
      RECT 51.4 3.865 51.41 4.085 ;
      RECT 51.39 3.868 51.4 4.058 ;
      RECT 51.715 4.295 51.94 4.465 ;
      RECT 51.045 3.107 51.215 3.56 ;
      RECT 51.045 3.107 51.305 3.526 ;
      RECT 51.045 3.107 51.335 3.51 ;
      RECT 51.045 3.107 51.365 3.483 ;
      RECT 51.301 3.085 51.38 3.465 ;
      RECT 51.08 3.092 51.385 3.45 ;
      RECT 51.08 3.1 51.395 3.413 ;
      RECT 51.04 3.127 51.395 3.385 ;
      RECT 51.025 3.14 51.395 3.35 ;
      RECT 51.045 3.115 51.415 3.34 ;
      RECT 51.02 3.18 51.415 3.31 ;
      RECT 51.02 3.21 51.42 3.293 ;
      RECT 51.015 3.24 51.42 3.28 ;
      RECT 51.08 3.089 51.38 3.465 ;
      RECT 51.215 3.086 51.301 3.544 ;
      RECT 51.166 3.087 51.38 3.465 ;
      RECT 51.31 4.747 51.355 4.94 ;
      RECT 51.3 4.717 51.31 4.94 ;
      RECT 51.295 4.702 51.3 4.94 ;
      RECT 51.255 4.612 51.295 4.94 ;
      RECT 51.25 4.525 51.255 4.94 ;
      RECT 51.24 4.495 51.25 4.94 ;
      RECT 51.235 4.455 51.24 4.94 ;
      RECT 51.225 4.417 51.235 4.94 ;
      RECT 51.22 4.382 51.225 4.94 ;
      RECT 51.2 4.335 51.22 4.94 ;
      RECT 51.185 4.26 51.2 4.94 ;
      RECT 51.18 4.215 51.185 4.935 ;
      RECT 51.175 4.195 51.18 4.908 ;
      RECT 51.17 4.175 51.175 4.893 ;
      RECT 51.165 4.15 51.17 4.873 ;
      RECT 51.16 4.128 51.165 4.858 ;
      RECT 51.155 4.106 51.16 4.84 ;
      RECT 51.15 4.085 51.155 4.83 ;
      RECT 51.14 4.057 51.15 4.8 ;
      RECT 51.13 4.02 51.14 4.768 ;
      RECT 51.12 3.98 51.13 4.735 ;
      RECT 51.11 3.958 51.12 4.705 ;
      RECT 51.08 3.91 51.11 4.637 ;
      RECT 51.065 3.87 51.08 4.564 ;
      RECT 51.055 3.87 51.065 4.53 ;
      RECT 51.05 3.87 51.055 4.505 ;
      RECT 51.045 3.87 51.05 4.49 ;
      RECT 51.04 3.87 51.045 4.468 ;
      RECT 51.035 3.87 51.04 4.455 ;
      RECT 51.02 3.87 51.035 4.42 ;
      RECT 51 3.87 51.02 4.36 ;
      RECT 50.99 3.87 51 4.31 ;
      RECT 50.97 3.87 50.99 4.258 ;
      RECT 50.95 3.87 50.97 4.215 ;
      RECT 50.94 3.87 50.95 4.203 ;
      RECT 50.91 3.87 50.94 4.19 ;
      RECT 50.88 3.891 50.91 4.17 ;
      RECT 50.87 3.919 50.88 4.15 ;
      RECT 50.855 3.936 50.87 4.118 ;
      RECT 50.85 3.95 50.855 4.085 ;
      RECT 50.845 3.958 50.85 4.058 ;
      RECT 50.84 3.966 50.845 4.02 ;
      RECT 50.845 4.49 50.85 4.825 ;
      RECT 50.81 4.477 50.845 4.824 ;
      RECT 50.74 4.417 50.81 4.823 ;
      RECT 50.66 4.36 50.74 4.822 ;
      RECT 50.525 4.32 50.66 4.821 ;
      RECT 50.525 4.507 50.86 4.81 ;
      RECT 50.485 4.507 50.86 4.8 ;
      RECT 50.485 4.525 50.865 4.795 ;
      RECT 50.485 4.615 50.87 4.785 ;
      RECT 50.48 4.31 50.645 4.765 ;
      RECT 50.475 4.31 50.645 4.508 ;
      RECT 50.475 4.467 50.84 4.508 ;
      RECT 50.475 4.455 50.835 4.508 ;
      RECT 49.605 7.305 49.775 8.775 ;
      RECT 49.605 8.6 49.78 8.77 ;
      RECT 49.235 3.035 49.405 4.225 ;
      RECT 49.235 3.035 49.705 3.205 ;
      RECT 49.235 9.255 49.705 9.425 ;
      RECT 49.235 8.235 49.405 9.425 ;
      RECT 48.245 3.035 48.415 4.225 ;
      RECT 48.245 3.035 48.715 3.205 ;
      RECT 48.245 9.255 48.715 9.425 ;
      RECT 48.245 8.235 48.415 9.425 ;
      RECT 46.395 3.93 46.565 5.16 ;
      RECT 46.45 2.15 46.62 4.1 ;
      RECT 46.395 1.87 46.565 2.32 ;
      RECT 46.395 10.14 46.565 10.59 ;
      RECT 46.45 8.36 46.62 10.31 ;
      RECT 46.395 7.3 46.565 8.53 ;
      RECT 45.875 1.87 46.045 5.16 ;
      RECT 45.875 3.37 46.28 3.7 ;
      RECT 45.875 2.53 46.28 2.86 ;
      RECT 45.875 7.3 46.045 10.59 ;
      RECT 45.875 9.6 46.28 9.93 ;
      RECT 45.875 8.76 46.28 9.09 ;
      RECT 43.21 3.27 43.94 3.51 ;
      RECT 43.752 3.065 43.94 3.51 ;
      RECT 43.58 3.077 43.955 3.504 ;
      RECT 43.495 3.092 43.975 3.489 ;
      RECT 43.495 3.107 43.98 3.479 ;
      RECT 43.45 3.127 43.995 3.471 ;
      RECT 43.427 3.162 44.01 3.425 ;
      RECT 43.341 3.185 44.015 3.385 ;
      RECT 43.341 3.203 44.025 3.355 ;
      RECT 43.21 3.272 44.03 3.318 ;
      RECT 43.255 3.215 44.025 3.355 ;
      RECT 43.341 3.167 44.01 3.425 ;
      RECT 43.427 3.136 43.995 3.471 ;
      RECT 43.45 3.117 43.98 3.479 ;
      RECT 43.495 3.09 43.955 3.504 ;
      RECT 43.58 3.072 43.94 3.51 ;
      RECT 43.666 3.066 43.94 3.51 ;
      RECT 43.752 3.061 43.885 3.51 ;
      RECT 43.838 3.056 43.885 3.51 ;
      RECT 43.53 3.954 43.7 4.34 ;
      RECT 43.525 3.954 43.7 4.335 ;
      RECT 43.5 3.954 43.7 4.3 ;
      RECT 43.5 3.982 43.71 4.29 ;
      RECT 43.48 3.982 43.71 4.25 ;
      RECT 43.475 3.982 43.71 4.223 ;
      RECT 43.475 4 43.715 4.215 ;
      RECT 43.42 4 43.715 4.15 ;
      RECT 43.42 4.017 43.725 4.133 ;
      RECT 43.41 4.017 43.725 4.073 ;
      RECT 43.41 4.034 43.73 4.07 ;
      RECT 43.405 3.87 43.575 4.048 ;
      RECT 43.405 3.904 43.661 4.048 ;
      RECT 43.4 4.67 43.405 4.683 ;
      RECT 43.395 4.565 43.4 4.688 ;
      RECT 43.37 4.425 43.395 4.703 ;
      RECT 43.335 4.376 43.37 4.735 ;
      RECT 43.33 4.344 43.335 4.755 ;
      RECT 43.325 4.335 43.33 4.755 ;
      RECT 43.245 4.3 43.325 4.755 ;
      RECT 43.182 4.27 43.245 4.755 ;
      RECT 43.096 4.258 43.182 4.755 ;
      RECT 43.01 4.244 43.096 4.755 ;
      RECT 42.93 4.231 43.01 4.741 ;
      RECT 42.895 4.223 42.93 4.721 ;
      RECT 42.885 4.22 42.895 4.712 ;
      RECT 42.855 4.215 42.885 4.699 ;
      RECT 42.805 4.19 42.855 4.675 ;
      RECT 42.791 4.164 42.805 4.657 ;
      RECT 42.705 4.124 42.791 4.633 ;
      RECT 42.66 4.072 42.705 4.602 ;
      RECT 42.65 4.047 42.66 4.589 ;
      RECT 42.645 3.828 42.65 3.85 ;
      RECT 42.64 4.03 42.65 4.585 ;
      RECT 42.64 3.826 42.645 3.94 ;
      RECT 42.63 3.822 42.64 4.581 ;
      RECT 42.586 3.82 42.63 4.569 ;
      RECT 42.5 3.82 42.586 4.54 ;
      RECT 42.47 3.82 42.5 4.513 ;
      RECT 42.455 3.82 42.47 4.501 ;
      RECT 42.415 3.832 42.455 4.486 ;
      RECT 42.395 3.851 42.415 4.465 ;
      RECT 42.385 3.861 42.395 4.449 ;
      RECT 42.375 3.867 42.385 4.438 ;
      RECT 42.355 3.877 42.375 4.421 ;
      RECT 42.35 3.886 42.355 4.408 ;
      RECT 42.345 3.89 42.35 4.358 ;
      RECT 42.335 3.896 42.345 4.275 ;
      RECT 42.33 3.9 42.335 4.189 ;
      RECT 42.325 3.92 42.33 4.126 ;
      RECT 42.32 3.943 42.325 4.073 ;
      RECT 42.315 3.961 42.32 4.018 ;
      RECT 42.925 3.78 43.095 4.04 ;
      RECT 43.095 3.745 43.14 4.026 ;
      RECT 43.056 3.747 43.145 4.009 ;
      RECT 42.945 3.764 43.231 3.98 ;
      RECT 42.945 3.779 43.235 3.952 ;
      RECT 42.945 3.76 43.145 4.009 ;
      RECT 42.97 3.748 43.095 4.04 ;
      RECT 43.056 3.746 43.14 4.026 ;
      RECT 42.11 3.135 42.28 3.625 ;
      RECT 42.11 3.135 42.315 3.605 ;
      RECT 42.245 3.055 42.355 3.565 ;
      RECT 42.226 3.059 42.375 3.535 ;
      RECT 42.14 3.067 42.395 3.518 ;
      RECT 42.14 3.073 42.4 3.508 ;
      RECT 42.14 3.082 42.42 3.496 ;
      RECT 42.115 3.107 42.45 3.474 ;
      RECT 42.115 3.127 42.455 3.454 ;
      RECT 42.11 3.14 42.465 3.434 ;
      RECT 42.11 3.207 42.47 3.415 ;
      RECT 42.11 3.34 42.475 3.402 ;
      RECT 42.105 3.145 42.465 3.235 ;
      RECT 42.115 3.102 42.42 3.496 ;
      RECT 42.226 3.057 42.355 3.565 ;
      RECT 42.1 4.81 42.4 5.065 ;
      RECT 42.185 4.776 42.4 5.065 ;
      RECT 42.185 4.779 42.405 4.925 ;
      RECT 42.12 4.8 42.405 4.925 ;
      RECT 42.155 4.79 42.4 5.065 ;
      RECT 42.15 4.795 42.405 4.925 ;
      RECT 42.185 4.774 42.386 5.065 ;
      RECT 42.271 4.765 42.386 5.065 ;
      RECT 42.271 4.759 42.3 5.065 ;
      RECT 41.76 4.4 41.77 4.89 ;
      RECT 41.42 4.335 41.43 4.635 ;
      RECT 41.935 4.507 41.94 4.726 ;
      RECT 41.925 4.487 41.935 4.743 ;
      RECT 41.915 4.467 41.925 4.773 ;
      RECT 41.91 4.457 41.915 4.788 ;
      RECT 41.905 4.453 41.91 4.793 ;
      RECT 41.89 4.445 41.905 4.8 ;
      RECT 41.85 4.425 41.89 4.825 ;
      RECT 41.825 4.407 41.85 4.858 ;
      RECT 41.82 4.405 41.825 4.871 ;
      RECT 41.8 4.402 41.82 4.875 ;
      RECT 41.77 4.4 41.8 4.885 ;
      RECT 41.7 4.402 41.76 4.886 ;
      RECT 41.68 4.402 41.7 4.88 ;
      RECT 41.655 4.4 41.68 4.877 ;
      RECT 41.62 4.395 41.655 4.873 ;
      RECT 41.6 4.389 41.62 4.86 ;
      RECT 41.59 4.386 41.6 4.848 ;
      RECT 41.57 4.383 41.59 4.833 ;
      RECT 41.55 4.379 41.57 4.815 ;
      RECT 41.545 4.376 41.55 4.805 ;
      RECT 41.54 4.375 41.545 4.803 ;
      RECT 41.53 4.372 41.54 4.795 ;
      RECT 41.52 4.366 41.53 4.778 ;
      RECT 41.51 4.36 41.52 4.76 ;
      RECT 41.5 4.354 41.51 4.748 ;
      RECT 41.49 4.348 41.5 4.728 ;
      RECT 41.485 4.344 41.49 4.713 ;
      RECT 41.48 4.342 41.485 4.705 ;
      RECT 41.475 4.34 41.48 4.698 ;
      RECT 41.47 4.338 41.475 4.688 ;
      RECT 41.465 4.336 41.47 4.682 ;
      RECT 41.455 4.335 41.465 4.672 ;
      RECT 41.445 4.335 41.455 4.663 ;
      RECT 41.43 4.335 41.445 4.648 ;
      RECT 41.39 4.335 41.42 4.632 ;
      RECT 41.37 4.337 41.39 4.627 ;
      RECT 41.365 4.342 41.37 4.625 ;
      RECT 41.335 4.35 41.365 4.623 ;
      RECT 41.305 4.365 41.335 4.622 ;
      RECT 41.26 4.387 41.305 4.627 ;
      RECT 41.255 4.402 41.26 4.631 ;
      RECT 41.24 4.407 41.255 4.633 ;
      RECT 41.235 4.411 41.24 4.635 ;
      RECT 41.175 4.434 41.235 4.644 ;
      RECT 41.155 4.46 41.175 4.657 ;
      RECT 41.145 4.467 41.155 4.661 ;
      RECT 41.13 4.474 41.145 4.664 ;
      RECT 41.11 4.484 41.13 4.667 ;
      RECT 41.105 4.492 41.11 4.67 ;
      RECT 41.06 4.497 41.105 4.677 ;
      RECT 41.05 4.5 41.06 4.684 ;
      RECT 41.04 4.5 41.05 4.688 ;
      RECT 41.005 4.502 41.04 4.7 ;
      RECT 40.985 4.505 41.005 4.713 ;
      RECT 40.945 4.508 40.985 4.724 ;
      RECT 40.93 4.51 40.945 4.737 ;
      RECT 40.92 4.51 40.93 4.742 ;
      RECT 40.895 4.511 40.92 4.75 ;
      RECT 40.885 4.513 40.895 4.755 ;
      RECT 40.88 4.514 40.885 4.758 ;
      RECT 40.855 4.512 40.88 4.761 ;
      RECT 40.84 4.51 40.855 4.762 ;
      RECT 40.82 4.507 40.84 4.764 ;
      RECT 40.8 4.502 40.82 4.764 ;
      RECT 40.74 4.497 40.8 4.761 ;
      RECT 40.705 4.472 40.74 4.757 ;
      RECT 40.695 4.449 40.705 4.755 ;
      RECT 40.665 4.426 40.695 4.755 ;
      RECT 40.655 4.405 40.665 4.755 ;
      RECT 40.63 4.387 40.655 4.753 ;
      RECT 40.615 4.365 40.63 4.75 ;
      RECT 40.6 4.347 40.615 4.748 ;
      RECT 40.58 4.337 40.6 4.746 ;
      RECT 40.565 4.332 40.58 4.745 ;
      RECT 40.55 4.33 40.565 4.744 ;
      RECT 40.52 4.331 40.55 4.742 ;
      RECT 40.5 4.334 40.52 4.74 ;
      RECT 40.443 4.338 40.5 4.74 ;
      RECT 40.357 4.347 40.443 4.74 ;
      RECT 40.271 4.358 40.357 4.74 ;
      RECT 40.185 4.369 40.271 4.74 ;
      RECT 40.165 4.376 40.185 4.748 ;
      RECT 40.155 4.379 40.165 4.755 ;
      RECT 40.09 4.384 40.155 4.773 ;
      RECT 40.06 4.391 40.09 4.798 ;
      RECT 40.05 4.394 40.06 4.805 ;
      RECT 40.005 4.398 40.05 4.81 ;
      RECT 39.975 4.403 40.005 4.815 ;
      RECT 39.974 4.405 39.975 4.815 ;
      RECT 39.888 4.411 39.974 4.815 ;
      RECT 39.802 4.422 39.888 4.815 ;
      RECT 39.716 4.434 39.802 4.815 ;
      RECT 39.63 4.445 39.716 4.815 ;
      RECT 39.615 4.452 39.63 4.81 ;
      RECT 39.61 4.454 39.615 4.804 ;
      RECT 39.59 4.465 39.61 4.799 ;
      RECT 39.58 4.483 39.59 4.793 ;
      RECT 39.575 4.495 39.58 4.593 ;
      RECT 41.87 3.248 41.89 3.335 ;
      RECT 41.865 3.183 41.87 3.367 ;
      RECT 41.855 3.15 41.865 3.372 ;
      RECT 41.85 3.13 41.855 3.378 ;
      RECT 41.82 3.13 41.85 3.395 ;
      RECT 41.771 3.13 41.82 3.431 ;
      RECT 41.685 3.13 41.771 3.489 ;
      RECT 41.656 3.14 41.685 3.538 ;
      RECT 41.57 3.182 41.656 3.591 ;
      RECT 41.55 3.22 41.57 3.638 ;
      RECT 41.525 3.237 41.55 3.658 ;
      RECT 41.515 3.251 41.525 3.678 ;
      RECT 41.51 3.257 41.515 3.688 ;
      RECT 41.505 3.261 41.51 3.695 ;
      RECT 41.455 3.281 41.505 3.7 ;
      RECT 41.39 3.325 41.455 3.7 ;
      RECT 41.365 3.375 41.39 3.7 ;
      RECT 41.355 3.405 41.365 3.7 ;
      RECT 41.35 3.432 41.355 3.7 ;
      RECT 41.345 3.45 41.35 3.7 ;
      RECT 41.335 3.492 41.345 3.7 ;
      RECT 41.685 4.05 41.855 4.225 ;
      RECT 41.625 3.878 41.685 4.213 ;
      RECT 41.615 3.871 41.625 4.196 ;
      RECT 41.57 4.05 41.855 4.176 ;
      RECT 41.551 4.05 41.855 4.154 ;
      RECT 41.465 4.05 41.855 4.119 ;
      RECT 41.445 3.87 41.615 4.075 ;
      RECT 41.445 4.017 41.85 4.075 ;
      RECT 41.445 3.965 41.825 4.075 ;
      RECT 41.445 3.92 41.79 4.075 ;
      RECT 41.445 3.902 41.755 4.075 ;
      RECT 41.445 3.892 41.75 4.075 ;
      RECT 41.095 7.3 41.265 10.59 ;
      RECT 41.095 9.6 41.5 9.93 ;
      RECT 41.095 8.76 41.5 9.09 ;
      RECT 41.165 4.85 41.355 5.075 ;
      RECT 41.155 4.851 41.36 5.07 ;
      RECT 41.155 4.853 41.37 5.05 ;
      RECT 41.155 4.857 41.375 5.035 ;
      RECT 41.155 4.844 41.325 5.07 ;
      RECT 41.155 4.847 41.35 5.07 ;
      RECT 41.165 4.843 41.325 5.075 ;
      RECT 41.251 4.841 41.325 5.075 ;
      RECT 40.875 4.092 41.045 4.33 ;
      RECT 40.875 4.092 41.131 4.244 ;
      RECT 40.875 4.092 41.135 4.154 ;
      RECT 40.925 3.865 41.145 4.133 ;
      RECT 40.92 3.882 41.15 4.106 ;
      RECT 40.885 4.04 41.15 4.106 ;
      RECT 40.905 3.89 41.045 4.33 ;
      RECT 40.895 3.972 41.155 4.089 ;
      RECT 40.89 4.02 41.155 4.089 ;
      RECT 40.895 3.93 41.15 4.106 ;
      RECT 40.92 3.867 41.145 4.133 ;
      RECT 40.485 3.842 40.655 4.04 ;
      RECT 40.485 3.842 40.7 4.015 ;
      RECT 40.555 3.785 40.725 3.973 ;
      RECT 40.53 3.8 40.725 3.973 ;
      RECT 40.145 3.846 40.175 4.04 ;
      RECT 40.14 3.818 40.145 4.04 ;
      RECT 40.11 3.792 40.14 4.042 ;
      RECT 40.085 3.75 40.11 4.045 ;
      RECT 40.075 3.722 40.085 4.047 ;
      RECT 40.04 3.702 40.075 4.049 ;
      RECT 39.975 3.687 40.04 4.055 ;
      RECT 39.925 3.685 39.975 4.061 ;
      RECT 39.902 3.687 39.925 4.066 ;
      RECT 39.816 3.698 39.902 4.072 ;
      RECT 39.73 3.716 39.816 4.082 ;
      RECT 39.715 3.727 39.73 4.088 ;
      RECT 39.645 3.75 39.715 4.094 ;
      RECT 39.59 3.782 39.645 4.102 ;
      RECT 39.55 3.805 39.59 4.108 ;
      RECT 39.536 3.818 39.55 4.111 ;
      RECT 39.45 3.84 39.536 4.117 ;
      RECT 39.435 3.865 39.45 4.123 ;
      RECT 39.395 3.88 39.435 4.127 ;
      RECT 39.345 3.895 39.395 4.132 ;
      RECT 39.32 3.902 39.345 4.136 ;
      RECT 39.26 3.897 39.32 4.14 ;
      RECT 39.245 3.888 39.26 4.144 ;
      RECT 39.175 3.878 39.245 4.14 ;
      RECT 39.15 3.87 39.17 4.13 ;
      RECT 39.091 3.87 39.15 4.108 ;
      RECT 39.005 3.87 39.091 4.065 ;
      RECT 39.17 3.87 39.175 4.135 ;
      RECT 39.865 3.101 40.035 3.435 ;
      RECT 39.835 3.101 40.035 3.43 ;
      RECT 39.775 3.068 39.835 3.418 ;
      RECT 39.775 3.124 40.045 3.413 ;
      RECT 39.75 3.124 40.045 3.407 ;
      RECT 39.745 3.065 39.775 3.404 ;
      RECT 39.73 3.071 39.865 3.402 ;
      RECT 39.725 3.079 39.95 3.39 ;
      RECT 39.725 3.131 40.06 3.343 ;
      RECT 39.71 3.087 39.95 3.338 ;
      RECT 39.71 3.157 40.07 3.279 ;
      RECT 39.68 3.107 40.035 3.24 ;
      RECT 39.68 3.197 40.08 3.236 ;
      RECT 39.73 3.076 39.95 3.402 ;
      RECT 39.07 3.406 39.125 3.67 ;
      RECT 39.07 3.406 39.19 3.669 ;
      RECT 39.07 3.406 39.215 3.668 ;
      RECT 39.07 3.406 39.28 3.667 ;
      RECT 39.215 3.372 39.295 3.666 ;
      RECT 39.03 3.416 39.44 3.665 ;
      RECT 39.07 3.413 39.44 3.665 ;
      RECT 39.03 3.421 39.445 3.658 ;
      RECT 39.015 3.423 39.445 3.657 ;
      RECT 39.015 3.43 39.45 3.653 ;
      RECT 38.995 3.429 39.445 3.649 ;
      RECT 38.995 3.437 39.455 3.648 ;
      RECT 38.99 3.434 39.45 3.644 ;
      RECT 38.99 3.447 39.465 3.643 ;
      RECT 38.975 3.437 39.455 3.642 ;
      RECT 38.94 3.45 39.465 3.635 ;
      RECT 39.125 3.405 39.435 3.665 ;
      RECT 39.125 3.39 39.385 3.665 ;
      RECT 39.19 3.377 39.32 3.665 ;
      RECT 38.735 4.466 38.75 4.859 ;
      RECT 38.7 4.471 38.75 4.858 ;
      RECT 38.735 4.47 38.795 4.857 ;
      RECT 38.68 4.481 38.795 4.856 ;
      RECT 38.695 4.477 38.795 4.856 ;
      RECT 38.66 4.487 38.87 4.853 ;
      RECT 38.66 4.506 38.915 4.851 ;
      RECT 38.66 4.513 38.92 4.848 ;
      RECT 38.645 4.49 38.87 4.845 ;
      RECT 38.625 4.495 38.87 4.838 ;
      RECT 38.62 4.499 38.87 4.834 ;
      RECT 38.62 4.516 38.93 4.833 ;
      RECT 38.6 4.51 38.915 4.829 ;
      RECT 38.6 4.519 38.935 4.823 ;
      RECT 38.595 4.525 38.935 4.595 ;
      RECT 38.66 4.485 38.795 4.853 ;
      RECT 38.535 3.848 38.735 4.16 ;
      RECT 38.61 3.826 38.735 4.16 ;
      RECT 38.55 3.845 38.74 4.145 ;
      RECT 38.52 3.856 38.74 4.143 ;
      RECT 38.535 3.851 38.745 4.109 ;
      RECT 38.52 3.955 38.75 4.076 ;
      RECT 38.55 3.827 38.735 4.16 ;
      RECT 38.61 3.805 38.71 4.16 ;
      RECT 38.635 3.802 38.71 4.16 ;
      RECT 38.635 3.797 38.655 4.16 ;
      RECT 38.04 3.865 38.215 4.04 ;
      RECT 38.035 3.865 38.215 4.038 ;
      RECT 38.01 3.865 38.215 4.033 ;
      RECT 37.955 3.845 38.125 4.023 ;
      RECT 37.955 3.852 38.19 4.023 ;
      RECT 38.04 4.532 38.055 4.715 ;
      RECT 38.03 4.51 38.04 4.715 ;
      RECT 38.015 4.49 38.03 4.715 ;
      RECT 38.005 4.465 38.015 4.715 ;
      RECT 37.975 4.43 38.005 4.715 ;
      RECT 37.94 4.37 37.975 4.715 ;
      RECT 37.935 4.332 37.94 4.715 ;
      RECT 37.885 4.283 37.935 4.715 ;
      RECT 37.875 4.233 37.885 4.703 ;
      RECT 37.86 4.212 37.875 4.663 ;
      RECT 37.84 4.18 37.86 4.613 ;
      RECT 37.815 4.136 37.84 4.553 ;
      RECT 37.81 4.108 37.815 4.508 ;
      RECT 37.805 4.099 37.81 4.494 ;
      RECT 37.8 4.092 37.805 4.481 ;
      RECT 37.795 4.087 37.8 4.47 ;
      RECT 37.79 4.072 37.795 4.46 ;
      RECT 37.785 4.05 37.79 4.447 ;
      RECT 37.775 4.01 37.785 4.422 ;
      RECT 37.75 3.94 37.775 4.378 ;
      RECT 37.745 3.88 37.75 4.343 ;
      RECT 37.73 3.86 37.745 4.31 ;
      RECT 37.725 3.86 37.73 4.285 ;
      RECT 37.695 3.86 37.725 4.24 ;
      RECT 37.65 3.86 37.695 4.18 ;
      RECT 37.575 3.86 37.65 4.128 ;
      RECT 37.57 3.86 37.575 4.093 ;
      RECT 37.565 3.86 37.57 4.083 ;
      RECT 37.56 3.86 37.565 4.063 ;
      RECT 37.825 3.08 37.995 3.55 ;
      RECT 37.77 3.073 37.965 3.534 ;
      RECT 37.77 3.087 38 3.533 ;
      RECT 37.755 3.088 38 3.514 ;
      RECT 37.75 3.106 38 3.5 ;
      RECT 37.755 3.089 38.005 3.498 ;
      RECT 37.74 3.12 38.005 3.483 ;
      RECT 37.755 3.095 38.01 3.468 ;
      RECT 37.735 3.135 38.01 3.465 ;
      RECT 37.75 3.107 38.015 3.45 ;
      RECT 37.75 3.119 38.02 3.43 ;
      RECT 37.735 3.135 38.025 3.413 ;
      RECT 37.735 3.145 38.03 3.268 ;
      RECT 37.73 3.145 38.03 3.225 ;
      RECT 37.73 3.16 38.035 3.203 ;
      RECT 37.825 3.07 37.965 3.55 ;
      RECT 37.825 3.068 37.935 3.55 ;
      RECT 37.911 3.065 37.935 3.55 ;
      RECT 37.57 4.732 37.575 4.778 ;
      RECT 37.56 4.58 37.57 4.802 ;
      RECT 37.555 4.425 37.56 4.827 ;
      RECT 37.54 4.387 37.555 4.838 ;
      RECT 37.535 4.37 37.54 4.845 ;
      RECT 37.525 4.358 37.535 4.852 ;
      RECT 37.52 4.349 37.525 4.854 ;
      RECT 37.515 4.347 37.52 4.858 ;
      RECT 37.47 4.338 37.515 4.873 ;
      RECT 37.465 4.33 37.47 4.887 ;
      RECT 37.46 4.327 37.465 4.891 ;
      RECT 37.445 4.322 37.46 4.899 ;
      RECT 37.39 4.312 37.445 4.91 ;
      RECT 37.355 4.3 37.39 4.911 ;
      RECT 37.346 4.295 37.355 4.905 ;
      RECT 37.26 4.295 37.346 4.895 ;
      RECT 37.23 4.295 37.26 4.873 ;
      RECT 37.22 4.295 37.225 4.853 ;
      RECT 37.215 4.295 37.22 4.815 ;
      RECT 37.21 4.295 37.215 4.773 ;
      RECT 37.205 4.295 37.21 4.733 ;
      RECT 37.2 4.295 37.205 4.663 ;
      RECT 37.19 4.295 37.2 4.585 ;
      RECT 37.185 4.295 37.19 4.485 ;
      RECT 37.225 4.295 37.23 4.855 ;
      RECT 36.72 4.377 36.81 4.855 ;
      RECT 36.705 4.38 36.825 4.853 ;
      RECT 36.72 4.379 36.825 4.853 ;
      RECT 36.685 4.386 36.85 4.843 ;
      RECT 36.705 4.38 36.85 4.843 ;
      RECT 36.67 4.392 36.85 4.831 ;
      RECT 36.705 4.383 36.9 4.824 ;
      RECT 36.656 4.4 36.9 4.822 ;
      RECT 36.685 4.39 36.91 4.81 ;
      RECT 36.656 4.411 36.94 4.801 ;
      RECT 36.57 4.435 36.94 4.795 ;
      RECT 36.57 4.448 36.98 4.778 ;
      RECT 36.565 4.47 36.98 4.771 ;
      RECT 36.535 4.485 36.98 4.761 ;
      RECT 36.53 4.496 36.98 4.751 ;
      RECT 36.5 4.509 36.98 4.742 ;
      RECT 36.485 4.527 36.98 4.731 ;
      RECT 36.46 4.54 36.98 4.721 ;
      RECT 36.72 4.376 36.73 4.855 ;
      RECT 36.766 3.8 36.805 4.045 ;
      RECT 36.68 3.8 36.815 4.043 ;
      RECT 36.565 3.825 36.815 4.04 ;
      RECT 36.565 3.825 36.82 4.038 ;
      RECT 36.565 3.825 36.835 4.033 ;
      RECT 36.671 3.8 36.85 4.013 ;
      RECT 36.585 3.808 36.85 4.013 ;
      RECT 36.255 3.16 36.425 3.595 ;
      RECT 36.245 3.194 36.425 3.578 ;
      RECT 36.325 3.13 36.495 3.565 ;
      RECT 36.23 3.205 36.495 3.543 ;
      RECT 36.325 3.14 36.5 3.533 ;
      RECT 36.255 3.192 36.53 3.518 ;
      RECT 36.215 3.218 36.53 3.503 ;
      RECT 36.215 3.26 36.54 3.483 ;
      RECT 36.21 3.285 36.545 3.465 ;
      RECT 36.21 3.295 36.55 3.45 ;
      RECT 36.205 3.232 36.53 3.448 ;
      RECT 36.205 3.305 36.555 3.433 ;
      RECT 36.2 3.242 36.53 3.43 ;
      RECT 36.195 3.326 36.56 3.413 ;
      RECT 36.195 3.358 36.565 3.393 ;
      RECT 36.19 3.272 36.54 3.385 ;
      RECT 36.195 3.257 36.53 3.413 ;
      RECT 36.21 3.227 36.53 3.465 ;
      RECT 36.055 3.814 36.28 4.07 ;
      RECT 36.055 3.847 36.3 4.06 ;
      RECT 36.02 3.847 36.3 4.058 ;
      RECT 36.02 3.86 36.305 4.048 ;
      RECT 36.02 3.88 36.315 4.04 ;
      RECT 36.02 3.977 36.32 4.033 ;
      RECT 36 3.725 36.13 4.023 ;
      RECT 35.955 3.88 36.315 3.965 ;
      RECT 35.945 3.725 36.13 3.91 ;
      RECT 35.945 3.757 36.216 3.91 ;
      RECT 35.91 4.287 35.93 4.465 ;
      RECT 35.875 4.24 35.91 4.465 ;
      RECT 35.86 4.18 35.875 4.465 ;
      RECT 35.835 4.127 35.86 4.465 ;
      RECT 35.82 4.08 35.835 4.465 ;
      RECT 35.8 4.057 35.82 4.465 ;
      RECT 35.775 4.022 35.8 4.465 ;
      RECT 35.765 3.868 35.775 4.465 ;
      RECT 35.735 3.863 35.765 4.456 ;
      RECT 35.73 3.86 35.735 4.446 ;
      RECT 35.715 3.86 35.73 4.42 ;
      RECT 35.71 3.86 35.715 4.383 ;
      RECT 35.685 3.86 35.71 4.335 ;
      RECT 35.665 3.86 35.685 4.26 ;
      RECT 35.655 3.86 35.665 4.22 ;
      RECT 35.65 3.86 35.655 4.195 ;
      RECT 35.645 3.86 35.65 4.178 ;
      RECT 35.64 3.86 35.645 4.16 ;
      RECT 35.635 3.861 35.64 4.15 ;
      RECT 35.625 3.863 35.635 4.118 ;
      RECT 35.615 3.865 35.625 4.085 ;
      RECT 35.605 3.868 35.615 4.058 ;
      RECT 35.93 4.295 36.155 4.465 ;
      RECT 35.26 3.107 35.43 3.56 ;
      RECT 35.26 3.107 35.52 3.526 ;
      RECT 35.26 3.107 35.55 3.51 ;
      RECT 35.26 3.107 35.58 3.483 ;
      RECT 35.516 3.085 35.595 3.465 ;
      RECT 35.295 3.092 35.6 3.45 ;
      RECT 35.295 3.1 35.61 3.413 ;
      RECT 35.255 3.127 35.61 3.385 ;
      RECT 35.24 3.14 35.61 3.35 ;
      RECT 35.26 3.115 35.63 3.34 ;
      RECT 35.235 3.18 35.63 3.31 ;
      RECT 35.235 3.21 35.635 3.293 ;
      RECT 35.23 3.24 35.635 3.28 ;
      RECT 35.295 3.089 35.595 3.465 ;
      RECT 35.43 3.086 35.516 3.544 ;
      RECT 35.381 3.087 35.595 3.465 ;
      RECT 35.525 4.747 35.57 4.94 ;
      RECT 35.515 4.717 35.525 4.94 ;
      RECT 35.51 4.702 35.515 4.94 ;
      RECT 35.47 4.612 35.51 4.94 ;
      RECT 35.465 4.525 35.47 4.94 ;
      RECT 35.455 4.495 35.465 4.94 ;
      RECT 35.45 4.455 35.455 4.94 ;
      RECT 35.44 4.417 35.45 4.94 ;
      RECT 35.435 4.382 35.44 4.94 ;
      RECT 35.415 4.335 35.435 4.94 ;
      RECT 35.4 4.26 35.415 4.94 ;
      RECT 35.395 4.215 35.4 4.935 ;
      RECT 35.39 4.195 35.395 4.908 ;
      RECT 35.385 4.175 35.39 4.893 ;
      RECT 35.38 4.15 35.385 4.873 ;
      RECT 35.375 4.128 35.38 4.858 ;
      RECT 35.37 4.106 35.375 4.84 ;
      RECT 35.365 4.085 35.37 4.83 ;
      RECT 35.355 4.057 35.365 4.8 ;
      RECT 35.345 4.02 35.355 4.768 ;
      RECT 35.335 3.98 35.345 4.735 ;
      RECT 35.325 3.958 35.335 4.705 ;
      RECT 35.295 3.91 35.325 4.637 ;
      RECT 35.28 3.87 35.295 4.564 ;
      RECT 35.27 3.87 35.28 4.53 ;
      RECT 35.265 3.87 35.27 4.505 ;
      RECT 35.26 3.87 35.265 4.49 ;
      RECT 35.255 3.87 35.26 4.468 ;
      RECT 35.25 3.87 35.255 4.455 ;
      RECT 35.235 3.87 35.25 4.42 ;
      RECT 35.215 3.87 35.235 4.36 ;
      RECT 35.205 3.87 35.215 4.31 ;
      RECT 35.185 3.87 35.205 4.258 ;
      RECT 35.165 3.87 35.185 4.215 ;
      RECT 35.155 3.87 35.165 4.203 ;
      RECT 35.125 3.87 35.155 4.19 ;
      RECT 35.095 3.891 35.125 4.17 ;
      RECT 35.085 3.919 35.095 4.15 ;
      RECT 35.07 3.936 35.085 4.118 ;
      RECT 35.065 3.95 35.07 4.085 ;
      RECT 35.06 3.958 35.065 4.058 ;
      RECT 35.055 3.966 35.06 4.02 ;
      RECT 35.06 4.49 35.065 4.825 ;
      RECT 35.025 4.477 35.06 4.824 ;
      RECT 34.955 4.417 35.025 4.823 ;
      RECT 34.875 4.36 34.955 4.822 ;
      RECT 34.74 4.32 34.875 4.821 ;
      RECT 34.74 4.507 35.075 4.81 ;
      RECT 34.7 4.507 35.075 4.8 ;
      RECT 34.7 4.525 35.08 4.795 ;
      RECT 34.7 4.615 35.085 4.785 ;
      RECT 34.695 4.31 34.86 4.765 ;
      RECT 34.69 4.31 34.86 4.508 ;
      RECT 34.69 4.467 35.055 4.508 ;
      RECT 34.69 4.455 35.05 4.508 ;
      RECT 33.83 7.305 34 8.775 ;
      RECT 33.83 8.6 34.005 8.77 ;
      RECT 33.46 3.035 33.63 4.225 ;
      RECT 33.46 3.035 33.93 3.205 ;
      RECT 33.46 9.255 33.93 9.425 ;
      RECT 33.46 8.235 33.63 9.425 ;
      RECT 32.47 3.035 32.64 4.225 ;
      RECT 32.47 3.035 32.94 3.205 ;
      RECT 32.47 9.255 32.94 9.425 ;
      RECT 32.47 8.235 32.64 9.425 ;
      RECT 30.62 3.93 30.79 5.16 ;
      RECT 30.675 2.15 30.845 4.1 ;
      RECT 30.62 1.87 30.79 2.32 ;
      RECT 30.62 10.14 30.79 10.59 ;
      RECT 30.675 8.36 30.845 10.31 ;
      RECT 30.62 7.3 30.79 8.53 ;
      RECT 30.1 1.87 30.27 5.16 ;
      RECT 30.1 3.37 30.505 3.7 ;
      RECT 30.1 2.53 30.505 2.86 ;
      RECT 30.1 7.3 30.27 10.59 ;
      RECT 30.1 9.6 30.505 9.93 ;
      RECT 30.1 8.76 30.505 9.09 ;
      RECT 27.435 3.27 28.165 3.51 ;
      RECT 27.977 3.065 28.165 3.51 ;
      RECT 27.805 3.077 28.18 3.504 ;
      RECT 27.72 3.092 28.2 3.489 ;
      RECT 27.72 3.107 28.205 3.479 ;
      RECT 27.675 3.127 28.22 3.471 ;
      RECT 27.652 3.162 28.235 3.425 ;
      RECT 27.566 3.185 28.24 3.385 ;
      RECT 27.566 3.203 28.25 3.355 ;
      RECT 27.435 3.272 28.255 3.318 ;
      RECT 27.48 3.215 28.25 3.355 ;
      RECT 27.566 3.167 28.235 3.425 ;
      RECT 27.652 3.136 28.22 3.471 ;
      RECT 27.675 3.117 28.205 3.479 ;
      RECT 27.72 3.09 28.18 3.504 ;
      RECT 27.805 3.072 28.165 3.51 ;
      RECT 27.891 3.066 28.165 3.51 ;
      RECT 27.977 3.061 28.11 3.51 ;
      RECT 28.063 3.056 28.11 3.51 ;
      RECT 27.755 3.954 27.925 4.34 ;
      RECT 27.75 3.954 27.925 4.335 ;
      RECT 27.725 3.954 27.925 4.3 ;
      RECT 27.725 3.982 27.935 4.29 ;
      RECT 27.705 3.982 27.935 4.25 ;
      RECT 27.7 3.982 27.935 4.223 ;
      RECT 27.7 4 27.94 4.215 ;
      RECT 27.645 4 27.94 4.15 ;
      RECT 27.645 4.017 27.95 4.133 ;
      RECT 27.635 4.017 27.95 4.073 ;
      RECT 27.635 4.034 27.955 4.07 ;
      RECT 27.63 3.87 27.8 4.048 ;
      RECT 27.63 3.904 27.886 4.048 ;
      RECT 27.625 4.67 27.63 4.683 ;
      RECT 27.62 4.565 27.625 4.688 ;
      RECT 27.595 4.425 27.62 4.703 ;
      RECT 27.56 4.376 27.595 4.735 ;
      RECT 27.555 4.344 27.56 4.755 ;
      RECT 27.55 4.335 27.555 4.755 ;
      RECT 27.47 4.3 27.55 4.755 ;
      RECT 27.407 4.27 27.47 4.755 ;
      RECT 27.321 4.258 27.407 4.755 ;
      RECT 27.235 4.244 27.321 4.755 ;
      RECT 27.155 4.231 27.235 4.741 ;
      RECT 27.12 4.223 27.155 4.721 ;
      RECT 27.11 4.22 27.12 4.712 ;
      RECT 27.08 4.215 27.11 4.699 ;
      RECT 27.03 4.19 27.08 4.675 ;
      RECT 27.016 4.164 27.03 4.657 ;
      RECT 26.93 4.124 27.016 4.633 ;
      RECT 26.885 4.072 26.93 4.602 ;
      RECT 26.875 4.047 26.885 4.589 ;
      RECT 26.87 3.828 26.875 3.85 ;
      RECT 26.865 4.03 26.875 4.585 ;
      RECT 26.865 3.826 26.87 3.94 ;
      RECT 26.855 3.822 26.865 4.581 ;
      RECT 26.811 3.82 26.855 4.569 ;
      RECT 26.725 3.82 26.811 4.54 ;
      RECT 26.695 3.82 26.725 4.513 ;
      RECT 26.68 3.82 26.695 4.501 ;
      RECT 26.64 3.832 26.68 4.486 ;
      RECT 26.62 3.851 26.64 4.465 ;
      RECT 26.61 3.861 26.62 4.449 ;
      RECT 26.6 3.867 26.61 4.438 ;
      RECT 26.58 3.877 26.6 4.421 ;
      RECT 26.575 3.886 26.58 4.408 ;
      RECT 26.57 3.89 26.575 4.358 ;
      RECT 26.56 3.896 26.57 4.275 ;
      RECT 26.555 3.9 26.56 4.189 ;
      RECT 26.55 3.92 26.555 4.126 ;
      RECT 26.545 3.943 26.55 4.073 ;
      RECT 26.54 3.961 26.545 4.018 ;
      RECT 27.15 3.78 27.32 4.04 ;
      RECT 27.32 3.745 27.365 4.026 ;
      RECT 27.281 3.747 27.37 4.009 ;
      RECT 27.17 3.764 27.456 3.98 ;
      RECT 27.17 3.779 27.46 3.952 ;
      RECT 27.17 3.76 27.37 4.009 ;
      RECT 27.195 3.748 27.32 4.04 ;
      RECT 27.281 3.746 27.365 4.026 ;
      RECT 26.335 3.135 26.505 3.625 ;
      RECT 26.335 3.135 26.54 3.605 ;
      RECT 26.47 3.055 26.58 3.565 ;
      RECT 26.451 3.059 26.6 3.535 ;
      RECT 26.365 3.067 26.62 3.518 ;
      RECT 26.365 3.073 26.625 3.508 ;
      RECT 26.365 3.082 26.645 3.496 ;
      RECT 26.34 3.107 26.675 3.474 ;
      RECT 26.34 3.127 26.68 3.454 ;
      RECT 26.335 3.14 26.69 3.434 ;
      RECT 26.335 3.207 26.695 3.415 ;
      RECT 26.335 3.34 26.7 3.402 ;
      RECT 26.33 3.145 26.69 3.235 ;
      RECT 26.34 3.102 26.645 3.496 ;
      RECT 26.451 3.057 26.58 3.565 ;
      RECT 26.325 4.81 26.625 5.065 ;
      RECT 26.41 4.776 26.625 5.065 ;
      RECT 26.41 4.779 26.63 4.925 ;
      RECT 26.345 4.8 26.63 4.925 ;
      RECT 26.38 4.79 26.625 5.065 ;
      RECT 26.375 4.795 26.63 4.925 ;
      RECT 26.41 4.774 26.611 5.065 ;
      RECT 26.496 4.765 26.611 5.065 ;
      RECT 26.496 4.759 26.525 5.065 ;
      RECT 25.985 4.4 25.995 4.89 ;
      RECT 25.645 4.335 25.655 4.635 ;
      RECT 26.16 4.507 26.165 4.726 ;
      RECT 26.15 4.487 26.16 4.743 ;
      RECT 26.14 4.467 26.15 4.773 ;
      RECT 26.135 4.457 26.14 4.788 ;
      RECT 26.13 4.453 26.135 4.793 ;
      RECT 26.115 4.445 26.13 4.8 ;
      RECT 26.075 4.425 26.115 4.825 ;
      RECT 26.05 4.407 26.075 4.858 ;
      RECT 26.045 4.405 26.05 4.871 ;
      RECT 26.025 4.402 26.045 4.875 ;
      RECT 25.995 4.4 26.025 4.885 ;
      RECT 25.925 4.402 25.985 4.886 ;
      RECT 25.905 4.402 25.925 4.88 ;
      RECT 25.88 4.4 25.905 4.877 ;
      RECT 25.845 4.395 25.88 4.873 ;
      RECT 25.825 4.389 25.845 4.86 ;
      RECT 25.815 4.386 25.825 4.848 ;
      RECT 25.795 4.383 25.815 4.833 ;
      RECT 25.775 4.379 25.795 4.815 ;
      RECT 25.77 4.376 25.775 4.805 ;
      RECT 25.765 4.375 25.77 4.803 ;
      RECT 25.755 4.372 25.765 4.795 ;
      RECT 25.745 4.366 25.755 4.778 ;
      RECT 25.735 4.36 25.745 4.76 ;
      RECT 25.725 4.354 25.735 4.748 ;
      RECT 25.715 4.348 25.725 4.728 ;
      RECT 25.71 4.344 25.715 4.713 ;
      RECT 25.705 4.342 25.71 4.705 ;
      RECT 25.7 4.34 25.705 4.698 ;
      RECT 25.695 4.338 25.7 4.688 ;
      RECT 25.69 4.336 25.695 4.682 ;
      RECT 25.68 4.335 25.69 4.672 ;
      RECT 25.67 4.335 25.68 4.663 ;
      RECT 25.655 4.335 25.67 4.648 ;
      RECT 25.615 4.335 25.645 4.632 ;
      RECT 25.595 4.337 25.615 4.627 ;
      RECT 25.59 4.342 25.595 4.625 ;
      RECT 25.56 4.35 25.59 4.623 ;
      RECT 25.53 4.365 25.56 4.622 ;
      RECT 25.485 4.387 25.53 4.627 ;
      RECT 25.48 4.402 25.485 4.631 ;
      RECT 25.465 4.407 25.48 4.633 ;
      RECT 25.46 4.411 25.465 4.635 ;
      RECT 25.4 4.434 25.46 4.644 ;
      RECT 25.38 4.46 25.4 4.657 ;
      RECT 25.37 4.467 25.38 4.661 ;
      RECT 25.355 4.474 25.37 4.664 ;
      RECT 25.335 4.484 25.355 4.667 ;
      RECT 25.33 4.492 25.335 4.67 ;
      RECT 25.285 4.497 25.33 4.677 ;
      RECT 25.275 4.5 25.285 4.684 ;
      RECT 25.265 4.5 25.275 4.688 ;
      RECT 25.23 4.502 25.265 4.7 ;
      RECT 25.21 4.505 25.23 4.713 ;
      RECT 25.17 4.508 25.21 4.724 ;
      RECT 25.155 4.51 25.17 4.737 ;
      RECT 25.145 4.51 25.155 4.742 ;
      RECT 25.12 4.511 25.145 4.75 ;
      RECT 25.11 4.513 25.12 4.755 ;
      RECT 25.105 4.514 25.11 4.758 ;
      RECT 25.08 4.512 25.105 4.761 ;
      RECT 25.065 4.51 25.08 4.762 ;
      RECT 25.045 4.507 25.065 4.764 ;
      RECT 25.025 4.502 25.045 4.764 ;
      RECT 24.965 4.497 25.025 4.761 ;
      RECT 24.93 4.472 24.965 4.757 ;
      RECT 24.92 4.449 24.93 4.755 ;
      RECT 24.89 4.426 24.92 4.755 ;
      RECT 24.88 4.405 24.89 4.755 ;
      RECT 24.855 4.387 24.88 4.753 ;
      RECT 24.84 4.365 24.855 4.75 ;
      RECT 24.825 4.347 24.84 4.748 ;
      RECT 24.805 4.337 24.825 4.746 ;
      RECT 24.79 4.332 24.805 4.745 ;
      RECT 24.775 4.33 24.79 4.744 ;
      RECT 24.745 4.331 24.775 4.742 ;
      RECT 24.725 4.334 24.745 4.74 ;
      RECT 24.668 4.338 24.725 4.74 ;
      RECT 24.582 4.347 24.668 4.74 ;
      RECT 24.496 4.358 24.582 4.74 ;
      RECT 24.41 4.369 24.496 4.74 ;
      RECT 24.39 4.376 24.41 4.748 ;
      RECT 24.38 4.379 24.39 4.755 ;
      RECT 24.315 4.384 24.38 4.773 ;
      RECT 24.285 4.391 24.315 4.798 ;
      RECT 24.275 4.394 24.285 4.805 ;
      RECT 24.23 4.398 24.275 4.81 ;
      RECT 24.2 4.403 24.23 4.815 ;
      RECT 24.199 4.405 24.2 4.815 ;
      RECT 24.113 4.411 24.199 4.815 ;
      RECT 24.027 4.422 24.113 4.815 ;
      RECT 23.941 4.434 24.027 4.815 ;
      RECT 23.855 4.445 23.941 4.815 ;
      RECT 23.84 4.452 23.855 4.81 ;
      RECT 23.835 4.454 23.84 4.804 ;
      RECT 23.815 4.465 23.835 4.799 ;
      RECT 23.805 4.483 23.815 4.793 ;
      RECT 23.8 4.495 23.805 4.593 ;
      RECT 26.095 3.248 26.115 3.335 ;
      RECT 26.09 3.183 26.095 3.367 ;
      RECT 26.08 3.15 26.09 3.372 ;
      RECT 26.075 3.13 26.08 3.378 ;
      RECT 26.045 3.13 26.075 3.395 ;
      RECT 25.996 3.13 26.045 3.431 ;
      RECT 25.91 3.13 25.996 3.489 ;
      RECT 25.881 3.14 25.91 3.538 ;
      RECT 25.795 3.182 25.881 3.591 ;
      RECT 25.775 3.22 25.795 3.638 ;
      RECT 25.75 3.237 25.775 3.658 ;
      RECT 25.74 3.251 25.75 3.678 ;
      RECT 25.735 3.257 25.74 3.688 ;
      RECT 25.73 3.261 25.735 3.695 ;
      RECT 25.68 3.281 25.73 3.7 ;
      RECT 25.615 3.325 25.68 3.7 ;
      RECT 25.59 3.375 25.615 3.7 ;
      RECT 25.58 3.405 25.59 3.7 ;
      RECT 25.575 3.432 25.58 3.7 ;
      RECT 25.57 3.45 25.575 3.7 ;
      RECT 25.56 3.492 25.57 3.7 ;
      RECT 25.91 4.05 26.08 4.225 ;
      RECT 25.85 3.878 25.91 4.213 ;
      RECT 25.84 3.871 25.85 4.196 ;
      RECT 25.795 4.05 26.08 4.176 ;
      RECT 25.776 4.05 26.08 4.154 ;
      RECT 25.69 4.05 26.08 4.119 ;
      RECT 25.67 3.87 25.84 4.075 ;
      RECT 25.67 4.017 26.075 4.075 ;
      RECT 25.67 3.965 26.05 4.075 ;
      RECT 25.67 3.92 26.015 4.075 ;
      RECT 25.67 3.902 25.98 4.075 ;
      RECT 25.67 3.892 25.975 4.075 ;
      RECT 25.32 7.3 25.49 10.59 ;
      RECT 25.32 9.6 25.725 9.93 ;
      RECT 25.32 8.76 25.725 9.09 ;
      RECT 25.39 4.85 25.58 5.075 ;
      RECT 25.38 4.851 25.585 5.07 ;
      RECT 25.38 4.853 25.595 5.05 ;
      RECT 25.38 4.857 25.6 5.035 ;
      RECT 25.38 4.844 25.55 5.07 ;
      RECT 25.38 4.847 25.575 5.07 ;
      RECT 25.39 4.843 25.55 5.075 ;
      RECT 25.476 4.841 25.55 5.075 ;
      RECT 25.1 4.092 25.27 4.33 ;
      RECT 25.1 4.092 25.356 4.244 ;
      RECT 25.1 4.092 25.36 4.154 ;
      RECT 25.15 3.865 25.37 4.133 ;
      RECT 25.145 3.882 25.375 4.106 ;
      RECT 25.11 4.04 25.375 4.106 ;
      RECT 25.13 3.89 25.27 4.33 ;
      RECT 25.12 3.972 25.38 4.089 ;
      RECT 25.115 4.02 25.38 4.089 ;
      RECT 25.12 3.93 25.375 4.106 ;
      RECT 25.145 3.867 25.37 4.133 ;
      RECT 24.71 3.842 24.88 4.04 ;
      RECT 24.71 3.842 24.925 4.015 ;
      RECT 24.78 3.785 24.95 3.973 ;
      RECT 24.755 3.8 24.95 3.973 ;
      RECT 24.37 3.846 24.4 4.04 ;
      RECT 24.365 3.818 24.37 4.04 ;
      RECT 24.335 3.792 24.365 4.042 ;
      RECT 24.31 3.75 24.335 4.045 ;
      RECT 24.3 3.722 24.31 4.047 ;
      RECT 24.265 3.702 24.3 4.049 ;
      RECT 24.2 3.687 24.265 4.055 ;
      RECT 24.15 3.685 24.2 4.061 ;
      RECT 24.127 3.687 24.15 4.066 ;
      RECT 24.041 3.698 24.127 4.072 ;
      RECT 23.955 3.716 24.041 4.082 ;
      RECT 23.94 3.727 23.955 4.088 ;
      RECT 23.87 3.75 23.94 4.094 ;
      RECT 23.815 3.782 23.87 4.102 ;
      RECT 23.775 3.805 23.815 4.108 ;
      RECT 23.761 3.818 23.775 4.111 ;
      RECT 23.675 3.84 23.761 4.117 ;
      RECT 23.66 3.865 23.675 4.123 ;
      RECT 23.62 3.88 23.66 4.127 ;
      RECT 23.57 3.895 23.62 4.132 ;
      RECT 23.545 3.902 23.57 4.136 ;
      RECT 23.485 3.897 23.545 4.14 ;
      RECT 23.47 3.888 23.485 4.144 ;
      RECT 23.4 3.878 23.47 4.14 ;
      RECT 23.375 3.87 23.395 4.13 ;
      RECT 23.316 3.87 23.375 4.108 ;
      RECT 23.23 3.87 23.316 4.065 ;
      RECT 23.395 3.87 23.4 4.135 ;
      RECT 24.09 3.101 24.26 3.435 ;
      RECT 24.06 3.101 24.26 3.43 ;
      RECT 24 3.068 24.06 3.418 ;
      RECT 24 3.124 24.27 3.413 ;
      RECT 23.975 3.124 24.27 3.407 ;
      RECT 23.97 3.065 24 3.404 ;
      RECT 23.955 3.071 24.09 3.402 ;
      RECT 23.95 3.079 24.175 3.39 ;
      RECT 23.95 3.131 24.285 3.343 ;
      RECT 23.935 3.087 24.175 3.338 ;
      RECT 23.935 3.157 24.295 3.279 ;
      RECT 23.905 3.107 24.26 3.24 ;
      RECT 23.905 3.197 24.305 3.236 ;
      RECT 23.955 3.076 24.175 3.402 ;
      RECT 23.295 3.406 23.35 3.67 ;
      RECT 23.295 3.406 23.415 3.669 ;
      RECT 23.295 3.406 23.44 3.668 ;
      RECT 23.295 3.406 23.505 3.667 ;
      RECT 23.44 3.372 23.52 3.666 ;
      RECT 23.255 3.416 23.665 3.665 ;
      RECT 23.295 3.413 23.665 3.665 ;
      RECT 23.255 3.421 23.67 3.658 ;
      RECT 23.24 3.423 23.67 3.657 ;
      RECT 23.24 3.43 23.675 3.653 ;
      RECT 23.22 3.429 23.67 3.649 ;
      RECT 23.22 3.437 23.68 3.648 ;
      RECT 23.215 3.434 23.675 3.644 ;
      RECT 23.215 3.447 23.69 3.643 ;
      RECT 23.2 3.437 23.68 3.642 ;
      RECT 23.165 3.45 23.69 3.635 ;
      RECT 23.35 3.405 23.66 3.665 ;
      RECT 23.35 3.39 23.61 3.665 ;
      RECT 23.415 3.377 23.545 3.665 ;
      RECT 22.96 4.466 22.975 4.859 ;
      RECT 22.925 4.471 22.975 4.858 ;
      RECT 22.96 4.47 23.02 4.857 ;
      RECT 22.905 4.481 23.02 4.856 ;
      RECT 22.92 4.477 23.02 4.856 ;
      RECT 22.885 4.487 23.095 4.853 ;
      RECT 22.885 4.506 23.14 4.851 ;
      RECT 22.885 4.513 23.145 4.848 ;
      RECT 22.87 4.49 23.095 4.845 ;
      RECT 22.85 4.495 23.095 4.838 ;
      RECT 22.845 4.499 23.095 4.834 ;
      RECT 22.845 4.516 23.155 4.833 ;
      RECT 22.825 4.51 23.14 4.829 ;
      RECT 22.825 4.519 23.16 4.823 ;
      RECT 22.82 4.525 23.16 4.595 ;
      RECT 22.885 4.485 23.02 4.853 ;
      RECT 22.76 3.848 22.96 4.16 ;
      RECT 22.835 3.826 22.96 4.16 ;
      RECT 22.775 3.845 22.965 4.145 ;
      RECT 22.745 3.856 22.965 4.143 ;
      RECT 22.76 3.851 22.97 4.109 ;
      RECT 22.745 3.955 22.975 4.076 ;
      RECT 22.775 3.827 22.96 4.16 ;
      RECT 22.835 3.805 22.935 4.16 ;
      RECT 22.86 3.802 22.935 4.16 ;
      RECT 22.86 3.797 22.88 4.16 ;
      RECT 22.265 3.865 22.44 4.04 ;
      RECT 22.26 3.865 22.44 4.038 ;
      RECT 22.235 3.865 22.44 4.033 ;
      RECT 22.18 3.845 22.35 4.023 ;
      RECT 22.18 3.852 22.415 4.023 ;
      RECT 22.265 4.532 22.28 4.715 ;
      RECT 22.255 4.51 22.265 4.715 ;
      RECT 22.24 4.49 22.255 4.715 ;
      RECT 22.23 4.465 22.24 4.715 ;
      RECT 22.2 4.43 22.23 4.715 ;
      RECT 22.165 4.37 22.2 4.715 ;
      RECT 22.16 4.332 22.165 4.715 ;
      RECT 22.11 4.283 22.16 4.715 ;
      RECT 22.1 4.233 22.11 4.703 ;
      RECT 22.085 4.212 22.1 4.663 ;
      RECT 22.065 4.18 22.085 4.613 ;
      RECT 22.04 4.136 22.065 4.553 ;
      RECT 22.035 4.108 22.04 4.508 ;
      RECT 22.03 4.099 22.035 4.494 ;
      RECT 22.025 4.092 22.03 4.481 ;
      RECT 22.02 4.087 22.025 4.47 ;
      RECT 22.015 4.072 22.02 4.46 ;
      RECT 22.01 4.05 22.015 4.447 ;
      RECT 22 4.01 22.01 4.422 ;
      RECT 21.975 3.94 22 4.378 ;
      RECT 21.97 3.88 21.975 4.343 ;
      RECT 21.955 3.86 21.97 4.31 ;
      RECT 21.95 3.86 21.955 4.285 ;
      RECT 21.92 3.86 21.95 4.24 ;
      RECT 21.875 3.86 21.92 4.18 ;
      RECT 21.8 3.86 21.875 4.128 ;
      RECT 21.795 3.86 21.8 4.093 ;
      RECT 21.79 3.86 21.795 4.083 ;
      RECT 21.785 3.86 21.79 4.063 ;
      RECT 22.05 3.08 22.22 3.55 ;
      RECT 21.995 3.073 22.19 3.534 ;
      RECT 21.995 3.087 22.225 3.533 ;
      RECT 21.98 3.088 22.225 3.514 ;
      RECT 21.975 3.106 22.225 3.5 ;
      RECT 21.98 3.089 22.23 3.498 ;
      RECT 21.965 3.12 22.23 3.483 ;
      RECT 21.98 3.095 22.235 3.468 ;
      RECT 21.96 3.135 22.235 3.465 ;
      RECT 21.975 3.107 22.24 3.45 ;
      RECT 21.975 3.119 22.245 3.43 ;
      RECT 21.96 3.135 22.25 3.413 ;
      RECT 21.96 3.145 22.255 3.268 ;
      RECT 21.955 3.145 22.255 3.225 ;
      RECT 21.955 3.16 22.26 3.203 ;
      RECT 22.05 3.07 22.19 3.55 ;
      RECT 22.05 3.068 22.16 3.55 ;
      RECT 22.136 3.065 22.16 3.55 ;
      RECT 21.795 4.732 21.8 4.778 ;
      RECT 21.785 4.58 21.795 4.802 ;
      RECT 21.78 4.425 21.785 4.827 ;
      RECT 21.765 4.387 21.78 4.838 ;
      RECT 21.76 4.37 21.765 4.845 ;
      RECT 21.75 4.358 21.76 4.852 ;
      RECT 21.745 4.349 21.75 4.854 ;
      RECT 21.74 4.347 21.745 4.858 ;
      RECT 21.695 4.338 21.74 4.873 ;
      RECT 21.69 4.33 21.695 4.887 ;
      RECT 21.685 4.327 21.69 4.891 ;
      RECT 21.67 4.322 21.685 4.899 ;
      RECT 21.615 4.312 21.67 4.91 ;
      RECT 21.58 4.3 21.615 4.911 ;
      RECT 21.571 4.295 21.58 4.905 ;
      RECT 21.485 4.295 21.571 4.895 ;
      RECT 21.455 4.295 21.485 4.873 ;
      RECT 21.445 4.295 21.45 4.853 ;
      RECT 21.44 4.295 21.445 4.815 ;
      RECT 21.435 4.295 21.44 4.773 ;
      RECT 21.43 4.295 21.435 4.733 ;
      RECT 21.425 4.295 21.43 4.663 ;
      RECT 21.415 4.295 21.425 4.585 ;
      RECT 21.41 4.295 21.415 4.485 ;
      RECT 21.45 4.295 21.455 4.855 ;
      RECT 20.945 4.377 21.035 4.855 ;
      RECT 20.93 4.38 21.05 4.853 ;
      RECT 20.945 4.379 21.05 4.853 ;
      RECT 20.91 4.386 21.075 4.843 ;
      RECT 20.93 4.38 21.075 4.843 ;
      RECT 20.895 4.392 21.075 4.831 ;
      RECT 20.93 4.383 21.125 4.824 ;
      RECT 20.881 4.4 21.125 4.822 ;
      RECT 20.91 4.39 21.135 4.81 ;
      RECT 20.881 4.411 21.165 4.801 ;
      RECT 20.795 4.435 21.165 4.795 ;
      RECT 20.795 4.448 21.205 4.778 ;
      RECT 20.79 4.47 21.205 4.771 ;
      RECT 20.76 4.485 21.205 4.761 ;
      RECT 20.755 4.496 21.205 4.751 ;
      RECT 20.725 4.509 21.205 4.742 ;
      RECT 20.71 4.527 21.205 4.731 ;
      RECT 20.685 4.54 21.205 4.721 ;
      RECT 20.945 4.376 20.955 4.855 ;
      RECT 20.991 3.8 21.03 4.045 ;
      RECT 20.905 3.8 21.04 4.043 ;
      RECT 20.79 3.825 21.04 4.04 ;
      RECT 20.79 3.825 21.045 4.038 ;
      RECT 20.79 3.825 21.06 4.033 ;
      RECT 20.896 3.8 21.075 4.013 ;
      RECT 20.81 3.808 21.075 4.013 ;
      RECT 20.48 3.16 20.65 3.595 ;
      RECT 20.47 3.194 20.65 3.578 ;
      RECT 20.55 3.13 20.72 3.565 ;
      RECT 20.455 3.205 20.72 3.543 ;
      RECT 20.55 3.14 20.725 3.533 ;
      RECT 20.48 3.192 20.755 3.518 ;
      RECT 20.44 3.218 20.755 3.503 ;
      RECT 20.44 3.26 20.765 3.483 ;
      RECT 20.435 3.285 20.77 3.465 ;
      RECT 20.435 3.295 20.775 3.45 ;
      RECT 20.43 3.232 20.755 3.448 ;
      RECT 20.43 3.305 20.78 3.433 ;
      RECT 20.425 3.242 20.755 3.43 ;
      RECT 20.42 3.326 20.785 3.413 ;
      RECT 20.42 3.358 20.79 3.393 ;
      RECT 20.415 3.272 20.765 3.385 ;
      RECT 20.42 3.257 20.755 3.413 ;
      RECT 20.435 3.227 20.755 3.465 ;
      RECT 20.28 3.814 20.505 4.07 ;
      RECT 20.28 3.847 20.525 4.06 ;
      RECT 20.245 3.847 20.525 4.058 ;
      RECT 20.245 3.86 20.53 4.048 ;
      RECT 20.245 3.88 20.54 4.04 ;
      RECT 20.245 3.977 20.545 4.033 ;
      RECT 20.225 3.725 20.355 4.023 ;
      RECT 20.18 3.88 20.54 3.965 ;
      RECT 20.17 3.725 20.355 3.91 ;
      RECT 20.17 3.757 20.441 3.91 ;
      RECT 20.135 4.287 20.155 4.465 ;
      RECT 20.1 4.24 20.135 4.465 ;
      RECT 20.085 4.18 20.1 4.465 ;
      RECT 20.06 4.127 20.085 4.465 ;
      RECT 20.045 4.08 20.06 4.465 ;
      RECT 20.025 4.057 20.045 4.465 ;
      RECT 20 4.022 20.025 4.465 ;
      RECT 19.99 3.868 20 4.465 ;
      RECT 19.96 3.863 19.99 4.456 ;
      RECT 19.955 3.86 19.96 4.446 ;
      RECT 19.94 3.86 19.955 4.42 ;
      RECT 19.935 3.86 19.94 4.383 ;
      RECT 19.91 3.86 19.935 4.335 ;
      RECT 19.89 3.86 19.91 4.26 ;
      RECT 19.88 3.86 19.89 4.22 ;
      RECT 19.875 3.86 19.88 4.195 ;
      RECT 19.87 3.86 19.875 4.178 ;
      RECT 19.865 3.86 19.87 4.16 ;
      RECT 19.86 3.861 19.865 4.15 ;
      RECT 19.85 3.863 19.86 4.118 ;
      RECT 19.84 3.865 19.85 4.085 ;
      RECT 19.83 3.868 19.84 4.058 ;
      RECT 20.155 4.295 20.38 4.465 ;
      RECT 19.485 3.107 19.655 3.56 ;
      RECT 19.485 3.107 19.745 3.526 ;
      RECT 19.485 3.107 19.775 3.51 ;
      RECT 19.485 3.107 19.805 3.483 ;
      RECT 19.741 3.085 19.82 3.465 ;
      RECT 19.52 3.092 19.825 3.45 ;
      RECT 19.52 3.1 19.835 3.413 ;
      RECT 19.48 3.127 19.835 3.385 ;
      RECT 19.465 3.14 19.835 3.35 ;
      RECT 19.485 3.115 19.855 3.34 ;
      RECT 19.46 3.18 19.855 3.31 ;
      RECT 19.46 3.21 19.86 3.293 ;
      RECT 19.455 3.24 19.86 3.28 ;
      RECT 19.52 3.089 19.82 3.465 ;
      RECT 19.655 3.086 19.741 3.544 ;
      RECT 19.606 3.087 19.82 3.465 ;
      RECT 19.75 4.747 19.795 4.94 ;
      RECT 19.74 4.717 19.75 4.94 ;
      RECT 19.735 4.702 19.74 4.94 ;
      RECT 19.695 4.612 19.735 4.94 ;
      RECT 19.69 4.525 19.695 4.94 ;
      RECT 19.68 4.495 19.69 4.94 ;
      RECT 19.675 4.455 19.68 4.94 ;
      RECT 19.665 4.417 19.675 4.94 ;
      RECT 19.66 4.382 19.665 4.94 ;
      RECT 19.64 4.335 19.66 4.94 ;
      RECT 19.625 4.26 19.64 4.94 ;
      RECT 19.62 4.215 19.625 4.935 ;
      RECT 19.615 4.195 19.62 4.908 ;
      RECT 19.61 4.175 19.615 4.893 ;
      RECT 19.605 4.15 19.61 4.873 ;
      RECT 19.6 4.128 19.605 4.858 ;
      RECT 19.595 4.106 19.6 4.84 ;
      RECT 19.59 4.085 19.595 4.83 ;
      RECT 19.58 4.057 19.59 4.8 ;
      RECT 19.57 4.02 19.58 4.768 ;
      RECT 19.56 3.98 19.57 4.735 ;
      RECT 19.55 3.958 19.56 4.705 ;
      RECT 19.52 3.91 19.55 4.637 ;
      RECT 19.505 3.87 19.52 4.564 ;
      RECT 19.495 3.87 19.505 4.53 ;
      RECT 19.49 3.87 19.495 4.505 ;
      RECT 19.485 3.87 19.49 4.49 ;
      RECT 19.48 3.87 19.485 4.468 ;
      RECT 19.475 3.87 19.48 4.455 ;
      RECT 19.46 3.87 19.475 4.42 ;
      RECT 19.44 3.87 19.46 4.36 ;
      RECT 19.43 3.87 19.44 4.31 ;
      RECT 19.41 3.87 19.43 4.258 ;
      RECT 19.39 3.87 19.41 4.215 ;
      RECT 19.38 3.87 19.39 4.203 ;
      RECT 19.35 3.87 19.38 4.19 ;
      RECT 19.32 3.891 19.35 4.17 ;
      RECT 19.31 3.919 19.32 4.15 ;
      RECT 19.295 3.936 19.31 4.118 ;
      RECT 19.29 3.95 19.295 4.085 ;
      RECT 19.285 3.958 19.29 4.058 ;
      RECT 19.28 3.966 19.285 4.02 ;
      RECT 19.285 4.49 19.29 4.825 ;
      RECT 19.25 4.477 19.285 4.824 ;
      RECT 19.18 4.417 19.25 4.823 ;
      RECT 19.1 4.36 19.18 4.822 ;
      RECT 18.965 4.32 19.1 4.821 ;
      RECT 18.965 4.507 19.3 4.81 ;
      RECT 18.925 4.507 19.3 4.8 ;
      RECT 18.925 4.525 19.305 4.795 ;
      RECT 18.925 4.615 19.31 4.785 ;
      RECT 18.92 4.31 19.085 4.765 ;
      RECT 18.915 4.31 19.085 4.508 ;
      RECT 18.915 4.467 19.28 4.508 ;
      RECT 18.915 4.455 19.275 4.508 ;
      RECT 18.05 7.305 18.22 8.775 ;
      RECT 18.05 8.6 18.225 8.77 ;
      RECT 17.68 3.035 17.85 4.225 ;
      RECT 17.68 3.035 18.15 3.205 ;
      RECT 17.68 9.255 18.15 9.425 ;
      RECT 17.68 8.235 17.85 9.425 ;
      RECT 16.69 3.035 16.86 4.225 ;
      RECT 16.69 3.035 17.16 3.205 ;
      RECT 16.69 9.255 17.16 9.425 ;
      RECT 16.69 8.235 16.86 9.425 ;
      RECT 14.84 3.93 15.01 5.16 ;
      RECT 14.895 2.15 15.065 4.1 ;
      RECT 14.84 1.87 15.01 2.32 ;
      RECT 14.84 10.14 15.01 10.59 ;
      RECT 14.895 8.36 15.065 10.31 ;
      RECT 14.84 7.3 15.01 8.53 ;
      RECT 14.32 1.87 14.49 5.16 ;
      RECT 14.32 3.37 14.725 3.7 ;
      RECT 14.32 2.53 14.725 2.86 ;
      RECT 14.32 7.3 14.49 10.59 ;
      RECT 14.32 9.6 14.725 9.93 ;
      RECT 14.32 8.76 14.725 9.09 ;
      RECT 11.655 3.27 12.385 3.51 ;
      RECT 12.197 3.065 12.385 3.51 ;
      RECT 12.025 3.077 12.4 3.504 ;
      RECT 11.94 3.092 12.42 3.489 ;
      RECT 11.94 3.107 12.425 3.479 ;
      RECT 11.895 3.127 12.44 3.471 ;
      RECT 11.872 3.162 12.455 3.425 ;
      RECT 11.786 3.185 12.46 3.385 ;
      RECT 11.786 3.203 12.47 3.355 ;
      RECT 11.655 3.272 12.475 3.318 ;
      RECT 11.7 3.215 12.47 3.355 ;
      RECT 11.786 3.167 12.455 3.425 ;
      RECT 11.872 3.136 12.44 3.471 ;
      RECT 11.895 3.117 12.425 3.479 ;
      RECT 11.94 3.09 12.4 3.504 ;
      RECT 12.025 3.072 12.385 3.51 ;
      RECT 12.111 3.066 12.385 3.51 ;
      RECT 12.197 3.061 12.33 3.51 ;
      RECT 12.283 3.056 12.33 3.51 ;
      RECT 11.975 3.954 12.145 4.34 ;
      RECT 11.97 3.954 12.145 4.335 ;
      RECT 11.945 3.954 12.145 4.3 ;
      RECT 11.945 3.982 12.155 4.29 ;
      RECT 11.925 3.982 12.155 4.25 ;
      RECT 11.92 3.982 12.155 4.223 ;
      RECT 11.92 4 12.16 4.215 ;
      RECT 11.865 4 12.16 4.15 ;
      RECT 11.865 4.017 12.17 4.133 ;
      RECT 11.855 4.017 12.17 4.073 ;
      RECT 11.855 4.034 12.175 4.07 ;
      RECT 11.85 3.87 12.02 4.048 ;
      RECT 11.85 3.904 12.106 4.048 ;
      RECT 11.845 4.67 11.85 4.683 ;
      RECT 11.84 4.565 11.845 4.688 ;
      RECT 11.815 4.425 11.84 4.703 ;
      RECT 11.78 4.376 11.815 4.735 ;
      RECT 11.775 4.344 11.78 4.755 ;
      RECT 11.77 4.335 11.775 4.755 ;
      RECT 11.69 4.3 11.77 4.755 ;
      RECT 11.627 4.27 11.69 4.755 ;
      RECT 11.541 4.258 11.627 4.755 ;
      RECT 11.455 4.244 11.541 4.755 ;
      RECT 11.375 4.231 11.455 4.741 ;
      RECT 11.34 4.223 11.375 4.721 ;
      RECT 11.33 4.22 11.34 4.712 ;
      RECT 11.3 4.215 11.33 4.699 ;
      RECT 11.25 4.19 11.3 4.675 ;
      RECT 11.236 4.164 11.25 4.657 ;
      RECT 11.15 4.124 11.236 4.633 ;
      RECT 11.105 4.072 11.15 4.602 ;
      RECT 11.095 4.047 11.105 4.589 ;
      RECT 11.09 3.828 11.095 3.85 ;
      RECT 11.085 4.03 11.095 4.585 ;
      RECT 11.085 3.826 11.09 3.94 ;
      RECT 11.075 3.822 11.085 4.581 ;
      RECT 11.031 3.82 11.075 4.569 ;
      RECT 10.945 3.82 11.031 4.54 ;
      RECT 10.915 3.82 10.945 4.513 ;
      RECT 10.9 3.82 10.915 4.501 ;
      RECT 10.86 3.832 10.9 4.486 ;
      RECT 10.84 3.851 10.86 4.465 ;
      RECT 10.83 3.861 10.84 4.449 ;
      RECT 10.82 3.867 10.83 4.438 ;
      RECT 10.8 3.877 10.82 4.421 ;
      RECT 10.795 3.886 10.8 4.408 ;
      RECT 10.79 3.89 10.795 4.358 ;
      RECT 10.78 3.896 10.79 4.275 ;
      RECT 10.775 3.9 10.78 4.189 ;
      RECT 10.77 3.92 10.775 4.126 ;
      RECT 10.765 3.943 10.77 4.073 ;
      RECT 10.76 3.961 10.765 4.018 ;
      RECT 11.37 3.78 11.54 4.04 ;
      RECT 11.54 3.745 11.585 4.026 ;
      RECT 11.501 3.747 11.59 4.009 ;
      RECT 11.39 3.764 11.676 3.98 ;
      RECT 11.39 3.779 11.68 3.952 ;
      RECT 11.39 3.76 11.59 4.009 ;
      RECT 11.415 3.748 11.54 4.04 ;
      RECT 11.501 3.746 11.585 4.026 ;
      RECT 10.555 3.135 10.725 3.625 ;
      RECT 10.555 3.135 10.76 3.605 ;
      RECT 10.69 3.055 10.8 3.565 ;
      RECT 10.671 3.059 10.82 3.535 ;
      RECT 10.585 3.067 10.84 3.518 ;
      RECT 10.585 3.073 10.845 3.508 ;
      RECT 10.585 3.082 10.865 3.496 ;
      RECT 10.56 3.107 10.895 3.474 ;
      RECT 10.56 3.127 10.9 3.454 ;
      RECT 10.555 3.14 10.91 3.434 ;
      RECT 10.555 3.207 10.915 3.415 ;
      RECT 10.555 3.34 10.92 3.402 ;
      RECT 10.55 3.145 10.91 3.235 ;
      RECT 10.56 3.102 10.865 3.496 ;
      RECT 10.671 3.057 10.8 3.565 ;
      RECT 10.545 4.81 10.845 5.065 ;
      RECT 10.63 4.776 10.845 5.065 ;
      RECT 10.63 4.779 10.85 4.925 ;
      RECT 10.565 4.8 10.85 4.925 ;
      RECT 10.6 4.79 10.845 5.065 ;
      RECT 10.595 4.795 10.85 4.925 ;
      RECT 10.63 4.774 10.831 5.065 ;
      RECT 10.716 4.765 10.831 5.065 ;
      RECT 10.716 4.759 10.745 5.065 ;
      RECT 10.205 4.4 10.215 4.89 ;
      RECT 9.865 4.335 9.875 4.635 ;
      RECT 10.38 4.507 10.385 4.726 ;
      RECT 10.37 4.487 10.38 4.743 ;
      RECT 10.36 4.467 10.37 4.773 ;
      RECT 10.355 4.457 10.36 4.788 ;
      RECT 10.35 4.453 10.355 4.793 ;
      RECT 10.335 4.445 10.35 4.8 ;
      RECT 10.295 4.425 10.335 4.825 ;
      RECT 10.27 4.407 10.295 4.858 ;
      RECT 10.265 4.405 10.27 4.871 ;
      RECT 10.245 4.402 10.265 4.875 ;
      RECT 10.215 4.4 10.245 4.885 ;
      RECT 10.145 4.402 10.205 4.886 ;
      RECT 10.125 4.402 10.145 4.88 ;
      RECT 10.1 4.4 10.125 4.877 ;
      RECT 10.065 4.395 10.1 4.873 ;
      RECT 10.045 4.389 10.065 4.86 ;
      RECT 10.035 4.386 10.045 4.848 ;
      RECT 10.015 4.383 10.035 4.833 ;
      RECT 9.995 4.379 10.015 4.815 ;
      RECT 9.99 4.376 9.995 4.805 ;
      RECT 9.985 4.375 9.99 4.803 ;
      RECT 9.975 4.372 9.985 4.795 ;
      RECT 9.965 4.366 9.975 4.778 ;
      RECT 9.955 4.36 9.965 4.76 ;
      RECT 9.945 4.354 9.955 4.748 ;
      RECT 9.935 4.348 9.945 4.728 ;
      RECT 9.93 4.344 9.935 4.713 ;
      RECT 9.925 4.342 9.93 4.705 ;
      RECT 9.92 4.34 9.925 4.698 ;
      RECT 9.915 4.338 9.92 4.688 ;
      RECT 9.91 4.336 9.915 4.682 ;
      RECT 9.9 4.335 9.91 4.672 ;
      RECT 9.89 4.335 9.9 4.663 ;
      RECT 9.875 4.335 9.89 4.648 ;
      RECT 9.835 4.335 9.865 4.632 ;
      RECT 9.815 4.337 9.835 4.627 ;
      RECT 9.81 4.342 9.815 4.625 ;
      RECT 9.78 4.35 9.81 4.623 ;
      RECT 9.75 4.365 9.78 4.622 ;
      RECT 9.705 4.387 9.75 4.627 ;
      RECT 9.7 4.402 9.705 4.631 ;
      RECT 9.685 4.407 9.7 4.633 ;
      RECT 9.68 4.411 9.685 4.635 ;
      RECT 9.62 4.434 9.68 4.644 ;
      RECT 9.6 4.46 9.62 4.657 ;
      RECT 9.59 4.467 9.6 4.661 ;
      RECT 9.575 4.474 9.59 4.664 ;
      RECT 9.555 4.484 9.575 4.667 ;
      RECT 9.55 4.492 9.555 4.67 ;
      RECT 9.505 4.497 9.55 4.677 ;
      RECT 9.495 4.5 9.505 4.684 ;
      RECT 9.485 4.5 9.495 4.688 ;
      RECT 9.45 4.502 9.485 4.7 ;
      RECT 9.43 4.505 9.45 4.713 ;
      RECT 9.39 4.508 9.43 4.724 ;
      RECT 9.375 4.51 9.39 4.737 ;
      RECT 9.365 4.51 9.375 4.742 ;
      RECT 9.34 4.511 9.365 4.75 ;
      RECT 9.33 4.513 9.34 4.755 ;
      RECT 9.325 4.514 9.33 4.758 ;
      RECT 9.3 4.512 9.325 4.761 ;
      RECT 9.285 4.51 9.3 4.762 ;
      RECT 9.265 4.507 9.285 4.764 ;
      RECT 9.245 4.502 9.265 4.764 ;
      RECT 9.185 4.497 9.245 4.761 ;
      RECT 9.15 4.472 9.185 4.757 ;
      RECT 9.14 4.449 9.15 4.755 ;
      RECT 9.11 4.426 9.14 4.755 ;
      RECT 9.1 4.405 9.11 4.755 ;
      RECT 9.075 4.387 9.1 4.753 ;
      RECT 9.06 4.365 9.075 4.75 ;
      RECT 9.045 4.347 9.06 4.748 ;
      RECT 9.025 4.337 9.045 4.746 ;
      RECT 9.01 4.332 9.025 4.745 ;
      RECT 8.995 4.33 9.01 4.744 ;
      RECT 8.965 4.331 8.995 4.742 ;
      RECT 8.945 4.334 8.965 4.74 ;
      RECT 8.888 4.338 8.945 4.74 ;
      RECT 8.802 4.347 8.888 4.74 ;
      RECT 8.716 4.358 8.802 4.74 ;
      RECT 8.63 4.369 8.716 4.74 ;
      RECT 8.61 4.376 8.63 4.748 ;
      RECT 8.6 4.379 8.61 4.755 ;
      RECT 8.535 4.384 8.6 4.773 ;
      RECT 8.505 4.391 8.535 4.798 ;
      RECT 8.495 4.394 8.505 4.805 ;
      RECT 8.45 4.398 8.495 4.81 ;
      RECT 8.42 4.403 8.45 4.815 ;
      RECT 8.419 4.405 8.42 4.815 ;
      RECT 8.333 4.411 8.419 4.815 ;
      RECT 8.247 4.422 8.333 4.815 ;
      RECT 8.161 4.434 8.247 4.815 ;
      RECT 8.075 4.445 8.161 4.815 ;
      RECT 8.06 4.452 8.075 4.81 ;
      RECT 8.055 4.454 8.06 4.804 ;
      RECT 8.035 4.465 8.055 4.799 ;
      RECT 8.025 4.483 8.035 4.793 ;
      RECT 8.02 4.495 8.025 4.593 ;
      RECT 10.315 3.248 10.335 3.335 ;
      RECT 10.31 3.183 10.315 3.367 ;
      RECT 10.3 3.15 10.31 3.372 ;
      RECT 10.295 3.13 10.3 3.378 ;
      RECT 10.265 3.13 10.295 3.395 ;
      RECT 10.216 3.13 10.265 3.431 ;
      RECT 10.13 3.13 10.216 3.489 ;
      RECT 10.101 3.14 10.13 3.538 ;
      RECT 10.015 3.182 10.101 3.591 ;
      RECT 9.995 3.22 10.015 3.638 ;
      RECT 9.97 3.237 9.995 3.658 ;
      RECT 9.96 3.251 9.97 3.678 ;
      RECT 9.955 3.257 9.96 3.688 ;
      RECT 9.95 3.261 9.955 3.695 ;
      RECT 9.9 3.281 9.95 3.7 ;
      RECT 9.835 3.325 9.9 3.7 ;
      RECT 9.81 3.375 9.835 3.7 ;
      RECT 9.8 3.405 9.81 3.7 ;
      RECT 9.795 3.432 9.8 3.7 ;
      RECT 9.79 3.45 9.795 3.7 ;
      RECT 9.78 3.492 9.79 3.7 ;
      RECT 10.13 4.05 10.3 4.225 ;
      RECT 10.07 3.878 10.13 4.213 ;
      RECT 10.06 3.871 10.07 4.196 ;
      RECT 10.015 4.05 10.3 4.176 ;
      RECT 9.996 4.05 10.3 4.154 ;
      RECT 9.91 4.05 10.3 4.119 ;
      RECT 9.89 3.87 10.06 4.075 ;
      RECT 9.89 4.017 10.295 4.075 ;
      RECT 9.89 3.965 10.27 4.075 ;
      RECT 9.89 3.92 10.235 4.075 ;
      RECT 9.89 3.902 10.2 4.075 ;
      RECT 9.89 3.892 10.195 4.075 ;
      RECT 9.54 7.3 9.71 10.59 ;
      RECT 9.54 9.6 9.945 9.93 ;
      RECT 9.54 8.76 9.945 9.09 ;
      RECT 9.61 4.85 9.8 5.075 ;
      RECT 9.6 4.851 9.805 5.07 ;
      RECT 9.6 4.853 9.815 5.05 ;
      RECT 9.6 4.857 9.82 5.035 ;
      RECT 9.6 4.844 9.77 5.07 ;
      RECT 9.6 4.847 9.795 5.07 ;
      RECT 9.61 4.843 9.77 5.075 ;
      RECT 9.696 4.841 9.77 5.075 ;
      RECT 9.32 4.092 9.49 4.33 ;
      RECT 9.32 4.092 9.576 4.244 ;
      RECT 9.32 4.092 9.58 4.154 ;
      RECT 9.37 3.865 9.59 4.133 ;
      RECT 9.365 3.882 9.595 4.106 ;
      RECT 9.33 4.04 9.595 4.106 ;
      RECT 9.35 3.89 9.49 4.33 ;
      RECT 9.34 3.972 9.6 4.089 ;
      RECT 9.335 4.02 9.6 4.089 ;
      RECT 9.34 3.93 9.595 4.106 ;
      RECT 9.365 3.867 9.59 4.133 ;
      RECT 8.93 3.842 9.1 4.04 ;
      RECT 8.93 3.842 9.145 4.015 ;
      RECT 9 3.785 9.17 3.973 ;
      RECT 8.975 3.8 9.17 3.973 ;
      RECT 8.59 3.846 8.62 4.04 ;
      RECT 8.585 3.818 8.59 4.04 ;
      RECT 8.555 3.792 8.585 4.042 ;
      RECT 8.53 3.75 8.555 4.045 ;
      RECT 8.52 3.722 8.53 4.047 ;
      RECT 8.485 3.702 8.52 4.049 ;
      RECT 8.42 3.687 8.485 4.055 ;
      RECT 8.37 3.685 8.42 4.061 ;
      RECT 8.347 3.687 8.37 4.066 ;
      RECT 8.261 3.698 8.347 4.072 ;
      RECT 8.175 3.716 8.261 4.082 ;
      RECT 8.16 3.727 8.175 4.088 ;
      RECT 8.09 3.75 8.16 4.094 ;
      RECT 8.035 3.782 8.09 4.102 ;
      RECT 7.995 3.805 8.035 4.108 ;
      RECT 7.981 3.818 7.995 4.111 ;
      RECT 7.895 3.84 7.981 4.117 ;
      RECT 7.88 3.865 7.895 4.123 ;
      RECT 7.84 3.88 7.88 4.127 ;
      RECT 7.79 3.895 7.84 4.132 ;
      RECT 7.765 3.902 7.79 4.136 ;
      RECT 7.705 3.897 7.765 4.14 ;
      RECT 7.69 3.888 7.705 4.144 ;
      RECT 7.62 3.878 7.69 4.14 ;
      RECT 7.595 3.87 7.615 4.13 ;
      RECT 7.536 3.87 7.595 4.108 ;
      RECT 7.45 3.87 7.536 4.065 ;
      RECT 7.615 3.87 7.62 4.135 ;
      RECT 8.31 3.101 8.48 3.435 ;
      RECT 8.28 3.101 8.48 3.43 ;
      RECT 8.22 3.068 8.28 3.418 ;
      RECT 8.22 3.124 8.49 3.413 ;
      RECT 8.195 3.124 8.49 3.407 ;
      RECT 8.19 3.065 8.22 3.404 ;
      RECT 8.175 3.071 8.31 3.402 ;
      RECT 8.17 3.079 8.395 3.39 ;
      RECT 8.17 3.131 8.505 3.343 ;
      RECT 8.155 3.087 8.395 3.338 ;
      RECT 8.155 3.157 8.515 3.279 ;
      RECT 8.125 3.107 8.48 3.24 ;
      RECT 8.125 3.197 8.525 3.236 ;
      RECT 8.175 3.076 8.395 3.402 ;
      RECT 7.515 3.406 7.57 3.67 ;
      RECT 7.515 3.406 7.635 3.669 ;
      RECT 7.515 3.406 7.66 3.668 ;
      RECT 7.515 3.406 7.725 3.667 ;
      RECT 7.66 3.372 7.74 3.666 ;
      RECT 7.475 3.416 7.885 3.665 ;
      RECT 7.515 3.413 7.885 3.665 ;
      RECT 7.475 3.421 7.89 3.658 ;
      RECT 7.46 3.423 7.89 3.657 ;
      RECT 7.46 3.43 7.895 3.653 ;
      RECT 7.44 3.429 7.89 3.649 ;
      RECT 7.44 3.437 7.9 3.648 ;
      RECT 7.435 3.434 7.895 3.644 ;
      RECT 7.435 3.447 7.91 3.643 ;
      RECT 7.42 3.437 7.9 3.642 ;
      RECT 7.385 3.45 7.91 3.635 ;
      RECT 7.57 3.405 7.88 3.665 ;
      RECT 7.57 3.39 7.83 3.665 ;
      RECT 7.635 3.377 7.765 3.665 ;
      RECT 7.18 4.466 7.195 4.859 ;
      RECT 7.145 4.471 7.195 4.858 ;
      RECT 7.18 4.47 7.24 4.857 ;
      RECT 7.125 4.481 7.24 4.856 ;
      RECT 7.14 4.477 7.24 4.856 ;
      RECT 7.105 4.487 7.315 4.853 ;
      RECT 7.105 4.506 7.36 4.851 ;
      RECT 7.105 4.513 7.365 4.848 ;
      RECT 7.09 4.49 7.315 4.845 ;
      RECT 7.07 4.495 7.315 4.838 ;
      RECT 7.065 4.499 7.315 4.834 ;
      RECT 7.065 4.516 7.375 4.833 ;
      RECT 7.045 4.51 7.36 4.829 ;
      RECT 7.045 4.519 7.38 4.823 ;
      RECT 7.04 4.525 7.38 4.595 ;
      RECT 7.105 4.485 7.24 4.853 ;
      RECT 6.98 3.848 7.18 4.16 ;
      RECT 7.055 3.826 7.18 4.16 ;
      RECT 6.995 3.845 7.185 4.145 ;
      RECT 6.965 3.856 7.185 4.143 ;
      RECT 6.98 3.851 7.19 4.109 ;
      RECT 6.965 3.955 7.195 4.076 ;
      RECT 6.995 3.827 7.18 4.16 ;
      RECT 7.055 3.805 7.155 4.16 ;
      RECT 7.08 3.802 7.155 4.16 ;
      RECT 7.08 3.797 7.1 4.16 ;
      RECT 6.485 3.865 6.66 4.04 ;
      RECT 6.48 3.865 6.66 4.038 ;
      RECT 6.455 3.865 6.66 4.033 ;
      RECT 6.4 3.845 6.57 4.023 ;
      RECT 6.4 3.852 6.635 4.023 ;
      RECT 6.485 4.532 6.5 4.715 ;
      RECT 6.475 4.51 6.485 4.715 ;
      RECT 6.46 4.49 6.475 4.715 ;
      RECT 6.45 4.465 6.46 4.715 ;
      RECT 6.42 4.43 6.45 4.715 ;
      RECT 6.385 4.37 6.42 4.715 ;
      RECT 6.38 4.332 6.385 4.715 ;
      RECT 6.33 4.283 6.38 4.715 ;
      RECT 6.32 4.233 6.33 4.703 ;
      RECT 6.305 4.212 6.32 4.663 ;
      RECT 6.285 4.18 6.305 4.613 ;
      RECT 6.26 4.136 6.285 4.553 ;
      RECT 6.255 4.108 6.26 4.508 ;
      RECT 6.25 4.099 6.255 4.494 ;
      RECT 6.245 4.092 6.25 4.481 ;
      RECT 6.24 4.087 6.245 4.47 ;
      RECT 6.235 4.072 6.24 4.46 ;
      RECT 6.23 4.05 6.235 4.447 ;
      RECT 6.22 4.01 6.23 4.422 ;
      RECT 6.195 3.94 6.22 4.378 ;
      RECT 6.19 3.88 6.195 4.343 ;
      RECT 6.175 3.86 6.19 4.31 ;
      RECT 6.17 3.86 6.175 4.285 ;
      RECT 6.14 3.86 6.17 4.24 ;
      RECT 6.095 3.86 6.14 4.18 ;
      RECT 6.02 3.86 6.095 4.128 ;
      RECT 6.015 3.86 6.02 4.093 ;
      RECT 6.01 3.86 6.015 4.083 ;
      RECT 6.005 3.86 6.01 4.063 ;
      RECT 6.27 3.08 6.44 3.55 ;
      RECT 6.215 3.073 6.41 3.534 ;
      RECT 6.215 3.087 6.445 3.533 ;
      RECT 6.2 3.088 6.445 3.514 ;
      RECT 6.195 3.106 6.445 3.5 ;
      RECT 6.2 3.089 6.45 3.498 ;
      RECT 6.185 3.12 6.45 3.483 ;
      RECT 6.2 3.095 6.455 3.468 ;
      RECT 6.18 3.135 6.455 3.465 ;
      RECT 6.195 3.107 6.46 3.45 ;
      RECT 6.195 3.119 6.465 3.43 ;
      RECT 6.18 3.135 6.47 3.413 ;
      RECT 6.18 3.145 6.475 3.268 ;
      RECT 6.175 3.145 6.475 3.225 ;
      RECT 6.175 3.16 6.48 3.203 ;
      RECT 6.27 3.07 6.41 3.55 ;
      RECT 6.27 3.068 6.38 3.55 ;
      RECT 6.356 3.065 6.38 3.55 ;
      RECT 6.015 4.732 6.02 4.778 ;
      RECT 6.005 4.58 6.015 4.802 ;
      RECT 6 4.425 6.005 4.827 ;
      RECT 5.985 4.387 6 4.838 ;
      RECT 5.98 4.37 5.985 4.845 ;
      RECT 5.97 4.358 5.98 4.852 ;
      RECT 5.965 4.349 5.97 4.854 ;
      RECT 5.96 4.347 5.965 4.858 ;
      RECT 5.915 4.338 5.96 4.873 ;
      RECT 5.91 4.33 5.915 4.887 ;
      RECT 5.905 4.327 5.91 4.891 ;
      RECT 5.89 4.322 5.905 4.899 ;
      RECT 5.835 4.312 5.89 4.91 ;
      RECT 5.8 4.3 5.835 4.911 ;
      RECT 5.791 4.295 5.8 4.905 ;
      RECT 5.705 4.295 5.791 4.895 ;
      RECT 5.675 4.295 5.705 4.873 ;
      RECT 5.665 4.295 5.67 4.853 ;
      RECT 5.66 4.295 5.665 4.815 ;
      RECT 5.655 4.295 5.66 4.773 ;
      RECT 5.65 4.295 5.655 4.733 ;
      RECT 5.645 4.295 5.65 4.663 ;
      RECT 5.635 4.295 5.645 4.585 ;
      RECT 5.63 4.295 5.635 4.485 ;
      RECT 5.67 4.295 5.675 4.855 ;
      RECT 5.165 4.377 5.255 4.855 ;
      RECT 5.15 4.38 5.27 4.853 ;
      RECT 5.165 4.379 5.27 4.853 ;
      RECT 5.13 4.386 5.295 4.843 ;
      RECT 5.15 4.38 5.295 4.843 ;
      RECT 5.115 4.392 5.295 4.831 ;
      RECT 5.15 4.383 5.345 4.824 ;
      RECT 5.101 4.4 5.345 4.822 ;
      RECT 5.13 4.39 5.355 4.81 ;
      RECT 5.101 4.411 5.385 4.801 ;
      RECT 5.015 4.435 5.385 4.795 ;
      RECT 5.015 4.448 5.425 4.778 ;
      RECT 5.01 4.47 5.425 4.771 ;
      RECT 4.98 4.485 5.425 4.761 ;
      RECT 4.975 4.496 5.425 4.751 ;
      RECT 4.945 4.509 5.425 4.742 ;
      RECT 4.93 4.527 5.425 4.731 ;
      RECT 4.905 4.54 5.425 4.721 ;
      RECT 5.165 4.376 5.175 4.855 ;
      RECT 5.211 3.8 5.25 4.045 ;
      RECT 5.125 3.8 5.26 4.043 ;
      RECT 5.01 3.825 5.26 4.04 ;
      RECT 5.01 3.825 5.265 4.038 ;
      RECT 5.01 3.825 5.28 4.033 ;
      RECT 5.116 3.8 5.295 4.013 ;
      RECT 5.03 3.808 5.295 4.013 ;
      RECT 4.7 3.16 4.87 3.595 ;
      RECT 4.69 3.194 4.87 3.578 ;
      RECT 4.77 3.13 4.94 3.565 ;
      RECT 4.675 3.205 4.94 3.543 ;
      RECT 4.77 3.14 4.945 3.533 ;
      RECT 4.7 3.192 4.975 3.518 ;
      RECT 4.66 3.218 4.975 3.503 ;
      RECT 4.66 3.26 4.985 3.483 ;
      RECT 4.655 3.285 4.99 3.465 ;
      RECT 4.655 3.295 4.995 3.45 ;
      RECT 4.65 3.232 4.975 3.448 ;
      RECT 4.65 3.305 5 3.433 ;
      RECT 4.645 3.242 4.975 3.43 ;
      RECT 4.64 3.326 5.005 3.413 ;
      RECT 4.64 3.358 5.01 3.393 ;
      RECT 4.635 3.272 4.985 3.385 ;
      RECT 4.64 3.257 4.975 3.413 ;
      RECT 4.655 3.227 4.975 3.465 ;
      RECT 4.5 3.814 4.725 4.07 ;
      RECT 4.5 3.847 4.745 4.06 ;
      RECT 4.465 3.847 4.745 4.058 ;
      RECT 4.465 3.86 4.75 4.048 ;
      RECT 4.465 3.88 4.76 4.04 ;
      RECT 4.465 3.977 4.765 4.033 ;
      RECT 4.445 3.725 4.575 4.023 ;
      RECT 4.4 3.88 4.76 3.965 ;
      RECT 4.39 3.725 4.575 3.91 ;
      RECT 4.39 3.757 4.661 3.91 ;
      RECT 4.355 4.287 4.375 4.465 ;
      RECT 4.32 4.24 4.355 4.465 ;
      RECT 4.305 4.18 4.32 4.465 ;
      RECT 4.28 4.127 4.305 4.465 ;
      RECT 4.265 4.08 4.28 4.465 ;
      RECT 4.245 4.057 4.265 4.465 ;
      RECT 4.22 4.022 4.245 4.465 ;
      RECT 4.21 3.868 4.22 4.465 ;
      RECT 4.18 3.863 4.21 4.456 ;
      RECT 4.175 3.86 4.18 4.446 ;
      RECT 4.16 3.86 4.175 4.42 ;
      RECT 4.155 3.86 4.16 4.383 ;
      RECT 4.13 3.86 4.155 4.335 ;
      RECT 4.11 3.86 4.13 4.26 ;
      RECT 4.1 3.86 4.11 4.22 ;
      RECT 4.095 3.86 4.1 4.195 ;
      RECT 4.09 3.86 4.095 4.178 ;
      RECT 4.085 3.86 4.09 4.16 ;
      RECT 4.08 3.861 4.085 4.15 ;
      RECT 4.07 3.863 4.08 4.118 ;
      RECT 4.06 3.865 4.07 4.085 ;
      RECT 4.05 3.868 4.06 4.058 ;
      RECT 4.375 4.295 4.6 4.465 ;
      RECT 3.705 3.107 3.875 3.56 ;
      RECT 3.705 3.107 3.965 3.526 ;
      RECT 3.705 3.107 3.995 3.51 ;
      RECT 3.705 3.107 4.025 3.483 ;
      RECT 3.961 3.085 4.04 3.465 ;
      RECT 3.74 3.092 4.045 3.45 ;
      RECT 3.74 3.1 4.055 3.413 ;
      RECT 3.7 3.127 4.055 3.385 ;
      RECT 3.685 3.14 4.055 3.35 ;
      RECT 3.705 3.115 4.075 3.34 ;
      RECT 3.68 3.18 4.075 3.31 ;
      RECT 3.68 3.21 4.08 3.293 ;
      RECT 3.675 3.24 4.08 3.28 ;
      RECT 3.74 3.089 4.04 3.465 ;
      RECT 3.875 3.086 3.961 3.544 ;
      RECT 3.826 3.087 4.04 3.465 ;
      RECT 3.97 4.747 4.015 4.94 ;
      RECT 3.96 4.717 3.97 4.94 ;
      RECT 3.955 4.702 3.96 4.94 ;
      RECT 3.915 4.612 3.955 4.94 ;
      RECT 3.91 4.525 3.915 4.94 ;
      RECT 3.9 4.495 3.91 4.94 ;
      RECT 3.895 4.455 3.9 4.94 ;
      RECT 3.885 4.417 3.895 4.94 ;
      RECT 3.88 4.382 3.885 4.94 ;
      RECT 3.86 4.335 3.88 4.94 ;
      RECT 3.845 4.26 3.86 4.94 ;
      RECT 3.84 4.215 3.845 4.935 ;
      RECT 3.835 4.195 3.84 4.908 ;
      RECT 3.83 4.175 3.835 4.893 ;
      RECT 3.825 4.15 3.83 4.873 ;
      RECT 3.82 4.128 3.825 4.858 ;
      RECT 3.815 4.106 3.82 4.84 ;
      RECT 3.81 4.085 3.815 4.83 ;
      RECT 3.8 4.057 3.81 4.8 ;
      RECT 3.79 4.02 3.8 4.768 ;
      RECT 3.78 3.98 3.79 4.735 ;
      RECT 3.77 3.958 3.78 4.705 ;
      RECT 3.74 3.91 3.77 4.637 ;
      RECT 3.725 3.87 3.74 4.564 ;
      RECT 3.715 3.87 3.725 4.53 ;
      RECT 3.71 3.87 3.715 4.505 ;
      RECT 3.705 3.87 3.71 4.49 ;
      RECT 3.7 3.87 3.705 4.468 ;
      RECT 3.695 3.87 3.7 4.455 ;
      RECT 3.68 3.87 3.695 4.42 ;
      RECT 3.66 3.87 3.68 4.36 ;
      RECT 3.65 3.87 3.66 4.31 ;
      RECT 3.63 3.87 3.65 4.258 ;
      RECT 3.61 3.87 3.63 4.215 ;
      RECT 3.6 3.87 3.61 4.203 ;
      RECT 3.57 3.87 3.6 4.19 ;
      RECT 3.54 3.891 3.57 4.17 ;
      RECT 3.53 3.919 3.54 4.15 ;
      RECT 3.515 3.936 3.53 4.118 ;
      RECT 3.51 3.95 3.515 4.085 ;
      RECT 3.505 3.958 3.51 4.058 ;
      RECT 3.5 3.966 3.505 4.02 ;
      RECT 3.505 4.49 3.51 4.825 ;
      RECT 3.47 4.477 3.505 4.824 ;
      RECT 3.4 4.417 3.47 4.823 ;
      RECT 3.32 4.36 3.4 4.822 ;
      RECT 3.185 4.32 3.32 4.821 ;
      RECT 3.185 4.507 3.52 4.81 ;
      RECT 3.145 4.507 3.52 4.8 ;
      RECT 3.145 4.525 3.525 4.795 ;
      RECT 3.145 4.615 3.53 4.785 ;
      RECT 3.14 4.31 3.305 4.765 ;
      RECT 3.135 4.31 3.305 4.508 ;
      RECT 3.135 4.467 3.5 4.508 ;
      RECT 3.135 4.455 3.495 4.508 ;
      RECT 2.03 7.3 2.2 10.59 ;
      RECT 1.985 7.29 2.155 7.35 ;
      RECT 1.17 10.14 1.34 10.59 ;
      RECT 1.225 8.36 1.395 10.31 ;
      RECT 1.17 7.3 1.34 8.53 ;
      RECT 0.65 7.3 0.82 10.59 ;
      RECT 0.65 9.6 1.055 9.93 ;
      RECT 0.65 8.76 1.055 9.09 ;
      RECT 81.175 10.085 81.345 10.595 ;
      RECT 80.185 1.865 80.355 2.375 ;
      RECT 80.185 3.685 80.355 5.155 ;
      RECT 80.185 7.305 80.355 8.775 ;
      RECT 80.185 10.085 80.355 10.595 ;
      RECT 78.825 1.87 78.995 5.16 ;
      RECT 78.825 7.3 78.995 10.59 ;
      RECT 78.395 1.87 78.565 2.38 ;
      RECT 78.395 2.95 78.565 5.16 ;
      RECT 78.395 7.3 78.565 9.51 ;
      RECT 78.395 10.08 78.565 10.59 ;
      RECT 76.005 4.145 76.375 4.515 ;
      RECT 74.045 7.3 74.215 10.59 ;
      RECT 73.615 7.3 73.785 9.51 ;
      RECT 73.615 10.08 73.785 10.59 ;
      RECT 65.39 10.085 65.56 10.595 ;
      RECT 64.4 1.865 64.57 2.375 ;
      RECT 64.4 3.685 64.57 5.155 ;
      RECT 64.4 7.305 64.57 8.775 ;
      RECT 64.4 10.085 64.57 10.595 ;
      RECT 63.04 1.87 63.21 5.16 ;
      RECT 63.04 7.3 63.21 10.59 ;
      RECT 62.61 1.87 62.78 2.38 ;
      RECT 62.61 2.95 62.78 5.16 ;
      RECT 62.61 7.3 62.78 9.51 ;
      RECT 62.61 10.08 62.78 10.59 ;
      RECT 60.22 4.145 60.59 4.515 ;
      RECT 58.26 7.3 58.43 10.59 ;
      RECT 57.83 7.3 58 9.51 ;
      RECT 57.83 10.08 58 10.59 ;
      RECT 49.605 10.085 49.775 10.595 ;
      RECT 48.615 1.865 48.785 2.375 ;
      RECT 48.615 3.685 48.785 5.155 ;
      RECT 48.615 7.305 48.785 8.775 ;
      RECT 48.615 10.085 48.785 10.595 ;
      RECT 47.255 1.87 47.425 5.16 ;
      RECT 47.255 7.3 47.425 10.59 ;
      RECT 46.825 1.87 46.995 2.38 ;
      RECT 46.825 2.95 46.995 5.16 ;
      RECT 46.825 7.3 46.995 9.51 ;
      RECT 46.825 10.08 46.995 10.59 ;
      RECT 44.435 4.145 44.805 4.515 ;
      RECT 42.475 7.3 42.645 10.59 ;
      RECT 42.045 7.3 42.215 9.51 ;
      RECT 42.045 10.08 42.215 10.59 ;
      RECT 33.83 10.085 34 10.595 ;
      RECT 32.84 1.865 33.01 2.375 ;
      RECT 32.84 3.685 33.01 5.155 ;
      RECT 32.84 7.305 33.01 8.775 ;
      RECT 32.84 10.085 33.01 10.595 ;
      RECT 31.48 1.87 31.65 5.16 ;
      RECT 31.48 7.3 31.65 10.59 ;
      RECT 31.05 1.87 31.22 2.38 ;
      RECT 31.05 2.95 31.22 5.16 ;
      RECT 31.05 7.3 31.22 9.51 ;
      RECT 31.05 10.08 31.22 10.59 ;
      RECT 28.66 4.145 29.03 4.515 ;
      RECT 26.7 7.3 26.87 10.59 ;
      RECT 26.27 7.3 26.44 9.51 ;
      RECT 26.27 10.08 26.44 10.59 ;
      RECT 18.05 10.085 18.22 10.595 ;
      RECT 17.06 1.865 17.23 2.375 ;
      RECT 17.06 3.685 17.23 5.155 ;
      RECT 17.06 7.305 17.23 8.775 ;
      RECT 17.06 10.085 17.23 10.595 ;
      RECT 15.7 1.87 15.87 5.16 ;
      RECT 15.7 7.3 15.87 10.59 ;
      RECT 15.27 1.87 15.44 2.38 ;
      RECT 15.27 2.95 15.44 5.16 ;
      RECT 15.27 7.3 15.44 9.51 ;
      RECT 15.27 10.08 15.44 10.59 ;
      RECT 12.88 4.145 13.25 4.515 ;
      RECT 10.92 7.3 11.09 10.59 ;
      RECT 10.49 7.3 10.66 9.51 ;
      RECT 10.49 10.08 10.66 10.59 ;
      RECT 1.6 7.3 1.77 9.51 ;
      RECT 1.6 10.08 1.77 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r2
  CLASS BLOCK ;
  ORIGIN -9.41 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r2 ;
  SIZE 81.775 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 27.51 1.865 27.68 2.375 ;
        RECT 27.51 3.685 27.68 5.155 ;
      LAYER met1 ;
        RECT 27.45 3.655 27.74 3.885 ;
        RECT 27.45 2.175 27.74 2.405 ;
        RECT 27.51 2.175 27.68 3.885 ;
      LAYER mcon ;
        RECT 27.51 3.685 27.68 3.855 ;
        RECT 27.51 2.205 27.68 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 43.29 1.865 43.46 2.375 ;
        RECT 43.29 3.685 43.46 5.155 ;
      LAYER met1 ;
        RECT 43.23 3.655 43.52 3.885 ;
        RECT 43.23 2.175 43.52 2.405 ;
        RECT 43.29 2.175 43.46 3.885 ;
      LAYER mcon ;
        RECT 43.29 3.685 43.46 3.855 ;
        RECT 43.29 2.205 43.46 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 59.065 1.865 59.235 2.375 ;
        RECT 59.065 3.685 59.235 5.155 ;
      LAYER met1 ;
        RECT 59.005 3.655 59.295 3.885 ;
        RECT 59.005 2.175 59.295 2.405 ;
        RECT 59.065 2.175 59.235 3.885 ;
      LAYER mcon ;
        RECT 59.065 3.685 59.235 3.855 ;
        RECT 59.065 2.205 59.235 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 74.85 1.865 75.02 2.375 ;
        RECT 74.85 3.685 75.02 5.155 ;
      LAYER met1 ;
        RECT 74.79 3.655 75.08 3.885 ;
        RECT 74.79 2.175 75.08 2.405 ;
        RECT 74.85 2.175 75.02 3.885 ;
      LAYER mcon ;
        RECT 74.85 3.685 75.02 3.855 ;
        RECT 74.85 2.205 75.02 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 90.635 1.865 90.805 2.375 ;
        RECT 90.635 3.685 90.805 5.155 ;
      LAYER met1 ;
        RECT 90.575 3.655 90.865 3.885 ;
        RECT 90.575 2.175 90.865 2.405 ;
        RECT 90.635 2.175 90.805 3.885 ;
      LAYER mcon ;
        RECT 90.635 3.685 90.805 3.855 ;
        RECT 90.635 2.205 90.805 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 23.275 8.14 23.625 8.49 ;
        RECT 23.27 4 23.62 4.35 ;
        RECT 23.345 4 23.52 8.49 ;
      LAYER li1 ;
        RECT 23.36 2.955 23.53 4.23 ;
        RECT 23.36 8.23 23.53 9.505 ;
        RECT 18.58 8.23 18.75 9.505 ;
      LAYER met1 ;
        RECT 23.27 4.06 23.76 4.23 ;
        RECT 23.27 4 23.62 4.35 ;
        RECT 18.52 8.23 23.76 8.4 ;
        RECT 23.275 8.14 23.625 8.49 ;
        RECT 18.52 8.2 18.81 8.43 ;
      LAYER via1 ;
        RECT 23.37 4.1 23.52 4.25 ;
        RECT 23.375 8.24 23.525 8.39 ;
      LAYER mcon ;
        RECT 18.58 8.23 18.75 8.4 ;
        RECT 23.36 8.23 23.53 8.4 ;
        RECT 23.36 4.06 23.53 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 39.055 8.14 39.405 8.49 ;
        RECT 39.05 4 39.4 4.35 ;
        RECT 39.125 4 39.3 8.49 ;
      LAYER li1 ;
        RECT 39.14 2.955 39.31 4.23 ;
        RECT 39.14 8.23 39.31 9.505 ;
        RECT 34.36 8.23 34.53 9.505 ;
      LAYER met1 ;
        RECT 39.05 4.06 39.54 4.23 ;
        RECT 39.05 4 39.4 4.35 ;
        RECT 34.3 8.23 39.54 8.4 ;
        RECT 39.055 8.14 39.405 8.49 ;
        RECT 34.3 8.2 34.59 8.43 ;
      LAYER via1 ;
        RECT 39.15 4.1 39.3 4.25 ;
        RECT 39.155 8.24 39.305 8.39 ;
      LAYER mcon ;
        RECT 34.36 8.23 34.53 8.4 ;
        RECT 39.14 8.23 39.31 8.4 ;
        RECT 39.14 4.06 39.31 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 54.83 8.14 55.18 8.49 ;
        RECT 54.825 4 55.175 4.35 ;
        RECT 54.9 4 55.075 8.49 ;
      LAYER li1 ;
        RECT 54.915 2.955 55.085 4.23 ;
        RECT 54.915 8.23 55.085 9.505 ;
        RECT 50.135 8.23 50.305 9.505 ;
      LAYER met1 ;
        RECT 54.825 4.06 55.315 4.23 ;
        RECT 54.825 4 55.175 4.35 ;
        RECT 50.075 8.23 55.315 8.4 ;
        RECT 54.83 8.14 55.18 8.49 ;
        RECT 50.075 8.2 50.365 8.43 ;
      LAYER via1 ;
        RECT 54.925 4.1 55.075 4.25 ;
        RECT 54.93 8.24 55.08 8.39 ;
      LAYER mcon ;
        RECT 50.135 8.23 50.305 8.4 ;
        RECT 54.915 8.23 55.085 8.4 ;
        RECT 54.915 4.06 55.085 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 70.615 8.14 70.965 8.49 ;
        RECT 70.61 4 70.96 4.35 ;
        RECT 70.685 4 70.86 8.49 ;
      LAYER li1 ;
        RECT 70.7 2.955 70.87 4.23 ;
        RECT 70.7 8.23 70.87 9.505 ;
        RECT 65.92 8.23 66.09 9.505 ;
      LAYER met1 ;
        RECT 70.61 4.06 71.1 4.23 ;
        RECT 70.61 4 70.96 4.35 ;
        RECT 65.86 8.23 71.1 8.4 ;
        RECT 70.615 8.14 70.965 8.49 ;
        RECT 65.86 8.2 66.15 8.43 ;
      LAYER via1 ;
        RECT 70.71 4.1 70.86 4.25 ;
        RECT 70.715 8.24 70.865 8.39 ;
      LAYER mcon ;
        RECT 65.92 8.23 66.09 8.4 ;
        RECT 70.7 8.23 70.87 8.4 ;
        RECT 70.7 4.06 70.87 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 86.4 8.14 86.75 8.49 ;
        RECT 86.395 4 86.745 4.35 ;
        RECT 86.47 4 86.645 8.49 ;
      LAYER li1 ;
        RECT 86.485 2.955 86.655 4.23 ;
        RECT 86.485 8.23 86.655 9.505 ;
        RECT 81.705 8.23 81.875 9.505 ;
      LAYER met1 ;
        RECT 86.395 4.06 86.885 4.23 ;
        RECT 86.395 4 86.745 4.35 ;
        RECT 81.645 8.23 86.885 8.4 ;
        RECT 86.4 8.14 86.75 8.49 ;
        RECT 81.645 8.2 81.935 8.43 ;
      LAYER via1 ;
        RECT 86.495 4.1 86.645 4.25 ;
        RECT 86.5 8.24 86.65 8.39 ;
      LAYER mcon ;
        RECT 81.705 8.23 81.875 8.4 ;
        RECT 86.485 8.23 86.655 8.4 ;
        RECT 86.485 4.06 86.655 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 9.705 8.23 9.875 9.505 ;
      LAYER met1 ;
        RECT 9.585 8.23 10.105 8.4 ;
        RECT 9.585 8.2 9.935 8.43 ;
      LAYER mcon ;
        RECT 9.705 8.23 9.875 8.4 ;
    END
  END start
  OBS
    LAYER met3 ;
      RECT 82.975 9.325 83.345 9.695 ;
      RECT 83.015 9.005 83.345 9.695 ;
      RECT 83.015 9.005 85.805 9.31 ;
      RECT 85.5 4.145 85.805 9.31 ;
      RECT 85.465 4.145 85.835 4.515 ;
      RECT 84.725 2.11 85.03 5.315 ;
      RECT 84.475 4.27 85.03 5 ;
      RECT 84.685 2.11 85.055 2.48 ;
      RECT 80.835 3.145 81.165 4.04 ;
      RECT 79.955 3.31 80.285 4.04 ;
      RECT 80.83 3.145 81.2 3.945 ;
      RECT 83.995 3.145 84.325 3.875 ;
      RECT 83.955 3.03 84.135 3.68 ;
      RECT 79.965 3.145 84.325 3.515 ;
      RECT 80.455 4.83 80.785 5.16 ;
      RECT 79.25 4.845 80.785 5.145 ;
      RECT 79.25 3.725 79.55 5.145 ;
      RECT 78.995 3.71 79.325 4.04 ;
      RECT 67.19 9.325 67.56 9.695 ;
      RECT 67.23 9.005 67.56 9.695 ;
      RECT 67.23 9.005 70.02 9.31 ;
      RECT 69.715 4.145 70.02 9.31 ;
      RECT 69.68 4.145 70.05 4.515 ;
      RECT 68.94 2.11 69.245 5.315 ;
      RECT 68.69 4.27 69.245 5 ;
      RECT 68.9 2.11 69.27 2.48 ;
      RECT 65.05 3.145 65.38 4.04 ;
      RECT 64.17 3.31 64.5 4.04 ;
      RECT 65.045 3.145 65.415 3.945 ;
      RECT 68.21 3.145 68.54 3.875 ;
      RECT 68.17 3.03 68.35 3.68 ;
      RECT 64.18 3.145 68.54 3.515 ;
      RECT 64.67 4.83 65 5.16 ;
      RECT 63.465 4.845 65 5.145 ;
      RECT 63.465 3.725 63.765 5.145 ;
      RECT 63.21 3.71 63.54 4.04 ;
      RECT 51.405 9.325 51.775 9.695 ;
      RECT 51.445 9.005 51.775 9.695 ;
      RECT 51.445 9.005 54.235 9.31 ;
      RECT 53.93 4.145 54.235 9.31 ;
      RECT 53.895 4.145 54.265 4.515 ;
      RECT 53.155 2.11 53.46 5.315 ;
      RECT 52.905 4.27 53.46 5 ;
      RECT 53.115 2.11 53.485 2.48 ;
      RECT 49.265 3.145 49.595 4.04 ;
      RECT 48.385 3.31 48.715 4.04 ;
      RECT 49.26 3.145 49.63 3.945 ;
      RECT 52.425 3.145 52.755 3.875 ;
      RECT 52.385 3.03 52.565 3.68 ;
      RECT 48.395 3.145 52.755 3.515 ;
      RECT 48.885 4.83 49.215 5.16 ;
      RECT 47.68 4.845 49.215 5.145 ;
      RECT 47.68 3.725 47.98 5.145 ;
      RECT 47.425 3.71 47.755 4.04 ;
      RECT 35.63 9.325 36 9.695 ;
      RECT 35.67 9.005 36 9.695 ;
      RECT 35.67 9.005 38.46 9.31 ;
      RECT 38.155 4.145 38.46 9.31 ;
      RECT 38.12 4.145 38.49 4.515 ;
      RECT 37.38 2.11 37.685 5.315 ;
      RECT 37.13 4.27 37.685 5 ;
      RECT 37.34 2.11 37.71 2.48 ;
      RECT 33.49 3.145 33.82 4.04 ;
      RECT 32.61 3.31 32.94 4.04 ;
      RECT 33.485 3.145 33.855 3.945 ;
      RECT 36.65 3.145 36.98 3.875 ;
      RECT 36.61 3.03 36.79 3.68 ;
      RECT 32.62 3.145 36.98 3.515 ;
      RECT 33.11 4.83 33.44 5.16 ;
      RECT 31.905 4.845 33.44 5.145 ;
      RECT 31.905 3.725 32.205 5.145 ;
      RECT 31.65 3.71 31.98 4.04 ;
      RECT 19.85 9.325 20.22 9.695 ;
      RECT 19.89 9.005 20.22 9.695 ;
      RECT 19.89 9.005 22.68 9.31 ;
      RECT 22.375 4.145 22.68 9.31 ;
      RECT 22.34 4.145 22.71 4.515 ;
      RECT 21.6 2.11 21.905 5.315 ;
      RECT 21.35 4.27 21.905 5 ;
      RECT 21.56 2.11 21.93 2.48 ;
      RECT 17.71 3.145 18.04 4.04 ;
      RECT 16.83 3.31 17.16 4.04 ;
      RECT 17.705 3.145 18.075 3.945 ;
      RECT 20.87 3.145 21.2 3.875 ;
      RECT 20.83 3.03 21.01 3.68 ;
      RECT 16.84 3.145 21.2 3.515 ;
      RECT 17.33 4.83 17.66 5.16 ;
      RECT 16.125 4.845 17.66 5.145 ;
      RECT 16.125 3.725 16.425 5.145 ;
      RECT 15.87 3.71 16.2 4.04 ;
      RECT 82.395 3.87 82.725 4.6 ;
      RECT 78.275 3.71 78.605 4.44 ;
      RECT 77.275 3.15 77.605 3.88 ;
      RECT 75.835 3.87 76.165 4.6 ;
      RECT 66.61 3.87 66.94 4.6 ;
      RECT 62.49 3.71 62.82 4.44 ;
      RECT 61.49 3.15 61.82 3.88 ;
      RECT 60.05 3.87 60.38 4.6 ;
      RECT 50.825 3.87 51.155 4.6 ;
      RECT 46.705 3.71 47.035 4.44 ;
      RECT 45.705 3.15 46.035 3.88 ;
      RECT 44.265 3.87 44.595 4.6 ;
      RECT 35.05 3.87 35.38 4.6 ;
      RECT 30.93 3.71 31.26 4.44 ;
      RECT 29.93 3.15 30.26 3.88 ;
      RECT 28.49 3.87 28.82 4.6 ;
      RECT 19.27 3.87 19.6 4.6 ;
      RECT 15.15 3.71 15.48 4.44 ;
      RECT 14.15 3.15 14.48 3.88 ;
      RECT 12.71 3.87 13.04 4.6 ;
      RECT 9.415 0 10.22 0.38 ;
      RECT 9.415 10.785 10.22 11.165 ;
    LAYER via2 ;
      RECT 85.55 4.23 85.75 4.43 ;
      RECT 84.77 2.195 84.97 2.395 ;
      RECT 84.54 4.335 84.74 4.535 ;
      RECT 84.06 3.61 84.26 3.81 ;
      RECT 83.06 9.41 83.26 9.61 ;
      RECT 82.46 4.335 82.66 4.535 ;
      RECT 80.9 3.775 81.1 3.975 ;
      RECT 80.52 4.895 80.72 5.095 ;
      RECT 80.02 3.775 80.22 3.975 ;
      RECT 79.06 3.775 79.26 3.975 ;
      RECT 78.34 3.775 78.54 3.975 ;
      RECT 77.34 3.215 77.54 3.415 ;
      RECT 75.9 4.335 76.1 4.535 ;
      RECT 69.765 4.23 69.965 4.43 ;
      RECT 68.985 2.195 69.185 2.395 ;
      RECT 68.755 4.335 68.955 4.535 ;
      RECT 68.275 3.61 68.475 3.81 ;
      RECT 67.275 9.41 67.475 9.61 ;
      RECT 66.675 4.335 66.875 4.535 ;
      RECT 65.115 3.775 65.315 3.975 ;
      RECT 64.735 4.895 64.935 5.095 ;
      RECT 64.235 3.775 64.435 3.975 ;
      RECT 63.275 3.775 63.475 3.975 ;
      RECT 62.555 3.775 62.755 3.975 ;
      RECT 61.555 3.215 61.755 3.415 ;
      RECT 60.115 4.335 60.315 4.535 ;
      RECT 53.98 4.23 54.18 4.43 ;
      RECT 53.2 2.195 53.4 2.395 ;
      RECT 52.97 4.335 53.17 4.535 ;
      RECT 52.49 3.61 52.69 3.81 ;
      RECT 51.49 9.41 51.69 9.61 ;
      RECT 50.89 4.335 51.09 4.535 ;
      RECT 49.33 3.775 49.53 3.975 ;
      RECT 48.95 4.895 49.15 5.095 ;
      RECT 48.45 3.775 48.65 3.975 ;
      RECT 47.49 3.775 47.69 3.975 ;
      RECT 46.77 3.775 46.97 3.975 ;
      RECT 45.77 3.215 45.97 3.415 ;
      RECT 44.33 4.335 44.53 4.535 ;
      RECT 38.205 4.23 38.405 4.43 ;
      RECT 37.425 2.195 37.625 2.395 ;
      RECT 37.195 4.335 37.395 4.535 ;
      RECT 36.715 3.61 36.915 3.81 ;
      RECT 35.715 9.41 35.915 9.61 ;
      RECT 35.115 4.335 35.315 4.535 ;
      RECT 33.555 3.775 33.755 3.975 ;
      RECT 33.175 4.895 33.375 5.095 ;
      RECT 32.675 3.775 32.875 3.975 ;
      RECT 31.715 3.775 31.915 3.975 ;
      RECT 30.995 3.775 31.195 3.975 ;
      RECT 29.995 3.215 30.195 3.415 ;
      RECT 28.555 4.335 28.755 4.535 ;
      RECT 22.425 4.23 22.625 4.43 ;
      RECT 21.645 2.195 21.845 2.395 ;
      RECT 21.415 4.335 21.615 4.535 ;
      RECT 20.935 3.61 21.135 3.81 ;
      RECT 19.935 9.41 20.135 9.61 ;
      RECT 19.335 4.335 19.535 4.535 ;
      RECT 17.775 3.775 17.975 3.975 ;
      RECT 17.395 4.895 17.595 5.095 ;
      RECT 16.895 3.775 17.095 3.975 ;
      RECT 15.935 3.775 16.135 3.975 ;
      RECT 15.215 3.775 15.415 3.975 ;
      RECT 14.215 3.215 14.415 3.415 ;
      RECT 12.775 4.335 12.975 4.535 ;
      RECT 9.695 0.09 9.895 0.29 ;
      RECT 9.695 10.875 9.895 11.075 ;
    LAYER met2 ;
      RECT 10.64 10.685 90.81 10.855 ;
      RECT 90.64 9.56 90.81 10.855 ;
      RECT 10.64 8.54 10.81 10.855 ;
      RECT 90.61 9.56 90.96 9.91 ;
      RECT 10.58 8.54 10.87 8.89 ;
      RECT 87.45 8.505 87.77 8.83 ;
      RECT 87.48 7.98 87.65 8.83 ;
      RECT 87.48 7.98 87.655 8.33 ;
      RECT 87.48 7.98 88.455 8.155 ;
      RECT 88.28 3.26 88.455 8.155 ;
      RECT 88.225 3.26 88.575 3.61 ;
      RECT 88.25 8.94 88.575 9.265 ;
      RECT 87.135 9.03 88.575 9.2 ;
      RECT 87.135 3.69 87.295 9.2 ;
      RECT 87.45 3.66 87.77 3.98 ;
      RECT 87.135 3.69 87.77 3.86 ;
      RECT 75.86 4.295 76.14 4.575 ;
      RECT 75.83 4.295 76.14 4.56 ;
      RECT 75.825 4.295 76.14 4.558 ;
      RECT 75.82 2.625 75.99 4.552 ;
      RECT 75.815 4.262 76.085 4.545 ;
      RECT 75.81 4.295 76.14 4.538 ;
      RECT 75.78 4.265 76.085 4.525 ;
      RECT 75.78 4.292 76.105 4.525 ;
      RECT 75.78 4.282 76.1 4.525 ;
      RECT 75.78 4.267 76.095 4.525 ;
      RECT 75.82 4.257 76.085 4.552 ;
      RECT 75.82 4.252 76.075 4.552 ;
      RECT 75.82 4.251 76.06 4.552 ;
      RECT 85.79 2.635 86.14 2.985 ;
      RECT 85.785 2.635 86.14 2.89 ;
      RECT 75.82 2.625 86.03 2.795 ;
      RECT 85.465 4.145 85.835 4.515 ;
      RECT 85.55 3.53 85.72 4.515 ;
      RECT 81.57 3.75 81.805 4.01 ;
      RECT 84.715 3.53 84.88 3.79 ;
      RECT 84.62 3.52 84.635 3.79 ;
      RECT 84.715 3.53 85.72 3.71 ;
      RECT 83.22 3.09 83.26 3.23 ;
      RECT 84.635 3.525 84.715 3.79 ;
      RECT 84.58 3.52 84.62 3.756 ;
      RECT 84.566 3.52 84.58 3.756 ;
      RECT 84.48 3.525 84.566 3.758 ;
      RECT 84.435 3.532 84.48 3.76 ;
      RECT 84.405 3.532 84.435 3.762 ;
      RECT 84.38 3.527 84.405 3.764 ;
      RECT 84.35 3.523 84.38 3.773 ;
      RECT 84.34 3.52 84.35 3.785 ;
      RECT 84.335 3.52 84.34 3.793 ;
      RECT 84.33 3.52 84.335 3.798 ;
      RECT 84.32 3.519 84.33 3.808 ;
      RECT 84.315 3.518 84.32 3.818 ;
      RECT 84.3 3.517 84.315 3.823 ;
      RECT 84.272 3.514 84.3 3.85 ;
      RECT 84.186 3.506 84.272 3.85 ;
      RECT 84.1 3.495 84.186 3.85 ;
      RECT 84.06 3.48 84.1 3.85 ;
      RECT 84.02 3.454 84.06 3.85 ;
      RECT 84.015 3.436 84.02 3.662 ;
      RECT 84.005 3.432 84.015 3.652 ;
      RECT 83.99 3.422 84.005 3.639 ;
      RECT 83.97 3.406 83.99 3.624 ;
      RECT 83.955 3.391 83.97 3.609 ;
      RECT 83.945 3.38 83.955 3.599 ;
      RECT 83.92 3.364 83.945 3.588 ;
      RECT 83.915 3.351 83.92 3.578 ;
      RECT 83.91 3.347 83.915 3.573 ;
      RECT 83.855 3.333 83.91 3.551 ;
      RECT 83.816 3.314 83.855 3.515 ;
      RECT 83.73 3.288 83.816 3.468 ;
      RECT 83.726 3.27 83.73 3.434 ;
      RECT 83.64 3.251 83.726 3.412 ;
      RECT 83.635 3.233 83.64 3.39 ;
      RECT 83.63 3.231 83.635 3.388 ;
      RECT 83.62 3.23 83.63 3.383 ;
      RECT 83.56 3.217 83.62 3.369 ;
      RECT 83.515 3.195 83.56 3.348 ;
      RECT 83.455 3.172 83.515 3.327 ;
      RECT 83.391 3.147 83.455 3.302 ;
      RECT 83.305 3.117 83.391 3.271 ;
      RECT 83.29 3.097 83.305 3.25 ;
      RECT 83.26 3.092 83.29 3.241 ;
      RECT 83.207 3.09 83.22 3.23 ;
      RECT 83.121 3.09 83.207 3.232 ;
      RECT 83.035 3.09 83.121 3.234 ;
      RECT 83.015 3.09 83.035 3.238 ;
      RECT 82.97 3.092 83.015 3.249 ;
      RECT 82.93 3.102 82.97 3.265 ;
      RECT 82.926 3.111 82.93 3.273 ;
      RECT 82.84 3.131 82.926 3.289 ;
      RECT 82.83 3.15 82.84 3.307 ;
      RECT 82.825 3.152 82.83 3.31 ;
      RECT 82.815 3.156 82.825 3.313 ;
      RECT 82.795 3.161 82.815 3.323 ;
      RECT 82.765 3.171 82.795 3.343 ;
      RECT 82.76 3.178 82.765 3.357 ;
      RECT 82.75 3.182 82.76 3.364 ;
      RECT 82.735 3.19 82.75 3.375 ;
      RECT 82.725 3.2 82.735 3.386 ;
      RECT 82.715 3.207 82.725 3.394 ;
      RECT 82.69 3.22 82.715 3.409 ;
      RECT 82.626 3.256 82.69 3.448 ;
      RECT 82.54 3.319 82.626 3.512 ;
      RECT 82.505 3.37 82.54 3.565 ;
      RECT 82.5 3.387 82.505 3.582 ;
      RECT 82.485 3.396 82.5 3.589 ;
      RECT 82.465 3.411 82.485 3.603 ;
      RECT 82.46 3.422 82.465 3.613 ;
      RECT 82.44 3.435 82.46 3.623 ;
      RECT 82.435 3.445 82.44 3.633 ;
      RECT 82.42 3.45 82.435 3.642 ;
      RECT 82.41 3.46 82.42 3.653 ;
      RECT 82.38 3.477 82.41 3.67 ;
      RECT 82.37 3.495 82.38 3.688 ;
      RECT 82.355 3.506 82.37 3.699 ;
      RECT 82.315 3.53 82.355 3.715 ;
      RECT 82.28 3.564 82.315 3.732 ;
      RECT 82.25 3.587 82.28 3.744 ;
      RECT 82.235 3.597 82.25 3.753 ;
      RECT 82.195 3.607 82.235 3.764 ;
      RECT 82.175 3.618 82.195 3.776 ;
      RECT 82.17 3.622 82.175 3.783 ;
      RECT 82.155 3.626 82.17 3.788 ;
      RECT 82.145 3.631 82.155 3.793 ;
      RECT 82.14 3.634 82.145 3.796 ;
      RECT 82.11 3.64 82.14 3.803 ;
      RECT 82.075 3.65 82.11 3.817 ;
      RECT 82.015 3.665 82.075 3.837 ;
      RECT 81.96 3.685 82.015 3.861 ;
      RECT 81.931 3.7 81.96 3.879 ;
      RECT 81.845 3.72 81.931 3.904 ;
      RECT 81.84 3.735 81.845 3.924 ;
      RECT 81.83 3.738 81.84 3.925 ;
      RECT 81.805 3.745 81.83 4.01 ;
      RECT 84.5 4.238 84.78 4.575 ;
      RECT 84.5 4.248 84.785 4.533 ;
      RECT 84.5 4.257 84.79 4.43 ;
      RECT 84.5 4.272 84.795 4.298 ;
      RECT 84.5 4.1 84.76 4.575 ;
      RECT 74.8 8.94 75.15 9.29 ;
      RECT 83.625 8.895 83.975 9.245 ;
      RECT 74.8 8.97 83.975 9.17 ;
      RECT 82.22 4.98 82.23 5.17 ;
      RECT 80.48 4.855 80.76 5.135 ;
      RECT 83.525 3.795 83.53 4.28 ;
      RECT 83.42 3.795 83.48 4.055 ;
      RECT 83.745 4.765 83.75 4.84 ;
      RECT 83.735 4.632 83.745 4.875 ;
      RECT 83.725 4.467 83.735 4.896 ;
      RECT 83.72 4.337 83.725 4.912 ;
      RECT 83.71 4.227 83.72 4.928 ;
      RECT 83.705 4.126 83.71 4.945 ;
      RECT 83.7 4.108 83.705 4.955 ;
      RECT 83.695 4.09 83.7 4.965 ;
      RECT 83.685 4.065 83.695 4.98 ;
      RECT 83.68 4.045 83.685 4.995 ;
      RECT 83.66 3.795 83.68 5.02 ;
      RECT 83.645 3.795 83.66 5.053 ;
      RECT 83.615 3.795 83.645 5.075 ;
      RECT 83.595 3.795 83.615 5.089 ;
      RECT 83.575 3.795 83.595 4.605 ;
      RECT 83.59 4.672 83.595 5.094 ;
      RECT 83.585 4.702 83.59 5.096 ;
      RECT 83.58 4.715 83.585 5.099 ;
      RECT 83.575 4.725 83.58 5.103 ;
      RECT 83.57 3.795 83.575 4.523 ;
      RECT 83.57 4.735 83.575 5.105 ;
      RECT 83.565 3.795 83.57 4.5 ;
      RECT 83.555 4.757 83.57 5.105 ;
      RECT 83.55 3.795 83.565 4.445 ;
      RECT 83.545 4.782 83.555 5.105 ;
      RECT 83.545 3.795 83.55 4.39 ;
      RECT 83.535 3.795 83.545 4.338 ;
      RECT 83.54 4.795 83.545 5.106 ;
      RECT 83.535 4.807 83.54 5.107 ;
      RECT 83.53 3.795 83.535 4.298 ;
      RECT 83.53 4.82 83.535 5.108 ;
      RECT 83.515 4.835 83.53 5.109 ;
      RECT 83.52 3.795 83.525 4.26 ;
      RECT 83.515 3.795 83.52 4.225 ;
      RECT 83.51 3.795 83.515 4.2 ;
      RECT 83.505 4.862 83.515 5.111 ;
      RECT 83.5 3.795 83.51 4.158 ;
      RECT 83.5 4.88 83.505 5.112 ;
      RECT 83.495 3.795 83.5 4.118 ;
      RECT 83.495 4.887 83.5 5.113 ;
      RECT 83.49 3.795 83.495 4.09 ;
      RECT 83.485 4.905 83.495 5.114 ;
      RECT 83.48 3.795 83.49 4.07 ;
      RECT 83.475 4.925 83.485 5.116 ;
      RECT 83.465 4.942 83.475 5.117 ;
      RECT 83.43 4.965 83.465 5.12 ;
      RECT 83.375 4.983 83.43 5.126 ;
      RECT 83.289 4.991 83.375 5.135 ;
      RECT 83.203 5.002 83.289 5.146 ;
      RECT 83.117 5.012 83.203 5.157 ;
      RECT 83.031 5.022 83.117 5.169 ;
      RECT 82.945 5.032 83.031 5.18 ;
      RECT 82.925 5.038 82.945 5.186 ;
      RECT 82.845 5.04 82.925 5.19 ;
      RECT 82.84 5.039 82.845 5.195 ;
      RECT 82.832 5.038 82.84 5.195 ;
      RECT 82.746 5.034 82.832 5.193 ;
      RECT 82.66 5.026 82.746 5.19 ;
      RECT 82.574 5.017 82.66 5.186 ;
      RECT 82.488 5.009 82.574 5.183 ;
      RECT 82.402 5.001 82.488 5.179 ;
      RECT 82.316 4.992 82.402 5.176 ;
      RECT 82.23 4.984 82.316 5.172 ;
      RECT 82.175 4.977 82.22 5.17 ;
      RECT 82.09 4.97 82.175 5.168 ;
      RECT 82.016 4.962 82.09 5.164 ;
      RECT 81.93 4.954 82.016 5.161 ;
      RECT 81.927 4.95 81.93 5.159 ;
      RECT 81.841 4.946 81.927 5.158 ;
      RECT 81.755 4.938 81.841 5.155 ;
      RECT 81.67 4.933 81.755 5.152 ;
      RECT 81.584 4.93 81.67 5.149 ;
      RECT 81.498 4.928 81.584 5.146 ;
      RECT 81.412 4.925 81.498 5.143 ;
      RECT 81.326 4.922 81.412 5.14 ;
      RECT 81.24 4.919 81.326 5.137 ;
      RECT 81.164 4.917 81.24 5.134 ;
      RECT 81.078 4.914 81.164 5.131 ;
      RECT 80.992 4.911 81.078 5.129 ;
      RECT 80.906 4.909 80.992 5.126 ;
      RECT 80.82 4.906 80.906 5.123 ;
      RECT 80.76 4.897 80.82 5.121 ;
      RECT 83.27 4.515 83.345 4.775 ;
      RECT 83.25 4.495 83.255 4.775 ;
      RECT 82.57 4.28 82.675 4.575 ;
      RECT 77.015 4.255 77.085 4.515 ;
      RECT 82.91 4.13 82.915 4.501 ;
      RECT 82.9 4.185 82.905 4.501 ;
      RECT 83.205 3.355 83.265 3.615 ;
      RECT 83.26 4.51 83.27 4.775 ;
      RECT 83.255 4.5 83.26 4.775 ;
      RECT 83.175 4.447 83.25 4.775 ;
      RECT 83.2 3.355 83.205 3.635 ;
      RECT 83.19 3.355 83.2 3.655 ;
      RECT 83.175 3.355 83.19 3.685 ;
      RECT 83.16 3.355 83.175 3.728 ;
      RECT 83.155 4.39 83.175 4.775 ;
      RECT 83.145 3.355 83.16 3.765 ;
      RECT 83.14 4.37 83.155 4.775 ;
      RECT 83.14 3.355 83.145 3.788 ;
      RECT 83.13 3.355 83.14 3.813 ;
      RECT 83.1 4.337 83.14 4.775 ;
      RECT 83.105 3.355 83.13 3.863 ;
      RECT 83.1 3.355 83.105 3.918 ;
      RECT 83.095 3.355 83.1 3.96 ;
      RECT 83.085 4.3 83.1 4.775 ;
      RECT 83.09 3.355 83.095 4.003 ;
      RECT 83.085 3.355 83.09 4.068 ;
      RECT 83.08 3.355 83.085 4.09 ;
      RECT 83.08 4.288 83.085 4.64 ;
      RECT 83.075 3.355 83.08 4.158 ;
      RECT 83.075 4.28 83.08 4.623 ;
      RECT 83.07 3.355 83.075 4.203 ;
      RECT 83.065 4.262 83.075 4.6 ;
      RECT 83.065 3.355 83.07 4.24 ;
      RECT 83.055 3.355 83.065 4.58 ;
      RECT 83.05 3.355 83.055 4.563 ;
      RECT 83.045 3.355 83.05 4.548 ;
      RECT 83.04 3.355 83.045 4.533 ;
      RECT 83.02 3.355 83.04 4.523 ;
      RECT 83.015 3.355 83.02 4.513 ;
      RECT 83.005 3.355 83.015 4.509 ;
      RECT 83 3.632 83.005 4.508 ;
      RECT 82.995 3.655 83 4.507 ;
      RECT 82.99 3.685 82.995 4.506 ;
      RECT 82.985 3.712 82.99 4.505 ;
      RECT 82.98 3.74 82.985 4.505 ;
      RECT 82.975 3.767 82.98 4.505 ;
      RECT 82.97 3.787 82.975 4.505 ;
      RECT 82.965 3.815 82.97 4.505 ;
      RECT 82.955 3.857 82.965 4.505 ;
      RECT 82.945 3.902 82.955 4.504 ;
      RECT 82.94 3.955 82.945 4.503 ;
      RECT 82.935 3.987 82.94 4.502 ;
      RECT 82.93 4.007 82.935 4.501 ;
      RECT 82.925 4.045 82.93 4.501 ;
      RECT 82.92 4.067 82.925 4.501 ;
      RECT 82.915 4.092 82.92 4.501 ;
      RECT 82.905 4.157 82.91 4.501 ;
      RECT 82.89 4.217 82.9 4.501 ;
      RECT 82.875 4.227 82.89 4.501 ;
      RECT 82.855 4.237 82.875 4.501 ;
      RECT 82.825 4.242 82.855 4.498 ;
      RECT 82.765 4.252 82.825 4.495 ;
      RECT 82.745 4.261 82.765 4.5 ;
      RECT 82.72 4.267 82.745 4.513 ;
      RECT 82.7 4.272 82.72 4.528 ;
      RECT 82.675 4.277 82.7 4.575 ;
      RECT 82.546 4.279 82.57 4.575 ;
      RECT 82.46 4.274 82.546 4.575 ;
      RECT 82.42 4.271 82.46 4.575 ;
      RECT 82.37 4.273 82.42 4.555 ;
      RECT 82.34 4.277 82.37 4.555 ;
      RECT 82.261 4.287 82.34 4.555 ;
      RECT 82.175 4.302 82.261 4.556 ;
      RECT 82.125 4.312 82.175 4.557 ;
      RECT 82.117 4.315 82.125 4.557 ;
      RECT 82.031 4.317 82.117 4.558 ;
      RECT 81.945 4.321 82.031 4.558 ;
      RECT 81.859 4.325 81.945 4.559 ;
      RECT 81.773 4.328 81.859 4.56 ;
      RECT 81.687 4.332 81.773 4.56 ;
      RECT 81.601 4.336 81.687 4.561 ;
      RECT 81.515 4.339 81.601 4.562 ;
      RECT 81.429 4.343 81.515 4.562 ;
      RECT 81.343 4.347 81.429 4.563 ;
      RECT 81.257 4.351 81.343 4.564 ;
      RECT 81.171 4.354 81.257 4.564 ;
      RECT 81.085 4.358 81.171 4.565 ;
      RECT 81.055 4.36 81.085 4.565 ;
      RECT 80.969 4.363 81.055 4.566 ;
      RECT 80.883 4.367 80.969 4.567 ;
      RECT 80.797 4.371 80.883 4.568 ;
      RECT 80.711 4.374 80.797 4.568 ;
      RECT 80.625 4.378 80.711 4.569 ;
      RECT 80.59 4.383 80.625 4.57 ;
      RECT 80.535 4.393 80.59 4.577 ;
      RECT 80.51 4.405 80.535 4.587 ;
      RECT 80.475 4.418 80.51 4.595 ;
      RECT 80.435 4.435 80.475 4.618 ;
      RECT 80.415 4.448 80.435 4.645 ;
      RECT 80.385 4.46 80.415 4.673 ;
      RECT 80.38 4.468 80.385 4.693 ;
      RECT 80.375 4.471 80.38 4.703 ;
      RECT 80.325 4.483 80.375 4.737 ;
      RECT 80.315 4.498 80.325 4.77 ;
      RECT 80.305 4.504 80.315 4.783 ;
      RECT 80.295 4.511 80.305 4.795 ;
      RECT 80.27 4.524 80.295 4.813 ;
      RECT 80.255 4.539 80.27 4.835 ;
      RECT 80.245 4.547 80.255 4.851 ;
      RECT 80.23 4.556 80.245 4.866 ;
      RECT 80.22 4.566 80.23 4.88 ;
      RECT 80.201 4.579 80.22 4.897 ;
      RECT 80.115 4.624 80.201 4.962 ;
      RECT 80.1 4.669 80.115 5.02 ;
      RECT 80.095 4.678 80.1 5.033 ;
      RECT 80.085 4.685 80.095 5.038 ;
      RECT 80.08 4.69 80.085 5.042 ;
      RECT 80.06 4.7 80.08 5.049 ;
      RECT 80.035 4.72 80.06 5.063 ;
      RECT 80 4.745 80.035 5.083 ;
      RECT 79.985 4.768 80 5.098 ;
      RECT 79.975 4.778 79.985 5.103 ;
      RECT 79.965 4.786 79.975 5.11 ;
      RECT 79.955 4.795 79.965 5.116 ;
      RECT 79.935 4.807 79.955 5.118 ;
      RECT 79.925 4.82 79.935 5.12 ;
      RECT 79.9 4.835 79.925 5.123 ;
      RECT 79.88 4.852 79.9 5.127 ;
      RECT 79.84 4.88 79.88 5.133 ;
      RECT 79.775 4.927 79.84 5.142 ;
      RECT 79.76 4.96 79.775 5.15 ;
      RECT 79.755 4.967 79.76 5.152 ;
      RECT 79.705 4.992 79.755 5.157 ;
      RECT 79.69 5.016 79.705 5.164 ;
      RECT 79.64 5.021 79.69 5.165 ;
      RECT 79.554 5.025 79.64 5.165 ;
      RECT 79.468 5.025 79.554 5.165 ;
      RECT 79.382 5.025 79.468 5.166 ;
      RECT 79.296 5.025 79.382 5.166 ;
      RECT 79.21 5.025 79.296 5.166 ;
      RECT 79.144 5.025 79.21 5.166 ;
      RECT 79.058 5.025 79.144 5.167 ;
      RECT 78.972 5.025 79.058 5.167 ;
      RECT 78.886 5.026 78.972 5.168 ;
      RECT 78.8 5.026 78.886 5.168 ;
      RECT 78.714 5.026 78.8 5.168 ;
      RECT 78.628 5.026 78.714 5.169 ;
      RECT 78.542 5.026 78.628 5.169 ;
      RECT 78.456 5.027 78.542 5.17 ;
      RECT 78.37 5.027 78.456 5.17 ;
      RECT 78.35 5.027 78.37 5.17 ;
      RECT 78.264 5.027 78.35 5.17 ;
      RECT 78.178 5.027 78.264 5.17 ;
      RECT 78.092 5.028 78.178 5.17 ;
      RECT 78.006 5.028 78.092 5.17 ;
      RECT 77.92 5.028 78.006 5.17 ;
      RECT 77.834 5.029 77.92 5.17 ;
      RECT 77.748 5.029 77.834 5.17 ;
      RECT 77.662 5.029 77.748 5.17 ;
      RECT 77.576 5.029 77.662 5.17 ;
      RECT 77.49 5.03 77.576 5.17 ;
      RECT 77.44 5.027 77.49 5.17 ;
      RECT 77.43 5.025 77.44 5.169 ;
      RECT 77.426 5.025 77.43 5.168 ;
      RECT 77.34 5.02 77.426 5.163 ;
      RECT 77.318 5.013 77.34 5.157 ;
      RECT 77.232 5.004 77.318 5.151 ;
      RECT 77.146 4.991 77.232 5.142 ;
      RECT 77.06 4.977 77.146 5.132 ;
      RECT 77.015 4.967 77.06 5.125 ;
      RECT 76.995 4.255 77.015 4.533 ;
      RECT 76.995 4.96 77.015 5.121 ;
      RECT 76.965 4.255 76.995 4.555 ;
      RECT 76.955 4.927 76.995 5.118 ;
      RECT 76.95 4.255 76.965 4.575 ;
      RECT 76.95 4.892 76.955 5.116 ;
      RECT 76.945 4.255 76.95 4.7 ;
      RECT 76.945 4.852 76.95 5.116 ;
      RECT 76.935 4.255 76.945 5.116 ;
      RECT 76.86 4.255 76.935 5.11 ;
      RECT 76.83 4.255 76.86 5.1 ;
      RECT 76.825 4.255 76.83 5.092 ;
      RECT 76.82 4.297 76.825 5.085 ;
      RECT 76.81 4.366 76.82 5.076 ;
      RECT 76.805 4.436 76.81 5.028 ;
      RECT 76.8 4.5 76.805 4.925 ;
      RECT 76.795 4.535 76.8 4.88 ;
      RECT 76.793 4.572 76.795 4.772 ;
      RECT 76.79 4.58 76.793 4.765 ;
      RECT 76.785 4.645 76.79 4.708 ;
      RECT 80.86 3.735 81.14 4.015 ;
      RECT 80.85 3.735 81.14 3.878 ;
      RECT 80.805 3.6 81.065 3.86 ;
      RECT 80.805 3.715 81.12 3.86 ;
      RECT 80.805 3.685 81.115 3.86 ;
      RECT 80.805 3.672 81.105 3.86 ;
      RECT 80.805 3.662 81.1 3.86 ;
      RECT 76.78 3.645 77.04 3.905 ;
      RECT 80.55 3.195 80.81 3.455 ;
      RECT 80.54 3.22 80.81 3.415 ;
      RECT 80.535 3.22 80.54 3.414 ;
      RECT 80.465 3.215 80.535 3.406 ;
      RECT 80.38 3.202 80.465 3.389 ;
      RECT 80.376 3.194 80.38 3.379 ;
      RECT 80.29 3.187 80.376 3.369 ;
      RECT 80.281 3.179 80.29 3.359 ;
      RECT 80.195 3.172 80.281 3.347 ;
      RECT 80.175 3.163 80.195 3.333 ;
      RECT 80.12 3.158 80.175 3.325 ;
      RECT 80.11 3.152 80.12 3.319 ;
      RECT 80.09 3.15 80.11 3.315 ;
      RECT 80.082 3.149 80.09 3.311 ;
      RECT 79.996 3.141 80.082 3.3 ;
      RECT 79.91 3.127 79.996 3.28 ;
      RECT 79.85 3.115 79.91 3.265 ;
      RECT 79.84 3.11 79.85 3.26 ;
      RECT 79.79 3.11 79.84 3.262 ;
      RECT 79.743 3.112 79.79 3.266 ;
      RECT 79.657 3.119 79.743 3.271 ;
      RECT 79.571 3.127 79.657 3.277 ;
      RECT 79.485 3.136 79.571 3.283 ;
      RECT 79.426 3.142 79.485 3.288 ;
      RECT 79.34 3.147 79.426 3.294 ;
      RECT 79.265 3.152 79.34 3.3 ;
      RECT 79.226 3.154 79.265 3.305 ;
      RECT 79.14 3.151 79.226 3.31 ;
      RECT 79.055 3.149 79.14 3.317 ;
      RECT 79.023 3.148 79.055 3.32 ;
      RECT 78.937 3.147 79.023 3.321 ;
      RECT 78.851 3.146 78.937 3.322 ;
      RECT 78.765 3.145 78.851 3.322 ;
      RECT 78.679 3.144 78.765 3.323 ;
      RECT 78.593 3.143 78.679 3.324 ;
      RECT 78.507 3.142 78.593 3.325 ;
      RECT 78.421 3.141 78.507 3.325 ;
      RECT 78.335 3.14 78.421 3.326 ;
      RECT 78.285 3.14 78.335 3.327 ;
      RECT 78.271 3.141 78.285 3.327 ;
      RECT 78.185 3.148 78.271 3.328 ;
      RECT 78.111 3.159 78.185 3.329 ;
      RECT 78.025 3.168 78.111 3.33 ;
      RECT 77.99 3.175 78.025 3.345 ;
      RECT 77.965 3.178 77.99 3.375 ;
      RECT 77.94 3.187 77.965 3.404 ;
      RECT 77.93 3.198 77.94 3.424 ;
      RECT 77.92 3.206 77.93 3.438 ;
      RECT 77.915 3.212 77.92 3.448 ;
      RECT 77.89 3.229 77.915 3.465 ;
      RECT 77.875 3.251 77.89 3.493 ;
      RECT 77.845 3.277 77.875 3.523 ;
      RECT 77.825 3.306 77.845 3.553 ;
      RECT 77.82 3.321 77.825 3.57 ;
      RECT 77.8 3.336 77.82 3.585 ;
      RECT 77.79 3.354 77.8 3.603 ;
      RECT 77.78 3.365 77.79 3.618 ;
      RECT 77.73 3.397 77.78 3.644 ;
      RECT 77.725 3.427 77.73 3.664 ;
      RECT 77.715 3.44 77.725 3.67 ;
      RECT 77.706 3.45 77.715 3.678 ;
      RECT 77.695 3.461 77.706 3.686 ;
      RECT 77.69 3.471 77.695 3.692 ;
      RECT 77.675 3.492 77.69 3.699 ;
      RECT 77.66 3.522 77.675 3.707 ;
      RECT 77.625 3.552 77.66 3.713 ;
      RECT 77.6 3.57 77.625 3.72 ;
      RECT 77.55 3.578 77.6 3.729 ;
      RECT 77.525 3.583 77.55 3.738 ;
      RECT 77.47 3.589 77.525 3.748 ;
      RECT 77.465 3.594 77.47 3.756 ;
      RECT 77.451 3.597 77.465 3.758 ;
      RECT 77.365 3.609 77.451 3.77 ;
      RECT 77.355 3.621 77.365 3.783 ;
      RECT 77.27 3.634 77.355 3.795 ;
      RECT 77.226 3.651 77.27 3.809 ;
      RECT 77.14 3.668 77.226 3.825 ;
      RECT 77.11 3.682 77.14 3.839 ;
      RECT 77.1 3.687 77.11 3.844 ;
      RECT 77.04 3.69 77.1 3.853 ;
      RECT 79.93 3.96 80.19 4.22 ;
      RECT 79.93 3.96 80.21 4.073 ;
      RECT 79.93 3.96 80.235 4.04 ;
      RECT 79.93 3.96 80.24 4.02 ;
      RECT 79.98 3.735 80.26 4.015 ;
      RECT 79.535 4.47 79.795 4.73 ;
      RECT 79.525 4.327 79.72 4.668 ;
      RECT 79.52 4.435 79.735 4.66 ;
      RECT 79.515 4.485 79.795 4.65 ;
      RECT 79.505 4.562 79.795 4.635 ;
      RECT 79.525 4.41 79.735 4.668 ;
      RECT 79.535 4.285 79.72 4.73 ;
      RECT 79.535 4.18 79.7 4.73 ;
      RECT 79.545 4.167 79.7 4.73 ;
      RECT 79.545 4.125 79.69 4.73 ;
      RECT 79.55 4.05 79.69 4.73 ;
      RECT 79.58 3.7 79.69 4.73 ;
      RECT 79.585 3.43 79.71 4.053 ;
      RECT 79.555 4.005 79.71 4.053 ;
      RECT 79.57 3.807 79.69 4.73 ;
      RECT 79.56 3.917 79.71 4.053 ;
      RECT 79.585 3.43 79.725 3.91 ;
      RECT 79.585 3.43 79.745 3.785 ;
      RECT 79.55 3.43 79.81 3.69 ;
      RECT 79.02 3.735 79.3 4.015 ;
      RECT 79.005 3.735 79.3 3.995 ;
      RECT 77.06 4.6 77.32 4.86 ;
      RECT 78.845 4.455 79.105 4.715 ;
      RECT 78.825 4.475 79.105 4.69 ;
      RECT 78.782 4.475 78.825 4.689 ;
      RECT 78.696 4.476 78.782 4.686 ;
      RECT 78.61 4.477 78.696 4.682 ;
      RECT 78.535 4.479 78.61 4.679 ;
      RECT 78.512 4.48 78.535 4.677 ;
      RECT 78.426 4.481 78.512 4.675 ;
      RECT 78.34 4.482 78.426 4.672 ;
      RECT 78.316 4.483 78.34 4.67 ;
      RECT 78.23 4.485 78.316 4.667 ;
      RECT 78.145 4.487 78.23 4.668 ;
      RECT 78.088 4.488 78.145 4.674 ;
      RECT 78.002 4.49 78.088 4.684 ;
      RECT 77.916 4.493 78.002 4.697 ;
      RECT 77.83 4.495 77.916 4.709 ;
      RECT 77.816 4.496 77.83 4.716 ;
      RECT 77.73 4.497 77.816 4.724 ;
      RECT 77.69 4.499 77.73 4.733 ;
      RECT 77.681 4.5 77.69 4.736 ;
      RECT 77.595 4.508 77.681 4.742 ;
      RECT 77.575 4.517 77.595 4.75 ;
      RECT 77.49 4.532 77.575 4.758 ;
      RECT 77.43 4.555 77.49 4.769 ;
      RECT 77.42 4.567 77.43 4.774 ;
      RECT 77.38 4.577 77.42 4.778 ;
      RECT 77.325 4.594 77.38 4.786 ;
      RECT 77.32 4.604 77.325 4.79 ;
      RECT 78.386 3.735 78.445 4.132 ;
      RECT 78.3 3.735 78.505 4.123 ;
      RECT 78.295 3.765 78.505 4.118 ;
      RECT 78.261 3.765 78.505 4.116 ;
      RECT 78.175 3.765 78.505 4.11 ;
      RECT 78.13 3.765 78.525 4.088 ;
      RECT 78.13 3.765 78.545 4.043 ;
      RECT 78.09 3.765 78.545 4.033 ;
      RECT 78.3 3.735 78.58 4.015 ;
      RECT 78.035 3.735 78.295 3.995 ;
      RECT 77.22 3.215 77.48 3.475 ;
      RECT 77.3 3.175 77.58 3.455 ;
      RECT 71.665 8.505 71.985 8.83 ;
      RECT 71.695 7.98 71.865 8.83 ;
      RECT 71.695 7.98 71.87 8.33 ;
      RECT 71.695 7.98 72.67 8.155 ;
      RECT 72.495 3.26 72.67 8.155 ;
      RECT 72.44 3.26 72.79 3.61 ;
      RECT 72.465 8.94 72.79 9.265 ;
      RECT 71.35 9.03 72.79 9.2 ;
      RECT 71.35 3.69 71.51 9.2 ;
      RECT 71.665 3.66 71.985 3.98 ;
      RECT 71.35 3.69 71.985 3.86 ;
      RECT 60.075 4.295 60.355 4.575 ;
      RECT 60.045 4.295 60.355 4.56 ;
      RECT 60.04 4.295 60.355 4.558 ;
      RECT 60.035 2.625 60.205 4.552 ;
      RECT 60.03 4.262 60.3 4.545 ;
      RECT 60.025 4.295 60.355 4.538 ;
      RECT 59.995 4.265 60.3 4.525 ;
      RECT 59.995 4.292 60.32 4.525 ;
      RECT 59.995 4.282 60.315 4.525 ;
      RECT 59.995 4.267 60.31 4.525 ;
      RECT 60.035 4.257 60.3 4.552 ;
      RECT 60.035 4.252 60.29 4.552 ;
      RECT 60.035 4.251 60.275 4.552 ;
      RECT 70.005 2.635 70.355 2.985 ;
      RECT 70 2.635 70.355 2.89 ;
      RECT 60.035 2.625 70.245 2.795 ;
      RECT 69.68 4.145 70.05 4.515 ;
      RECT 69.765 3.53 69.935 4.515 ;
      RECT 65.785 3.75 66.02 4.01 ;
      RECT 68.93 3.53 69.095 3.79 ;
      RECT 68.835 3.52 68.85 3.79 ;
      RECT 68.93 3.53 69.935 3.71 ;
      RECT 67.435 3.09 67.475 3.23 ;
      RECT 68.85 3.525 68.93 3.79 ;
      RECT 68.795 3.52 68.835 3.756 ;
      RECT 68.781 3.52 68.795 3.756 ;
      RECT 68.695 3.525 68.781 3.758 ;
      RECT 68.65 3.532 68.695 3.76 ;
      RECT 68.62 3.532 68.65 3.762 ;
      RECT 68.595 3.527 68.62 3.764 ;
      RECT 68.565 3.523 68.595 3.773 ;
      RECT 68.555 3.52 68.565 3.785 ;
      RECT 68.55 3.52 68.555 3.793 ;
      RECT 68.545 3.52 68.55 3.798 ;
      RECT 68.535 3.519 68.545 3.808 ;
      RECT 68.53 3.518 68.535 3.818 ;
      RECT 68.515 3.517 68.53 3.823 ;
      RECT 68.487 3.514 68.515 3.85 ;
      RECT 68.401 3.506 68.487 3.85 ;
      RECT 68.315 3.495 68.401 3.85 ;
      RECT 68.275 3.48 68.315 3.85 ;
      RECT 68.235 3.454 68.275 3.85 ;
      RECT 68.23 3.436 68.235 3.662 ;
      RECT 68.22 3.432 68.23 3.652 ;
      RECT 68.205 3.422 68.22 3.639 ;
      RECT 68.185 3.406 68.205 3.624 ;
      RECT 68.17 3.391 68.185 3.609 ;
      RECT 68.16 3.38 68.17 3.599 ;
      RECT 68.135 3.364 68.16 3.588 ;
      RECT 68.13 3.351 68.135 3.578 ;
      RECT 68.125 3.347 68.13 3.573 ;
      RECT 68.07 3.333 68.125 3.551 ;
      RECT 68.031 3.314 68.07 3.515 ;
      RECT 67.945 3.288 68.031 3.468 ;
      RECT 67.941 3.27 67.945 3.434 ;
      RECT 67.855 3.251 67.941 3.412 ;
      RECT 67.85 3.233 67.855 3.39 ;
      RECT 67.845 3.231 67.85 3.388 ;
      RECT 67.835 3.23 67.845 3.383 ;
      RECT 67.775 3.217 67.835 3.369 ;
      RECT 67.73 3.195 67.775 3.348 ;
      RECT 67.67 3.172 67.73 3.327 ;
      RECT 67.606 3.147 67.67 3.302 ;
      RECT 67.52 3.117 67.606 3.271 ;
      RECT 67.505 3.097 67.52 3.25 ;
      RECT 67.475 3.092 67.505 3.241 ;
      RECT 67.422 3.09 67.435 3.23 ;
      RECT 67.336 3.09 67.422 3.232 ;
      RECT 67.25 3.09 67.336 3.234 ;
      RECT 67.23 3.09 67.25 3.238 ;
      RECT 67.185 3.092 67.23 3.249 ;
      RECT 67.145 3.102 67.185 3.265 ;
      RECT 67.141 3.111 67.145 3.273 ;
      RECT 67.055 3.131 67.141 3.289 ;
      RECT 67.045 3.15 67.055 3.307 ;
      RECT 67.04 3.152 67.045 3.31 ;
      RECT 67.03 3.156 67.04 3.313 ;
      RECT 67.01 3.161 67.03 3.323 ;
      RECT 66.98 3.171 67.01 3.343 ;
      RECT 66.975 3.178 66.98 3.357 ;
      RECT 66.965 3.182 66.975 3.364 ;
      RECT 66.95 3.19 66.965 3.375 ;
      RECT 66.94 3.2 66.95 3.386 ;
      RECT 66.93 3.207 66.94 3.394 ;
      RECT 66.905 3.22 66.93 3.409 ;
      RECT 66.841 3.256 66.905 3.448 ;
      RECT 66.755 3.319 66.841 3.512 ;
      RECT 66.72 3.37 66.755 3.565 ;
      RECT 66.715 3.387 66.72 3.582 ;
      RECT 66.7 3.396 66.715 3.589 ;
      RECT 66.68 3.411 66.7 3.603 ;
      RECT 66.675 3.422 66.68 3.613 ;
      RECT 66.655 3.435 66.675 3.623 ;
      RECT 66.65 3.445 66.655 3.633 ;
      RECT 66.635 3.45 66.65 3.642 ;
      RECT 66.625 3.46 66.635 3.653 ;
      RECT 66.595 3.477 66.625 3.67 ;
      RECT 66.585 3.495 66.595 3.688 ;
      RECT 66.57 3.506 66.585 3.699 ;
      RECT 66.53 3.53 66.57 3.715 ;
      RECT 66.495 3.564 66.53 3.732 ;
      RECT 66.465 3.587 66.495 3.744 ;
      RECT 66.45 3.597 66.465 3.753 ;
      RECT 66.41 3.607 66.45 3.764 ;
      RECT 66.39 3.618 66.41 3.776 ;
      RECT 66.385 3.622 66.39 3.783 ;
      RECT 66.37 3.626 66.385 3.788 ;
      RECT 66.36 3.631 66.37 3.793 ;
      RECT 66.355 3.634 66.36 3.796 ;
      RECT 66.325 3.64 66.355 3.803 ;
      RECT 66.29 3.65 66.325 3.817 ;
      RECT 66.23 3.665 66.29 3.837 ;
      RECT 66.175 3.685 66.23 3.861 ;
      RECT 66.146 3.7 66.175 3.879 ;
      RECT 66.06 3.72 66.146 3.904 ;
      RECT 66.055 3.735 66.06 3.924 ;
      RECT 66.045 3.738 66.055 3.925 ;
      RECT 66.02 3.745 66.045 4.01 ;
      RECT 68.715 4.238 68.995 4.575 ;
      RECT 68.715 4.248 69 4.533 ;
      RECT 68.715 4.257 69.005 4.43 ;
      RECT 68.715 4.272 69.01 4.298 ;
      RECT 68.715 4.1 68.975 4.575 ;
      RECT 59.015 8.94 59.365 9.29 ;
      RECT 67.84 8.895 68.19 9.245 ;
      RECT 59.015 8.97 68.19 9.17 ;
      RECT 66.435 4.98 66.445 5.17 ;
      RECT 64.695 4.855 64.975 5.135 ;
      RECT 67.74 3.795 67.745 4.28 ;
      RECT 67.635 3.795 67.695 4.055 ;
      RECT 67.96 4.765 67.965 4.84 ;
      RECT 67.95 4.632 67.96 4.875 ;
      RECT 67.94 4.467 67.95 4.896 ;
      RECT 67.935 4.337 67.94 4.912 ;
      RECT 67.925 4.227 67.935 4.928 ;
      RECT 67.92 4.126 67.925 4.945 ;
      RECT 67.915 4.108 67.92 4.955 ;
      RECT 67.91 4.09 67.915 4.965 ;
      RECT 67.9 4.065 67.91 4.98 ;
      RECT 67.895 4.045 67.9 4.995 ;
      RECT 67.875 3.795 67.895 5.02 ;
      RECT 67.86 3.795 67.875 5.053 ;
      RECT 67.83 3.795 67.86 5.075 ;
      RECT 67.81 3.795 67.83 5.089 ;
      RECT 67.79 3.795 67.81 4.605 ;
      RECT 67.805 4.672 67.81 5.094 ;
      RECT 67.8 4.702 67.805 5.096 ;
      RECT 67.795 4.715 67.8 5.099 ;
      RECT 67.79 4.725 67.795 5.103 ;
      RECT 67.785 3.795 67.79 4.523 ;
      RECT 67.785 4.735 67.79 5.105 ;
      RECT 67.78 3.795 67.785 4.5 ;
      RECT 67.77 4.757 67.785 5.105 ;
      RECT 67.765 3.795 67.78 4.445 ;
      RECT 67.76 4.782 67.77 5.105 ;
      RECT 67.76 3.795 67.765 4.39 ;
      RECT 67.75 3.795 67.76 4.338 ;
      RECT 67.755 4.795 67.76 5.106 ;
      RECT 67.75 4.807 67.755 5.107 ;
      RECT 67.745 3.795 67.75 4.298 ;
      RECT 67.745 4.82 67.75 5.108 ;
      RECT 67.73 4.835 67.745 5.109 ;
      RECT 67.735 3.795 67.74 4.26 ;
      RECT 67.73 3.795 67.735 4.225 ;
      RECT 67.725 3.795 67.73 4.2 ;
      RECT 67.72 4.862 67.73 5.111 ;
      RECT 67.715 3.795 67.725 4.158 ;
      RECT 67.715 4.88 67.72 5.112 ;
      RECT 67.71 3.795 67.715 4.118 ;
      RECT 67.71 4.887 67.715 5.113 ;
      RECT 67.705 3.795 67.71 4.09 ;
      RECT 67.7 4.905 67.71 5.114 ;
      RECT 67.695 3.795 67.705 4.07 ;
      RECT 67.69 4.925 67.7 5.116 ;
      RECT 67.68 4.942 67.69 5.117 ;
      RECT 67.645 4.965 67.68 5.12 ;
      RECT 67.59 4.983 67.645 5.126 ;
      RECT 67.504 4.991 67.59 5.135 ;
      RECT 67.418 5.002 67.504 5.146 ;
      RECT 67.332 5.012 67.418 5.157 ;
      RECT 67.246 5.022 67.332 5.169 ;
      RECT 67.16 5.032 67.246 5.18 ;
      RECT 67.14 5.038 67.16 5.186 ;
      RECT 67.06 5.04 67.14 5.19 ;
      RECT 67.055 5.039 67.06 5.195 ;
      RECT 67.047 5.038 67.055 5.195 ;
      RECT 66.961 5.034 67.047 5.193 ;
      RECT 66.875 5.026 66.961 5.19 ;
      RECT 66.789 5.017 66.875 5.186 ;
      RECT 66.703 5.009 66.789 5.183 ;
      RECT 66.617 5.001 66.703 5.179 ;
      RECT 66.531 4.992 66.617 5.176 ;
      RECT 66.445 4.984 66.531 5.172 ;
      RECT 66.39 4.977 66.435 5.17 ;
      RECT 66.305 4.97 66.39 5.168 ;
      RECT 66.231 4.962 66.305 5.164 ;
      RECT 66.145 4.954 66.231 5.161 ;
      RECT 66.142 4.95 66.145 5.159 ;
      RECT 66.056 4.946 66.142 5.158 ;
      RECT 65.97 4.938 66.056 5.155 ;
      RECT 65.885 4.933 65.97 5.152 ;
      RECT 65.799 4.93 65.885 5.149 ;
      RECT 65.713 4.928 65.799 5.146 ;
      RECT 65.627 4.925 65.713 5.143 ;
      RECT 65.541 4.922 65.627 5.14 ;
      RECT 65.455 4.919 65.541 5.137 ;
      RECT 65.379 4.917 65.455 5.134 ;
      RECT 65.293 4.914 65.379 5.131 ;
      RECT 65.207 4.911 65.293 5.129 ;
      RECT 65.121 4.909 65.207 5.126 ;
      RECT 65.035 4.906 65.121 5.123 ;
      RECT 64.975 4.897 65.035 5.121 ;
      RECT 67.485 4.515 67.56 4.775 ;
      RECT 67.465 4.495 67.47 4.775 ;
      RECT 66.785 4.28 66.89 4.575 ;
      RECT 61.23 4.255 61.3 4.515 ;
      RECT 67.125 4.13 67.13 4.501 ;
      RECT 67.115 4.185 67.12 4.501 ;
      RECT 67.42 3.355 67.48 3.615 ;
      RECT 67.475 4.51 67.485 4.775 ;
      RECT 67.47 4.5 67.475 4.775 ;
      RECT 67.39 4.447 67.465 4.775 ;
      RECT 67.415 3.355 67.42 3.635 ;
      RECT 67.405 3.355 67.415 3.655 ;
      RECT 67.39 3.355 67.405 3.685 ;
      RECT 67.375 3.355 67.39 3.728 ;
      RECT 67.37 4.39 67.39 4.775 ;
      RECT 67.36 3.355 67.375 3.765 ;
      RECT 67.355 4.37 67.37 4.775 ;
      RECT 67.355 3.355 67.36 3.788 ;
      RECT 67.345 3.355 67.355 3.813 ;
      RECT 67.315 4.337 67.355 4.775 ;
      RECT 67.32 3.355 67.345 3.863 ;
      RECT 67.315 3.355 67.32 3.918 ;
      RECT 67.31 3.355 67.315 3.96 ;
      RECT 67.3 4.3 67.315 4.775 ;
      RECT 67.305 3.355 67.31 4.003 ;
      RECT 67.3 3.355 67.305 4.068 ;
      RECT 67.295 3.355 67.3 4.09 ;
      RECT 67.295 4.288 67.3 4.64 ;
      RECT 67.29 3.355 67.295 4.158 ;
      RECT 67.29 4.28 67.295 4.623 ;
      RECT 67.285 3.355 67.29 4.203 ;
      RECT 67.28 4.262 67.29 4.6 ;
      RECT 67.28 3.355 67.285 4.24 ;
      RECT 67.27 3.355 67.28 4.58 ;
      RECT 67.265 3.355 67.27 4.563 ;
      RECT 67.26 3.355 67.265 4.548 ;
      RECT 67.255 3.355 67.26 4.533 ;
      RECT 67.235 3.355 67.255 4.523 ;
      RECT 67.23 3.355 67.235 4.513 ;
      RECT 67.22 3.355 67.23 4.509 ;
      RECT 67.215 3.632 67.22 4.508 ;
      RECT 67.21 3.655 67.215 4.507 ;
      RECT 67.205 3.685 67.21 4.506 ;
      RECT 67.2 3.712 67.205 4.505 ;
      RECT 67.195 3.74 67.2 4.505 ;
      RECT 67.19 3.767 67.195 4.505 ;
      RECT 67.185 3.787 67.19 4.505 ;
      RECT 67.18 3.815 67.185 4.505 ;
      RECT 67.17 3.857 67.18 4.505 ;
      RECT 67.16 3.902 67.17 4.504 ;
      RECT 67.155 3.955 67.16 4.503 ;
      RECT 67.15 3.987 67.155 4.502 ;
      RECT 67.145 4.007 67.15 4.501 ;
      RECT 67.14 4.045 67.145 4.501 ;
      RECT 67.135 4.067 67.14 4.501 ;
      RECT 67.13 4.092 67.135 4.501 ;
      RECT 67.12 4.157 67.125 4.501 ;
      RECT 67.105 4.217 67.115 4.501 ;
      RECT 67.09 4.227 67.105 4.501 ;
      RECT 67.07 4.237 67.09 4.501 ;
      RECT 67.04 4.242 67.07 4.498 ;
      RECT 66.98 4.252 67.04 4.495 ;
      RECT 66.96 4.261 66.98 4.5 ;
      RECT 66.935 4.267 66.96 4.513 ;
      RECT 66.915 4.272 66.935 4.528 ;
      RECT 66.89 4.277 66.915 4.575 ;
      RECT 66.761 4.279 66.785 4.575 ;
      RECT 66.675 4.274 66.761 4.575 ;
      RECT 66.635 4.271 66.675 4.575 ;
      RECT 66.585 4.273 66.635 4.555 ;
      RECT 66.555 4.277 66.585 4.555 ;
      RECT 66.476 4.287 66.555 4.555 ;
      RECT 66.39 4.302 66.476 4.556 ;
      RECT 66.34 4.312 66.39 4.557 ;
      RECT 66.332 4.315 66.34 4.557 ;
      RECT 66.246 4.317 66.332 4.558 ;
      RECT 66.16 4.321 66.246 4.558 ;
      RECT 66.074 4.325 66.16 4.559 ;
      RECT 65.988 4.328 66.074 4.56 ;
      RECT 65.902 4.332 65.988 4.56 ;
      RECT 65.816 4.336 65.902 4.561 ;
      RECT 65.73 4.339 65.816 4.562 ;
      RECT 65.644 4.343 65.73 4.562 ;
      RECT 65.558 4.347 65.644 4.563 ;
      RECT 65.472 4.351 65.558 4.564 ;
      RECT 65.386 4.354 65.472 4.564 ;
      RECT 65.3 4.358 65.386 4.565 ;
      RECT 65.27 4.36 65.3 4.565 ;
      RECT 65.184 4.363 65.27 4.566 ;
      RECT 65.098 4.367 65.184 4.567 ;
      RECT 65.012 4.371 65.098 4.568 ;
      RECT 64.926 4.374 65.012 4.568 ;
      RECT 64.84 4.378 64.926 4.569 ;
      RECT 64.805 4.383 64.84 4.57 ;
      RECT 64.75 4.393 64.805 4.577 ;
      RECT 64.725 4.405 64.75 4.587 ;
      RECT 64.69 4.418 64.725 4.595 ;
      RECT 64.65 4.435 64.69 4.618 ;
      RECT 64.63 4.448 64.65 4.645 ;
      RECT 64.6 4.46 64.63 4.673 ;
      RECT 64.595 4.468 64.6 4.693 ;
      RECT 64.59 4.471 64.595 4.703 ;
      RECT 64.54 4.483 64.59 4.737 ;
      RECT 64.53 4.498 64.54 4.77 ;
      RECT 64.52 4.504 64.53 4.783 ;
      RECT 64.51 4.511 64.52 4.795 ;
      RECT 64.485 4.524 64.51 4.813 ;
      RECT 64.47 4.539 64.485 4.835 ;
      RECT 64.46 4.547 64.47 4.851 ;
      RECT 64.445 4.556 64.46 4.866 ;
      RECT 64.435 4.566 64.445 4.88 ;
      RECT 64.416 4.579 64.435 4.897 ;
      RECT 64.33 4.624 64.416 4.962 ;
      RECT 64.315 4.669 64.33 5.02 ;
      RECT 64.31 4.678 64.315 5.033 ;
      RECT 64.3 4.685 64.31 5.038 ;
      RECT 64.295 4.69 64.3 5.042 ;
      RECT 64.275 4.7 64.295 5.049 ;
      RECT 64.25 4.72 64.275 5.063 ;
      RECT 64.215 4.745 64.25 5.083 ;
      RECT 64.2 4.768 64.215 5.098 ;
      RECT 64.19 4.778 64.2 5.103 ;
      RECT 64.18 4.786 64.19 5.11 ;
      RECT 64.17 4.795 64.18 5.116 ;
      RECT 64.15 4.807 64.17 5.118 ;
      RECT 64.14 4.82 64.15 5.12 ;
      RECT 64.115 4.835 64.14 5.123 ;
      RECT 64.095 4.852 64.115 5.127 ;
      RECT 64.055 4.88 64.095 5.133 ;
      RECT 63.99 4.927 64.055 5.142 ;
      RECT 63.975 4.96 63.99 5.15 ;
      RECT 63.97 4.967 63.975 5.152 ;
      RECT 63.92 4.992 63.97 5.157 ;
      RECT 63.905 5.016 63.92 5.164 ;
      RECT 63.855 5.021 63.905 5.165 ;
      RECT 63.769 5.025 63.855 5.165 ;
      RECT 63.683 5.025 63.769 5.165 ;
      RECT 63.597 5.025 63.683 5.166 ;
      RECT 63.511 5.025 63.597 5.166 ;
      RECT 63.425 5.025 63.511 5.166 ;
      RECT 63.359 5.025 63.425 5.166 ;
      RECT 63.273 5.025 63.359 5.167 ;
      RECT 63.187 5.025 63.273 5.167 ;
      RECT 63.101 5.026 63.187 5.168 ;
      RECT 63.015 5.026 63.101 5.168 ;
      RECT 62.929 5.026 63.015 5.168 ;
      RECT 62.843 5.026 62.929 5.169 ;
      RECT 62.757 5.026 62.843 5.169 ;
      RECT 62.671 5.027 62.757 5.17 ;
      RECT 62.585 5.027 62.671 5.17 ;
      RECT 62.565 5.027 62.585 5.17 ;
      RECT 62.479 5.027 62.565 5.17 ;
      RECT 62.393 5.027 62.479 5.17 ;
      RECT 62.307 5.028 62.393 5.17 ;
      RECT 62.221 5.028 62.307 5.17 ;
      RECT 62.135 5.028 62.221 5.17 ;
      RECT 62.049 5.029 62.135 5.17 ;
      RECT 61.963 5.029 62.049 5.17 ;
      RECT 61.877 5.029 61.963 5.17 ;
      RECT 61.791 5.029 61.877 5.17 ;
      RECT 61.705 5.03 61.791 5.17 ;
      RECT 61.655 5.027 61.705 5.17 ;
      RECT 61.645 5.025 61.655 5.169 ;
      RECT 61.641 5.025 61.645 5.168 ;
      RECT 61.555 5.02 61.641 5.163 ;
      RECT 61.533 5.013 61.555 5.157 ;
      RECT 61.447 5.004 61.533 5.151 ;
      RECT 61.361 4.991 61.447 5.142 ;
      RECT 61.275 4.977 61.361 5.132 ;
      RECT 61.23 4.967 61.275 5.125 ;
      RECT 61.21 4.255 61.23 4.533 ;
      RECT 61.21 4.96 61.23 5.121 ;
      RECT 61.18 4.255 61.21 4.555 ;
      RECT 61.17 4.927 61.21 5.118 ;
      RECT 61.165 4.255 61.18 4.575 ;
      RECT 61.165 4.892 61.17 5.116 ;
      RECT 61.16 4.255 61.165 4.7 ;
      RECT 61.16 4.852 61.165 5.116 ;
      RECT 61.15 4.255 61.16 5.116 ;
      RECT 61.075 4.255 61.15 5.11 ;
      RECT 61.045 4.255 61.075 5.1 ;
      RECT 61.04 4.255 61.045 5.092 ;
      RECT 61.035 4.297 61.04 5.085 ;
      RECT 61.025 4.366 61.035 5.076 ;
      RECT 61.02 4.436 61.025 5.028 ;
      RECT 61.015 4.5 61.02 4.925 ;
      RECT 61.01 4.535 61.015 4.88 ;
      RECT 61.008 4.572 61.01 4.772 ;
      RECT 61.005 4.58 61.008 4.765 ;
      RECT 61 4.645 61.005 4.708 ;
      RECT 65.075 3.735 65.355 4.015 ;
      RECT 65.065 3.735 65.355 3.878 ;
      RECT 65.02 3.6 65.28 3.86 ;
      RECT 65.02 3.715 65.335 3.86 ;
      RECT 65.02 3.685 65.33 3.86 ;
      RECT 65.02 3.672 65.32 3.86 ;
      RECT 65.02 3.662 65.315 3.86 ;
      RECT 60.995 3.645 61.255 3.905 ;
      RECT 64.765 3.195 65.025 3.455 ;
      RECT 64.755 3.22 65.025 3.415 ;
      RECT 64.75 3.22 64.755 3.414 ;
      RECT 64.68 3.215 64.75 3.406 ;
      RECT 64.595 3.202 64.68 3.389 ;
      RECT 64.591 3.194 64.595 3.379 ;
      RECT 64.505 3.187 64.591 3.369 ;
      RECT 64.496 3.179 64.505 3.359 ;
      RECT 64.41 3.172 64.496 3.347 ;
      RECT 64.39 3.163 64.41 3.333 ;
      RECT 64.335 3.158 64.39 3.325 ;
      RECT 64.325 3.152 64.335 3.319 ;
      RECT 64.305 3.15 64.325 3.315 ;
      RECT 64.297 3.149 64.305 3.311 ;
      RECT 64.211 3.141 64.297 3.3 ;
      RECT 64.125 3.127 64.211 3.28 ;
      RECT 64.065 3.115 64.125 3.265 ;
      RECT 64.055 3.11 64.065 3.26 ;
      RECT 64.005 3.11 64.055 3.262 ;
      RECT 63.958 3.112 64.005 3.266 ;
      RECT 63.872 3.119 63.958 3.271 ;
      RECT 63.786 3.127 63.872 3.277 ;
      RECT 63.7 3.136 63.786 3.283 ;
      RECT 63.641 3.142 63.7 3.288 ;
      RECT 63.555 3.147 63.641 3.294 ;
      RECT 63.48 3.152 63.555 3.3 ;
      RECT 63.441 3.154 63.48 3.305 ;
      RECT 63.355 3.151 63.441 3.31 ;
      RECT 63.27 3.149 63.355 3.317 ;
      RECT 63.238 3.148 63.27 3.32 ;
      RECT 63.152 3.147 63.238 3.321 ;
      RECT 63.066 3.146 63.152 3.322 ;
      RECT 62.98 3.145 63.066 3.322 ;
      RECT 62.894 3.144 62.98 3.323 ;
      RECT 62.808 3.143 62.894 3.324 ;
      RECT 62.722 3.142 62.808 3.325 ;
      RECT 62.636 3.141 62.722 3.325 ;
      RECT 62.55 3.14 62.636 3.326 ;
      RECT 62.5 3.14 62.55 3.327 ;
      RECT 62.486 3.141 62.5 3.327 ;
      RECT 62.4 3.148 62.486 3.328 ;
      RECT 62.326 3.159 62.4 3.329 ;
      RECT 62.24 3.168 62.326 3.33 ;
      RECT 62.205 3.175 62.24 3.345 ;
      RECT 62.18 3.178 62.205 3.375 ;
      RECT 62.155 3.187 62.18 3.404 ;
      RECT 62.145 3.198 62.155 3.424 ;
      RECT 62.135 3.206 62.145 3.438 ;
      RECT 62.13 3.212 62.135 3.448 ;
      RECT 62.105 3.229 62.13 3.465 ;
      RECT 62.09 3.251 62.105 3.493 ;
      RECT 62.06 3.277 62.09 3.523 ;
      RECT 62.04 3.306 62.06 3.553 ;
      RECT 62.035 3.321 62.04 3.57 ;
      RECT 62.015 3.336 62.035 3.585 ;
      RECT 62.005 3.354 62.015 3.603 ;
      RECT 61.995 3.365 62.005 3.618 ;
      RECT 61.945 3.397 61.995 3.644 ;
      RECT 61.94 3.427 61.945 3.664 ;
      RECT 61.93 3.44 61.94 3.67 ;
      RECT 61.921 3.45 61.93 3.678 ;
      RECT 61.91 3.461 61.921 3.686 ;
      RECT 61.905 3.471 61.91 3.692 ;
      RECT 61.89 3.492 61.905 3.699 ;
      RECT 61.875 3.522 61.89 3.707 ;
      RECT 61.84 3.552 61.875 3.713 ;
      RECT 61.815 3.57 61.84 3.72 ;
      RECT 61.765 3.578 61.815 3.729 ;
      RECT 61.74 3.583 61.765 3.738 ;
      RECT 61.685 3.589 61.74 3.748 ;
      RECT 61.68 3.594 61.685 3.756 ;
      RECT 61.666 3.597 61.68 3.758 ;
      RECT 61.58 3.609 61.666 3.77 ;
      RECT 61.57 3.621 61.58 3.783 ;
      RECT 61.485 3.634 61.57 3.795 ;
      RECT 61.441 3.651 61.485 3.809 ;
      RECT 61.355 3.668 61.441 3.825 ;
      RECT 61.325 3.682 61.355 3.839 ;
      RECT 61.315 3.687 61.325 3.844 ;
      RECT 61.255 3.69 61.315 3.853 ;
      RECT 64.145 3.96 64.405 4.22 ;
      RECT 64.145 3.96 64.425 4.073 ;
      RECT 64.145 3.96 64.45 4.04 ;
      RECT 64.145 3.96 64.455 4.02 ;
      RECT 64.195 3.735 64.475 4.015 ;
      RECT 63.75 4.47 64.01 4.73 ;
      RECT 63.74 4.327 63.935 4.668 ;
      RECT 63.735 4.435 63.95 4.66 ;
      RECT 63.73 4.485 64.01 4.65 ;
      RECT 63.72 4.562 64.01 4.635 ;
      RECT 63.74 4.41 63.95 4.668 ;
      RECT 63.75 4.285 63.935 4.73 ;
      RECT 63.75 4.18 63.915 4.73 ;
      RECT 63.76 4.167 63.915 4.73 ;
      RECT 63.76 4.125 63.905 4.73 ;
      RECT 63.765 4.05 63.905 4.73 ;
      RECT 63.795 3.7 63.905 4.73 ;
      RECT 63.8 3.43 63.925 4.053 ;
      RECT 63.77 4.005 63.925 4.053 ;
      RECT 63.785 3.807 63.905 4.73 ;
      RECT 63.775 3.917 63.925 4.053 ;
      RECT 63.8 3.43 63.94 3.91 ;
      RECT 63.8 3.43 63.96 3.785 ;
      RECT 63.765 3.43 64.025 3.69 ;
      RECT 63.235 3.735 63.515 4.015 ;
      RECT 63.22 3.735 63.515 3.995 ;
      RECT 61.275 4.6 61.535 4.86 ;
      RECT 63.06 4.455 63.32 4.715 ;
      RECT 63.04 4.475 63.32 4.69 ;
      RECT 62.997 4.475 63.04 4.689 ;
      RECT 62.911 4.476 62.997 4.686 ;
      RECT 62.825 4.477 62.911 4.682 ;
      RECT 62.75 4.479 62.825 4.679 ;
      RECT 62.727 4.48 62.75 4.677 ;
      RECT 62.641 4.481 62.727 4.675 ;
      RECT 62.555 4.482 62.641 4.672 ;
      RECT 62.531 4.483 62.555 4.67 ;
      RECT 62.445 4.485 62.531 4.667 ;
      RECT 62.36 4.487 62.445 4.668 ;
      RECT 62.303 4.488 62.36 4.674 ;
      RECT 62.217 4.49 62.303 4.684 ;
      RECT 62.131 4.493 62.217 4.697 ;
      RECT 62.045 4.495 62.131 4.709 ;
      RECT 62.031 4.496 62.045 4.716 ;
      RECT 61.945 4.497 62.031 4.724 ;
      RECT 61.905 4.499 61.945 4.733 ;
      RECT 61.896 4.5 61.905 4.736 ;
      RECT 61.81 4.508 61.896 4.742 ;
      RECT 61.79 4.517 61.81 4.75 ;
      RECT 61.705 4.532 61.79 4.758 ;
      RECT 61.645 4.555 61.705 4.769 ;
      RECT 61.635 4.567 61.645 4.774 ;
      RECT 61.595 4.577 61.635 4.778 ;
      RECT 61.54 4.594 61.595 4.786 ;
      RECT 61.535 4.604 61.54 4.79 ;
      RECT 62.601 3.735 62.66 4.132 ;
      RECT 62.515 3.735 62.72 4.123 ;
      RECT 62.51 3.765 62.72 4.118 ;
      RECT 62.476 3.765 62.72 4.116 ;
      RECT 62.39 3.765 62.72 4.11 ;
      RECT 62.345 3.765 62.74 4.088 ;
      RECT 62.345 3.765 62.76 4.043 ;
      RECT 62.305 3.765 62.76 4.033 ;
      RECT 62.515 3.735 62.795 4.015 ;
      RECT 62.25 3.735 62.51 3.995 ;
      RECT 61.435 3.215 61.695 3.475 ;
      RECT 61.515 3.175 61.795 3.455 ;
      RECT 55.88 8.505 56.2 8.83 ;
      RECT 55.91 7.98 56.08 8.83 ;
      RECT 55.91 7.98 56.085 8.33 ;
      RECT 55.91 7.98 56.885 8.155 ;
      RECT 56.71 3.26 56.885 8.155 ;
      RECT 56.655 3.26 57.005 3.61 ;
      RECT 56.68 8.94 57.005 9.265 ;
      RECT 55.565 9.03 57.005 9.2 ;
      RECT 55.565 3.69 55.725 9.2 ;
      RECT 55.88 3.66 56.2 3.98 ;
      RECT 55.565 3.69 56.2 3.86 ;
      RECT 44.29 4.295 44.57 4.575 ;
      RECT 44.26 4.295 44.57 4.56 ;
      RECT 44.255 4.295 44.57 4.558 ;
      RECT 44.25 2.625 44.42 4.552 ;
      RECT 44.245 4.262 44.515 4.545 ;
      RECT 44.24 4.295 44.57 4.538 ;
      RECT 44.21 4.265 44.515 4.525 ;
      RECT 44.21 4.292 44.535 4.525 ;
      RECT 44.21 4.282 44.53 4.525 ;
      RECT 44.21 4.267 44.525 4.525 ;
      RECT 44.25 4.257 44.515 4.552 ;
      RECT 44.25 4.252 44.505 4.552 ;
      RECT 44.25 4.251 44.49 4.552 ;
      RECT 54.22 2.635 54.57 2.985 ;
      RECT 54.215 2.635 54.57 2.89 ;
      RECT 44.25 2.625 54.46 2.795 ;
      RECT 53.895 4.145 54.265 4.515 ;
      RECT 53.98 3.53 54.15 4.515 ;
      RECT 50 3.75 50.235 4.01 ;
      RECT 53.145 3.53 53.31 3.79 ;
      RECT 53.05 3.52 53.065 3.79 ;
      RECT 53.145 3.53 54.15 3.71 ;
      RECT 51.65 3.09 51.69 3.23 ;
      RECT 53.065 3.525 53.145 3.79 ;
      RECT 53.01 3.52 53.05 3.756 ;
      RECT 52.996 3.52 53.01 3.756 ;
      RECT 52.91 3.525 52.996 3.758 ;
      RECT 52.865 3.532 52.91 3.76 ;
      RECT 52.835 3.532 52.865 3.762 ;
      RECT 52.81 3.527 52.835 3.764 ;
      RECT 52.78 3.523 52.81 3.773 ;
      RECT 52.77 3.52 52.78 3.785 ;
      RECT 52.765 3.52 52.77 3.793 ;
      RECT 52.76 3.52 52.765 3.798 ;
      RECT 52.75 3.519 52.76 3.808 ;
      RECT 52.745 3.518 52.75 3.818 ;
      RECT 52.73 3.517 52.745 3.823 ;
      RECT 52.702 3.514 52.73 3.85 ;
      RECT 52.616 3.506 52.702 3.85 ;
      RECT 52.53 3.495 52.616 3.85 ;
      RECT 52.49 3.48 52.53 3.85 ;
      RECT 52.45 3.454 52.49 3.85 ;
      RECT 52.445 3.436 52.45 3.662 ;
      RECT 52.435 3.432 52.445 3.652 ;
      RECT 52.42 3.422 52.435 3.639 ;
      RECT 52.4 3.406 52.42 3.624 ;
      RECT 52.385 3.391 52.4 3.609 ;
      RECT 52.375 3.38 52.385 3.599 ;
      RECT 52.35 3.364 52.375 3.588 ;
      RECT 52.345 3.351 52.35 3.578 ;
      RECT 52.34 3.347 52.345 3.573 ;
      RECT 52.285 3.333 52.34 3.551 ;
      RECT 52.246 3.314 52.285 3.515 ;
      RECT 52.16 3.288 52.246 3.468 ;
      RECT 52.156 3.27 52.16 3.434 ;
      RECT 52.07 3.251 52.156 3.412 ;
      RECT 52.065 3.233 52.07 3.39 ;
      RECT 52.06 3.231 52.065 3.388 ;
      RECT 52.05 3.23 52.06 3.383 ;
      RECT 51.99 3.217 52.05 3.369 ;
      RECT 51.945 3.195 51.99 3.348 ;
      RECT 51.885 3.172 51.945 3.327 ;
      RECT 51.821 3.147 51.885 3.302 ;
      RECT 51.735 3.117 51.821 3.271 ;
      RECT 51.72 3.097 51.735 3.25 ;
      RECT 51.69 3.092 51.72 3.241 ;
      RECT 51.637 3.09 51.65 3.23 ;
      RECT 51.551 3.09 51.637 3.232 ;
      RECT 51.465 3.09 51.551 3.234 ;
      RECT 51.445 3.09 51.465 3.238 ;
      RECT 51.4 3.092 51.445 3.249 ;
      RECT 51.36 3.102 51.4 3.265 ;
      RECT 51.356 3.111 51.36 3.273 ;
      RECT 51.27 3.131 51.356 3.289 ;
      RECT 51.26 3.15 51.27 3.307 ;
      RECT 51.255 3.152 51.26 3.31 ;
      RECT 51.245 3.156 51.255 3.313 ;
      RECT 51.225 3.161 51.245 3.323 ;
      RECT 51.195 3.171 51.225 3.343 ;
      RECT 51.19 3.178 51.195 3.357 ;
      RECT 51.18 3.182 51.19 3.364 ;
      RECT 51.165 3.19 51.18 3.375 ;
      RECT 51.155 3.2 51.165 3.386 ;
      RECT 51.145 3.207 51.155 3.394 ;
      RECT 51.12 3.22 51.145 3.409 ;
      RECT 51.056 3.256 51.12 3.448 ;
      RECT 50.97 3.319 51.056 3.512 ;
      RECT 50.935 3.37 50.97 3.565 ;
      RECT 50.93 3.387 50.935 3.582 ;
      RECT 50.915 3.396 50.93 3.589 ;
      RECT 50.895 3.411 50.915 3.603 ;
      RECT 50.89 3.422 50.895 3.613 ;
      RECT 50.87 3.435 50.89 3.623 ;
      RECT 50.865 3.445 50.87 3.633 ;
      RECT 50.85 3.45 50.865 3.642 ;
      RECT 50.84 3.46 50.85 3.653 ;
      RECT 50.81 3.477 50.84 3.67 ;
      RECT 50.8 3.495 50.81 3.688 ;
      RECT 50.785 3.506 50.8 3.699 ;
      RECT 50.745 3.53 50.785 3.715 ;
      RECT 50.71 3.564 50.745 3.732 ;
      RECT 50.68 3.587 50.71 3.744 ;
      RECT 50.665 3.597 50.68 3.753 ;
      RECT 50.625 3.607 50.665 3.764 ;
      RECT 50.605 3.618 50.625 3.776 ;
      RECT 50.6 3.622 50.605 3.783 ;
      RECT 50.585 3.626 50.6 3.788 ;
      RECT 50.575 3.631 50.585 3.793 ;
      RECT 50.57 3.634 50.575 3.796 ;
      RECT 50.54 3.64 50.57 3.803 ;
      RECT 50.505 3.65 50.54 3.817 ;
      RECT 50.445 3.665 50.505 3.837 ;
      RECT 50.39 3.685 50.445 3.861 ;
      RECT 50.361 3.7 50.39 3.879 ;
      RECT 50.275 3.72 50.361 3.904 ;
      RECT 50.27 3.735 50.275 3.924 ;
      RECT 50.26 3.738 50.27 3.925 ;
      RECT 50.235 3.745 50.26 4.01 ;
      RECT 52.93 4.238 53.21 4.575 ;
      RECT 52.93 4.248 53.215 4.533 ;
      RECT 52.93 4.257 53.22 4.43 ;
      RECT 52.93 4.272 53.225 4.298 ;
      RECT 52.93 4.1 53.19 4.575 ;
      RECT 43.285 8.945 43.635 9.295 ;
      RECT 52.11 8.9 52.46 9.25 ;
      RECT 43.285 8.975 52.46 9.175 ;
      RECT 50.65 4.98 50.66 5.17 ;
      RECT 48.91 4.855 49.19 5.135 ;
      RECT 51.955 3.795 51.96 4.28 ;
      RECT 51.85 3.795 51.91 4.055 ;
      RECT 52.175 4.765 52.18 4.84 ;
      RECT 52.165 4.632 52.175 4.875 ;
      RECT 52.155 4.467 52.165 4.896 ;
      RECT 52.15 4.337 52.155 4.912 ;
      RECT 52.14 4.227 52.15 4.928 ;
      RECT 52.135 4.126 52.14 4.945 ;
      RECT 52.13 4.108 52.135 4.955 ;
      RECT 52.125 4.09 52.13 4.965 ;
      RECT 52.115 4.065 52.125 4.98 ;
      RECT 52.11 4.045 52.115 4.995 ;
      RECT 52.09 3.795 52.11 5.02 ;
      RECT 52.075 3.795 52.09 5.053 ;
      RECT 52.045 3.795 52.075 5.075 ;
      RECT 52.025 3.795 52.045 5.089 ;
      RECT 52.005 3.795 52.025 4.605 ;
      RECT 52.02 4.672 52.025 5.094 ;
      RECT 52.015 4.702 52.02 5.096 ;
      RECT 52.01 4.715 52.015 5.099 ;
      RECT 52.005 4.725 52.01 5.103 ;
      RECT 52 3.795 52.005 4.523 ;
      RECT 52 4.735 52.005 5.105 ;
      RECT 51.995 3.795 52 4.5 ;
      RECT 51.985 4.757 52 5.105 ;
      RECT 51.98 3.795 51.995 4.445 ;
      RECT 51.975 4.782 51.985 5.105 ;
      RECT 51.975 3.795 51.98 4.39 ;
      RECT 51.965 3.795 51.975 4.338 ;
      RECT 51.97 4.795 51.975 5.106 ;
      RECT 51.965 4.807 51.97 5.107 ;
      RECT 51.96 3.795 51.965 4.298 ;
      RECT 51.96 4.82 51.965 5.108 ;
      RECT 51.945 4.835 51.96 5.109 ;
      RECT 51.95 3.795 51.955 4.26 ;
      RECT 51.945 3.795 51.95 4.225 ;
      RECT 51.94 3.795 51.945 4.2 ;
      RECT 51.935 4.862 51.945 5.111 ;
      RECT 51.93 3.795 51.94 4.158 ;
      RECT 51.93 4.88 51.935 5.112 ;
      RECT 51.925 3.795 51.93 4.118 ;
      RECT 51.925 4.887 51.93 5.113 ;
      RECT 51.92 3.795 51.925 4.09 ;
      RECT 51.915 4.905 51.925 5.114 ;
      RECT 51.91 3.795 51.92 4.07 ;
      RECT 51.905 4.925 51.915 5.116 ;
      RECT 51.895 4.942 51.905 5.117 ;
      RECT 51.86 4.965 51.895 5.12 ;
      RECT 51.805 4.983 51.86 5.126 ;
      RECT 51.719 4.991 51.805 5.135 ;
      RECT 51.633 5.002 51.719 5.146 ;
      RECT 51.547 5.012 51.633 5.157 ;
      RECT 51.461 5.022 51.547 5.169 ;
      RECT 51.375 5.032 51.461 5.18 ;
      RECT 51.355 5.038 51.375 5.186 ;
      RECT 51.275 5.04 51.355 5.19 ;
      RECT 51.27 5.039 51.275 5.195 ;
      RECT 51.262 5.038 51.27 5.195 ;
      RECT 51.176 5.034 51.262 5.193 ;
      RECT 51.09 5.026 51.176 5.19 ;
      RECT 51.004 5.017 51.09 5.186 ;
      RECT 50.918 5.009 51.004 5.183 ;
      RECT 50.832 5.001 50.918 5.179 ;
      RECT 50.746 4.992 50.832 5.176 ;
      RECT 50.66 4.984 50.746 5.172 ;
      RECT 50.605 4.977 50.65 5.17 ;
      RECT 50.52 4.97 50.605 5.168 ;
      RECT 50.446 4.962 50.52 5.164 ;
      RECT 50.36 4.954 50.446 5.161 ;
      RECT 50.357 4.95 50.36 5.159 ;
      RECT 50.271 4.946 50.357 5.158 ;
      RECT 50.185 4.938 50.271 5.155 ;
      RECT 50.1 4.933 50.185 5.152 ;
      RECT 50.014 4.93 50.1 5.149 ;
      RECT 49.928 4.928 50.014 5.146 ;
      RECT 49.842 4.925 49.928 5.143 ;
      RECT 49.756 4.922 49.842 5.14 ;
      RECT 49.67 4.919 49.756 5.137 ;
      RECT 49.594 4.917 49.67 5.134 ;
      RECT 49.508 4.914 49.594 5.131 ;
      RECT 49.422 4.911 49.508 5.129 ;
      RECT 49.336 4.909 49.422 5.126 ;
      RECT 49.25 4.906 49.336 5.123 ;
      RECT 49.19 4.897 49.25 5.121 ;
      RECT 51.7 4.515 51.775 4.775 ;
      RECT 51.68 4.495 51.685 4.775 ;
      RECT 51 4.28 51.105 4.575 ;
      RECT 45.445 4.255 45.515 4.515 ;
      RECT 51.34 4.13 51.345 4.501 ;
      RECT 51.33 4.185 51.335 4.501 ;
      RECT 51.635 3.355 51.695 3.615 ;
      RECT 51.69 4.51 51.7 4.775 ;
      RECT 51.685 4.5 51.69 4.775 ;
      RECT 51.605 4.447 51.68 4.775 ;
      RECT 51.63 3.355 51.635 3.635 ;
      RECT 51.62 3.355 51.63 3.655 ;
      RECT 51.605 3.355 51.62 3.685 ;
      RECT 51.59 3.355 51.605 3.728 ;
      RECT 51.585 4.39 51.605 4.775 ;
      RECT 51.575 3.355 51.59 3.765 ;
      RECT 51.57 4.37 51.585 4.775 ;
      RECT 51.57 3.355 51.575 3.788 ;
      RECT 51.56 3.355 51.57 3.813 ;
      RECT 51.53 4.337 51.57 4.775 ;
      RECT 51.535 3.355 51.56 3.863 ;
      RECT 51.53 3.355 51.535 3.918 ;
      RECT 51.525 3.355 51.53 3.96 ;
      RECT 51.515 4.3 51.53 4.775 ;
      RECT 51.52 3.355 51.525 4.003 ;
      RECT 51.515 3.355 51.52 4.068 ;
      RECT 51.51 3.355 51.515 4.09 ;
      RECT 51.51 4.288 51.515 4.64 ;
      RECT 51.505 3.355 51.51 4.158 ;
      RECT 51.505 4.28 51.51 4.623 ;
      RECT 51.5 3.355 51.505 4.203 ;
      RECT 51.495 4.262 51.505 4.6 ;
      RECT 51.495 3.355 51.5 4.24 ;
      RECT 51.485 3.355 51.495 4.58 ;
      RECT 51.48 3.355 51.485 4.563 ;
      RECT 51.475 3.355 51.48 4.548 ;
      RECT 51.47 3.355 51.475 4.533 ;
      RECT 51.45 3.355 51.47 4.523 ;
      RECT 51.445 3.355 51.45 4.513 ;
      RECT 51.435 3.355 51.445 4.509 ;
      RECT 51.43 3.632 51.435 4.508 ;
      RECT 51.425 3.655 51.43 4.507 ;
      RECT 51.42 3.685 51.425 4.506 ;
      RECT 51.415 3.712 51.42 4.505 ;
      RECT 51.41 3.74 51.415 4.505 ;
      RECT 51.405 3.767 51.41 4.505 ;
      RECT 51.4 3.787 51.405 4.505 ;
      RECT 51.395 3.815 51.4 4.505 ;
      RECT 51.385 3.857 51.395 4.505 ;
      RECT 51.375 3.902 51.385 4.504 ;
      RECT 51.37 3.955 51.375 4.503 ;
      RECT 51.365 3.987 51.37 4.502 ;
      RECT 51.36 4.007 51.365 4.501 ;
      RECT 51.355 4.045 51.36 4.501 ;
      RECT 51.35 4.067 51.355 4.501 ;
      RECT 51.345 4.092 51.35 4.501 ;
      RECT 51.335 4.157 51.34 4.501 ;
      RECT 51.32 4.217 51.33 4.501 ;
      RECT 51.305 4.227 51.32 4.501 ;
      RECT 51.285 4.237 51.305 4.501 ;
      RECT 51.255 4.242 51.285 4.498 ;
      RECT 51.195 4.252 51.255 4.495 ;
      RECT 51.175 4.261 51.195 4.5 ;
      RECT 51.15 4.267 51.175 4.513 ;
      RECT 51.13 4.272 51.15 4.528 ;
      RECT 51.105 4.277 51.13 4.575 ;
      RECT 50.976 4.279 51 4.575 ;
      RECT 50.89 4.274 50.976 4.575 ;
      RECT 50.85 4.271 50.89 4.575 ;
      RECT 50.8 4.273 50.85 4.555 ;
      RECT 50.77 4.277 50.8 4.555 ;
      RECT 50.691 4.287 50.77 4.555 ;
      RECT 50.605 4.302 50.691 4.556 ;
      RECT 50.555 4.312 50.605 4.557 ;
      RECT 50.547 4.315 50.555 4.557 ;
      RECT 50.461 4.317 50.547 4.558 ;
      RECT 50.375 4.321 50.461 4.558 ;
      RECT 50.289 4.325 50.375 4.559 ;
      RECT 50.203 4.328 50.289 4.56 ;
      RECT 50.117 4.332 50.203 4.56 ;
      RECT 50.031 4.336 50.117 4.561 ;
      RECT 49.945 4.339 50.031 4.562 ;
      RECT 49.859 4.343 49.945 4.562 ;
      RECT 49.773 4.347 49.859 4.563 ;
      RECT 49.687 4.351 49.773 4.564 ;
      RECT 49.601 4.354 49.687 4.564 ;
      RECT 49.515 4.358 49.601 4.565 ;
      RECT 49.485 4.36 49.515 4.565 ;
      RECT 49.399 4.363 49.485 4.566 ;
      RECT 49.313 4.367 49.399 4.567 ;
      RECT 49.227 4.371 49.313 4.568 ;
      RECT 49.141 4.374 49.227 4.568 ;
      RECT 49.055 4.378 49.141 4.569 ;
      RECT 49.02 4.383 49.055 4.57 ;
      RECT 48.965 4.393 49.02 4.577 ;
      RECT 48.94 4.405 48.965 4.587 ;
      RECT 48.905 4.418 48.94 4.595 ;
      RECT 48.865 4.435 48.905 4.618 ;
      RECT 48.845 4.448 48.865 4.645 ;
      RECT 48.815 4.46 48.845 4.673 ;
      RECT 48.81 4.468 48.815 4.693 ;
      RECT 48.805 4.471 48.81 4.703 ;
      RECT 48.755 4.483 48.805 4.737 ;
      RECT 48.745 4.498 48.755 4.77 ;
      RECT 48.735 4.504 48.745 4.783 ;
      RECT 48.725 4.511 48.735 4.795 ;
      RECT 48.7 4.524 48.725 4.813 ;
      RECT 48.685 4.539 48.7 4.835 ;
      RECT 48.675 4.547 48.685 4.851 ;
      RECT 48.66 4.556 48.675 4.866 ;
      RECT 48.65 4.566 48.66 4.88 ;
      RECT 48.631 4.579 48.65 4.897 ;
      RECT 48.545 4.624 48.631 4.962 ;
      RECT 48.53 4.669 48.545 5.02 ;
      RECT 48.525 4.678 48.53 5.033 ;
      RECT 48.515 4.685 48.525 5.038 ;
      RECT 48.51 4.69 48.515 5.042 ;
      RECT 48.49 4.7 48.51 5.049 ;
      RECT 48.465 4.72 48.49 5.063 ;
      RECT 48.43 4.745 48.465 5.083 ;
      RECT 48.415 4.768 48.43 5.098 ;
      RECT 48.405 4.778 48.415 5.103 ;
      RECT 48.395 4.786 48.405 5.11 ;
      RECT 48.385 4.795 48.395 5.116 ;
      RECT 48.365 4.807 48.385 5.118 ;
      RECT 48.355 4.82 48.365 5.12 ;
      RECT 48.33 4.835 48.355 5.123 ;
      RECT 48.31 4.852 48.33 5.127 ;
      RECT 48.27 4.88 48.31 5.133 ;
      RECT 48.205 4.927 48.27 5.142 ;
      RECT 48.19 4.96 48.205 5.15 ;
      RECT 48.185 4.967 48.19 5.152 ;
      RECT 48.135 4.992 48.185 5.157 ;
      RECT 48.12 5.016 48.135 5.164 ;
      RECT 48.07 5.021 48.12 5.165 ;
      RECT 47.984 5.025 48.07 5.165 ;
      RECT 47.898 5.025 47.984 5.165 ;
      RECT 47.812 5.025 47.898 5.166 ;
      RECT 47.726 5.025 47.812 5.166 ;
      RECT 47.64 5.025 47.726 5.166 ;
      RECT 47.574 5.025 47.64 5.166 ;
      RECT 47.488 5.025 47.574 5.167 ;
      RECT 47.402 5.025 47.488 5.167 ;
      RECT 47.316 5.026 47.402 5.168 ;
      RECT 47.23 5.026 47.316 5.168 ;
      RECT 47.144 5.026 47.23 5.168 ;
      RECT 47.058 5.026 47.144 5.169 ;
      RECT 46.972 5.026 47.058 5.169 ;
      RECT 46.886 5.027 46.972 5.17 ;
      RECT 46.8 5.027 46.886 5.17 ;
      RECT 46.78 5.027 46.8 5.17 ;
      RECT 46.694 5.027 46.78 5.17 ;
      RECT 46.608 5.027 46.694 5.17 ;
      RECT 46.522 5.028 46.608 5.17 ;
      RECT 46.436 5.028 46.522 5.17 ;
      RECT 46.35 5.028 46.436 5.17 ;
      RECT 46.264 5.029 46.35 5.17 ;
      RECT 46.178 5.029 46.264 5.17 ;
      RECT 46.092 5.029 46.178 5.17 ;
      RECT 46.006 5.029 46.092 5.17 ;
      RECT 45.92 5.03 46.006 5.17 ;
      RECT 45.87 5.027 45.92 5.17 ;
      RECT 45.86 5.025 45.87 5.169 ;
      RECT 45.856 5.025 45.86 5.168 ;
      RECT 45.77 5.02 45.856 5.163 ;
      RECT 45.748 5.013 45.77 5.157 ;
      RECT 45.662 5.004 45.748 5.151 ;
      RECT 45.576 4.991 45.662 5.142 ;
      RECT 45.49 4.977 45.576 5.132 ;
      RECT 45.445 4.967 45.49 5.125 ;
      RECT 45.425 4.255 45.445 4.533 ;
      RECT 45.425 4.96 45.445 5.121 ;
      RECT 45.395 4.255 45.425 4.555 ;
      RECT 45.385 4.927 45.425 5.118 ;
      RECT 45.38 4.255 45.395 4.575 ;
      RECT 45.38 4.892 45.385 5.116 ;
      RECT 45.375 4.255 45.38 4.7 ;
      RECT 45.375 4.852 45.38 5.116 ;
      RECT 45.365 4.255 45.375 5.116 ;
      RECT 45.29 4.255 45.365 5.11 ;
      RECT 45.26 4.255 45.29 5.1 ;
      RECT 45.255 4.255 45.26 5.092 ;
      RECT 45.25 4.297 45.255 5.085 ;
      RECT 45.24 4.366 45.25 5.076 ;
      RECT 45.235 4.436 45.24 5.028 ;
      RECT 45.23 4.5 45.235 4.925 ;
      RECT 45.225 4.535 45.23 4.88 ;
      RECT 45.223 4.572 45.225 4.772 ;
      RECT 45.22 4.58 45.223 4.765 ;
      RECT 45.215 4.645 45.22 4.708 ;
      RECT 49.29 3.735 49.57 4.015 ;
      RECT 49.28 3.735 49.57 3.878 ;
      RECT 49.235 3.6 49.495 3.86 ;
      RECT 49.235 3.715 49.55 3.86 ;
      RECT 49.235 3.685 49.545 3.86 ;
      RECT 49.235 3.672 49.535 3.86 ;
      RECT 49.235 3.662 49.53 3.86 ;
      RECT 45.21 3.645 45.47 3.905 ;
      RECT 48.98 3.195 49.24 3.455 ;
      RECT 48.97 3.22 49.24 3.415 ;
      RECT 48.965 3.22 48.97 3.414 ;
      RECT 48.895 3.215 48.965 3.406 ;
      RECT 48.81 3.202 48.895 3.389 ;
      RECT 48.806 3.194 48.81 3.379 ;
      RECT 48.72 3.187 48.806 3.369 ;
      RECT 48.711 3.179 48.72 3.359 ;
      RECT 48.625 3.172 48.711 3.347 ;
      RECT 48.605 3.163 48.625 3.333 ;
      RECT 48.55 3.158 48.605 3.325 ;
      RECT 48.54 3.152 48.55 3.319 ;
      RECT 48.52 3.15 48.54 3.315 ;
      RECT 48.512 3.149 48.52 3.311 ;
      RECT 48.426 3.141 48.512 3.3 ;
      RECT 48.34 3.127 48.426 3.28 ;
      RECT 48.28 3.115 48.34 3.265 ;
      RECT 48.27 3.11 48.28 3.26 ;
      RECT 48.22 3.11 48.27 3.262 ;
      RECT 48.173 3.112 48.22 3.266 ;
      RECT 48.087 3.119 48.173 3.271 ;
      RECT 48.001 3.127 48.087 3.277 ;
      RECT 47.915 3.136 48.001 3.283 ;
      RECT 47.856 3.142 47.915 3.288 ;
      RECT 47.77 3.147 47.856 3.294 ;
      RECT 47.695 3.152 47.77 3.3 ;
      RECT 47.656 3.154 47.695 3.305 ;
      RECT 47.57 3.151 47.656 3.31 ;
      RECT 47.485 3.149 47.57 3.317 ;
      RECT 47.453 3.148 47.485 3.32 ;
      RECT 47.367 3.147 47.453 3.321 ;
      RECT 47.281 3.146 47.367 3.322 ;
      RECT 47.195 3.145 47.281 3.322 ;
      RECT 47.109 3.144 47.195 3.323 ;
      RECT 47.023 3.143 47.109 3.324 ;
      RECT 46.937 3.142 47.023 3.325 ;
      RECT 46.851 3.141 46.937 3.325 ;
      RECT 46.765 3.14 46.851 3.326 ;
      RECT 46.715 3.14 46.765 3.327 ;
      RECT 46.701 3.141 46.715 3.327 ;
      RECT 46.615 3.148 46.701 3.328 ;
      RECT 46.541 3.159 46.615 3.329 ;
      RECT 46.455 3.168 46.541 3.33 ;
      RECT 46.42 3.175 46.455 3.345 ;
      RECT 46.395 3.178 46.42 3.375 ;
      RECT 46.37 3.187 46.395 3.404 ;
      RECT 46.36 3.198 46.37 3.424 ;
      RECT 46.35 3.206 46.36 3.438 ;
      RECT 46.345 3.212 46.35 3.448 ;
      RECT 46.32 3.229 46.345 3.465 ;
      RECT 46.305 3.251 46.32 3.493 ;
      RECT 46.275 3.277 46.305 3.523 ;
      RECT 46.255 3.306 46.275 3.553 ;
      RECT 46.25 3.321 46.255 3.57 ;
      RECT 46.23 3.336 46.25 3.585 ;
      RECT 46.22 3.354 46.23 3.603 ;
      RECT 46.21 3.365 46.22 3.618 ;
      RECT 46.16 3.397 46.21 3.644 ;
      RECT 46.155 3.427 46.16 3.664 ;
      RECT 46.145 3.44 46.155 3.67 ;
      RECT 46.136 3.45 46.145 3.678 ;
      RECT 46.125 3.461 46.136 3.686 ;
      RECT 46.12 3.471 46.125 3.692 ;
      RECT 46.105 3.492 46.12 3.699 ;
      RECT 46.09 3.522 46.105 3.707 ;
      RECT 46.055 3.552 46.09 3.713 ;
      RECT 46.03 3.57 46.055 3.72 ;
      RECT 45.98 3.578 46.03 3.729 ;
      RECT 45.955 3.583 45.98 3.738 ;
      RECT 45.9 3.589 45.955 3.748 ;
      RECT 45.895 3.594 45.9 3.756 ;
      RECT 45.881 3.597 45.895 3.758 ;
      RECT 45.795 3.609 45.881 3.77 ;
      RECT 45.785 3.621 45.795 3.783 ;
      RECT 45.7 3.634 45.785 3.795 ;
      RECT 45.656 3.651 45.7 3.809 ;
      RECT 45.57 3.668 45.656 3.825 ;
      RECT 45.54 3.682 45.57 3.839 ;
      RECT 45.53 3.687 45.54 3.844 ;
      RECT 45.47 3.69 45.53 3.853 ;
      RECT 48.36 3.96 48.62 4.22 ;
      RECT 48.36 3.96 48.64 4.073 ;
      RECT 48.36 3.96 48.665 4.04 ;
      RECT 48.36 3.96 48.67 4.02 ;
      RECT 48.41 3.735 48.69 4.015 ;
      RECT 47.965 4.47 48.225 4.73 ;
      RECT 47.955 4.327 48.15 4.668 ;
      RECT 47.95 4.435 48.165 4.66 ;
      RECT 47.945 4.485 48.225 4.65 ;
      RECT 47.935 4.562 48.225 4.635 ;
      RECT 47.955 4.41 48.165 4.668 ;
      RECT 47.965 4.285 48.15 4.73 ;
      RECT 47.965 4.18 48.13 4.73 ;
      RECT 47.975 4.167 48.13 4.73 ;
      RECT 47.975 4.125 48.12 4.73 ;
      RECT 47.98 4.05 48.12 4.73 ;
      RECT 48.01 3.7 48.12 4.73 ;
      RECT 48.015 3.43 48.14 4.053 ;
      RECT 47.985 4.005 48.14 4.053 ;
      RECT 48 3.807 48.12 4.73 ;
      RECT 47.99 3.917 48.14 4.053 ;
      RECT 48.015 3.43 48.155 3.91 ;
      RECT 48.015 3.43 48.175 3.785 ;
      RECT 47.98 3.43 48.24 3.69 ;
      RECT 47.45 3.735 47.73 4.015 ;
      RECT 47.435 3.735 47.73 3.995 ;
      RECT 45.49 4.6 45.75 4.86 ;
      RECT 47.275 4.455 47.535 4.715 ;
      RECT 47.255 4.475 47.535 4.69 ;
      RECT 47.212 4.475 47.255 4.689 ;
      RECT 47.126 4.476 47.212 4.686 ;
      RECT 47.04 4.477 47.126 4.682 ;
      RECT 46.965 4.479 47.04 4.679 ;
      RECT 46.942 4.48 46.965 4.677 ;
      RECT 46.856 4.481 46.942 4.675 ;
      RECT 46.77 4.482 46.856 4.672 ;
      RECT 46.746 4.483 46.77 4.67 ;
      RECT 46.66 4.485 46.746 4.667 ;
      RECT 46.575 4.487 46.66 4.668 ;
      RECT 46.518 4.488 46.575 4.674 ;
      RECT 46.432 4.49 46.518 4.684 ;
      RECT 46.346 4.493 46.432 4.697 ;
      RECT 46.26 4.495 46.346 4.709 ;
      RECT 46.246 4.496 46.26 4.716 ;
      RECT 46.16 4.497 46.246 4.724 ;
      RECT 46.12 4.499 46.16 4.733 ;
      RECT 46.111 4.5 46.12 4.736 ;
      RECT 46.025 4.508 46.111 4.742 ;
      RECT 46.005 4.517 46.025 4.75 ;
      RECT 45.92 4.532 46.005 4.758 ;
      RECT 45.86 4.555 45.92 4.769 ;
      RECT 45.85 4.567 45.86 4.774 ;
      RECT 45.81 4.577 45.85 4.778 ;
      RECT 45.755 4.594 45.81 4.786 ;
      RECT 45.75 4.604 45.755 4.79 ;
      RECT 46.816 3.735 46.875 4.132 ;
      RECT 46.73 3.735 46.935 4.123 ;
      RECT 46.725 3.765 46.935 4.118 ;
      RECT 46.691 3.765 46.935 4.116 ;
      RECT 46.605 3.765 46.935 4.11 ;
      RECT 46.56 3.765 46.955 4.088 ;
      RECT 46.56 3.765 46.975 4.043 ;
      RECT 46.52 3.765 46.975 4.033 ;
      RECT 46.73 3.735 47.01 4.015 ;
      RECT 46.465 3.735 46.725 3.995 ;
      RECT 45.65 3.215 45.91 3.475 ;
      RECT 45.73 3.175 46.01 3.455 ;
      RECT 40.105 8.505 40.425 8.83 ;
      RECT 40.135 7.98 40.305 8.83 ;
      RECT 40.135 7.98 40.31 8.33 ;
      RECT 40.135 7.98 41.11 8.155 ;
      RECT 40.935 3.26 41.11 8.155 ;
      RECT 40.88 3.26 41.23 3.61 ;
      RECT 40.905 8.94 41.23 9.265 ;
      RECT 39.79 9.03 41.23 9.2 ;
      RECT 39.79 3.69 39.95 9.2 ;
      RECT 40.105 3.66 40.425 3.98 ;
      RECT 39.79 3.69 40.425 3.86 ;
      RECT 28.515 4.295 28.795 4.575 ;
      RECT 28.485 4.295 28.795 4.56 ;
      RECT 28.48 4.295 28.795 4.558 ;
      RECT 28.475 2.625 28.645 4.552 ;
      RECT 28.47 4.262 28.74 4.545 ;
      RECT 28.465 4.295 28.795 4.538 ;
      RECT 28.435 4.265 28.74 4.525 ;
      RECT 28.435 4.292 28.76 4.525 ;
      RECT 28.435 4.282 28.755 4.525 ;
      RECT 28.435 4.267 28.75 4.525 ;
      RECT 28.475 4.257 28.74 4.552 ;
      RECT 28.475 4.252 28.73 4.552 ;
      RECT 28.475 4.251 28.715 4.552 ;
      RECT 38.445 2.635 38.795 2.985 ;
      RECT 38.44 2.635 38.795 2.89 ;
      RECT 28.475 2.625 38.685 2.795 ;
      RECT 38.12 4.145 38.49 4.515 ;
      RECT 38.205 3.53 38.375 4.515 ;
      RECT 34.225 3.75 34.46 4.01 ;
      RECT 37.37 3.53 37.535 3.79 ;
      RECT 37.275 3.52 37.29 3.79 ;
      RECT 37.37 3.53 38.375 3.71 ;
      RECT 35.875 3.09 35.915 3.23 ;
      RECT 37.29 3.525 37.37 3.79 ;
      RECT 37.235 3.52 37.275 3.756 ;
      RECT 37.221 3.52 37.235 3.756 ;
      RECT 37.135 3.525 37.221 3.758 ;
      RECT 37.09 3.532 37.135 3.76 ;
      RECT 37.06 3.532 37.09 3.762 ;
      RECT 37.035 3.527 37.06 3.764 ;
      RECT 37.005 3.523 37.035 3.773 ;
      RECT 36.995 3.52 37.005 3.785 ;
      RECT 36.99 3.52 36.995 3.793 ;
      RECT 36.985 3.52 36.99 3.798 ;
      RECT 36.975 3.519 36.985 3.808 ;
      RECT 36.97 3.518 36.975 3.818 ;
      RECT 36.955 3.517 36.97 3.823 ;
      RECT 36.927 3.514 36.955 3.85 ;
      RECT 36.841 3.506 36.927 3.85 ;
      RECT 36.755 3.495 36.841 3.85 ;
      RECT 36.715 3.48 36.755 3.85 ;
      RECT 36.675 3.454 36.715 3.85 ;
      RECT 36.67 3.436 36.675 3.662 ;
      RECT 36.66 3.432 36.67 3.652 ;
      RECT 36.645 3.422 36.66 3.639 ;
      RECT 36.625 3.406 36.645 3.624 ;
      RECT 36.61 3.391 36.625 3.609 ;
      RECT 36.6 3.38 36.61 3.599 ;
      RECT 36.575 3.364 36.6 3.588 ;
      RECT 36.57 3.351 36.575 3.578 ;
      RECT 36.565 3.347 36.57 3.573 ;
      RECT 36.51 3.333 36.565 3.551 ;
      RECT 36.471 3.314 36.51 3.515 ;
      RECT 36.385 3.288 36.471 3.468 ;
      RECT 36.381 3.27 36.385 3.434 ;
      RECT 36.295 3.251 36.381 3.412 ;
      RECT 36.29 3.233 36.295 3.39 ;
      RECT 36.285 3.231 36.29 3.388 ;
      RECT 36.275 3.23 36.285 3.383 ;
      RECT 36.215 3.217 36.275 3.369 ;
      RECT 36.17 3.195 36.215 3.348 ;
      RECT 36.11 3.172 36.17 3.327 ;
      RECT 36.046 3.147 36.11 3.302 ;
      RECT 35.96 3.117 36.046 3.271 ;
      RECT 35.945 3.097 35.96 3.25 ;
      RECT 35.915 3.092 35.945 3.241 ;
      RECT 35.862 3.09 35.875 3.23 ;
      RECT 35.776 3.09 35.862 3.232 ;
      RECT 35.69 3.09 35.776 3.234 ;
      RECT 35.67 3.09 35.69 3.238 ;
      RECT 35.625 3.092 35.67 3.249 ;
      RECT 35.585 3.102 35.625 3.265 ;
      RECT 35.581 3.111 35.585 3.273 ;
      RECT 35.495 3.131 35.581 3.289 ;
      RECT 35.485 3.15 35.495 3.307 ;
      RECT 35.48 3.152 35.485 3.31 ;
      RECT 35.47 3.156 35.48 3.313 ;
      RECT 35.45 3.161 35.47 3.323 ;
      RECT 35.42 3.171 35.45 3.343 ;
      RECT 35.415 3.178 35.42 3.357 ;
      RECT 35.405 3.182 35.415 3.364 ;
      RECT 35.39 3.19 35.405 3.375 ;
      RECT 35.38 3.2 35.39 3.386 ;
      RECT 35.37 3.207 35.38 3.394 ;
      RECT 35.345 3.22 35.37 3.409 ;
      RECT 35.281 3.256 35.345 3.448 ;
      RECT 35.195 3.319 35.281 3.512 ;
      RECT 35.16 3.37 35.195 3.565 ;
      RECT 35.155 3.387 35.16 3.582 ;
      RECT 35.14 3.396 35.155 3.589 ;
      RECT 35.12 3.411 35.14 3.603 ;
      RECT 35.115 3.422 35.12 3.613 ;
      RECT 35.095 3.435 35.115 3.623 ;
      RECT 35.09 3.445 35.095 3.633 ;
      RECT 35.075 3.45 35.09 3.642 ;
      RECT 35.065 3.46 35.075 3.653 ;
      RECT 35.035 3.477 35.065 3.67 ;
      RECT 35.025 3.495 35.035 3.688 ;
      RECT 35.01 3.506 35.025 3.699 ;
      RECT 34.97 3.53 35.01 3.715 ;
      RECT 34.935 3.564 34.97 3.732 ;
      RECT 34.905 3.587 34.935 3.744 ;
      RECT 34.89 3.597 34.905 3.753 ;
      RECT 34.85 3.607 34.89 3.764 ;
      RECT 34.83 3.618 34.85 3.776 ;
      RECT 34.825 3.622 34.83 3.783 ;
      RECT 34.81 3.626 34.825 3.788 ;
      RECT 34.8 3.631 34.81 3.793 ;
      RECT 34.795 3.634 34.8 3.796 ;
      RECT 34.765 3.64 34.795 3.803 ;
      RECT 34.73 3.65 34.765 3.817 ;
      RECT 34.67 3.665 34.73 3.837 ;
      RECT 34.615 3.685 34.67 3.861 ;
      RECT 34.586 3.7 34.615 3.879 ;
      RECT 34.5 3.72 34.586 3.904 ;
      RECT 34.495 3.735 34.5 3.924 ;
      RECT 34.485 3.738 34.495 3.925 ;
      RECT 34.46 3.745 34.485 4.01 ;
      RECT 37.155 4.238 37.435 4.575 ;
      RECT 37.155 4.248 37.44 4.533 ;
      RECT 37.155 4.257 37.445 4.43 ;
      RECT 37.155 4.272 37.45 4.298 ;
      RECT 37.155 4.1 37.415 4.575 ;
      RECT 27.505 8.94 27.855 9.29 ;
      RECT 36.33 8.895 36.68 9.245 ;
      RECT 27.505 8.97 36.68 9.17 ;
      RECT 34.875 4.98 34.885 5.17 ;
      RECT 33.135 4.855 33.415 5.135 ;
      RECT 36.18 3.795 36.185 4.28 ;
      RECT 36.075 3.795 36.135 4.055 ;
      RECT 36.4 4.765 36.405 4.84 ;
      RECT 36.39 4.632 36.4 4.875 ;
      RECT 36.38 4.467 36.39 4.896 ;
      RECT 36.375 4.337 36.38 4.912 ;
      RECT 36.365 4.227 36.375 4.928 ;
      RECT 36.36 4.126 36.365 4.945 ;
      RECT 36.355 4.108 36.36 4.955 ;
      RECT 36.35 4.09 36.355 4.965 ;
      RECT 36.34 4.065 36.35 4.98 ;
      RECT 36.335 4.045 36.34 4.995 ;
      RECT 36.315 3.795 36.335 5.02 ;
      RECT 36.3 3.795 36.315 5.053 ;
      RECT 36.27 3.795 36.3 5.075 ;
      RECT 36.25 3.795 36.27 5.089 ;
      RECT 36.23 3.795 36.25 4.605 ;
      RECT 36.245 4.672 36.25 5.094 ;
      RECT 36.24 4.702 36.245 5.096 ;
      RECT 36.235 4.715 36.24 5.099 ;
      RECT 36.23 4.725 36.235 5.103 ;
      RECT 36.225 3.795 36.23 4.523 ;
      RECT 36.225 4.735 36.23 5.105 ;
      RECT 36.22 3.795 36.225 4.5 ;
      RECT 36.21 4.757 36.225 5.105 ;
      RECT 36.205 3.795 36.22 4.445 ;
      RECT 36.2 4.782 36.21 5.105 ;
      RECT 36.2 3.795 36.205 4.39 ;
      RECT 36.19 3.795 36.2 4.338 ;
      RECT 36.195 4.795 36.2 5.106 ;
      RECT 36.19 4.807 36.195 5.107 ;
      RECT 36.185 3.795 36.19 4.298 ;
      RECT 36.185 4.82 36.19 5.108 ;
      RECT 36.17 4.835 36.185 5.109 ;
      RECT 36.175 3.795 36.18 4.26 ;
      RECT 36.17 3.795 36.175 4.225 ;
      RECT 36.165 3.795 36.17 4.2 ;
      RECT 36.16 4.862 36.17 5.111 ;
      RECT 36.155 3.795 36.165 4.158 ;
      RECT 36.155 4.88 36.16 5.112 ;
      RECT 36.15 3.795 36.155 4.118 ;
      RECT 36.15 4.887 36.155 5.113 ;
      RECT 36.145 3.795 36.15 4.09 ;
      RECT 36.14 4.905 36.15 5.114 ;
      RECT 36.135 3.795 36.145 4.07 ;
      RECT 36.13 4.925 36.14 5.116 ;
      RECT 36.12 4.942 36.13 5.117 ;
      RECT 36.085 4.965 36.12 5.12 ;
      RECT 36.03 4.983 36.085 5.126 ;
      RECT 35.944 4.991 36.03 5.135 ;
      RECT 35.858 5.002 35.944 5.146 ;
      RECT 35.772 5.012 35.858 5.157 ;
      RECT 35.686 5.022 35.772 5.169 ;
      RECT 35.6 5.032 35.686 5.18 ;
      RECT 35.58 5.038 35.6 5.186 ;
      RECT 35.5 5.04 35.58 5.19 ;
      RECT 35.495 5.039 35.5 5.195 ;
      RECT 35.487 5.038 35.495 5.195 ;
      RECT 35.401 5.034 35.487 5.193 ;
      RECT 35.315 5.026 35.401 5.19 ;
      RECT 35.229 5.017 35.315 5.186 ;
      RECT 35.143 5.009 35.229 5.183 ;
      RECT 35.057 5.001 35.143 5.179 ;
      RECT 34.971 4.992 35.057 5.176 ;
      RECT 34.885 4.984 34.971 5.172 ;
      RECT 34.83 4.977 34.875 5.17 ;
      RECT 34.745 4.97 34.83 5.168 ;
      RECT 34.671 4.962 34.745 5.164 ;
      RECT 34.585 4.954 34.671 5.161 ;
      RECT 34.582 4.95 34.585 5.159 ;
      RECT 34.496 4.946 34.582 5.158 ;
      RECT 34.41 4.938 34.496 5.155 ;
      RECT 34.325 4.933 34.41 5.152 ;
      RECT 34.239 4.93 34.325 5.149 ;
      RECT 34.153 4.928 34.239 5.146 ;
      RECT 34.067 4.925 34.153 5.143 ;
      RECT 33.981 4.922 34.067 5.14 ;
      RECT 33.895 4.919 33.981 5.137 ;
      RECT 33.819 4.917 33.895 5.134 ;
      RECT 33.733 4.914 33.819 5.131 ;
      RECT 33.647 4.911 33.733 5.129 ;
      RECT 33.561 4.909 33.647 5.126 ;
      RECT 33.475 4.906 33.561 5.123 ;
      RECT 33.415 4.897 33.475 5.121 ;
      RECT 35.925 4.515 36 4.775 ;
      RECT 35.905 4.495 35.91 4.775 ;
      RECT 35.225 4.28 35.33 4.575 ;
      RECT 29.67 4.255 29.74 4.515 ;
      RECT 35.565 4.13 35.57 4.501 ;
      RECT 35.555 4.185 35.56 4.501 ;
      RECT 35.86 3.355 35.92 3.615 ;
      RECT 35.915 4.51 35.925 4.775 ;
      RECT 35.91 4.5 35.915 4.775 ;
      RECT 35.83 4.447 35.905 4.775 ;
      RECT 35.855 3.355 35.86 3.635 ;
      RECT 35.845 3.355 35.855 3.655 ;
      RECT 35.83 3.355 35.845 3.685 ;
      RECT 35.815 3.355 35.83 3.728 ;
      RECT 35.81 4.39 35.83 4.775 ;
      RECT 35.8 3.355 35.815 3.765 ;
      RECT 35.795 4.37 35.81 4.775 ;
      RECT 35.795 3.355 35.8 3.788 ;
      RECT 35.785 3.355 35.795 3.813 ;
      RECT 35.755 4.337 35.795 4.775 ;
      RECT 35.76 3.355 35.785 3.863 ;
      RECT 35.755 3.355 35.76 3.918 ;
      RECT 35.75 3.355 35.755 3.96 ;
      RECT 35.74 4.3 35.755 4.775 ;
      RECT 35.745 3.355 35.75 4.003 ;
      RECT 35.74 3.355 35.745 4.068 ;
      RECT 35.735 3.355 35.74 4.09 ;
      RECT 35.735 4.288 35.74 4.64 ;
      RECT 35.73 3.355 35.735 4.158 ;
      RECT 35.73 4.28 35.735 4.623 ;
      RECT 35.725 3.355 35.73 4.203 ;
      RECT 35.72 4.262 35.73 4.6 ;
      RECT 35.72 3.355 35.725 4.24 ;
      RECT 35.71 3.355 35.72 4.58 ;
      RECT 35.705 3.355 35.71 4.563 ;
      RECT 35.7 3.355 35.705 4.548 ;
      RECT 35.695 3.355 35.7 4.533 ;
      RECT 35.675 3.355 35.695 4.523 ;
      RECT 35.67 3.355 35.675 4.513 ;
      RECT 35.66 3.355 35.67 4.509 ;
      RECT 35.655 3.632 35.66 4.508 ;
      RECT 35.65 3.655 35.655 4.507 ;
      RECT 35.645 3.685 35.65 4.506 ;
      RECT 35.64 3.712 35.645 4.505 ;
      RECT 35.635 3.74 35.64 4.505 ;
      RECT 35.63 3.767 35.635 4.505 ;
      RECT 35.625 3.787 35.63 4.505 ;
      RECT 35.62 3.815 35.625 4.505 ;
      RECT 35.61 3.857 35.62 4.505 ;
      RECT 35.6 3.902 35.61 4.504 ;
      RECT 35.595 3.955 35.6 4.503 ;
      RECT 35.59 3.987 35.595 4.502 ;
      RECT 35.585 4.007 35.59 4.501 ;
      RECT 35.58 4.045 35.585 4.501 ;
      RECT 35.575 4.067 35.58 4.501 ;
      RECT 35.57 4.092 35.575 4.501 ;
      RECT 35.56 4.157 35.565 4.501 ;
      RECT 35.545 4.217 35.555 4.501 ;
      RECT 35.53 4.227 35.545 4.501 ;
      RECT 35.51 4.237 35.53 4.501 ;
      RECT 35.48 4.242 35.51 4.498 ;
      RECT 35.42 4.252 35.48 4.495 ;
      RECT 35.4 4.261 35.42 4.5 ;
      RECT 35.375 4.267 35.4 4.513 ;
      RECT 35.355 4.272 35.375 4.528 ;
      RECT 35.33 4.277 35.355 4.575 ;
      RECT 35.201 4.279 35.225 4.575 ;
      RECT 35.115 4.274 35.201 4.575 ;
      RECT 35.075 4.271 35.115 4.575 ;
      RECT 35.025 4.273 35.075 4.555 ;
      RECT 34.995 4.277 35.025 4.555 ;
      RECT 34.916 4.287 34.995 4.555 ;
      RECT 34.83 4.302 34.916 4.556 ;
      RECT 34.78 4.312 34.83 4.557 ;
      RECT 34.772 4.315 34.78 4.557 ;
      RECT 34.686 4.317 34.772 4.558 ;
      RECT 34.6 4.321 34.686 4.558 ;
      RECT 34.514 4.325 34.6 4.559 ;
      RECT 34.428 4.328 34.514 4.56 ;
      RECT 34.342 4.332 34.428 4.56 ;
      RECT 34.256 4.336 34.342 4.561 ;
      RECT 34.17 4.339 34.256 4.562 ;
      RECT 34.084 4.343 34.17 4.562 ;
      RECT 33.998 4.347 34.084 4.563 ;
      RECT 33.912 4.351 33.998 4.564 ;
      RECT 33.826 4.354 33.912 4.564 ;
      RECT 33.74 4.358 33.826 4.565 ;
      RECT 33.71 4.36 33.74 4.565 ;
      RECT 33.624 4.363 33.71 4.566 ;
      RECT 33.538 4.367 33.624 4.567 ;
      RECT 33.452 4.371 33.538 4.568 ;
      RECT 33.366 4.374 33.452 4.568 ;
      RECT 33.28 4.378 33.366 4.569 ;
      RECT 33.245 4.383 33.28 4.57 ;
      RECT 33.19 4.393 33.245 4.577 ;
      RECT 33.165 4.405 33.19 4.587 ;
      RECT 33.13 4.418 33.165 4.595 ;
      RECT 33.09 4.435 33.13 4.618 ;
      RECT 33.07 4.448 33.09 4.645 ;
      RECT 33.04 4.46 33.07 4.673 ;
      RECT 33.035 4.468 33.04 4.693 ;
      RECT 33.03 4.471 33.035 4.703 ;
      RECT 32.98 4.483 33.03 4.737 ;
      RECT 32.97 4.498 32.98 4.77 ;
      RECT 32.96 4.504 32.97 4.783 ;
      RECT 32.95 4.511 32.96 4.795 ;
      RECT 32.925 4.524 32.95 4.813 ;
      RECT 32.91 4.539 32.925 4.835 ;
      RECT 32.9 4.547 32.91 4.851 ;
      RECT 32.885 4.556 32.9 4.866 ;
      RECT 32.875 4.566 32.885 4.88 ;
      RECT 32.856 4.579 32.875 4.897 ;
      RECT 32.77 4.624 32.856 4.962 ;
      RECT 32.755 4.669 32.77 5.02 ;
      RECT 32.75 4.678 32.755 5.033 ;
      RECT 32.74 4.685 32.75 5.038 ;
      RECT 32.735 4.69 32.74 5.042 ;
      RECT 32.715 4.7 32.735 5.049 ;
      RECT 32.69 4.72 32.715 5.063 ;
      RECT 32.655 4.745 32.69 5.083 ;
      RECT 32.64 4.768 32.655 5.098 ;
      RECT 32.63 4.778 32.64 5.103 ;
      RECT 32.62 4.786 32.63 5.11 ;
      RECT 32.61 4.795 32.62 5.116 ;
      RECT 32.59 4.807 32.61 5.118 ;
      RECT 32.58 4.82 32.59 5.12 ;
      RECT 32.555 4.835 32.58 5.123 ;
      RECT 32.535 4.852 32.555 5.127 ;
      RECT 32.495 4.88 32.535 5.133 ;
      RECT 32.43 4.927 32.495 5.142 ;
      RECT 32.415 4.96 32.43 5.15 ;
      RECT 32.41 4.967 32.415 5.152 ;
      RECT 32.36 4.992 32.41 5.157 ;
      RECT 32.345 5.016 32.36 5.164 ;
      RECT 32.295 5.021 32.345 5.165 ;
      RECT 32.209 5.025 32.295 5.165 ;
      RECT 32.123 5.025 32.209 5.165 ;
      RECT 32.037 5.025 32.123 5.166 ;
      RECT 31.951 5.025 32.037 5.166 ;
      RECT 31.865 5.025 31.951 5.166 ;
      RECT 31.799 5.025 31.865 5.166 ;
      RECT 31.713 5.025 31.799 5.167 ;
      RECT 31.627 5.025 31.713 5.167 ;
      RECT 31.541 5.026 31.627 5.168 ;
      RECT 31.455 5.026 31.541 5.168 ;
      RECT 31.369 5.026 31.455 5.168 ;
      RECT 31.283 5.026 31.369 5.169 ;
      RECT 31.197 5.026 31.283 5.169 ;
      RECT 31.111 5.027 31.197 5.17 ;
      RECT 31.025 5.027 31.111 5.17 ;
      RECT 31.005 5.027 31.025 5.17 ;
      RECT 30.919 5.027 31.005 5.17 ;
      RECT 30.833 5.027 30.919 5.17 ;
      RECT 30.747 5.028 30.833 5.17 ;
      RECT 30.661 5.028 30.747 5.17 ;
      RECT 30.575 5.028 30.661 5.17 ;
      RECT 30.489 5.029 30.575 5.17 ;
      RECT 30.403 5.029 30.489 5.17 ;
      RECT 30.317 5.029 30.403 5.17 ;
      RECT 30.231 5.029 30.317 5.17 ;
      RECT 30.145 5.03 30.231 5.17 ;
      RECT 30.095 5.027 30.145 5.17 ;
      RECT 30.085 5.025 30.095 5.169 ;
      RECT 30.081 5.025 30.085 5.168 ;
      RECT 29.995 5.02 30.081 5.163 ;
      RECT 29.973 5.013 29.995 5.157 ;
      RECT 29.887 5.004 29.973 5.151 ;
      RECT 29.801 4.991 29.887 5.142 ;
      RECT 29.715 4.977 29.801 5.132 ;
      RECT 29.67 4.967 29.715 5.125 ;
      RECT 29.65 4.255 29.67 4.533 ;
      RECT 29.65 4.96 29.67 5.121 ;
      RECT 29.62 4.255 29.65 4.555 ;
      RECT 29.61 4.927 29.65 5.118 ;
      RECT 29.605 4.255 29.62 4.575 ;
      RECT 29.605 4.892 29.61 5.116 ;
      RECT 29.6 4.255 29.605 4.7 ;
      RECT 29.6 4.852 29.605 5.116 ;
      RECT 29.59 4.255 29.6 5.116 ;
      RECT 29.515 4.255 29.59 5.11 ;
      RECT 29.485 4.255 29.515 5.1 ;
      RECT 29.48 4.255 29.485 5.092 ;
      RECT 29.475 4.297 29.48 5.085 ;
      RECT 29.465 4.366 29.475 5.076 ;
      RECT 29.46 4.436 29.465 5.028 ;
      RECT 29.455 4.5 29.46 4.925 ;
      RECT 29.45 4.535 29.455 4.88 ;
      RECT 29.448 4.572 29.45 4.772 ;
      RECT 29.445 4.58 29.448 4.765 ;
      RECT 29.44 4.645 29.445 4.708 ;
      RECT 33.515 3.735 33.795 4.015 ;
      RECT 33.505 3.735 33.795 3.878 ;
      RECT 33.46 3.6 33.72 3.86 ;
      RECT 33.46 3.715 33.775 3.86 ;
      RECT 33.46 3.685 33.77 3.86 ;
      RECT 33.46 3.672 33.76 3.86 ;
      RECT 33.46 3.662 33.755 3.86 ;
      RECT 29.435 3.645 29.695 3.905 ;
      RECT 33.205 3.195 33.465 3.455 ;
      RECT 33.195 3.22 33.465 3.415 ;
      RECT 33.19 3.22 33.195 3.414 ;
      RECT 33.12 3.215 33.19 3.406 ;
      RECT 33.035 3.202 33.12 3.389 ;
      RECT 33.031 3.194 33.035 3.379 ;
      RECT 32.945 3.187 33.031 3.369 ;
      RECT 32.936 3.179 32.945 3.359 ;
      RECT 32.85 3.172 32.936 3.347 ;
      RECT 32.83 3.163 32.85 3.333 ;
      RECT 32.775 3.158 32.83 3.325 ;
      RECT 32.765 3.152 32.775 3.319 ;
      RECT 32.745 3.15 32.765 3.315 ;
      RECT 32.737 3.149 32.745 3.311 ;
      RECT 32.651 3.141 32.737 3.3 ;
      RECT 32.565 3.127 32.651 3.28 ;
      RECT 32.505 3.115 32.565 3.265 ;
      RECT 32.495 3.11 32.505 3.26 ;
      RECT 32.445 3.11 32.495 3.262 ;
      RECT 32.398 3.112 32.445 3.266 ;
      RECT 32.312 3.119 32.398 3.271 ;
      RECT 32.226 3.127 32.312 3.277 ;
      RECT 32.14 3.136 32.226 3.283 ;
      RECT 32.081 3.142 32.14 3.288 ;
      RECT 31.995 3.147 32.081 3.294 ;
      RECT 31.92 3.152 31.995 3.3 ;
      RECT 31.881 3.154 31.92 3.305 ;
      RECT 31.795 3.151 31.881 3.31 ;
      RECT 31.71 3.149 31.795 3.317 ;
      RECT 31.678 3.148 31.71 3.32 ;
      RECT 31.592 3.147 31.678 3.321 ;
      RECT 31.506 3.146 31.592 3.322 ;
      RECT 31.42 3.145 31.506 3.322 ;
      RECT 31.334 3.144 31.42 3.323 ;
      RECT 31.248 3.143 31.334 3.324 ;
      RECT 31.162 3.142 31.248 3.325 ;
      RECT 31.076 3.141 31.162 3.325 ;
      RECT 30.99 3.14 31.076 3.326 ;
      RECT 30.94 3.14 30.99 3.327 ;
      RECT 30.926 3.141 30.94 3.327 ;
      RECT 30.84 3.148 30.926 3.328 ;
      RECT 30.766 3.159 30.84 3.329 ;
      RECT 30.68 3.168 30.766 3.33 ;
      RECT 30.645 3.175 30.68 3.345 ;
      RECT 30.62 3.178 30.645 3.375 ;
      RECT 30.595 3.187 30.62 3.404 ;
      RECT 30.585 3.198 30.595 3.424 ;
      RECT 30.575 3.206 30.585 3.438 ;
      RECT 30.57 3.212 30.575 3.448 ;
      RECT 30.545 3.229 30.57 3.465 ;
      RECT 30.53 3.251 30.545 3.493 ;
      RECT 30.5 3.277 30.53 3.523 ;
      RECT 30.48 3.306 30.5 3.553 ;
      RECT 30.475 3.321 30.48 3.57 ;
      RECT 30.455 3.336 30.475 3.585 ;
      RECT 30.445 3.354 30.455 3.603 ;
      RECT 30.435 3.365 30.445 3.618 ;
      RECT 30.385 3.397 30.435 3.644 ;
      RECT 30.38 3.427 30.385 3.664 ;
      RECT 30.37 3.44 30.38 3.67 ;
      RECT 30.361 3.45 30.37 3.678 ;
      RECT 30.35 3.461 30.361 3.686 ;
      RECT 30.345 3.471 30.35 3.692 ;
      RECT 30.33 3.492 30.345 3.699 ;
      RECT 30.315 3.522 30.33 3.707 ;
      RECT 30.28 3.552 30.315 3.713 ;
      RECT 30.255 3.57 30.28 3.72 ;
      RECT 30.205 3.578 30.255 3.729 ;
      RECT 30.18 3.583 30.205 3.738 ;
      RECT 30.125 3.589 30.18 3.748 ;
      RECT 30.12 3.594 30.125 3.756 ;
      RECT 30.106 3.597 30.12 3.758 ;
      RECT 30.02 3.609 30.106 3.77 ;
      RECT 30.01 3.621 30.02 3.783 ;
      RECT 29.925 3.634 30.01 3.795 ;
      RECT 29.881 3.651 29.925 3.809 ;
      RECT 29.795 3.668 29.881 3.825 ;
      RECT 29.765 3.682 29.795 3.839 ;
      RECT 29.755 3.687 29.765 3.844 ;
      RECT 29.695 3.69 29.755 3.853 ;
      RECT 32.585 3.96 32.845 4.22 ;
      RECT 32.585 3.96 32.865 4.073 ;
      RECT 32.585 3.96 32.89 4.04 ;
      RECT 32.585 3.96 32.895 4.02 ;
      RECT 32.635 3.735 32.915 4.015 ;
      RECT 32.19 4.47 32.45 4.73 ;
      RECT 32.18 4.327 32.375 4.668 ;
      RECT 32.175 4.435 32.39 4.66 ;
      RECT 32.17 4.485 32.45 4.65 ;
      RECT 32.16 4.562 32.45 4.635 ;
      RECT 32.18 4.41 32.39 4.668 ;
      RECT 32.19 4.285 32.375 4.73 ;
      RECT 32.19 4.18 32.355 4.73 ;
      RECT 32.2 4.167 32.355 4.73 ;
      RECT 32.2 4.125 32.345 4.73 ;
      RECT 32.205 4.05 32.345 4.73 ;
      RECT 32.235 3.7 32.345 4.73 ;
      RECT 32.24 3.43 32.365 4.053 ;
      RECT 32.21 4.005 32.365 4.053 ;
      RECT 32.225 3.807 32.345 4.73 ;
      RECT 32.215 3.917 32.365 4.053 ;
      RECT 32.24 3.43 32.38 3.91 ;
      RECT 32.24 3.43 32.4 3.785 ;
      RECT 32.205 3.43 32.465 3.69 ;
      RECT 31.675 3.735 31.955 4.015 ;
      RECT 31.66 3.735 31.955 3.995 ;
      RECT 29.715 4.6 29.975 4.86 ;
      RECT 31.5 4.455 31.76 4.715 ;
      RECT 31.48 4.475 31.76 4.69 ;
      RECT 31.437 4.475 31.48 4.689 ;
      RECT 31.351 4.476 31.437 4.686 ;
      RECT 31.265 4.477 31.351 4.682 ;
      RECT 31.19 4.479 31.265 4.679 ;
      RECT 31.167 4.48 31.19 4.677 ;
      RECT 31.081 4.481 31.167 4.675 ;
      RECT 30.995 4.482 31.081 4.672 ;
      RECT 30.971 4.483 30.995 4.67 ;
      RECT 30.885 4.485 30.971 4.667 ;
      RECT 30.8 4.487 30.885 4.668 ;
      RECT 30.743 4.488 30.8 4.674 ;
      RECT 30.657 4.49 30.743 4.684 ;
      RECT 30.571 4.493 30.657 4.697 ;
      RECT 30.485 4.495 30.571 4.709 ;
      RECT 30.471 4.496 30.485 4.716 ;
      RECT 30.385 4.497 30.471 4.724 ;
      RECT 30.345 4.499 30.385 4.733 ;
      RECT 30.336 4.5 30.345 4.736 ;
      RECT 30.25 4.508 30.336 4.742 ;
      RECT 30.23 4.517 30.25 4.75 ;
      RECT 30.145 4.532 30.23 4.758 ;
      RECT 30.085 4.555 30.145 4.769 ;
      RECT 30.075 4.567 30.085 4.774 ;
      RECT 30.035 4.577 30.075 4.778 ;
      RECT 29.98 4.594 30.035 4.786 ;
      RECT 29.975 4.604 29.98 4.79 ;
      RECT 31.041 3.735 31.1 4.132 ;
      RECT 30.955 3.735 31.16 4.123 ;
      RECT 30.95 3.765 31.16 4.118 ;
      RECT 30.916 3.765 31.16 4.116 ;
      RECT 30.83 3.765 31.16 4.11 ;
      RECT 30.785 3.765 31.18 4.088 ;
      RECT 30.785 3.765 31.2 4.043 ;
      RECT 30.745 3.765 31.2 4.033 ;
      RECT 30.955 3.735 31.235 4.015 ;
      RECT 30.69 3.735 30.95 3.995 ;
      RECT 29.875 3.215 30.135 3.475 ;
      RECT 29.955 3.175 30.235 3.455 ;
      RECT 24.325 8.505 24.645 8.83 ;
      RECT 24.355 7.98 24.525 8.83 ;
      RECT 24.355 7.98 24.53 8.33 ;
      RECT 24.355 7.98 25.33 8.155 ;
      RECT 25.155 3.26 25.33 8.155 ;
      RECT 25.1 3.26 25.45 3.61 ;
      RECT 25.125 8.94 25.45 9.265 ;
      RECT 24.01 9.03 25.45 9.2 ;
      RECT 24.01 3.69 24.17 9.2 ;
      RECT 24.325 3.66 24.645 3.98 ;
      RECT 24.01 3.69 24.645 3.86 ;
      RECT 12.735 4.295 13.015 4.575 ;
      RECT 12.705 4.295 13.015 4.56 ;
      RECT 12.7 4.295 13.015 4.558 ;
      RECT 12.695 2.625 12.865 4.552 ;
      RECT 12.69 4.262 12.96 4.545 ;
      RECT 12.685 4.295 13.015 4.538 ;
      RECT 12.655 4.265 12.96 4.525 ;
      RECT 12.655 4.292 12.98 4.525 ;
      RECT 12.655 4.282 12.975 4.525 ;
      RECT 12.655 4.267 12.97 4.525 ;
      RECT 12.695 4.257 12.96 4.552 ;
      RECT 12.695 4.252 12.95 4.552 ;
      RECT 12.695 4.251 12.935 4.552 ;
      RECT 22.665 2.635 23.015 2.985 ;
      RECT 22.66 2.635 23.015 2.89 ;
      RECT 12.695 2.625 22.905 2.795 ;
      RECT 22.34 4.145 22.71 4.515 ;
      RECT 22.425 3.53 22.595 4.515 ;
      RECT 18.445 3.75 18.68 4.01 ;
      RECT 21.59 3.53 21.755 3.79 ;
      RECT 21.495 3.52 21.51 3.79 ;
      RECT 21.59 3.53 22.595 3.71 ;
      RECT 20.095 3.09 20.135 3.23 ;
      RECT 21.51 3.525 21.59 3.79 ;
      RECT 21.455 3.52 21.495 3.756 ;
      RECT 21.441 3.52 21.455 3.756 ;
      RECT 21.355 3.525 21.441 3.758 ;
      RECT 21.31 3.532 21.355 3.76 ;
      RECT 21.28 3.532 21.31 3.762 ;
      RECT 21.255 3.527 21.28 3.764 ;
      RECT 21.225 3.523 21.255 3.773 ;
      RECT 21.215 3.52 21.225 3.785 ;
      RECT 21.21 3.52 21.215 3.793 ;
      RECT 21.205 3.52 21.21 3.798 ;
      RECT 21.195 3.519 21.205 3.808 ;
      RECT 21.19 3.518 21.195 3.818 ;
      RECT 21.175 3.517 21.19 3.823 ;
      RECT 21.147 3.514 21.175 3.85 ;
      RECT 21.061 3.506 21.147 3.85 ;
      RECT 20.975 3.495 21.061 3.85 ;
      RECT 20.935 3.48 20.975 3.85 ;
      RECT 20.895 3.454 20.935 3.85 ;
      RECT 20.89 3.436 20.895 3.662 ;
      RECT 20.88 3.432 20.89 3.652 ;
      RECT 20.865 3.422 20.88 3.639 ;
      RECT 20.845 3.406 20.865 3.624 ;
      RECT 20.83 3.391 20.845 3.609 ;
      RECT 20.82 3.38 20.83 3.599 ;
      RECT 20.795 3.364 20.82 3.588 ;
      RECT 20.79 3.351 20.795 3.578 ;
      RECT 20.785 3.347 20.79 3.573 ;
      RECT 20.73 3.333 20.785 3.551 ;
      RECT 20.691 3.314 20.73 3.515 ;
      RECT 20.605 3.288 20.691 3.468 ;
      RECT 20.601 3.27 20.605 3.434 ;
      RECT 20.515 3.251 20.601 3.412 ;
      RECT 20.51 3.233 20.515 3.39 ;
      RECT 20.505 3.231 20.51 3.388 ;
      RECT 20.495 3.23 20.505 3.383 ;
      RECT 20.435 3.217 20.495 3.369 ;
      RECT 20.39 3.195 20.435 3.348 ;
      RECT 20.33 3.172 20.39 3.327 ;
      RECT 20.266 3.147 20.33 3.302 ;
      RECT 20.18 3.117 20.266 3.271 ;
      RECT 20.165 3.097 20.18 3.25 ;
      RECT 20.135 3.092 20.165 3.241 ;
      RECT 20.082 3.09 20.095 3.23 ;
      RECT 19.996 3.09 20.082 3.232 ;
      RECT 19.91 3.09 19.996 3.234 ;
      RECT 19.89 3.09 19.91 3.238 ;
      RECT 19.845 3.092 19.89 3.249 ;
      RECT 19.805 3.102 19.845 3.265 ;
      RECT 19.801 3.111 19.805 3.273 ;
      RECT 19.715 3.131 19.801 3.289 ;
      RECT 19.705 3.15 19.715 3.307 ;
      RECT 19.7 3.152 19.705 3.31 ;
      RECT 19.69 3.156 19.7 3.313 ;
      RECT 19.67 3.161 19.69 3.323 ;
      RECT 19.64 3.171 19.67 3.343 ;
      RECT 19.635 3.178 19.64 3.357 ;
      RECT 19.625 3.182 19.635 3.364 ;
      RECT 19.61 3.19 19.625 3.375 ;
      RECT 19.6 3.2 19.61 3.386 ;
      RECT 19.59 3.207 19.6 3.394 ;
      RECT 19.565 3.22 19.59 3.409 ;
      RECT 19.501 3.256 19.565 3.448 ;
      RECT 19.415 3.319 19.501 3.512 ;
      RECT 19.38 3.37 19.415 3.565 ;
      RECT 19.375 3.387 19.38 3.582 ;
      RECT 19.36 3.396 19.375 3.589 ;
      RECT 19.34 3.411 19.36 3.603 ;
      RECT 19.335 3.422 19.34 3.613 ;
      RECT 19.315 3.435 19.335 3.623 ;
      RECT 19.31 3.445 19.315 3.633 ;
      RECT 19.295 3.45 19.31 3.642 ;
      RECT 19.285 3.46 19.295 3.653 ;
      RECT 19.255 3.477 19.285 3.67 ;
      RECT 19.245 3.495 19.255 3.688 ;
      RECT 19.23 3.506 19.245 3.699 ;
      RECT 19.19 3.53 19.23 3.715 ;
      RECT 19.155 3.564 19.19 3.732 ;
      RECT 19.125 3.587 19.155 3.744 ;
      RECT 19.11 3.597 19.125 3.753 ;
      RECT 19.07 3.607 19.11 3.764 ;
      RECT 19.05 3.618 19.07 3.776 ;
      RECT 19.045 3.622 19.05 3.783 ;
      RECT 19.03 3.626 19.045 3.788 ;
      RECT 19.02 3.631 19.03 3.793 ;
      RECT 19.015 3.634 19.02 3.796 ;
      RECT 18.985 3.64 19.015 3.803 ;
      RECT 18.95 3.65 18.985 3.817 ;
      RECT 18.89 3.665 18.95 3.837 ;
      RECT 18.835 3.685 18.89 3.861 ;
      RECT 18.806 3.7 18.835 3.879 ;
      RECT 18.72 3.72 18.806 3.904 ;
      RECT 18.715 3.735 18.72 3.924 ;
      RECT 18.705 3.738 18.715 3.925 ;
      RECT 18.68 3.745 18.705 4.01 ;
      RECT 21.375 4.238 21.655 4.575 ;
      RECT 21.375 4.248 21.66 4.533 ;
      RECT 21.375 4.257 21.665 4.43 ;
      RECT 21.375 4.272 21.67 4.298 ;
      RECT 21.375 4.1 21.635 4.575 ;
      RECT 10.955 9.28 11.245 9.63 ;
      RECT 10.955 9.34 12.37 9.51 ;
      RECT 12.2 8.97 12.37 9.51 ;
      RECT 20.52 8.89 20.87 9.24 ;
      RECT 12.2 8.97 20.87 9.14 ;
      RECT 19.095 4.98 19.105 5.17 ;
      RECT 17.355 4.855 17.635 5.135 ;
      RECT 20.4 3.795 20.405 4.28 ;
      RECT 20.295 3.795 20.355 4.055 ;
      RECT 20.62 4.765 20.625 4.84 ;
      RECT 20.61 4.632 20.62 4.875 ;
      RECT 20.6 4.467 20.61 4.896 ;
      RECT 20.595 4.337 20.6 4.912 ;
      RECT 20.585 4.227 20.595 4.928 ;
      RECT 20.58 4.126 20.585 4.945 ;
      RECT 20.575 4.108 20.58 4.955 ;
      RECT 20.57 4.09 20.575 4.965 ;
      RECT 20.56 4.065 20.57 4.98 ;
      RECT 20.555 4.045 20.56 4.995 ;
      RECT 20.535 3.795 20.555 5.02 ;
      RECT 20.52 3.795 20.535 5.053 ;
      RECT 20.49 3.795 20.52 5.075 ;
      RECT 20.47 3.795 20.49 5.089 ;
      RECT 20.45 3.795 20.47 4.605 ;
      RECT 20.465 4.672 20.47 5.094 ;
      RECT 20.46 4.702 20.465 5.096 ;
      RECT 20.455 4.715 20.46 5.099 ;
      RECT 20.45 4.725 20.455 5.103 ;
      RECT 20.445 3.795 20.45 4.523 ;
      RECT 20.445 4.735 20.45 5.105 ;
      RECT 20.44 3.795 20.445 4.5 ;
      RECT 20.43 4.757 20.445 5.105 ;
      RECT 20.425 3.795 20.44 4.445 ;
      RECT 20.42 4.782 20.43 5.105 ;
      RECT 20.42 3.795 20.425 4.39 ;
      RECT 20.41 3.795 20.42 4.338 ;
      RECT 20.415 4.795 20.42 5.106 ;
      RECT 20.41 4.807 20.415 5.107 ;
      RECT 20.405 3.795 20.41 4.298 ;
      RECT 20.405 4.82 20.41 5.108 ;
      RECT 20.39 4.835 20.405 5.109 ;
      RECT 20.395 3.795 20.4 4.26 ;
      RECT 20.39 3.795 20.395 4.225 ;
      RECT 20.385 3.795 20.39 4.2 ;
      RECT 20.38 4.862 20.39 5.111 ;
      RECT 20.375 3.795 20.385 4.158 ;
      RECT 20.375 4.88 20.38 5.112 ;
      RECT 20.37 3.795 20.375 4.118 ;
      RECT 20.37 4.887 20.375 5.113 ;
      RECT 20.365 3.795 20.37 4.09 ;
      RECT 20.36 4.905 20.37 5.114 ;
      RECT 20.355 3.795 20.365 4.07 ;
      RECT 20.35 4.925 20.36 5.116 ;
      RECT 20.34 4.942 20.35 5.117 ;
      RECT 20.305 4.965 20.34 5.12 ;
      RECT 20.25 4.983 20.305 5.126 ;
      RECT 20.164 4.991 20.25 5.135 ;
      RECT 20.078 5.002 20.164 5.146 ;
      RECT 19.992 5.012 20.078 5.157 ;
      RECT 19.906 5.022 19.992 5.169 ;
      RECT 19.82 5.032 19.906 5.18 ;
      RECT 19.8 5.038 19.82 5.186 ;
      RECT 19.72 5.04 19.8 5.19 ;
      RECT 19.715 5.039 19.72 5.195 ;
      RECT 19.707 5.038 19.715 5.195 ;
      RECT 19.621 5.034 19.707 5.193 ;
      RECT 19.535 5.026 19.621 5.19 ;
      RECT 19.449 5.017 19.535 5.186 ;
      RECT 19.363 5.009 19.449 5.183 ;
      RECT 19.277 5.001 19.363 5.179 ;
      RECT 19.191 4.992 19.277 5.176 ;
      RECT 19.105 4.984 19.191 5.172 ;
      RECT 19.05 4.977 19.095 5.17 ;
      RECT 18.965 4.97 19.05 5.168 ;
      RECT 18.891 4.962 18.965 5.164 ;
      RECT 18.805 4.954 18.891 5.161 ;
      RECT 18.802 4.95 18.805 5.159 ;
      RECT 18.716 4.946 18.802 5.158 ;
      RECT 18.63 4.938 18.716 5.155 ;
      RECT 18.545 4.933 18.63 5.152 ;
      RECT 18.459 4.93 18.545 5.149 ;
      RECT 18.373 4.928 18.459 5.146 ;
      RECT 18.287 4.925 18.373 5.143 ;
      RECT 18.201 4.922 18.287 5.14 ;
      RECT 18.115 4.919 18.201 5.137 ;
      RECT 18.039 4.917 18.115 5.134 ;
      RECT 17.953 4.914 18.039 5.131 ;
      RECT 17.867 4.911 17.953 5.129 ;
      RECT 17.781 4.909 17.867 5.126 ;
      RECT 17.695 4.906 17.781 5.123 ;
      RECT 17.635 4.897 17.695 5.121 ;
      RECT 20.145 4.515 20.22 4.775 ;
      RECT 20.125 4.495 20.13 4.775 ;
      RECT 19.445 4.28 19.55 4.575 ;
      RECT 13.89 4.255 13.96 4.515 ;
      RECT 19.785 4.13 19.79 4.501 ;
      RECT 19.775 4.185 19.78 4.501 ;
      RECT 20.08 3.355 20.14 3.615 ;
      RECT 20.135 4.51 20.145 4.775 ;
      RECT 20.13 4.5 20.135 4.775 ;
      RECT 20.05 4.447 20.125 4.775 ;
      RECT 20.075 3.355 20.08 3.635 ;
      RECT 20.065 3.355 20.075 3.655 ;
      RECT 20.05 3.355 20.065 3.685 ;
      RECT 20.035 3.355 20.05 3.728 ;
      RECT 20.03 4.39 20.05 4.775 ;
      RECT 20.02 3.355 20.035 3.765 ;
      RECT 20.015 4.37 20.03 4.775 ;
      RECT 20.015 3.355 20.02 3.788 ;
      RECT 20.005 3.355 20.015 3.813 ;
      RECT 19.975 4.337 20.015 4.775 ;
      RECT 19.98 3.355 20.005 3.863 ;
      RECT 19.975 3.355 19.98 3.918 ;
      RECT 19.97 3.355 19.975 3.96 ;
      RECT 19.96 4.3 19.975 4.775 ;
      RECT 19.965 3.355 19.97 4.003 ;
      RECT 19.96 3.355 19.965 4.068 ;
      RECT 19.955 3.355 19.96 4.09 ;
      RECT 19.955 4.288 19.96 4.64 ;
      RECT 19.95 3.355 19.955 4.158 ;
      RECT 19.95 4.28 19.955 4.623 ;
      RECT 19.945 3.355 19.95 4.203 ;
      RECT 19.94 4.262 19.95 4.6 ;
      RECT 19.94 3.355 19.945 4.24 ;
      RECT 19.93 3.355 19.94 4.58 ;
      RECT 19.925 3.355 19.93 4.563 ;
      RECT 19.92 3.355 19.925 4.548 ;
      RECT 19.915 3.355 19.92 4.533 ;
      RECT 19.895 3.355 19.915 4.523 ;
      RECT 19.89 3.355 19.895 4.513 ;
      RECT 19.88 3.355 19.89 4.509 ;
      RECT 19.875 3.632 19.88 4.508 ;
      RECT 19.87 3.655 19.875 4.507 ;
      RECT 19.865 3.685 19.87 4.506 ;
      RECT 19.86 3.712 19.865 4.505 ;
      RECT 19.855 3.74 19.86 4.505 ;
      RECT 19.85 3.767 19.855 4.505 ;
      RECT 19.845 3.787 19.85 4.505 ;
      RECT 19.84 3.815 19.845 4.505 ;
      RECT 19.83 3.857 19.84 4.505 ;
      RECT 19.82 3.902 19.83 4.504 ;
      RECT 19.815 3.955 19.82 4.503 ;
      RECT 19.81 3.987 19.815 4.502 ;
      RECT 19.805 4.007 19.81 4.501 ;
      RECT 19.8 4.045 19.805 4.501 ;
      RECT 19.795 4.067 19.8 4.501 ;
      RECT 19.79 4.092 19.795 4.501 ;
      RECT 19.78 4.157 19.785 4.501 ;
      RECT 19.765 4.217 19.775 4.501 ;
      RECT 19.75 4.227 19.765 4.501 ;
      RECT 19.73 4.237 19.75 4.501 ;
      RECT 19.7 4.242 19.73 4.498 ;
      RECT 19.64 4.252 19.7 4.495 ;
      RECT 19.62 4.261 19.64 4.5 ;
      RECT 19.595 4.267 19.62 4.513 ;
      RECT 19.575 4.272 19.595 4.528 ;
      RECT 19.55 4.277 19.575 4.575 ;
      RECT 19.421 4.279 19.445 4.575 ;
      RECT 19.335 4.274 19.421 4.575 ;
      RECT 19.295 4.271 19.335 4.575 ;
      RECT 19.245 4.273 19.295 4.555 ;
      RECT 19.215 4.277 19.245 4.555 ;
      RECT 19.136 4.287 19.215 4.555 ;
      RECT 19.05 4.302 19.136 4.556 ;
      RECT 19 4.312 19.05 4.557 ;
      RECT 18.992 4.315 19 4.557 ;
      RECT 18.906 4.317 18.992 4.558 ;
      RECT 18.82 4.321 18.906 4.558 ;
      RECT 18.734 4.325 18.82 4.559 ;
      RECT 18.648 4.328 18.734 4.56 ;
      RECT 18.562 4.332 18.648 4.56 ;
      RECT 18.476 4.336 18.562 4.561 ;
      RECT 18.39 4.339 18.476 4.562 ;
      RECT 18.304 4.343 18.39 4.562 ;
      RECT 18.218 4.347 18.304 4.563 ;
      RECT 18.132 4.351 18.218 4.564 ;
      RECT 18.046 4.354 18.132 4.564 ;
      RECT 17.96 4.358 18.046 4.565 ;
      RECT 17.93 4.36 17.96 4.565 ;
      RECT 17.844 4.363 17.93 4.566 ;
      RECT 17.758 4.367 17.844 4.567 ;
      RECT 17.672 4.371 17.758 4.568 ;
      RECT 17.586 4.374 17.672 4.568 ;
      RECT 17.5 4.378 17.586 4.569 ;
      RECT 17.465 4.383 17.5 4.57 ;
      RECT 17.41 4.393 17.465 4.577 ;
      RECT 17.385 4.405 17.41 4.587 ;
      RECT 17.35 4.418 17.385 4.595 ;
      RECT 17.31 4.435 17.35 4.618 ;
      RECT 17.29 4.448 17.31 4.645 ;
      RECT 17.26 4.46 17.29 4.673 ;
      RECT 17.255 4.468 17.26 4.693 ;
      RECT 17.25 4.471 17.255 4.703 ;
      RECT 17.2 4.483 17.25 4.737 ;
      RECT 17.19 4.498 17.2 4.77 ;
      RECT 17.18 4.504 17.19 4.783 ;
      RECT 17.17 4.511 17.18 4.795 ;
      RECT 17.145 4.524 17.17 4.813 ;
      RECT 17.13 4.539 17.145 4.835 ;
      RECT 17.12 4.547 17.13 4.851 ;
      RECT 17.105 4.556 17.12 4.866 ;
      RECT 17.095 4.566 17.105 4.88 ;
      RECT 17.076 4.579 17.095 4.897 ;
      RECT 16.99 4.624 17.076 4.962 ;
      RECT 16.975 4.669 16.99 5.02 ;
      RECT 16.97 4.678 16.975 5.033 ;
      RECT 16.96 4.685 16.97 5.038 ;
      RECT 16.955 4.69 16.96 5.042 ;
      RECT 16.935 4.7 16.955 5.049 ;
      RECT 16.91 4.72 16.935 5.063 ;
      RECT 16.875 4.745 16.91 5.083 ;
      RECT 16.86 4.768 16.875 5.098 ;
      RECT 16.85 4.778 16.86 5.103 ;
      RECT 16.84 4.786 16.85 5.11 ;
      RECT 16.83 4.795 16.84 5.116 ;
      RECT 16.81 4.807 16.83 5.118 ;
      RECT 16.8 4.82 16.81 5.12 ;
      RECT 16.775 4.835 16.8 5.123 ;
      RECT 16.755 4.852 16.775 5.127 ;
      RECT 16.715 4.88 16.755 5.133 ;
      RECT 16.65 4.927 16.715 5.142 ;
      RECT 16.635 4.96 16.65 5.15 ;
      RECT 16.63 4.967 16.635 5.152 ;
      RECT 16.58 4.992 16.63 5.157 ;
      RECT 16.565 5.016 16.58 5.164 ;
      RECT 16.515 5.021 16.565 5.165 ;
      RECT 16.429 5.025 16.515 5.165 ;
      RECT 16.343 5.025 16.429 5.165 ;
      RECT 16.257 5.025 16.343 5.166 ;
      RECT 16.171 5.025 16.257 5.166 ;
      RECT 16.085 5.025 16.171 5.166 ;
      RECT 16.019 5.025 16.085 5.166 ;
      RECT 15.933 5.025 16.019 5.167 ;
      RECT 15.847 5.025 15.933 5.167 ;
      RECT 15.761 5.026 15.847 5.168 ;
      RECT 15.675 5.026 15.761 5.168 ;
      RECT 15.589 5.026 15.675 5.168 ;
      RECT 15.503 5.026 15.589 5.169 ;
      RECT 15.417 5.026 15.503 5.169 ;
      RECT 15.331 5.027 15.417 5.17 ;
      RECT 15.245 5.027 15.331 5.17 ;
      RECT 15.225 5.027 15.245 5.17 ;
      RECT 15.139 5.027 15.225 5.17 ;
      RECT 15.053 5.027 15.139 5.17 ;
      RECT 14.967 5.028 15.053 5.17 ;
      RECT 14.881 5.028 14.967 5.17 ;
      RECT 14.795 5.028 14.881 5.17 ;
      RECT 14.709 5.029 14.795 5.17 ;
      RECT 14.623 5.029 14.709 5.17 ;
      RECT 14.537 5.029 14.623 5.17 ;
      RECT 14.451 5.029 14.537 5.17 ;
      RECT 14.365 5.03 14.451 5.17 ;
      RECT 14.315 5.027 14.365 5.17 ;
      RECT 14.305 5.025 14.315 5.169 ;
      RECT 14.301 5.025 14.305 5.168 ;
      RECT 14.215 5.02 14.301 5.163 ;
      RECT 14.193 5.013 14.215 5.157 ;
      RECT 14.107 5.004 14.193 5.151 ;
      RECT 14.021 4.991 14.107 5.142 ;
      RECT 13.935 4.977 14.021 5.132 ;
      RECT 13.89 4.967 13.935 5.125 ;
      RECT 13.87 4.255 13.89 4.533 ;
      RECT 13.87 4.96 13.89 5.121 ;
      RECT 13.84 4.255 13.87 4.555 ;
      RECT 13.83 4.927 13.87 5.118 ;
      RECT 13.825 4.255 13.84 4.575 ;
      RECT 13.825 4.892 13.83 5.116 ;
      RECT 13.82 4.255 13.825 4.7 ;
      RECT 13.82 4.852 13.825 5.116 ;
      RECT 13.81 4.255 13.82 5.116 ;
      RECT 13.735 4.255 13.81 5.11 ;
      RECT 13.705 4.255 13.735 5.1 ;
      RECT 13.7 4.255 13.705 5.092 ;
      RECT 13.695 4.297 13.7 5.085 ;
      RECT 13.685 4.366 13.695 5.076 ;
      RECT 13.68 4.436 13.685 5.028 ;
      RECT 13.675 4.5 13.68 4.925 ;
      RECT 13.67 4.535 13.675 4.88 ;
      RECT 13.668 4.572 13.67 4.772 ;
      RECT 13.665 4.58 13.668 4.765 ;
      RECT 13.66 4.645 13.665 4.708 ;
      RECT 17.735 3.735 18.015 4.015 ;
      RECT 17.725 3.735 18.015 3.878 ;
      RECT 17.68 3.6 17.94 3.86 ;
      RECT 17.68 3.715 17.995 3.86 ;
      RECT 17.68 3.685 17.99 3.86 ;
      RECT 17.68 3.672 17.98 3.86 ;
      RECT 17.68 3.662 17.975 3.86 ;
      RECT 13.655 3.645 13.915 3.905 ;
      RECT 17.425 3.195 17.685 3.455 ;
      RECT 17.415 3.22 17.685 3.415 ;
      RECT 17.41 3.22 17.415 3.414 ;
      RECT 17.34 3.215 17.41 3.406 ;
      RECT 17.255 3.202 17.34 3.389 ;
      RECT 17.251 3.194 17.255 3.379 ;
      RECT 17.165 3.187 17.251 3.369 ;
      RECT 17.156 3.179 17.165 3.359 ;
      RECT 17.07 3.172 17.156 3.347 ;
      RECT 17.05 3.163 17.07 3.333 ;
      RECT 16.995 3.158 17.05 3.325 ;
      RECT 16.985 3.152 16.995 3.319 ;
      RECT 16.965 3.15 16.985 3.315 ;
      RECT 16.957 3.149 16.965 3.311 ;
      RECT 16.871 3.141 16.957 3.3 ;
      RECT 16.785 3.127 16.871 3.28 ;
      RECT 16.725 3.115 16.785 3.265 ;
      RECT 16.715 3.11 16.725 3.26 ;
      RECT 16.665 3.11 16.715 3.262 ;
      RECT 16.618 3.112 16.665 3.266 ;
      RECT 16.532 3.119 16.618 3.271 ;
      RECT 16.446 3.127 16.532 3.277 ;
      RECT 16.36 3.136 16.446 3.283 ;
      RECT 16.301 3.142 16.36 3.288 ;
      RECT 16.215 3.147 16.301 3.294 ;
      RECT 16.14 3.152 16.215 3.3 ;
      RECT 16.101 3.154 16.14 3.305 ;
      RECT 16.015 3.151 16.101 3.31 ;
      RECT 15.93 3.149 16.015 3.317 ;
      RECT 15.898 3.148 15.93 3.32 ;
      RECT 15.812 3.147 15.898 3.321 ;
      RECT 15.726 3.146 15.812 3.322 ;
      RECT 15.64 3.145 15.726 3.322 ;
      RECT 15.554 3.144 15.64 3.323 ;
      RECT 15.468 3.143 15.554 3.324 ;
      RECT 15.382 3.142 15.468 3.325 ;
      RECT 15.296 3.141 15.382 3.325 ;
      RECT 15.21 3.14 15.296 3.326 ;
      RECT 15.16 3.14 15.21 3.327 ;
      RECT 15.146 3.141 15.16 3.327 ;
      RECT 15.06 3.148 15.146 3.328 ;
      RECT 14.986 3.159 15.06 3.329 ;
      RECT 14.9 3.168 14.986 3.33 ;
      RECT 14.865 3.175 14.9 3.345 ;
      RECT 14.84 3.178 14.865 3.375 ;
      RECT 14.815 3.187 14.84 3.404 ;
      RECT 14.805 3.198 14.815 3.424 ;
      RECT 14.795 3.206 14.805 3.438 ;
      RECT 14.79 3.212 14.795 3.448 ;
      RECT 14.765 3.229 14.79 3.465 ;
      RECT 14.75 3.251 14.765 3.493 ;
      RECT 14.72 3.277 14.75 3.523 ;
      RECT 14.7 3.306 14.72 3.553 ;
      RECT 14.695 3.321 14.7 3.57 ;
      RECT 14.675 3.336 14.695 3.585 ;
      RECT 14.665 3.354 14.675 3.603 ;
      RECT 14.655 3.365 14.665 3.618 ;
      RECT 14.605 3.397 14.655 3.644 ;
      RECT 14.6 3.427 14.605 3.664 ;
      RECT 14.59 3.44 14.6 3.67 ;
      RECT 14.581 3.45 14.59 3.678 ;
      RECT 14.57 3.461 14.581 3.686 ;
      RECT 14.565 3.471 14.57 3.692 ;
      RECT 14.55 3.492 14.565 3.699 ;
      RECT 14.535 3.522 14.55 3.707 ;
      RECT 14.5 3.552 14.535 3.713 ;
      RECT 14.475 3.57 14.5 3.72 ;
      RECT 14.425 3.578 14.475 3.729 ;
      RECT 14.4 3.583 14.425 3.738 ;
      RECT 14.345 3.589 14.4 3.748 ;
      RECT 14.34 3.594 14.345 3.756 ;
      RECT 14.326 3.597 14.34 3.758 ;
      RECT 14.24 3.609 14.326 3.77 ;
      RECT 14.23 3.621 14.24 3.783 ;
      RECT 14.145 3.634 14.23 3.795 ;
      RECT 14.101 3.651 14.145 3.809 ;
      RECT 14.015 3.668 14.101 3.825 ;
      RECT 13.985 3.682 14.015 3.839 ;
      RECT 13.975 3.687 13.985 3.844 ;
      RECT 13.915 3.69 13.975 3.853 ;
      RECT 16.805 3.96 17.065 4.22 ;
      RECT 16.805 3.96 17.085 4.073 ;
      RECT 16.805 3.96 17.11 4.04 ;
      RECT 16.805 3.96 17.115 4.02 ;
      RECT 16.855 3.735 17.135 4.015 ;
      RECT 16.41 4.47 16.67 4.73 ;
      RECT 16.4 4.327 16.595 4.668 ;
      RECT 16.395 4.435 16.61 4.66 ;
      RECT 16.39 4.485 16.67 4.65 ;
      RECT 16.38 4.562 16.67 4.635 ;
      RECT 16.4 4.41 16.61 4.668 ;
      RECT 16.41 4.285 16.595 4.73 ;
      RECT 16.41 4.18 16.575 4.73 ;
      RECT 16.42 4.167 16.575 4.73 ;
      RECT 16.42 4.125 16.565 4.73 ;
      RECT 16.425 4.05 16.565 4.73 ;
      RECT 16.455 3.7 16.565 4.73 ;
      RECT 16.46 3.43 16.585 4.053 ;
      RECT 16.43 4.005 16.585 4.053 ;
      RECT 16.445 3.807 16.565 4.73 ;
      RECT 16.435 3.917 16.585 4.053 ;
      RECT 16.46 3.43 16.6 3.91 ;
      RECT 16.46 3.43 16.62 3.785 ;
      RECT 16.425 3.43 16.685 3.69 ;
      RECT 15.895 3.735 16.175 4.015 ;
      RECT 15.88 3.735 16.175 3.995 ;
      RECT 13.935 4.6 14.195 4.86 ;
      RECT 15.72 4.455 15.98 4.715 ;
      RECT 15.7 4.475 15.98 4.69 ;
      RECT 15.657 4.475 15.7 4.689 ;
      RECT 15.571 4.476 15.657 4.686 ;
      RECT 15.485 4.477 15.571 4.682 ;
      RECT 15.41 4.479 15.485 4.679 ;
      RECT 15.387 4.48 15.41 4.677 ;
      RECT 15.301 4.481 15.387 4.675 ;
      RECT 15.215 4.482 15.301 4.672 ;
      RECT 15.191 4.483 15.215 4.67 ;
      RECT 15.105 4.485 15.191 4.667 ;
      RECT 15.02 4.487 15.105 4.668 ;
      RECT 14.963 4.488 15.02 4.674 ;
      RECT 14.877 4.49 14.963 4.684 ;
      RECT 14.791 4.493 14.877 4.697 ;
      RECT 14.705 4.495 14.791 4.709 ;
      RECT 14.691 4.496 14.705 4.716 ;
      RECT 14.605 4.497 14.691 4.724 ;
      RECT 14.565 4.499 14.605 4.733 ;
      RECT 14.556 4.5 14.565 4.736 ;
      RECT 14.47 4.508 14.556 4.742 ;
      RECT 14.45 4.517 14.47 4.75 ;
      RECT 14.365 4.532 14.45 4.758 ;
      RECT 14.305 4.555 14.365 4.769 ;
      RECT 14.295 4.567 14.305 4.774 ;
      RECT 14.255 4.577 14.295 4.778 ;
      RECT 14.2 4.594 14.255 4.786 ;
      RECT 14.195 4.604 14.2 4.79 ;
      RECT 15.261 3.735 15.32 4.132 ;
      RECT 15.175 3.735 15.38 4.123 ;
      RECT 15.17 3.765 15.38 4.118 ;
      RECT 15.136 3.765 15.38 4.116 ;
      RECT 15.05 3.765 15.38 4.11 ;
      RECT 15.005 3.765 15.4 4.088 ;
      RECT 15.005 3.765 15.42 4.043 ;
      RECT 14.965 3.765 15.42 4.033 ;
      RECT 15.175 3.735 15.455 4.015 ;
      RECT 14.91 3.735 15.17 3.995 ;
      RECT 14.095 3.215 14.355 3.475 ;
      RECT 14.175 3.175 14.455 3.455 ;
      RECT 9.605 10.785 9.985 11.165 ;
      RECT 9.65 0 9.79 11.165 ;
      RECT 9.605 0 9.985 0.38 ;
      RECT 84.685 2.11 85.055 2.48 ;
      RECT 82.975 9.325 83.345 9.695 ;
      RECT 68.9 2.11 69.27 2.48 ;
      RECT 67.19 9.325 67.56 9.695 ;
      RECT 53.115 2.11 53.485 2.48 ;
      RECT 51.405 9.325 51.775 9.695 ;
      RECT 37.34 2.11 37.71 2.48 ;
      RECT 35.63 9.325 36 9.695 ;
      RECT 21.56 2.11 21.93 2.48 ;
      RECT 19.85 9.325 20.22 9.695 ;
    LAYER via1 ;
      RECT 90.71 9.66 90.86 9.81 ;
      RECT 88.34 9.025 88.49 9.175 ;
      RECT 88.325 3.36 88.475 3.51 ;
      RECT 87.535 3.745 87.685 3.895 ;
      RECT 87.535 8.61 87.685 8.76 ;
      RECT 85.89 2.735 86.04 2.885 ;
      RECT 85.575 4.255 85.725 4.405 ;
      RECT 84.795 2.22 84.945 2.37 ;
      RECT 84.675 3.585 84.825 3.735 ;
      RECT 84.555 4.155 84.705 4.305 ;
      RECT 83.725 8.995 83.875 9.145 ;
      RECT 83.475 3.85 83.625 4 ;
      RECT 83.14 4.57 83.29 4.72 ;
      RECT 83.085 9.435 83.235 9.585 ;
      RECT 83.06 3.41 83.21 3.56 ;
      RECT 81.625 3.805 81.775 3.955 ;
      RECT 80.86 3.655 81.01 3.805 ;
      RECT 80.605 3.25 80.755 3.4 ;
      RECT 79.985 4.015 80.135 4.165 ;
      RECT 79.605 3.485 79.755 3.635 ;
      RECT 79.59 4.525 79.74 4.675 ;
      RECT 79.06 3.79 79.21 3.94 ;
      RECT 78.9 4.51 79.05 4.66 ;
      RECT 78.09 3.79 78.24 3.94 ;
      RECT 77.275 3.27 77.425 3.42 ;
      RECT 77.115 4.655 77.265 4.805 ;
      RECT 76.88 4.31 77.03 4.46 ;
      RECT 76.835 3.7 76.985 3.85 ;
      RECT 75.835 4.32 75.985 4.47 ;
      RECT 74.9 9.04 75.05 9.19 ;
      RECT 72.555 9.025 72.705 9.175 ;
      RECT 72.54 3.36 72.69 3.51 ;
      RECT 71.75 3.745 71.9 3.895 ;
      RECT 71.75 8.61 71.9 8.76 ;
      RECT 70.105 2.735 70.255 2.885 ;
      RECT 69.79 4.255 69.94 4.405 ;
      RECT 69.01 2.22 69.16 2.37 ;
      RECT 68.89 3.585 69.04 3.735 ;
      RECT 68.77 4.155 68.92 4.305 ;
      RECT 67.94 8.995 68.09 9.145 ;
      RECT 67.69 3.85 67.84 4 ;
      RECT 67.355 4.57 67.505 4.72 ;
      RECT 67.3 9.435 67.45 9.585 ;
      RECT 67.275 3.41 67.425 3.56 ;
      RECT 65.84 3.805 65.99 3.955 ;
      RECT 65.075 3.655 65.225 3.805 ;
      RECT 64.82 3.25 64.97 3.4 ;
      RECT 64.2 4.015 64.35 4.165 ;
      RECT 63.82 3.485 63.97 3.635 ;
      RECT 63.805 4.525 63.955 4.675 ;
      RECT 63.275 3.79 63.425 3.94 ;
      RECT 63.115 4.51 63.265 4.66 ;
      RECT 62.305 3.79 62.455 3.94 ;
      RECT 61.49 3.27 61.64 3.42 ;
      RECT 61.33 4.655 61.48 4.805 ;
      RECT 61.095 4.31 61.245 4.46 ;
      RECT 61.05 3.7 61.2 3.85 ;
      RECT 60.05 4.32 60.2 4.47 ;
      RECT 59.115 9.04 59.265 9.19 ;
      RECT 56.77 9.025 56.92 9.175 ;
      RECT 56.755 3.36 56.905 3.51 ;
      RECT 55.965 3.745 56.115 3.895 ;
      RECT 55.965 8.61 56.115 8.76 ;
      RECT 54.32 2.735 54.47 2.885 ;
      RECT 54.005 4.255 54.155 4.405 ;
      RECT 53.225 2.22 53.375 2.37 ;
      RECT 53.105 3.585 53.255 3.735 ;
      RECT 52.985 4.155 53.135 4.305 ;
      RECT 52.21 9 52.36 9.15 ;
      RECT 51.905 3.85 52.055 4 ;
      RECT 51.57 4.57 51.72 4.72 ;
      RECT 51.515 9.435 51.665 9.585 ;
      RECT 51.49 3.41 51.64 3.56 ;
      RECT 50.055 3.805 50.205 3.955 ;
      RECT 49.29 3.655 49.44 3.805 ;
      RECT 49.035 3.25 49.185 3.4 ;
      RECT 48.415 4.015 48.565 4.165 ;
      RECT 48.035 3.485 48.185 3.635 ;
      RECT 48.02 4.525 48.17 4.675 ;
      RECT 47.49 3.79 47.64 3.94 ;
      RECT 47.33 4.51 47.48 4.66 ;
      RECT 46.52 3.79 46.67 3.94 ;
      RECT 45.705 3.27 45.855 3.42 ;
      RECT 45.545 4.655 45.695 4.805 ;
      RECT 45.31 4.31 45.46 4.46 ;
      RECT 45.265 3.7 45.415 3.85 ;
      RECT 44.265 4.32 44.415 4.47 ;
      RECT 43.385 9.045 43.535 9.195 ;
      RECT 40.995 9.025 41.145 9.175 ;
      RECT 40.98 3.36 41.13 3.51 ;
      RECT 40.19 3.745 40.34 3.895 ;
      RECT 40.19 8.61 40.34 8.76 ;
      RECT 38.545 2.735 38.695 2.885 ;
      RECT 38.23 4.255 38.38 4.405 ;
      RECT 37.45 2.22 37.6 2.37 ;
      RECT 37.33 3.585 37.48 3.735 ;
      RECT 37.21 4.155 37.36 4.305 ;
      RECT 36.43 8.995 36.58 9.145 ;
      RECT 36.13 3.85 36.28 4 ;
      RECT 35.795 4.57 35.945 4.72 ;
      RECT 35.74 9.435 35.89 9.585 ;
      RECT 35.715 3.41 35.865 3.56 ;
      RECT 34.28 3.805 34.43 3.955 ;
      RECT 33.515 3.655 33.665 3.805 ;
      RECT 33.26 3.25 33.41 3.4 ;
      RECT 32.64 4.015 32.79 4.165 ;
      RECT 32.26 3.485 32.41 3.635 ;
      RECT 32.245 4.525 32.395 4.675 ;
      RECT 31.715 3.79 31.865 3.94 ;
      RECT 31.555 4.51 31.705 4.66 ;
      RECT 30.745 3.79 30.895 3.94 ;
      RECT 29.93 3.27 30.08 3.42 ;
      RECT 29.77 4.655 29.92 4.805 ;
      RECT 29.535 4.31 29.685 4.46 ;
      RECT 29.49 3.7 29.64 3.85 ;
      RECT 28.49 4.32 28.64 4.47 ;
      RECT 27.605 9.04 27.755 9.19 ;
      RECT 25.215 9.025 25.365 9.175 ;
      RECT 25.2 3.36 25.35 3.51 ;
      RECT 24.41 3.745 24.56 3.895 ;
      RECT 24.41 8.61 24.56 8.76 ;
      RECT 22.765 2.735 22.915 2.885 ;
      RECT 22.45 4.255 22.6 4.405 ;
      RECT 21.67 2.22 21.82 2.37 ;
      RECT 21.55 3.585 21.7 3.735 ;
      RECT 21.43 4.155 21.58 4.305 ;
      RECT 20.62 8.99 20.77 9.14 ;
      RECT 20.35 3.85 20.5 4 ;
      RECT 20.015 4.57 20.165 4.72 ;
      RECT 19.96 9.435 20.11 9.585 ;
      RECT 19.935 3.41 20.085 3.56 ;
      RECT 18.5 3.805 18.65 3.955 ;
      RECT 17.735 3.655 17.885 3.805 ;
      RECT 17.48 3.25 17.63 3.4 ;
      RECT 16.86 4.015 17.01 4.165 ;
      RECT 16.48 3.485 16.63 3.635 ;
      RECT 16.465 4.525 16.615 4.675 ;
      RECT 15.935 3.79 16.085 3.94 ;
      RECT 15.775 4.51 15.925 4.66 ;
      RECT 14.965 3.79 15.115 3.94 ;
      RECT 14.15 3.27 14.3 3.42 ;
      RECT 13.99 4.655 14.14 4.805 ;
      RECT 13.755 4.31 13.905 4.46 ;
      RECT 13.71 3.7 13.86 3.85 ;
      RECT 12.71 4.32 12.86 4.47 ;
      RECT 11.025 9.38 11.175 9.53 ;
      RECT 10.65 8.64 10.8 8.79 ;
      RECT 9.72 0.115 9.87 0.265 ;
      RECT 9.72 10.9 9.87 11.05 ;
    LAYER met1 ;
      RECT 75.585 2.555 85.245 3.035 ;
      RECT 59.8 2.555 69.46 3.035 ;
      RECT 44.015 2.555 53.675 3.035 ;
      RECT 28.24 2.555 37.9 3.035 ;
      RECT 12.46 2.555 22.12 3.035 ;
      RECT 75.585 2.555 85.3 2.885 ;
      RECT 59.8 2.555 69.515 2.885 ;
      RECT 44.015 2.555 53.73 2.885 ;
      RECT 28.24 2.555 37.955 2.885 ;
      RECT 12.46 2.555 22.175 2.885 ;
      RECT 75.7 0 85.415 2.88 ;
      RECT 59.915 0 69.63 2.88 ;
      RECT 44.13 0 53.845 2.88 ;
      RECT 28.355 0 38.07 2.88 ;
      RECT 12.575 0 22.29 2.88 ;
      RECT 9.415 0 91.185 1.6 ;
      RECT 9.41 10.86 91.185 12.46 ;
      RECT 82.27 8.6 82.44 12.46 ;
      RECT 66.485 8.6 66.655 12.46 ;
      RECT 50.7 8.6 50.87 12.46 ;
      RECT 34.925 8.6 35.095 12.46 ;
      RECT 19.145 8.6 19.315 12.46 ;
      RECT 9.41 10.85 10.22 12.46 ;
      RECT 9.62 10.83 9.97 12.46 ;
      RECT 82.64 8.57 82.93 8.8 ;
      RECT 66.855 8.57 67.145 8.8 ;
      RECT 51.07 8.57 51.36 8.8 ;
      RECT 35.295 8.57 35.585 8.8 ;
      RECT 19.515 8.57 19.805 8.8 ;
      RECT 82.27 8.6 82.93 8.77 ;
      RECT 66.485 8.6 67.145 8.77 ;
      RECT 50.7 8.6 51.36 8.77 ;
      RECT 34.925 8.6 35.585 8.77 ;
      RECT 19.145 8.6 19.805 8.77 ;
      RECT 89.045 5.425 91.025 7.035 ;
      RECT 73.26 5.425 75.24 7.035 ;
      RECT 57.475 5.425 59.455 7.035 ;
      RECT 41.7 5.425 43.68 7.035 ;
      RECT 25.92 5.425 27.9 7.035 ;
      RECT 9.415 5.43 91.18 7.03 ;
      RECT 75.585 5.275 85.245 7.03 ;
      RECT 59.8 5.275 69.46 7.03 ;
      RECT 44.015 5.275 53.675 7.03 ;
      RECT 28.24 5.275 37.9 7.03 ;
      RECT 12.46 5.275 22.12 7.03 ;
      RECT 90.575 10.055 90.865 10.285 ;
      RECT 90.635 8.575 90.805 10.285 ;
      RECT 90.61 9.56 90.96 9.91 ;
      RECT 90.575 8.575 90.865 8.805 ;
      RECT 90.17 3.69 90.275 4.26 ;
      RECT 90.17 4.025 90.495 4.255 ;
      RECT 90.17 4.055 90.665 4.225 ;
      RECT 90.17 3.69 90.36 4.255 ;
      RECT 89.585 3.655 89.875 3.885 ;
      RECT 89.585 3.69 90.36 3.86 ;
      RECT 89.645 2.175 89.815 3.885 ;
      RECT 89.585 2.175 89.875 2.405 ;
      RECT 89.585 10.055 89.875 10.285 ;
      RECT 89.645 8.575 89.815 10.285 ;
      RECT 89.585 8.575 89.875 8.805 ;
      RECT 89.585 8.61 90.435 8.77 ;
      RECT 90.27 8.205 90.435 8.77 ;
      RECT 89.585 8.605 89.98 8.77 ;
      RECT 90.205 8.205 90.495 8.435 ;
      RECT 90.205 8.235 90.665 8.405 ;
      RECT 89.215 4.025 89.505 4.255 ;
      RECT 89.215 4.055 89.675 4.225 ;
      RECT 89.28 2.95 89.445 4.255 ;
      RECT 87.795 2.92 88.085 3.15 ;
      RECT 87.795 2.95 89.445 3.12 ;
      RECT 87.855 2.18 88.025 3.15 ;
      RECT 87.795 2.18 88.085 2.41 ;
      RECT 87.795 10.05 88.085 10.28 ;
      RECT 87.855 9.31 88.025 10.28 ;
      RECT 87.855 9.405 89.445 9.575 ;
      RECT 89.275 8.205 89.445 9.575 ;
      RECT 87.795 9.31 88.085 9.54 ;
      RECT 89.215 8.205 89.505 8.435 ;
      RECT 89.215 8.235 89.675 8.405 ;
      RECT 88.225 3.26 88.575 3.61 ;
      RECT 85.89 3.32 88.575 3.49 ;
      RECT 85.89 2.635 86.06 3.49 ;
      RECT 85.79 2.635 86.14 2.985 ;
      RECT 88.25 8.94 88.575 9.265 ;
      RECT 83.625 8.895 83.975 9.245 ;
      RECT 88.225 8.94 88.575 9.17 ;
      RECT 83.445 8.94 83.975 9.17 ;
      RECT 83.275 8.97 88.575 9.14 ;
      RECT 87.45 3.66 87.77 3.98 ;
      RECT 87.42 3.66 87.77 3.89 ;
      RECT 87.25 3.69 87.77 3.86 ;
      RECT 87.45 8.54 87.77 8.83 ;
      RECT 87.42 8.57 87.77 8.8 ;
      RECT 87.25 8.6 87.77 8.77 ;
      RECT 84.085 3.76 84.27 3.97 ;
      RECT 84.075 3.765 84.285 3.963 ;
      RECT 84.075 3.765 84.371 3.94 ;
      RECT 84.075 3.765 84.43 3.915 ;
      RECT 84.075 3.765 84.485 3.895 ;
      RECT 84.075 3.765 84.495 3.883 ;
      RECT 84.075 3.765 84.69 3.822 ;
      RECT 84.075 3.765 84.72 3.805 ;
      RECT 84.075 3.765 84.74 3.795 ;
      RECT 84.62 3.53 84.88 3.79 ;
      RECT 84.605 3.62 84.62 3.837 ;
      RECT 84.14 3.752 84.88 3.79 ;
      RECT 84.591 3.631 84.605 3.843 ;
      RECT 84.18 3.745 84.88 3.79 ;
      RECT 84.505 3.671 84.591 3.862 ;
      RECT 84.43 3.732 84.88 3.79 ;
      RECT 84.5 3.707 84.505 3.879 ;
      RECT 84.485 3.717 84.88 3.79 ;
      RECT 84.495 3.712 84.5 3.881 ;
      RECT 84.79 4.217 84.795 4.309 ;
      RECT 84.785 4.195 84.79 4.326 ;
      RECT 84.78 4.185 84.785 4.338 ;
      RECT 84.77 4.176 84.78 4.348 ;
      RECT 84.765 4.171 84.77 4.356 ;
      RECT 84.76 4.03 84.765 4.359 ;
      RECT 84.726 4.03 84.76 4.37 ;
      RECT 84.64 4.03 84.726 4.405 ;
      RECT 84.56 4.03 84.64 4.453 ;
      RECT 84.531 4.03 84.56 4.477 ;
      RECT 84.445 4.03 84.531 4.483 ;
      RECT 84.44 4.214 84.445 4.488 ;
      RECT 84.405 4.225 84.44 4.491 ;
      RECT 84.38 4.24 84.405 4.495 ;
      RECT 84.366 4.249 84.38 4.497 ;
      RECT 84.28 4.276 84.366 4.503 ;
      RECT 84.215 4.317 84.28 4.512 ;
      RECT 84.2 4.337 84.215 4.517 ;
      RECT 84.17 4.347 84.2 4.52 ;
      RECT 84.165 4.357 84.17 4.523 ;
      RECT 84.135 4.362 84.165 4.525 ;
      RECT 84.115 4.367 84.135 4.529 ;
      RECT 84.03 4.37 84.115 4.536 ;
      RECT 84.015 4.367 84.03 4.542 ;
      RECT 84.005 4.364 84.015 4.544 ;
      RECT 83.985 4.361 84.005 4.546 ;
      RECT 83.965 4.357 83.985 4.547 ;
      RECT 83.95 4.353 83.965 4.549 ;
      RECT 83.94 4.35 83.95 4.55 ;
      RECT 83.9 4.344 83.94 4.548 ;
      RECT 83.89 4.339 83.9 4.546 ;
      RECT 83.875 4.336 83.89 4.542 ;
      RECT 83.85 4.331 83.875 4.535 ;
      RECT 83.8 4.322 83.85 4.523 ;
      RECT 83.73 4.308 83.8 4.505 ;
      RECT 83.672 4.293 83.73 4.487 ;
      RECT 83.586 4.276 83.672 4.467 ;
      RECT 83.5 4.255 83.586 4.442 ;
      RECT 83.45 4.24 83.5 4.423 ;
      RECT 83.446 4.234 83.45 4.415 ;
      RECT 83.36 4.224 83.446 4.402 ;
      RECT 83.325 4.209 83.36 4.385 ;
      RECT 83.31 4.202 83.325 4.378 ;
      RECT 83.25 4.19 83.31 4.366 ;
      RECT 83.23 4.177 83.25 4.354 ;
      RECT 83.19 4.168 83.23 4.346 ;
      RECT 83.185 4.16 83.19 4.339 ;
      RECT 83.105 4.15 83.185 4.325 ;
      RECT 83.09 4.137 83.105 4.31 ;
      RECT 83.085 4.135 83.09 4.308 ;
      RECT 83.006 4.123 83.085 4.295 ;
      RECT 82.92 4.098 83.006 4.27 ;
      RECT 82.905 4.067 82.92 4.255 ;
      RECT 82.89 4.042 82.905 4.251 ;
      RECT 82.875 4.035 82.89 4.247 ;
      RECT 82.7 4.04 82.705 4.243 ;
      RECT 82.695 4.045 82.7 4.238 ;
      RECT 82.705 4.035 82.875 4.245 ;
      RECT 83.42 3.795 83.525 4.055 ;
      RECT 84.235 3.32 84.24 3.545 ;
      RECT 84.365 3.32 84.42 3.53 ;
      RECT 84.42 3.325 84.43 3.523 ;
      RECT 84.326 3.32 84.365 3.533 ;
      RECT 84.24 3.32 84.326 3.54 ;
      RECT 84.22 3.325 84.235 3.546 ;
      RECT 84.21 3.365 84.22 3.548 ;
      RECT 84.18 3.375 84.21 3.55 ;
      RECT 84.175 3.38 84.18 3.552 ;
      RECT 84.15 3.385 84.175 3.554 ;
      RECT 84.135 3.39 84.15 3.556 ;
      RECT 84.12 3.392 84.135 3.558 ;
      RECT 84.115 3.397 84.12 3.56 ;
      RECT 84.065 3.405 84.115 3.563 ;
      RECT 84.04 3.414 84.065 3.568 ;
      RECT 84.03 3.421 84.04 3.573 ;
      RECT 84.025 3.424 84.03 3.577 ;
      RECT 84.005 3.427 84.025 3.586 ;
      RECT 83.975 3.435 84.005 3.606 ;
      RECT 83.946 3.448 83.975 3.628 ;
      RECT 83.86 3.482 83.946 3.672 ;
      RECT 83.855 3.508 83.86 3.71 ;
      RECT 83.85 3.512 83.855 3.719 ;
      RECT 83.815 3.525 83.85 3.752 ;
      RECT 83.805 3.539 83.815 3.79 ;
      RECT 83.8 3.543 83.805 3.803 ;
      RECT 83.795 3.547 83.8 3.808 ;
      RECT 83.785 3.555 83.795 3.82 ;
      RECT 83.78 3.562 83.785 3.835 ;
      RECT 83.755 3.575 83.78 3.86 ;
      RECT 83.715 3.604 83.755 3.915 ;
      RECT 83.7 3.629 83.715 3.97 ;
      RECT 83.69 3.64 83.7 3.993 ;
      RECT 83.685 3.647 83.69 4.005 ;
      RECT 83.68 3.651 83.685 4.013 ;
      RECT 83.625 3.679 83.68 4.055 ;
      RECT 83.605 3.715 83.625 4.055 ;
      RECT 83.59 3.73 83.605 4.055 ;
      RECT 83.535 3.762 83.59 4.055 ;
      RECT 83.525 3.792 83.535 4.055 ;
      RECT 83.135 3.407 83.32 3.645 ;
      RECT 83.12 3.409 83.33 3.64 ;
      RECT 83.005 3.355 83.265 3.615 ;
      RECT 83 3.392 83.265 3.569 ;
      RECT 82.995 3.402 83.265 3.566 ;
      RECT 82.99 3.442 83.33 3.56 ;
      RECT 82.985 3.475 83.33 3.55 ;
      RECT 82.995 3.417 83.345 3.488 ;
      RECT 83.292 4.515 83.305 5.045 ;
      RECT 83.206 4.515 83.305 5.044 ;
      RECT 83.206 4.515 83.31 5.043 ;
      RECT 83.12 4.515 83.31 5.041 ;
      RECT 83.115 4.515 83.31 5.038 ;
      RECT 83.115 4.515 83.32 5.036 ;
      RECT 83.11 4.807 83.32 5.033 ;
      RECT 83.11 4.817 83.325 5.03 ;
      RECT 83.11 4.885 83.33 5.026 ;
      RECT 83.1 4.89 83.33 5.025 ;
      RECT 83.1 4.982 83.335 5.022 ;
      RECT 83.085 4.515 83.345 4.775 ;
      RECT 83.015 10.05 83.305 10.28 ;
      RECT 83.075 9.31 83.245 10.28 ;
      RECT 82.99 9.34 83.33 9.685 ;
      RECT 83.015 9.31 83.305 9.685 ;
      RECT 82.315 3.505 82.36 5.04 ;
      RECT 82.515 3.505 82.545 3.72 ;
      RECT 80.89 3.245 81.01 3.455 ;
      RECT 80.55 3.195 80.81 3.455 ;
      RECT 80.55 3.24 80.845 3.445 ;
      RECT 82.555 3.521 82.56 3.575 ;
      RECT 82.55 3.514 82.555 3.708 ;
      RECT 82.545 3.508 82.55 3.715 ;
      RECT 82.5 3.505 82.515 3.728 ;
      RECT 82.495 3.505 82.5 3.75 ;
      RECT 82.49 3.505 82.495 3.798 ;
      RECT 82.485 3.505 82.49 3.818 ;
      RECT 82.475 3.505 82.485 3.925 ;
      RECT 82.47 3.505 82.475 3.988 ;
      RECT 82.465 3.505 82.47 4.045 ;
      RECT 82.46 3.505 82.465 4.053 ;
      RECT 82.445 3.505 82.46 4.16 ;
      RECT 82.435 3.505 82.445 4.295 ;
      RECT 82.425 3.505 82.435 4.405 ;
      RECT 82.415 3.505 82.425 4.462 ;
      RECT 82.41 3.505 82.415 4.502 ;
      RECT 82.405 3.505 82.41 4.538 ;
      RECT 82.395 3.505 82.405 4.578 ;
      RECT 82.39 3.505 82.395 4.62 ;
      RECT 82.37 3.505 82.39 4.685 ;
      RECT 82.375 4.83 82.38 5.01 ;
      RECT 82.37 4.812 82.375 5.018 ;
      RECT 82.365 3.505 82.37 4.748 ;
      RECT 82.365 4.792 82.37 5.025 ;
      RECT 82.36 3.505 82.365 5.035 ;
      RECT 82.305 3.505 82.315 3.805 ;
      RECT 82.31 4.052 82.315 5.04 ;
      RECT 82.305 4.117 82.31 5.04 ;
      RECT 82.3 3.506 82.305 3.795 ;
      RECT 82.295 4.182 82.305 5.04 ;
      RECT 82.29 3.507 82.3 3.785 ;
      RECT 82.28 4.295 82.295 5.04 ;
      RECT 82.285 3.508 82.29 3.775 ;
      RECT 82.265 3.509 82.285 3.753 ;
      RECT 82.27 4.392 82.28 5.04 ;
      RECT 82.265 4.467 82.27 5.04 ;
      RECT 82.255 3.508 82.265 3.73 ;
      RECT 82.26 4.51 82.265 5.04 ;
      RECT 82.255 4.537 82.26 5.04 ;
      RECT 82.245 3.506 82.255 3.718 ;
      RECT 82.25 4.58 82.255 5.04 ;
      RECT 82.245 4.607 82.25 5.04 ;
      RECT 82.235 3.505 82.245 3.705 ;
      RECT 82.24 4.622 82.245 5.04 ;
      RECT 82.2 4.68 82.24 5.04 ;
      RECT 82.23 3.504 82.235 3.69 ;
      RECT 82.225 3.502 82.23 3.683 ;
      RECT 82.215 3.499 82.225 3.673 ;
      RECT 82.21 3.496 82.215 3.658 ;
      RECT 82.195 3.492 82.21 3.651 ;
      RECT 82.19 4.735 82.2 5.04 ;
      RECT 82.19 3.489 82.195 3.646 ;
      RECT 82.175 3.485 82.19 3.64 ;
      RECT 82.185 4.752 82.19 5.04 ;
      RECT 82.175 4.815 82.185 5.04 ;
      RECT 82.095 3.47 82.175 3.62 ;
      RECT 82.17 4.822 82.175 5.035 ;
      RECT 82.165 4.83 82.17 5.025 ;
      RECT 82.085 3.456 82.095 3.604 ;
      RECT 82.07 3.452 82.085 3.602 ;
      RECT 82.06 3.447 82.07 3.598 ;
      RECT 82.035 3.44 82.06 3.59 ;
      RECT 82.03 3.435 82.035 3.585 ;
      RECT 82.02 3.435 82.03 3.583 ;
      RECT 82.01 3.433 82.02 3.581 ;
      RECT 81.98 3.425 82.01 3.575 ;
      RECT 81.965 3.417 81.98 3.568 ;
      RECT 81.945 3.412 81.965 3.561 ;
      RECT 81.94 3.408 81.945 3.556 ;
      RECT 81.91 3.401 81.94 3.55 ;
      RECT 81.885 3.392 81.91 3.54 ;
      RECT 81.855 3.385 81.885 3.532 ;
      RECT 81.83 3.375 81.855 3.523 ;
      RECT 81.815 3.367 81.83 3.517 ;
      RECT 81.79 3.362 81.815 3.512 ;
      RECT 81.78 3.358 81.79 3.507 ;
      RECT 81.76 3.353 81.78 3.502 ;
      RECT 81.725 3.348 81.76 3.495 ;
      RECT 81.665 3.343 81.725 3.488 ;
      RECT 81.652 3.339 81.665 3.486 ;
      RECT 81.566 3.334 81.652 3.483 ;
      RECT 81.48 3.324 81.566 3.479 ;
      RECT 81.439 3.317 81.48 3.476 ;
      RECT 81.353 3.31 81.439 3.473 ;
      RECT 81.267 3.3 81.353 3.469 ;
      RECT 81.181 3.29 81.267 3.464 ;
      RECT 81.095 3.28 81.181 3.46 ;
      RECT 81.085 3.265 81.095 3.458 ;
      RECT 81.075 3.25 81.085 3.458 ;
      RECT 81.01 3.245 81.075 3.457 ;
      RECT 80.845 3.242 80.89 3.45 ;
      RECT 82.09 4.147 82.095 4.338 ;
      RECT 82.085 4.142 82.09 4.345 ;
      RECT 82.071 4.14 82.085 4.351 ;
      RECT 81.985 4.14 82.071 4.353 ;
      RECT 81.981 4.14 81.985 4.356 ;
      RECT 81.895 4.14 81.981 4.374 ;
      RECT 81.885 4.145 81.895 4.393 ;
      RECT 81.875 4.2 81.885 4.397 ;
      RECT 81.85 4.215 81.875 4.404 ;
      RECT 81.81 4.235 81.85 4.417 ;
      RECT 81.805 4.247 81.81 4.427 ;
      RECT 81.79 4.253 81.805 4.432 ;
      RECT 81.785 4.258 81.79 4.436 ;
      RECT 81.765 4.265 81.785 4.441 ;
      RECT 81.695 4.29 81.765 4.458 ;
      RECT 81.655 4.318 81.695 4.478 ;
      RECT 81.65 4.328 81.655 4.486 ;
      RECT 81.63 4.335 81.65 4.488 ;
      RECT 81.625 4.342 81.63 4.491 ;
      RECT 81.595 4.35 81.625 4.494 ;
      RECT 81.59 4.355 81.595 4.498 ;
      RECT 81.516 4.359 81.59 4.506 ;
      RECT 81.43 4.368 81.516 4.522 ;
      RECT 81.426 4.373 81.43 4.531 ;
      RECT 81.34 4.378 81.426 4.541 ;
      RECT 81.3 4.386 81.34 4.553 ;
      RECT 81.25 4.392 81.3 4.56 ;
      RECT 81.165 4.401 81.25 4.575 ;
      RECT 81.09 4.412 81.165 4.593 ;
      RECT 81.055 4.419 81.09 4.603 ;
      RECT 80.98 4.427 81.055 4.608 ;
      RECT 80.925 4.436 80.98 4.608 ;
      RECT 80.9 4.441 80.925 4.606 ;
      RECT 80.89 4.444 80.9 4.604 ;
      RECT 80.855 4.446 80.89 4.602 ;
      RECT 80.825 4.448 80.855 4.598 ;
      RECT 80.78 4.447 80.825 4.594 ;
      RECT 80.76 4.442 80.78 4.591 ;
      RECT 80.71 4.427 80.76 4.588 ;
      RECT 80.7 4.412 80.71 4.583 ;
      RECT 80.65 4.397 80.7 4.573 ;
      RECT 80.6 4.372 80.65 4.553 ;
      RECT 80.59 4.357 80.6 4.535 ;
      RECT 80.585 4.355 80.59 4.529 ;
      RECT 80.565 4.35 80.585 4.524 ;
      RECT 80.56 4.342 80.565 4.518 ;
      RECT 80.545 4.336 80.56 4.511 ;
      RECT 80.54 4.331 80.545 4.503 ;
      RECT 80.52 4.326 80.54 4.495 ;
      RECT 80.505 4.319 80.52 4.488 ;
      RECT 80.49 4.313 80.505 4.479 ;
      RECT 80.485 4.307 80.49 4.472 ;
      RECT 80.44 4.282 80.485 4.458 ;
      RECT 80.425 4.252 80.44 4.44 ;
      RECT 80.41 4.235 80.425 4.431 ;
      RECT 80.385 4.215 80.41 4.419 ;
      RECT 80.345 4.185 80.385 4.399 ;
      RECT 80.335 4.155 80.345 4.384 ;
      RECT 80.32 4.145 80.335 4.377 ;
      RECT 80.265 4.11 80.32 4.356 ;
      RECT 80.25 4.073 80.265 4.335 ;
      RECT 80.24 4.06 80.25 4.327 ;
      RECT 80.19 4.03 80.24 4.309 ;
      RECT 80.175 3.96 80.19 4.29 ;
      RECT 80.13 3.96 80.175 4.273 ;
      RECT 80.105 3.96 80.13 4.255 ;
      RECT 80.095 3.96 80.105 4.248 ;
      RECT 80.016 3.96 80.095 4.241 ;
      RECT 79.93 3.96 80.016 4.233 ;
      RECT 79.915 3.992 79.93 4.228 ;
      RECT 79.84 4.002 79.915 4.224 ;
      RECT 79.82 4.012 79.84 4.219 ;
      RECT 79.795 4.012 79.82 4.216 ;
      RECT 79.785 4.002 79.795 4.215 ;
      RECT 79.775 3.975 79.785 4.214 ;
      RECT 79.735 3.97 79.775 4.212 ;
      RECT 79.69 3.97 79.735 4.208 ;
      RECT 79.665 3.97 79.69 4.203 ;
      RECT 79.615 3.97 79.665 4.19 ;
      RECT 79.575 3.975 79.585 4.175 ;
      RECT 79.585 3.97 79.615 4.18 ;
      RECT 81.57 3.75 81.83 4.01 ;
      RECT 81.565 3.772 81.83 3.968 ;
      RECT 80.805 3.6 81.025 3.965 ;
      RECT 80.787 3.687 81.025 3.964 ;
      RECT 80.77 3.692 81.025 3.961 ;
      RECT 80.77 3.692 81.045 3.96 ;
      RECT 80.74 3.702 81.045 3.958 ;
      RECT 80.735 3.717 81.045 3.954 ;
      RECT 80.735 3.717 81.05 3.953 ;
      RECT 80.73 3.775 81.05 3.951 ;
      RECT 80.73 3.775 81.06 3.948 ;
      RECT 80.725 3.84 81.06 3.943 ;
      RECT 80.805 3.6 81.065 3.86 ;
      RECT 79.55 3.43 79.81 3.69 ;
      RECT 79.55 3.473 79.896 3.664 ;
      RECT 79.55 3.473 79.94 3.663 ;
      RECT 79.55 3.473 79.96 3.661 ;
      RECT 79.55 3.473 80.06 3.66 ;
      RECT 79.55 3.473 80.08 3.658 ;
      RECT 79.55 3.473 80.09 3.653 ;
      RECT 79.96 3.44 80.15 3.65 ;
      RECT 79.96 3.442 80.155 3.648 ;
      RECT 79.95 3.447 80.16 3.64 ;
      RECT 79.896 3.471 80.16 3.64 ;
      RECT 79.94 3.465 79.95 3.662 ;
      RECT 79.95 3.445 80.155 3.648 ;
      RECT 78.905 4.505 79.11 4.735 ;
      RECT 78.845 4.455 78.9 4.715 ;
      RECT 78.905 4.455 79.105 4.735 ;
      RECT 79.875 4.77 79.88 4.797 ;
      RECT 79.865 4.68 79.875 4.802 ;
      RECT 79.86 4.602 79.865 4.808 ;
      RECT 79.85 4.592 79.86 4.815 ;
      RECT 79.845 4.582 79.85 4.821 ;
      RECT 79.835 4.577 79.845 4.823 ;
      RECT 79.82 4.569 79.835 4.831 ;
      RECT 79.805 4.56 79.82 4.843 ;
      RECT 79.795 4.552 79.805 4.853 ;
      RECT 79.76 4.47 79.795 4.871 ;
      RECT 79.725 4.47 79.76 4.89 ;
      RECT 79.71 4.47 79.725 4.898 ;
      RECT 79.655 4.47 79.71 4.898 ;
      RECT 79.621 4.47 79.655 4.889 ;
      RECT 79.535 4.47 79.621 4.865 ;
      RECT 79.525 4.53 79.535 4.847 ;
      RECT 79.485 4.532 79.525 4.838 ;
      RECT 79.48 4.534 79.485 4.828 ;
      RECT 79.46 4.536 79.48 4.823 ;
      RECT 79.45 4.539 79.46 4.818 ;
      RECT 79.44 4.54 79.45 4.813 ;
      RECT 79.416 4.541 79.44 4.805 ;
      RECT 79.33 4.546 79.416 4.783 ;
      RECT 79.275 4.545 79.33 4.756 ;
      RECT 79.26 4.538 79.275 4.743 ;
      RECT 79.225 4.533 79.26 4.739 ;
      RECT 79.17 4.525 79.225 4.738 ;
      RECT 79.11 4.512 79.17 4.736 ;
      RECT 78.9 4.455 78.905 4.723 ;
      RECT 78.975 3.825 79.16 4.035 ;
      RECT 78.965 3.83 79.175 4.028 ;
      RECT 79.005 3.735 79.265 3.995 ;
      RECT 78.96 3.892 79.265 3.918 ;
      RECT 78.305 3.685 78.31 4.485 ;
      RECT 78.25 3.735 78.28 4.485 ;
      RECT 78.24 3.735 78.245 4.045 ;
      RECT 78.225 3.735 78.23 4.04 ;
      RECT 77.77 3.78 77.785 3.995 ;
      RECT 77.7 3.78 77.785 3.99 ;
      RECT 78.965 3.36 79.035 3.57 ;
      RECT 79.035 3.367 79.045 3.565 ;
      RECT 78.931 3.36 78.965 3.577 ;
      RECT 78.845 3.36 78.931 3.601 ;
      RECT 78.835 3.365 78.845 3.62 ;
      RECT 78.83 3.377 78.835 3.623 ;
      RECT 78.815 3.392 78.83 3.627 ;
      RECT 78.81 3.41 78.815 3.631 ;
      RECT 78.77 3.42 78.81 3.64 ;
      RECT 78.755 3.427 78.77 3.652 ;
      RECT 78.74 3.432 78.755 3.657 ;
      RECT 78.725 3.435 78.74 3.662 ;
      RECT 78.715 3.437 78.725 3.666 ;
      RECT 78.68 3.444 78.715 3.674 ;
      RECT 78.645 3.452 78.68 3.688 ;
      RECT 78.635 3.458 78.645 3.697 ;
      RECT 78.63 3.46 78.635 3.699 ;
      RECT 78.61 3.463 78.63 3.705 ;
      RECT 78.58 3.47 78.61 3.716 ;
      RECT 78.57 3.476 78.58 3.723 ;
      RECT 78.545 3.479 78.57 3.73 ;
      RECT 78.535 3.483 78.545 3.738 ;
      RECT 78.53 3.484 78.535 3.76 ;
      RECT 78.525 3.485 78.53 3.775 ;
      RECT 78.52 3.486 78.525 3.79 ;
      RECT 78.515 3.487 78.52 3.805 ;
      RECT 78.51 3.488 78.515 3.835 ;
      RECT 78.5 3.49 78.51 3.868 ;
      RECT 78.485 3.494 78.5 3.915 ;
      RECT 78.475 3.497 78.485 3.96 ;
      RECT 78.47 3.5 78.475 3.988 ;
      RECT 78.46 3.502 78.47 4.015 ;
      RECT 78.455 3.505 78.46 4.05 ;
      RECT 78.425 3.51 78.455 4.108 ;
      RECT 78.42 3.515 78.425 4.193 ;
      RECT 78.415 3.517 78.42 4.228 ;
      RECT 78.41 3.519 78.415 4.31 ;
      RECT 78.405 3.521 78.41 4.398 ;
      RECT 78.395 3.523 78.405 4.48 ;
      RECT 78.38 3.537 78.395 4.485 ;
      RECT 78.345 3.582 78.38 4.485 ;
      RECT 78.335 3.622 78.345 4.485 ;
      RECT 78.32 3.65 78.335 4.485 ;
      RECT 78.315 3.667 78.32 4.485 ;
      RECT 78.31 3.675 78.315 4.485 ;
      RECT 78.3 3.69 78.305 4.485 ;
      RECT 78.295 3.697 78.3 4.485 ;
      RECT 78.285 3.717 78.295 4.485 ;
      RECT 78.28 3.73 78.285 4.485 ;
      RECT 78.245 3.735 78.25 4.07 ;
      RECT 78.23 4.125 78.25 4.485 ;
      RECT 78.23 3.735 78.24 4.043 ;
      RECT 78.225 4.165 78.23 4.485 ;
      RECT 78.175 3.735 78.225 4.038 ;
      RECT 78.22 4.202 78.225 4.485 ;
      RECT 78.21 4.225 78.22 4.485 ;
      RECT 78.205 4.27 78.21 4.485 ;
      RECT 78.195 4.28 78.205 4.478 ;
      RECT 78.121 3.735 78.175 4.032 ;
      RECT 78.035 3.735 78.121 4.025 ;
      RECT 77.986 3.782 78.035 4.018 ;
      RECT 77.9 3.79 77.986 4.011 ;
      RECT 77.885 3.787 77.9 4.006 ;
      RECT 77.871 3.78 77.885 4.005 ;
      RECT 77.785 3.78 77.871 4 ;
      RECT 77.69 3.785 77.7 3.985 ;
      RECT 77.28 3.215 77.295 3.615 ;
      RECT 77.475 3.215 77.48 3.475 ;
      RECT 77.22 3.215 77.265 3.475 ;
      RECT 77.675 4.52 77.68 4.725 ;
      RECT 77.67 4.51 77.675 4.73 ;
      RECT 77.665 4.497 77.67 4.735 ;
      RECT 77.66 4.477 77.665 4.735 ;
      RECT 77.635 4.43 77.66 4.735 ;
      RECT 77.6 4.345 77.635 4.735 ;
      RECT 77.595 4.282 77.6 4.735 ;
      RECT 77.59 4.267 77.595 4.735 ;
      RECT 77.575 4.227 77.59 4.735 ;
      RECT 77.57 4.202 77.575 4.735 ;
      RECT 77.56 4.185 77.57 4.735 ;
      RECT 77.525 4.107 77.56 4.735 ;
      RECT 77.52 4.05 77.525 4.735 ;
      RECT 77.515 4.037 77.52 4.735 ;
      RECT 77.505 4.015 77.515 4.735 ;
      RECT 77.495 3.98 77.505 4.735 ;
      RECT 77.485 3.95 77.495 4.735 ;
      RECT 77.475 3.865 77.485 4.378 ;
      RECT 77.482 4.51 77.485 4.735 ;
      RECT 77.48 4.52 77.482 4.735 ;
      RECT 77.47 4.53 77.48 4.73 ;
      RECT 77.465 3.215 77.475 3.61 ;
      RECT 77.47 3.742 77.475 4.353 ;
      RECT 77.465 3.64 77.47 4.336 ;
      RECT 77.455 3.215 77.465 4.312 ;
      RECT 77.45 3.215 77.455 4.283 ;
      RECT 77.445 3.215 77.45 4.273 ;
      RECT 77.425 3.215 77.445 4.235 ;
      RECT 77.42 3.215 77.425 4.193 ;
      RECT 77.415 3.215 77.42 4.173 ;
      RECT 77.385 3.215 77.415 4.123 ;
      RECT 77.375 3.215 77.385 4.07 ;
      RECT 77.37 3.215 77.375 4.043 ;
      RECT 77.365 3.215 77.37 4.028 ;
      RECT 77.355 3.215 77.365 4.005 ;
      RECT 77.345 3.215 77.355 3.98 ;
      RECT 77.34 3.215 77.345 3.92 ;
      RECT 77.33 3.215 77.34 3.858 ;
      RECT 77.325 3.215 77.33 3.778 ;
      RECT 77.32 3.215 77.325 3.743 ;
      RECT 77.315 3.215 77.32 3.718 ;
      RECT 77.31 3.215 77.315 3.703 ;
      RECT 77.305 3.215 77.31 3.673 ;
      RECT 77.3 3.215 77.305 3.65 ;
      RECT 77.295 3.215 77.3 3.623 ;
      RECT 77.265 3.215 77.28 3.61 ;
      RECT 76.42 4.75 76.605 4.96 ;
      RECT 76.41 4.755 76.62 4.953 ;
      RECT 76.41 4.755 76.64 4.925 ;
      RECT 76.41 4.755 76.655 4.904 ;
      RECT 76.41 4.755 76.67 4.902 ;
      RECT 76.41 4.755 76.68 4.901 ;
      RECT 76.41 4.755 76.71 4.898 ;
      RECT 77.06 4.6 77.32 4.86 ;
      RECT 77.02 4.647 77.32 4.843 ;
      RECT 77.011 4.655 77.02 4.846 ;
      RECT 76.605 4.748 77.32 4.843 ;
      RECT 76.925 4.673 77.011 4.853 ;
      RECT 76.62 4.745 77.32 4.843 ;
      RECT 76.866 4.695 76.925 4.865 ;
      RECT 76.64 4.741 77.32 4.843 ;
      RECT 76.78 4.707 76.866 4.876 ;
      RECT 76.655 4.737 77.32 4.843 ;
      RECT 76.725 4.72 76.78 4.888 ;
      RECT 76.67 4.735 77.32 4.843 ;
      RECT 76.71 4.726 76.725 4.894 ;
      RECT 76.68 4.731 77.32 4.843 ;
      RECT 76.825 4.255 77.085 4.515 ;
      RECT 76.825 4.275 77.195 4.485 ;
      RECT 76.825 4.28 77.205 4.48 ;
      RECT 77.016 3.694 77.095 3.925 ;
      RECT 76.93 3.697 77.145 3.92 ;
      RECT 76.925 3.697 77.145 3.915 ;
      RECT 76.925 3.702 77.155 3.913 ;
      RECT 76.9 3.702 77.155 3.91 ;
      RECT 76.9 3.71 77.165 3.908 ;
      RECT 76.78 3.645 77.04 3.905 ;
      RECT 76.78 3.692 77.09 3.905 ;
      RECT 76.035 4.265 76.04 4.525 ;
      RECT 75.865 4.035 75.87 4.525 ;
      RECT 75.75 4.275 75.755 4.5 ;
      RECT 76.46 3.37 76.465 3.58 ;
      RECT 76.465 3.375 76.48 3.575 ;
      RECT 76.4 3.37 76.46 3.588 ;
      RECT 76.385 3.37 76.4 3.598 ;
      RECT 76.335 3.37 76.385 3.615 ;
      RECT 76.315 3.37 76.335 3.638 ;
      RECT 76.3 3.37 76.315 3.65 ;
      RECT 76.28 3.37 76.3 3.66 ;
      RECT 76.27 3.375 76.28 3.669 ;
      RECT 76.265 3.385 76.27 3.674 ;
      RECT 76.26 3.397 76.265 3.678 ;
      RECT 76.25 3.42 76.26 3.683 ;
      RECT 76.245 3.435 76.25 3.687 ;
      RECT 76.24 3.452 76.245 3.69 ;
      RECT 76.235 3.46 76.24 3.693 ;
      RECT 76.225 3.465 76.235 3.697 ;
      RECT 76.22 3.472 76.225 3.702 ;
      RECT 76.21 3.477 76.22 3.706 ;
      RECT 76.185 3.489 76.21 3.717 ;
      RECT 76.165 3.506 76.185 3.733 ;
      RECT 76.14 3.523 76.165 3.755 ;
      RECT 76.105 3.546 76.14 3.813 ;
      RECT 76.085 3.568 76.105 3.875 ;
      RECT 76.08 3.578 76.085 3.91 ;
      RECT 76.07 3.585 76.08 3.948 ;
      RECT 76.065 3.592 76.07 3.968 ;
      RECT 76.06 3.603 76.065 4.005 ;
      RECT 76.055 3.611 76.06 4.07 ;
      RECT 76.045 3.622 76.055 4.123 ;
      RECT 76.04 3.64 76.045 4.193 ;
      RECT 76.035 3.65 76.04 4.23 ;
      RECT 76.03 3.66 76.035 4.525 ;
      RECT 76.025 3.672 76.03 4.525 ;
      RECT 76.02 3.682 76.025 4.525 ;
      RECT 76.01 3.692 76.02 4.525 ;
      RECT 76 3.715 76.01 4.525 ;
      RECT 75.985 3.75 76 4.525 ;
      RECT 75.945 3.812 75.985 4.525 ;
      RECT 75.94 3.865 75.945 4.525 ;
      RECT 75.915 3.9 75.94 4.525 ;
      RECT 75.9 3.945 75.915 4.525 ;
      RECT 75.895 3.967 75.9 4.525 ;
      RECT 75.885 3.98 75.895 4.525 ;
      RECT 75.875 4.005 75.885 4.525 ;
      RECT 75.87 4.027 75.875 4.525 ;
      RECT 75.845 4.065 75.865 4.525 ;
      RECT 75.805 4.122 75.845 4.525 ;
      RECT 75.8 4.172 75.805 4.525 ;
      RECT 75.795 4.19 75.8 4.525 ;
      RECT 75.79 4.202 75.795 4.525 ;
      RECT 75.78 4.22 75.79 4.525 ;
      RECT 75.77 4.24 75.78 4.5 ;
      RECT 75.765 4.257 75.77 4.5 ;
      RECT 75.755 4.27 75.765 4.5 ;
      RECT 75.725 4.28 75.75 4.5 ;
      RECT 75.715 4.287 75.725 4.5 ;
      RECT 75.7 4.297 75.715 4.495 ;
      RECT 74.79 10.055 75.08 10.285 ;
      RECT 74.85 8.575 75.02 10.285 ;
      RECT 74.8 8.94 75.15 9.29 ;
      RECT 74.79 8.575 75.08 8.805 ;
      RECT 74.385 3.69 74.49 4.26 ;
      RECT 74.385 4.025 74.71 4.255 ;
      RECT 74.385 4.055 74.88 4.225 ;
      RECT 74.385 3.69 74.575 4.255 ;
      RECT 73.8 3.655 74.09 3.885 ;
      RECT 73.8 3.69 74.575 3.86 ;
      RECT 73.86 2.175 74.03 3.885 ;
      RECT 73.8 2.175 74.09 2.405 ;
      RECT 73.8 10.055 74.09 10.285 ;
      RECT 73.86 8.575 74.03 10.285 ;
      RECT 73.8 8.575 74.09 8.805 ;
      RECT 73.8 8.61 74.65 8.77 ;
      RECT 74.485 8.205 74.65 8.77 ;
      RECT 73.8 8.605 74.195 8.77 ;
      RECT 74.42 8.205 74.71 8.435 ;
      RECT 74.42 8.235 74.88 8.405 ;
      RECT 73.43 4.025 73.72 4.255 ;
      RECT 73.43 4.055 73.89 4.225 ;
      RECT 73.495 2.95 73.66 4.255 ;
      RECT 72.01 2.92 72.3 3.15 ;
      RECT 72.01 2.95 73.66 3.12 ;
      RECT 72.07 2.18 72.24 3.15 ;
      RECT 72.01 2.18 72.3 2.41 ;
      RECT 72.01 10.05 72.3 10.28 ;
      RECT 72.07 9.31 72.24 10.28 ;
      RECT 72.07 9.405 73.66 9.575 ;
      RECT 73.49 8.205 73.66 9.575 ;
      RECT 72.01 9.31 72.3 9.54 ;
      RECT 73.43 8.205 73.72 8.435 ;
      RECT 73.43 8.235 73.89 8.405 ;
      RECT 72.44 3.26 72.79 3.61 ;
      RECT 70.105 3.32 72.79 3.49 ;
      RECT 70.105 2.635 70.275 3.49 ;
      RECT 70.005 2.635 70.355 2.985 ;
      RECT 72.465 8.94 72.79 9.265 ;
      RECT 67.84 8.895 68.19 9.245 ;
      RECT 72.44 8.94 72.79 9.17 ;
      RECT 67.66 8.94 68.19 9.17 ;
      RECT 67.49 8.97 72.79 9.14 ;
      RECT 71.665 3.66 71.985 3.98 ;
      RECT 71.635 3.66 71.985 3.89 ;
      RECT 71.465 3.69 71.985 3.86 ;
      RECT 71.665 8.54 71.985 8.83 ;
      RECT 71.635 8.57 71.985 8.8 ;
      RECT 71.465 8.6 71.985 8.77 ;
      RECT 68.3 3.76 68.485 3.97 ;
      RECT 68.29 3.765 68.5 3.963 ;
      RECT 68.29 3.765 68.586 3.94 ;
      RECT 68.29 3.765 68.645 3.915 ;
      RECT 68.29 3.765 68.7 3.895 ;
      RECT 68.29 3.765 68.71 3.883 ;
      RECT 68.29 3.765 68.905 3.822 ;
      RECT 68.29 3.765 68.935 3.805 ;
      RECT 68.29 3.765 68.955 3.795 ;
      RECT 68.835 3.53 69.095 3.79 ;
      RECT 68.82 3.62 68.835 3.837 ;
      RECT 68.355 3.752 69.095 3.79 ;
      RECT 68.806 3.631 68.82 3.843 ;
      RECT 68.395 3.745 69.095 3.79 ;
      RECT 68.72 3.671 68.806 3.862 ;
      RECT 68.645 3.732 69.095 3.79 ;
      RECT 68.715 3.707 68.72 3.879 ;
      RECT 68.7 3.717 69.095 3.79 ;
      RECT 68.71 3.712 68.715 3.881 ;
      RECT 69.005 4.217 69.01 4.309 ;
      RECT 69 4.195 69.005 4.326 ;
      RECT 68.995 4.185 69 4.338 ;
      RECT 68.985 4.176 68.995 4.348 ;
      RECT 68.98 4.171 68.985 4.356 ;
      RECT 68.975 4.03 68.98 4.359 ;
      RECT 68.941 4.03 68.975 4.37 ;
      RECT 68.855 4.03 68.941 4.405 ;
      RECT 68.775 4.03 68.855 4.453 ;
      RECT 68.746 4.03 68.775 4.477 ;
      RECT 68.66 4.03 68.746 4.483 ;
      RECT 68.655 4.214 68.66 4.488 ;
      RECT 68.62 4.225 68.655 4.491 ;
      RECT 68.595 4.24 68.62 4.495 ;
      RECT 68.581 4.249 68.595 4.497 ;
      RECT 68.495 4.276 68.581 4.503 ;
      RECT 68.43 4.317 68.495 4.512 ;
      RECT 68.415 4.337 68.43 4.517 ;
      RECT 68.385 4.347 68.415 4.52 ;
      RECT 68.38 4.357 68.385 4.523 ;
      RECT 68.35 4.362 68.38 4.525 ;
      RECT 68.33 4.367 68.35 4.529 ;
      RECT 68.245 4.37 68.33 4.536 ;
      RECT 68.23 4.367 68.245 4.542 ;
      RECT 68.22 4.364 68.23 4.544 ;
      RECT 68.2 4.361 68.22 4.546 ;
      RECT 68.18 4.357 68.2 4.547 ;
      RECT 68.165 4.353 68.18 4.549 ;
      RECT 68.155 4.35 68.165 4.55 ;
      RECT 68.115 4.344 68.155 4.548 ;
      RECT 68.105 4.339 68.115 4.546 ;
      RECT 68.09 4.336 68.105 4.542 ;
      RECT 68.065 4.331 68.09 4.535 ;
      RECT 68.015 4.322 68.065 4.523 ;
      RECT 67.945 4.308 68.015 4.505 ;
      RECT 67.887 4.293 67.945 4.487 ;
      RECT 67.801 4.276 67.887 4.467 ;
      RECT 67.715 4.255 67.801 4.442 ;
      RECT 67.665 4.24 67.715 4.423 ;
      RECT 67.661 4.234 67.665 4.415 ;
      RECT 67.575 4.224 67.661 4.402 ;
      RECT 67.54 4.209 67.575 4.385 ;
      RECT 67.525 4.202 67.54 4.378 ;
      RECT 67.465 4.19 67.525 4.366 ;
      RECT 67.445 4.177 67.465 4.354 ;
      RECT 67.405 4.168 67.445 4.346 ;
      RECT 67.4 4.16 67.405 4.339 ;
      RECT 67.32 4.15 67.4 4.325 ;
      RECT 67.305 4.137 67.32 4.31 ;
      RECT 67.3 4.135 67.305 4.308 ;
      RECT 67.221 4.123 67.3 4.295 ;
      RECT 67.135 4.098 67.221 4.27 ;
      RECT 67.12 4.067 67.135 4.255 ;
      RECT 67.105 4.042 67.12 4.251 ;
      RECT 67.09 4.035 67.105 4.247 ;
      RECT 66.915 4.04 66.92 4.243 ;
      RECT 66.91 4.045 66.915 4.238 ;
      RECT 66.92 4.035 67.09 4.245 ;
      RECT 67.635 3.795 67.74 4.055 ;
      RECT 68.45 3.32 68.455 3.545 ;
      RECT 68.58 3.32 68.635 3.53 ;
      RECT 68.635 3.325 68.645 3.523 ;
      RECT 68.541 3.32 68.58 3.533 ;
      RECT 68.455 3.32 68.541 3.54 ;
      RECT 68.435 3.325 68.45 3.546 ;
      RECT 68.425 3.365 68.435 3.548 ;
      RECT 68.395 3.375 68.425 3.55 ;
      RECT 68.39 3.38 68.395 3.552 ;
      RECT 68.365 3.385 68.39 3.554 ;
      RECT 68.35 3.39 68.365 3.556 ;
      RECT 68.335 3.392 68.35 3.558 ;
      RECT 68.33 3.397 68.335 3.56 ;
      RECT 68.28 3.405 68.33 3.563 ;
      RECT 68.255 3.414 68.28 3.568 ;
      RECT 68.245 3.421 68.255 3.573 ;
      RECT 68.24 3.424 68.245 3.577 ;
      RECT 68.22 3.427 68.24 3.586 ;
      RECT 68.19 3.435 68.22 3.606 ;
      RECT 68.161 3.448 68.19 3.628 ;
      RECT 68.075 3.482 68.161 3.672 ;
      RECT 68.07 3.508 68.075 3.71 ;
      RECT 68.065 3.512 68.07 3.719 ;
      RECT 68.03 3.525 68.065 3.752 ;
      RECT 68.02 3.539 68.03 3.79 ;
      RECT 68.015 3.543 68.02 3.803 ;
      RECT 68.01 3.547 68.015 3.808 ;
      RECT 68 3.555 68.01 3.82 ;
      RECT 67.995 3.562 68 3.835 ;
      RECT 67.97 3.575 67.995 3.86 ;
      RECT 67.93 3.604 67.97 3.915 ;
      RECT 67.915 3.629 67.93 3.97 ;
      RECT 67.905 3.64 67.915 3.993 ;
      RECT 67.9 3.647 67.905 4.005 ;
      RECT 67.895 3.651 67.9 4.013 ;
      RECT 67.84 3.679 67.895 4.055 ;
      RECT 67.82 3.715 67.84 4.055 ;
      RECT 67.805 3.73 67.82 4.055 ;
      RECT 67.75 3.762 67.805 4.055 ;
      RECT 67.74 3.792 67.75 4.055 ;
      RECT 67.35 3.407 67.535 3.645 ;
      RECT 67.335 3.409 67.545 3.64 ;
      RECT 67.22 3.355 67.48 3.615 ;
      RECT 67.215 3.392 67.48 3.569 ;
      RECT 67.21 3.402 67.48 3.566 ;
      RECT 67.205 3.442 67.545 3.56 ;
      RECT 67.2 3.475 67.545 3.55 ;
      RECT 67.21 3.417 67.56 3.488 ;
      RECT 67.507 4.515 67.52 5.045 ;
      RECT 67.421 4.515 67.52 5.044 ;
      RECT 67.421 4.515 67.525 5.043 ;
      RECT 67.335 4.515 67.525 5.041 ;
      RECT 67.33 4.515 67.525 5.038 ;
      RECT 67.33 4.515 67.535 5.036 ;
      RECT 67.325 4.807 67.535 5.033 ;
      RECT 67.325 4.817 67.54 5.03 ;
      RECT 67.325 4.885 67.545 5.026 ;
      RECT 67.315 4.89 67.545 5.025 ;
      RECT 67.315 4.982 67.55 5.022 ;
      RECT 67.3 4.515 67.56 4.775 ;
      RECT 67.23 10.05 67.52 10.28 ;
      RECT 67.29 9.31 67.46 10.28 ;
      RECT 67.205 9.34 67.545 9.685 ;
      RECT 67.23 9.31 67.52 9.685 ;
      RECT 66.53 3.505 66.575 5.04 ;
      RECT 66.73 3.505 66.76 3.72 ;
      RECT 65.105 3.245 65.225 3.455 ;
      RECT 64.765 3.195 65.025 3.455 ;
      RECT 64.765 3.24 65.06 3.445 ;
      RECT 66.77 3.521 66.775 3.575 ;
      RECT 66.765 3.514 66.77 3.708 ;
      RECT 66.76 3.508 66.765 3.715 ;
      RECT 66.715 3.505 66.73 3.728 ;
      RECT 66.71 3.505 66.715 3.75 ;
      RECT 66.705 3.505 66.71 3.798 ;
      RECT 66.7 3.505 66.705 3.818 ;
      RECT 66.69 3.505 66.7 3.925 ;
      RECT 66.685 3.505 66.69 3.988 ;
      RECT 66.68 3.505 66.685 4.045 ;
      RECT 66.675 3.505 66.68 4.053 ;
      RECT 66.66 3.505 66.675 4.16 ;
      RECT 66.65 3.505 66.66 4.295 ;
      RECT 66.64 3.505 66.65 4.405 ;
      RECT 66.63 3.505 66.64 4.462 ;
      RECT 66.625 3.505 66.63 4.502 ;
      RECT 66.62 3.505 66.625 4.538 ;
      RECT 66.61 3.505 66.62 4.578 ;
      RECT 66.605 3.505 66.61 4.62 ;
      RECT 66.585 3.505 66.605 4.685 ;
      RECT 66.59 4.83 66.595 5.01 ;
      RECT 66.585 4.812 66.59 5.018 ;
      RECT 66.58 3.505 66.585 4.748 ;
      RECT 66.58 4.792 66.585 5.025 ;
      RECT 66.575 3.505 66.58 5.035 ;
      RECT 66.52 3.505 66.53 3.805 ;
      RECT 66.525 4.052 66.53 5.04 ;
      RECT 66.52 4.117 66.525 5.04 ;
      RECT 66.515 3.506 66.52 3.795 ;
      RECT 66.51 4.182 66.52 5.04 ;
      RECT 66.505 3.507 66.515 3.785 ;
      RECT 66.495 4.295 66.51 5.04 ;
      RECT 66.5 3.508 66.505 3.775 ;
      RECT 66.48 3.509 66.5 3.753 ;
      RECT 66.485 4.392 66.495 5.04 ;
      RECT 66.48 4.467 66.485 5.04 ;
      RECT 66.47 3.508 66.48 3.73 ;
      RECT 66.475 4.51 66.48 5.04 ;
      RECT 66.47 4.537 66.475 5.04 ;
      RECT 66.46 3.506 66.47 3.718 ;
      RECT 66.465 4.58 66.47 5.04 ;
      RECT 66.46 4.607 66.465 5.04 ;
      RECT 66.45 3.505 66.46 3.705 ;
      RECT 66.455 4.622 66.46 5.04 ;
      RECT 66.415 4.68 66.455 5.04 ;
      RECT 66.445 3.504 66.45 3.69 ;
      RECT 66.44 3.502 66.445 3.683 ;
      RECT 66.43 3.499 66.44 3.673 ;
      RECT 66.425 3.496 66.43 3.658 ;
      RECT 66.41 3.492 66.425 3.651 ;
      RECT 66.405 4.735 66.415 5.04 ;
      RECT 66.405 3.489 66.41 3.646 ;
      RECT 66.39 3.485 66.405 3.64 ;
      RECT 66.4 4.752 66.405 5.04 ;
      RECT 66.39 4.815 66.4 5.04 ;
      RECT 66.31 3.47 66.39 3.62 ;
      RECT 66.385 4.822 66.39 5.035 ;
      RECT 66.38 4.83 66.385 5.025 ;
      RECT 66.3 3.456 66.31 3.604 ;
      RECT 66.285 3.452 66.3 3.602 ;
      RECT 66.275 3.447 66.285 3.598 ;
      RECT 66.25 3.44 66.275 3.59 ;
      RECT 66.245 3.435 66.25 3.585 ;
      RECT 66.235 3.435 66.245 3.583 ;
      RECT 66.225 3.433 66.235 3.581 ;
      RECT 66.195 3.425 66.225 3.575 ;
      RECT 66.18 3.417 66.195 3.568 ;
      RECT 66.16 3.412 66.18 3.561 ;
      RECT 66.155 3.408 66.16 3.556 ;
      RECT 66.125 3.401 66.155 3.55 ;
      RECT 66.1 3.392 66.125 3.54 ;
      RECT 66.07 3.385 66.1 3.532 ;
      RECT 66.045 3.375 66.07 3.523 ;
      RECT 66.03 3.367 66.045 3.517 ;
      RECT 66.005 3.362 66.03 3.512 ;
      RECT 65.995 3.358 66.005 3.507 ;
      RECT 65.975 3.353 65.995 3.502 ;
      RECT 65.94 3.348 65.975 3.495 ;
      RECT 65.88 3.343 65.94 3.488 ;
      RECT 65.867 3.339 65.88 3.486 ;
      RECT 65.781 3.334 65.867 3.483 ;
      RECT 65.695 3.324 65.781 3.479 ;
      RECT 65.654 3.317 65.695 3.476 ;
      RECT 65.568 3.31 65.654 3.473 ;
      RECT 65.482 3.3 65.568 3.469 ;
      RECT 65.396 3.29 65.482 3.464 ;
      RECT 65.31 3.28 65.396 3.46 ;
      RECT 65.3 3.265 65.31 3.458 ;
      RECT 65.29 3.25 65.3 3.458 ;
      RECT 65.225 3.245 65.29 3.457 ;
      RECT 65.06 3.242 65.105 3.45 ;
      RECT 66.305 4.147 66.31 4.338 ;
      RECT 66.3 4.142 66.305 4.345 ;
      RECT 66.286 4.14 66.3 4.351 ;
      RECT 66.2 4.14 66.286 4.353 ;
      RECT 66.196 4.14 66.2 4.356 ;
      RECT 66.11 4.14 66.196 4.374 ;
      RECT 66.1 4.145 66.11 4.393 ;
      RECT 66.09 4.2 66.1 4.397 ;
      RECT 66.065 4.215 66.09 4.404 ;
      RECT 66.025 4.235 66.065 4.417 ;
      RECT 66.02 4.247 66.025 4.427 ;
      RECT 66.005 4.253 66.02 4.432 ;
      RECT 66 4.258 66.005 4.436 ;
      RECT 65.98 4.265 66 4.441 ;
      RECT 65.91 4.29 65.98 4.458 ;
      RECT 65.87 4.318 65.91 4.478 ;
      RECT 65.865 4.328 65.87 4.486 ;
      RECT 65.845 4.335 65.865 4.488 ;
      RECT 65.84 4.342 65.845 4.491 ;
      RECT 65.81 4.35 65.84 4.494 ;
      RECT 65.805 4.355 65.81 4.498 ;
      RECT 65.731 4.359 65.805 4.506 ;
      RECT 65.645 4.368 65.731 4.522 ;
      RECT 65.641 4.373 65.645 4.531 ;
      RECT 65.555 4.378 65.641 4.541 ;
      RECT 65.515 4.386 65.555 4.553 ;
      RECT 65.465 4.392 65.515 4.56 ;
      RECT 65.38 4.401 65.465 4.575 ;
      RECT 65.305 4.412 65.38 4.593 ;
      RECT 65.27 4.419 65.305 4.603 ;
      RECT 65.195 4.427 65.27 4.608 ;
      RECT 65.14 4.436 65.195 4.608 ;
      RECT 65.115 4.441 65.14 4.606 ;
      RECT 65.105 4.444 65.115 4.604 ;
      RECT 65.07 4.446 65.105 4.602 ;
      RECT 65.04 4.448 65.07 4.598 ;
      RECT 64.995 4.447 65.04 4.594 ;
      RECT 64.975 4.442 64.995 4.591 ;
      RECT 64.925 4.427 64.975 4.588 ;
      RECT 64.915 4.412 64.925 4.583 ;
      RECT 64.865 4.397 64.915 4.573 ;
      RECT 64.815 4.372 64.865 4.553 ;
      RECT 64.805 4.357 64.815 4.535 ;
      RECT 64.8 4.355 64.805 4.529 ;
      RECT 64.78 4.35 64.8 4.524 ;
      RECT 64.775 4.342 64.78 4.518 ;
      RECT 64.76 4.336 64.775 4.511 ;
      RECT 64.755 4.331 64.76 4.503 ;
      RECT 64.735 4.326 64.755 4.495 ;
      RECT 64.72 4.319 64.735 4.488 ;
      RECT 64.705 4.313 64.72 4.479 ;
      RECT 64.7 4.307 64.705 4.472 ;
      RECT 64.655 4.282 64.7 4.458 ;
      RECT 64.64 4.252 64.655 4.44 ;
      RECT 64.625 4.235 64.64 4.431 ;
      RECT 64.6 4.215 64.625 4.419 ;
      RECT 64.56 4.185 64.6 4.399 ;
      RECT 64.55 4.155 64.56 4.384 ;
      RECT 64.535 4.145 64.55 4.377 ;
      RECT 64.48 4.11 64.535 4.356 ;
      RECT 64.465 4.073 64.48 4.335 ;
      RECT 64.455 4.06 64.465 4.327 ;
      RECT 64.405 4.03 64.455 4.309 ;
      RECT 64.39 3.96 64.405 4.29 ;
      RECT 64.345 3.96 64.39 4.273 ;
      RECT 64.32 3.96 64.345 4.255 ;
      RECT 64.31 3.96 64.32 4.248 ;
      RECT 64.231 3.96 64.31 4.241 ;
      RECT 64.145 3.96 64.231 4.233 ;
      RECT 64.13 3.992 64.145 4.228 ;
      RECT 64.055 4.002 64.13 4.224 ;
      RECT 64.035 4.012 64.055 4.219 ;
      RECT 64.01 4.012 64.035 4.216 ;
      RECT 64 4.002 64.01 4.215 ;
      RECT 63.99 3.975 64 4.214 ;
      RECT 63.95 3.97 63.99 4.212 ;
      RECT 63.905 3.97 63.95 4.208 ;
      RECT 63.88 3.97 63.905 4.203 ;
      RECT 63.83 3.97 63.88 4.19 ;
      RECT 63.79 3.975 63.8 4.175 ;
      RECT 63.8 3.97 63.83 4.18 ;
      RECT 65.785 3.75 66.045 4.01 ;
      RECT 65.78 3.772 66.045 3.968 ;
      RECT 65.02 3.6 65.24 3.965 ;
      RECT 65.002 3.687 65.24 3.964 ;
      RECT 64.985 3.692 65.24 3.961 ;
      RECT 64.985 3.692 65.26 3.96 ;
      RECT 64.955 3.702 65.26 3.958 ;
      RECT 64.95 3.717 65.26 3.954 ;
      RECT 64.95 3.717 65.265 3.953 ;
      RECT 64.945 3.775 65.265 3.951 ;
      RECT 64.945 3.775 65.275 3.948 ;
      RECT 64.94 3.84 65.275 3.943 ;
      RECT 65.02 3.6 65.28 3.86 ;
      RECT 63.765 3.43 64.025 3.69 ;
      RECT 63.765 3.473 64.111 3.664 ;
      RECT 63.765 3.473 64.155 3.663 ;
      RECT 63.765 3.473 64.175 3.661 ;
      RECT 63.765 3.473 64.275 3.66 ;
      RECT 63.765 3.473 64.295 3.658 ;
      RECT 63.765 3.473 64.305 3.653 ;
      RECT 64.175 3.44 64.365 3.65 ;
      RECT 64.175 3.442 64.37 3.648 ;
      RECT 64.165 3.447 64.375 3.64 ;
      RECT 64.111 3.471 64.375 3.64 ;
      RECT 64.155 3.465 64.165 3.662 ;
      RECT 64.165 3.445 64.37 3.648 ;
      RECT 63.12 4.505 63.325 4.735 ;
      RECT 63.06 4.455 63.115 4.715 ;
      RECT 63.12 4.455 63.32 4.735 ;
      RECT 64.09 4.77 64.095 4.797 ;
      RECT 64.08 4.68 64.09 4.802 ;
      RECT 64.075 4.602 64.08 4.808 ;
      RECT 64.065 4.592 64.075 4.815 ;
      RECT 64.06 4.582 64.065 4.821 ;
      RECT 64.05 4.577 64.06 4.823 ;
      RECT 64.035 4.569 64.05 4.831 ;
      RECT 64.02 4.56 64.035 4.843 ;
      RECT 64.01 4.552 64.02 4.853 ;
      RECT 63.975 4.47 64.01 4.871 ;
      RECT 63.94 4.47 63.975 4.89 ;
      RECT 63.925 4.47 63.94 4.898 ;
      RECT 63.87 4.47 63.925 4.898 ;
      RECT 63.836 4.47 63.87 4.889 ;
      RECT 63.75 4.47 63.836 4.865 ;
      RECT 63.74 4.53 63.75 4.847 ;
      RECT 63.7 4.532 63.74 4.838 ;
      RECT 63.695 4.534 63.7 4.828 ;
      RECT 63.675 4.536 63.695 4.823 ;
      RECT 63.665 4.539 63.675 4.818 ;
      RECT 63.655 4.54 63.665 4.813 ;
      RECT 63.631 4.541 63.655 4.805 ;
      RECT 63.545 4.546 63.631 4.783 ;
      RECT 63.49 4.545 63.545 4.756 ;
      RECT 63.475 4.538 63.49 4.743 ;
      RECT 63.44 4.533 63.475 4.739 ;
      RECT 63.385 4.525 63.44 4.738 ;
      RECT 63.325 4.512 63.385 4.736 ;
      RECT 63.115 4.455 63.12 4.723 ;
      RECT 63.19 3.825 63.375 4.035 ;
      RECT 63.18 3.83 63.39 4.028 ;
      RECT 63.22 3.735 63.48 3.995 ;
      RECT 63.175 3.892 63.48 3.918 ;
      RECT 62.52 3.685 62.525 4.485 ;
      RECT 62.465 3.735 62.495 4.485 ;
      RECT 62.455 3.735 62.46 4.045 ;
      RECT 62.44 3.735 62.445 4.04 ;
      RECT 61.985 3.78 62 3.995 ;
      RECT 61.915 3.78 62 3.99 ;
      RECT 63.18 3.36 63.25 3.57 ;
      RECT 63.25 3.367 63.26 3.565 ;
      RECT 63.146 3.36 63.18 3.577 ;
      RECT 63.06 3.36 63.146 3.601 ;
      RECT 63.05 3.365 63.06 3.62 ;
      RECT 63.045 3.377 63.05 3.623 ;
      RECT 63.03 3.392 63.045 3.627 ;
      RECT 63.025 3.41 63.03 3.631 ;
      RECT 62.985 3.42 63.025 3.64 ;
      RECT 62.97 3.427 62.985 3.652 ;
      RECT 62.955 3.432 62.97 3.657 ;
      RECT 62.94 3.435 62.955 3.662 ;
      RECT 62.93 3.437 62.94 3.666 ;
      RECT 62.895 3.444 62.93 3.674 ;
      RECT 62.86 3.452 62.895 3.688 ;
      RECT 62.85 3.458 62.86 3.697 ;
      RECT 62.845 3.46 62.85 3.699 ;
      RECT 62.825 3.463 62.845 3.705 ;
      RECT 62.795 3.47 62.825 3.716 ;
      RECT 62.785 3.476 62.795 3.723 ;
      RECT 62.76 3.479 62.785 3.73 ;
      RECT 62.75 3.483 62.76 3.738 ;
      RECT 62.745 3.484 62.75 3.76 ;
      RECT 62.74 3.485 62.745 3.775 ;
      RECT 62.735 3.486 62.74 3.79 ;
      RECT 62.73 3.487 62.735 3.805 ;
      RECT 62.725 3.488 62.73 3.835 ;
      RECT 62.715 3.49 62.725 3.868 ;
      RECT 62.7 3.494 62.715 3.915 ;
      RECT 62.69 3.497 62.7 3.96 ;
      RECT 62.685 3.5 62.69 3.988 ;
      RECT 62.675 3.502 62.685 4.015 ;
      RECT 62.67 3.505 62.675 4.05 ;
      RECT 62.64 3.51 62.67 4.108 ;
      RECT 62.635 3.515 62.64 4.193 ;
      RECT 62.63 3.517 62.635 4.228 ;
      RECT 62.625 3.519 62.63 4.31 ;
      RECT 62.62 3.521 62.625 4.398 ;
      RECT 62.61 3.523 62.62 4.48 ;
      RECT 62.595 3.537 62.61 4.485 ;
      RECT 62.56 3.582 62.595 4.485 ;
      RECT 62.55 3.622 62.56 4.485 ;
      RECT 62.535 3.65 62.55 4.485 ;
      RECT 62.53 3.667 62.535 4.485 ;
      RECT 62.525 3.675 62.53 4.485 ;
      RECT 62.515 3.69 62.52 4.485 ;
      RECT 62.51 3.697 62.515 4.485 ;
      RECT 62.5 3.717 62.51 4.485 ;
      RECT 62.495 3.73 62.5 4.485 ;
      RECT 62.46 3.735 62.465 4.07 ;
      RECT 62.445 4.125 62.465 4.485 ;
      RECT 62.445 3.735 62.455 4.043 ;
      RECT 62.44 4.165 62.445 4.485 ;
      RECT 62.39 3.735 62.44 4.038 ;
      RECT 62.435 4.202 62.44 4.485 ;
      RECT 62.425 4.225 62.435 4.485 ;
      RECT 62.42 4.27 62.425 4.485 ;
      RECT 62.41 4.28 62.42 4.478 ;
      RECT 62.336 3.735 62.39 4.032 ;
      RECT 62.25 3.735 62.336 4.025 ;
      RECT 62.201 3.782 62.25 4.018 ;
      RECT 62.115 3.79 62.201 4.011 ;
      RECT 62.1 3.787 62.115 4.006 ;
      RECT 62.086 3.78 62.1 4.005 ;
      RECT 62 3.78 62.086 4 ;
      RECT 61.905 3.785 61.915 3.985 ;
      RECT 61.495 3.215 61.51 3.615 ;
      RECT 61.69 3.215 61.695 3.475 ;
      RECT 61.435 3.215 61.48 3.475 ;
      RECT 61.89 4.52 61.895 4.725 ;
      RECT 61.885 4.51 61.89 4.73 ;
      RECT 61.88 4.497 61.885 4.735 ;
      RECT 61.875 4.477 61.88 4.735 ;
      RECT 61.85 4.43 61.875 4.735 ;
      RECT 61.815 4.345 61.85 4.735 ;
      RECT 61.81 4.282 61.815 4.735 ;
      RECT 61.805 4.267 61.81 4.735 ;
      RECT 61.79 4.227 61.805 4.735 ;
      RECT 61.785 4.202 61.79 4.735 ;
      RECT 61.775 4.185 61.785 4.735 ;
      RECT 61.74 4.107 61.775 4.735 ;
      RECT 61.735 4.05 61.74 4.735 ;
      RECT 61.73 4.037 61.735 4.735 ;
      RECT 61.72 4.015 61.73 4.735 ;
      RECT 61.71 3.98 61.72 4.735 ;
      RECT 61.7 3.95 61.71 4.735 ;
      RECT 61.69 3.865 61.7 4.378 ;
      RECT 61.697 4.51 61.7 4.735 ;
      RECT 61.695 4.52 61.697 4.735 ;
      RECT 61.685 4.53 61.695 4.73 ;
      RECT 61.68 3.215 61.69 3.61 ;
      RECT 61.685 3.742 61.69 4.353 ;
      RECT 61.68 3.64 61.685 4.336 ;
      RECT 61.67 3.215 61.68 4.312 ;
      RECT 61.665 3.215 61.67 4.283 ;
      RECT 61.66 3.215 61.665 4.273 ;
      RECT 61.64 3.215 61.66 4.235 ;
      RECT 61.635 3.215 61.64 4.193 ;
      RECT 61.63 3.215 61.635 4.173 ;
      RECT 61.6 3.215 61.63 4.123 ;
      RECT 61.59 3.215 61.6 4.07 ;
      RECT 61.585 3.215 61.59 4.043 ;
      RECT 61.58 3.215 61.585 4.028 ;
      RECT 61.57 3.215 61.58 4.005 ;
      RECT 61.56 3.215 61.57 3.98 ;
      RECT 61.555 3.215 61.56 3.92 ;
      RECT 61.545 3.215 61.555 3.858 ;
      RECT 61.54 3.215 61.545 3.778 ;
      RECT 61.535 3.215 61.54 3.743 ;
      RECT 61.53 3.215 61.535 3.718 ;
      RECT 61.525 3.215 61.53 3.703 ;
      RECT 61.52 3.215 61.525 3.673 ;
      RECT 61.515 3.215 61.52 3.65 ;
      RECT 61.51 3.215 61.515 3.623 ;
      RECT 61.48 3.215 61.495 3.61 ;
      RECT 60.635 4.75 60.82 4.96 ;
      RECT 60.625 4.755 60.835 4.953 ;
      RECT 60.625 4.755 60.855 4.925 ;
      RECT 60.625 4.755 60.87 4.904 ;
      RECT 60.625 4.755 60.885 4.902 ;
      RECT 60.625 4.755 60.895 4.901 ;
      RECT 60.625 4.755 60.925 4.898 ;
      RECT 61.275 4.6 61.535 4.86 ;
      RECT 61.235 4.647 61.535 4.843 ;
      RECT 61.226 4.655 61.235 4.846 ;
      RECT 60.82 4.748 61.535 4.843 ;
      RECT 61.14 4.673 61.226 4.853 ;
      RECT 60.835 4.745 61.535 4.843 ;
      RECT 61.081 4.695 61.14 4.865 ;
      RECT 60.855 4.741 61.535 4.843 ;
      RECT 60.995 4.707 61.081 4.876 ;
      RECT 60.87 4.737 61.535 4.843 ;
      RECT 60.94 4.72 60.995 4.888 ;
      RECT 60.885 4.735 61.535 4.843 ;
      RECT 60.925 4.726 60.94 4.894 ;
      RECT 60.895 4.731 61.535 4.843 ;
      RECT 61.04 4.255 61.3 4.515 ;
      RECT 61.04 4.275 61.41 4.485 ;
      RECT 61.04 4.28 61.42 4.48 ;
      RECT 61.231 3.694 61.31 3.925 ;
      RECT 61.145 3.697 61.36 3.92 ;
      RECT 61.14 3.697 61.36 3.915 ;
      RECT 61.14 3.702 61.37 3.913 ;
      RECT 61.115 3.702 61.37 3.91 ;
      RECT 61.115 3.71 61.38 3.908 ;
      RECT 60.995 3.645 61.255 3.905 ;
      RECT 60.995 3.692 61.305 3.905 ;
      RECT 60.25 4.265 60.255 4.525 ;
      RECT 60.08 4.035 60.085 4.525 ;
      RECT 59.965 4.275 59.97 4.5 ;
      RECT 60.675 3.37 60.68 3.58 ;
      RECT 60.68 3.375 60.695 3.575 ;
      RECT 60.615 3.37 60.675 3.588 ;
      RECT 60.6 3.37 60.615 3.598 ;
      RECT 60.55 3.37 60.6 3.615 ;
      RECT 60.53 3.37 60.55 3.638 ;
      RECT 60.515 3.37 60.53 3.65 ;
      RECT 60.495 3.37 60.515 3.66 ;
      RECT 60.485 3.375 60.495 3.669 ;
      RECT 60.48 3.385 60.485 3.674 ;
      RECT 60.475 3.397 60.48 3.678 ;
      RECT 60.465 3.42 60.475 3.683 ;
      RECT 60.46 3.435 60.465 3.687 ;
      RECT 60.455 3.452 60.46 3.69 ;
      RECT 60.45 3.46 60.455 3.693 ;
      RECT 60.44 3.465 60.45 3.697 ;
      RECT 60.435 3.472 60.44 3.702 ;
      RECT 60.425 3.477 60.435 3.706 ;
      RECT 60.4 3.489 60.425 3.717 ;
      RECT 60.38 3.506 60.4 3.733 ;
      RECT 60.355 3.523 60.38 3.755 ;
      RECT 60.32 3.546 60.355 3.813 ;
      RECT 60.3 3.568 60.32 3.875 ;
      RECT 60.295 3.578 60.3 3.91 ;
      RECT 60.285 3.585 60.295 3.948 ;
      RECT 60.28 3.592 60.285 3.968 ;
      RECT 60.275 3.603 60.28 4.005 ;
      RECT 60.27 3.611 60.275 4.07 ;
      RECT 60.26 3.622 60.27 4.123 ;
      RECT 60.255 3.64 60.26 4.193 ;
      RECT 60.25 3.65 60.255 4.23 ;
      RECT 60.245 3.66 60.25 4.525 ;
      RECT 60.24 3.672 60.245 4.525 ;
      RECT 60.235 3.682 60.24 4.525 ;
      RECT 60.225 3.692 60.235 4.525 ;
      RECT 60.215 3.715 60.225 4.525 ;
      RECT 60.2 3.75 60.215 4.525 ;
      RECT 60.16 3.812 60.2 4.525 ;
      RECT 60.155 3.865 60.16 4.525 ;
      RECT 60.13 3.9 60.155 4.525 ;
      RECT 60.115 3.945 60.13 4.525 ;
      RECT 60.11 3.967 60.115 4.525 ;
      RECT 60.1 3.98 60.11 4.525 ;
      RECT 60.09 4.005 60.1 4.525 ;
      RECT 60.085 4.027 60.09 4.525 ;
      RECT 60.06 4.065 60.08 4.525 ;
      RECT 60.02 4.122 60.06 4.525 ;
      RECT 60.015 4.172 60.02 4.525 ;
      RECT 60.01 4.19 60.015 4.525 ;
      RECT 60.005 4.202 60.01 4.525 ;
      RECT 59.995 4.22 60.005 4.525 ;
      RECT 59.985 4.24 59.995 4.5 ;
      RECT 59.98 4.257 59.985 4.5 ;
      RECT 59.97 4.27 59.98 4.5 ;
      RECT 59.94 4.28 59.965 4.5 ;
      RECT 59.93 4.287 59.94 4.5 ;
      RECT 59.915 4.297 59.93 4.495 ;
      RECT 59.005 10.055 59.295 10.285 ;
      RECT 59.065 8.575 59.235 10.285 ;
      RECT 59.015 8.94 59.365 9.29 ;
      RECT 59.005 8.575 59.295 8.805 ;
      RECT 58.6 3.69 58.705 4.26 ;
      RECT 58.6 4.025 58.925 4.255 ;
      RECT 58.6 4.055 59.095 4.225 ;
      RECT 58.6 3.69 58.79 4.255 ;
      RECT 58.015 3.655 58.305 3.885 ;
      RECT 58.015 3.69 58.79 3.86 ;
      RECT 58.075 2.175 58.245 3.885 ;
      RECT 58.015 2.175 58.305 2.405 ;
      RECT 58.015 10.055 58.305 10.285 ;
      RECT 58.075 8.575 58.245 10.285 ;
      RECT 58.015 8.575 58.305 8.805 ;
      RECT 58.015 8.61 58.865 8.77 ;
      RECT 58.7 8.205 58.865 8.77 ;
      RECT 58.015 8.605 58.41 8.77 ;
      RECT 58.635 8.205 58.925 8.435 ;
      RECT 58.635 8.235 59.095 8.405 ;
      RECT 57.645 4.025 57.935 4.255 ;
      RECT 57.645 4.055 58.105 4.225 ;
      RECT 57.71 2.95 57.875 4.255 ;
      RECT 56.225 2.92 56.515 3.15 ;
      RECT 56.225 2.95 57.875 3.12 ;
      RECT 56.285 2.18 56.455 3.15 ;
      RECT 56.225 2.18 56.515 2.41 ;
      RECT 56.225 10.05 56.515 10.28 ;
      RECT 56.285 9.31 56.455 10.28 ;
      RECT 56.285 9.405 57.875 9.575 ;
      RECT 57.705 8.205 57.875 9.575 ;
      RECT 56.225 9.31 56.515 9.54 ;
      RECT 57.645 8.205 57.935 8.435 ;
      RECT 57.645 8.235 58.105 8.405 ;
      RECT 56.655 3.26 57.005 3.61 ;
      RECT 54.32 3.32 57.005 3.49 ;
      RECT 54.32 2.635 54.49 3.49 ;
      RECT 54.22 2.635 54.57 2.985 ;
      RECT 56.68 8.94 57.005 9.265 ;
      RECT 52.11 8.9 52.46 9.25 ;
      RECT 56.655 8.94 57.005 9.17 ;
      RECT 51.875 8.94 52.46 9.17 ;
      RECT 51.705 8.97 57.005 9.14 ;
      RECT 55.88 3.66 56.2 3.98 ;
      RECT 55.85 3.66 56.2 3.89 ;
      RECT 55.68 3.69 56.2 3.86 ;
      RECT 55.88 8.54 56.2 8.83 ;
      RECT 55.85 8.57 56.2 8.8 ;
      RECT 55.68 8.6 56.2 8.77 ;
      RECT 52.515 3.76 52.7 3.97 ;
      RECT 52.505 3.765 52.715 3.963 ;
      RECT 52.505 3.765 52.801 3.94 ;
      RECT 52.505 3.765 52.86 3.915 ;
      RECT 52.505 3.765 52.915 3.895 ;
      RECT 52.505 3.765 52.925 3.883 ;
      RECT 52.505 3.765 53.12 3.822 ;
      RECT 52.505 3.765 53.15 3.805 ;
      RECT 52.505 3.765 53.17 3.795 ;
      RECT 53.05 3.53 53.31 3.79 ;
      RECT 53.035 3.62 53.05 3.837 ;
      RECT 52.57 3.752 53.31 3.79 ;
      RECT 53.021 3.631 53.035 3.843 ;
      RECT 52.61 3.745 53.31 3.79 ;
      RECT 52.935 3.671 53.021 3.862 ;
      RECT 52.86 3.732 53.31 3.79 ;
      RECT 52.93 3.707 52.935 3.879 ;
      RECT 52.915 3.717 53.31 3.79 ;
      RECT 52.925 3.712 52.93 3.881 ;
      RECT 53.22 4.217 53.225 4.309 ;
      RECT 53.215 4.195 53.22 4.326 ;
      RECT 53.21 4.185 53.215 4.338 ;
      RECT 53.2 4.176 53.21 4.348 ;
      RECT 53.195 4.171 53.2 4.356 ;
      RECT 53.19 4.03 53.195 4.359 ;
      RECT 53.156 4.03 53.19 4.37 ;
      RECT 53.07 4.03 53.156 4.405 ;
      RECT 52.99 4.03 53.07 4.453 ;
      RECT 52.961 4.03 52.99 4.477 ;
      RECT 52.875 4.03 52.961 4.483 ;
      RECT 52.87 4.214 52.875 4.488 ;
      RECT 52.835 4.225 52.87 4.491 ;
      RECT 52.81 4.24 52.835 4.495 ;
      RECT 52.796 4.249 52.81 4.497 ;
      RECT 52.71 4.276 52.796 4.503 ;
      RECT 52.645 4.317 52.71 4.512 ;
      RECT 52.63 4.337 52.645 4.517 ;
      RECT 52.6 4.347 52.63 4.52 ;
      RECT 52.595 4.357 52.6 4.523 ;
      RECT 52.565 4.362 52.595 4.525 ;
      RECT 52.545 4.367 52.565 4.529 ;
      RECT 52.46 4.37 52.545 4.536 ;
      RECT 52.445 4.367 52.46 4.542 ;
      RECT 52.435 4.364 52.445 4.544 ;
      RECT 52.415 4.361 52.435 4.546 ;
      RECT 52.395 4.357 52.415 4.547 ;
      RECT 52.38 4.353 52.395 4.549 ;
      RECT 52.37 4.35 52.38 4.55 ;
      RECT 52.33 4.344 52.37 4.548 ;
      RECT 52.32 4.339 52.33 4.546 ;
      RECT 52.305 4.336 52.32 4.542 ;
      RECT 52.28 4.331 52.305 4.535 ;
      RECT 52.23 4.322 52.28 4.523 ;
      RECT 52.16 4.308 52.23 4.505 ;
      RECT 52.102 4.293 52.16 4.487 ;
      RECT 52.016 4.276 52.102 4.467 ;
      RECT 51.93 4.255 52.016 4.442 ;
      RECT 51.88 4.24 51.93 4.423 ;
      RECT 51.876 4.234 51.88 4.415 ;
      RECT 51.79 4.224 51.876 4.402 ;
      RECT 51.755 4.209 51.79 4.385 ;
      RECT 51.74 4.202 51.755 4.378 ;
      RECT 51.68 4.19 51.74 4.366 ;
      RECT 51.66 4.177 51.68 4.354 ;
      RECT 51.62 4.168 51.66 4.346 ;
      RECT 51.615 4.16 51.62 4.339 ;
      RECT 51.535 4.15 51.615 4.325 ;
      RECT 51.52 4.137 51.535 4.31 ;
      RECT 51.515 4.135 51.52 4.308 ;
      RECT 51.436 4.123 51.515 4.295 ;
      RECT 51.35 4.098 51.436 4.27 ;
      RECT 51.335 4.067 51.35 4.255 ;
      RECT 51.32 4.042 51.335 4.251 ;
      RECT 51.305 4.035 51.32 4.247 ;
      RECT 51.13 4.04 51.135 4.243 ;
      RECT 51.125 4.045 51.13 4.238 ;
      RECT 51.135 4.035 51.305 4.245 ;
      RECT 51.85 3.795 51.955 4.055 ;
      RECT 52.665 3.32 52.67 3.545 ;
      RECT 52.795 3.32 52.85 3.53 ;
      RECT 52.85 3.325 52.86 3.523 ;
      RECT 52.756 3.32 52.795 3.533 ;
      RECT 52.67 3.32 52.756 3.54 ;
      RECT 52.65 3.325 52.665 3.546 ;
      RECT 52.64 3.365 52.65 3.548 ;
      RECT 52.61 3.375 52.64 3.55 ;
      RECT 52.605 3.38 52.61 3.552 ;
      RECT 52.58 3.385 52.605 3.554 ;
      RECT 52.565 3.39 52.58 3.556 ;
      RECT 52.55 3.392 52.565 3.558 ;
      RECT 52.545 3.397 52.55 3.56 ;
      RECT 52.495 3.405 52.545 3.563 ;
      RECT 52.47 3.414 52.495 3.568 ;
      RECT 52.46 3.421 52.47 3.573 ;
      RECT 52.455 3.424 52.46 3.577 ;
      RECT 52.435 3.427 52.455 3.586 ;
      RECT 52.405 3.435 52.435 3.606 ;
      RECT 52.376 3.448 52.405 3.628 ;
      RECT 52.29 3.482 52.376 3.672 ;
      RECT 52.285 3.508 52.29 3.71 ;
      RECT 52.28 3.512 52.285 3.719 ;
      RECT 52.245 3.525 52.28 3.752 ;
      RECT 52.235 3.539 52.245 3.79 ;
      RECT 52.23 3.543 52.235 3.803 ;
      RECT 52.225 3.547 52.23 3.808 ;
      RECT 52.215 3.555 52.225 3.82 ;
      RECT 52.21 3.562 52.215 3.835 ;
      RECT 52.185 3.575 52.21 3.86 ;
      RECT 52.145 3.604 52.185 3.915 ;
      RECT 52.13 3.629 52.145 3.97 ;
      RECT 52.12 3.64 52.13 3.993 ;
      RECT 52.115 3.647 52.12 4.005 ;
      RECT 52.11 3.651 52.115 4.013 ;
      RECT 52.055 3.679 52.11 4.055 ;
      RECT 52.035 3.715 52.055 4.055 ;
      RECT 52.02 3.73 52.035 4.055 ;
      RECT 51.965 3.762 52.02 4.055 ;
      RECT 51.955 3.792 51.965 4.055 ;
      RECT 51.565 3.407 51.75 3.645 ;
      RECT 51.55 3.409 51.76 3.64 ;
      RECT 51.435 3.355 51.695 3.615 ;
      RECT 51.43 3.392 51.695 3.569 ;
      RECT 51.425 3.402 51.695 3.566 ;
      RECT 51.42 3.442 51.76 3.56 ;
      RECT 51.415 3.475 51.76 3.55 ;
      RECT 51.425 3.417 51.775 3.488 ;
      RECT 51.722 4.515 51.735 5.045 ;
      RECT 51.636 4.515 51.735 5.044 ;
      RECT 51.636 4.515 51.74 5.043 ;
      RECT 51.55 4.515 51.74 5.041 ;
      RECT 51.545 4.515 51.74 5.038 ;
      RECT 51.545 4.515 51.75 5.036 ;
      RECT 51.54 4.807 51.75 5.033 ;
      RECT 51.54 4.817 51.755 5.03 ;
      RECT 51.54 4.885 51.76 5.026 ;
      RECT 51.53 4.89 51.76 5.025 ;
      RECT 51.53 4.982 51.765 5.022 ;
      RECT 51.515 4.515 51.775 4.775 ;
      RECT 51.445 10.05 51.735 10.28 ;
      RECT 51.505 9.31 51.675 10.28 ;
      RECT 51.42 9.34 51.76 9.685 ;
      RECT 51.445 9.31 51.735 9.685 ;
      RECT 50.745 3.505 50.79 5.04 ;
      RECT 50.945 3.505 50.975 3.72 ;
      RECT 49.32 3.245 49.44 3.455 ;
      RECT 48.98 3.195 49.24 3.455 ;
      RECT 48.98 3.24 49.275 3.445 ;
      RECT 50.985 3.521 50.99 3.575 ;
      RECT 50.98 3.514 50.985 3.708 ;
      RECT 50.975 3.508 50.98 3.715 ;
      RECT 50.93 3.505 50.945 3.728 ;
      RECT 50.925 3.505 50.93 3.75 ;
      RECT 50.92 3.505 50.925 3.798 ;
      RECT 50.915 3.505 50.92 3.818 ;
      RECT 50.905 3.505 50.915 3.925 ;
      RECT 50.9 3.505 50.905 3.988 ;
      RECT 50.895 3.505 50.9 4.045 ;
      RECT 50.89 3.505 50.895 4.053 ;
      RECT 50.875 3.505 50.89 4.16 ;
      RECT 50.865 3.505 50.875 4.295 ;
      RECT 50.855 3.505 50.865 4.405 ;
      RECT 50.845 3.505 50.855 4.462 ;
      RECT 50.84 3.505 50.845 4.502 ;
      RECT 50.835 3.505 50.84 4.538 ;
      RECT 50.825 3.505 50.835 4.578 ;
      RECT 50.82 3.505 50.825 4.62 ;
      RECT 50.8 3.505 50.82 4.685 ;
      RECT 50.805 4.83 50.81 5.01 ;
      RECT 50.8 4.812 50.805 5.018 ;
      RECT 50.795 3.505 50.8 4.748 ;
      RECT 50.795 4.792 50.8 5.025 ;
      RECT 50.79 3.505 50.795 5.035 ;
      RECT 50.735 3.505 50.745 3.805 ;
      RECT 50.74 4.052 50.745 5.04 ;
      RECT 50.735 4.117 50.74 5.04 ;
      RECT 50.73 3.506 50.735 3.795 ;
      RECT 50.725 4.182 50.735 5.04 ;
      RECT 50.72 3.507 50.73 3.785 ;
      RECT 50.71 4.295 50.725 5.04 ;
      RECT 50.715 3.508 50.72 3.775 ;
      RECT 50.695 3.509 50.715 3.753 ;
      RECT 50.7 4.392 50.71 5.04 ;
      RECT 50.695 4.467 50.7 5.04 ;
      RECT 50.685 3.508 50.695 3.73 ;
      RECT 50.69 4.51 50.695 5.04 ;
      RECT 50.685 4.537 50.69 5.04 ;
      RECT 50.675 3.506 50.685 3.718 ;
      RECT 50.68 4.58 50.685 5.04 ;
      RECT 50.675 4.607 50.68 5.04 ;
      RECT 50.665 3.505 50.675 3.705 ;
      RECT 50.67 4.622 50.675 5.04 ;
      RECT 50.63 4.68 50.67 5.04 ;
      RECT 50.66 3.504 50.665 3.69 ;
      RECT 50.655 3.502 50.66 3.683 ;
      RECT 50.645 3.499 50.655 3.673 ;
      RECT 50.64 3.496 50.645 3.658 ;
      RECT 50.625 3.492 50.64 3.651 ;
      RECT 50.62 4.735 50.63 5.04 ;
      RECT 50.62 3.489 50.625 3.646 ;
      RECT 50.605 3.485 50.62 3.64 ;
      RECT 50.615 4.752 50.62 5.04 ;
      RECT 50.605 4.815 50.615 5.04 ;
      RECT 50.525 3.47 50.605 3.62 ;
      RECT 50.6 4.822 50.605 5.035 ;
      RECT 50.595 4.83 50.6 5.025 ;
      RECT 50.515 3.456 50.525 3.604 ;
      RECT 50.5 3.452 50.515 3.602 ;
      RECT 50.49 3.447 50.5 3.598 ;
      RECT 50.465 3.44 50.49 3.59 ;
      RECT 50.46 3.435 50.465 3.585 ;
      RECT 50.45 3.435 50.46 3.583 ;
      RECT 50.44 3.433 50.45 3.581 ;
      RECT 50.41 3.425 50.44 3.575 ;
      RECT 50.395 3.417 50.41 3.568 ;
      RECT 50.375 3.412 50.395 3.561 ;
      RECT 50.37 3.408 50.375 3.556 ;
      RECT 50.34 3.401 50.37 3.55 ;
      RECT 50.315 3.392 50.34 3.54 ;
      RECT 50.285 3.385 50.315 3.532 ;
      RECT 50.26 3.375 50.285 3.523 ;
      RECT 50.245 3.367 50.26 3.517 ;
      RECT 50.22 3.362 50.245 3.512 ;
      RECT 50.21 3.358 50.22 3.507 ;
      RECT 50.19 3.353 50.21 3.502 ;
      RECT 50.155 3.348 50.19 3.495 ;
      RECT 50.095 3.343 50.155 3.488 ;
      RECT 50.082 3.339 50.095 3.486 ;
      RECT 49.996 3.334 50.082 3.483 ;
      RECT 49.91 3.324 49.996 3.479 ;
      RECT 49.869 3.317 49.91 3.476 ;
      RECT 49.783 3.31 49.869 3.473 ;
      RECT 49.697 3.3 49.783 3.469 ;
      RECT 49.611 3.29 49.697 3.464 ;
      RECT 49.525 3.28 49.611 3.46 ;
      RECT 49.515 3.265 49.525 3.458 ;
      RECT 49.505 3.25 49.515 3.458 ;
      RECT 49.44 3.245 49.505 3.457 ;
      RECT 49.275 3.242 49.32 3.45 ;
      RECT 50.52 4.147 50.525 4.338 ;
      RECT 50.515 4.142 50.52 4.345 ;
      RECT 50.501 4.14 50.515 4.351 ;
      RECT 50.415 4.14 50.501 4.353 ;
      RECT 50.411 4.14 50.415 4.356 ;
      RECT 50.325 4.14 50.411 4.374 ;
      RECT 50.315 4.145 50.325 4.393 ;
      RECT 50.305 4.2 50.315 4.397 ;
      RECT 50.28 4.215 50.305 4.404 ;
      RECT 50.24 4.235 50.28 4.417 ;
      RECT 50.235 4.247 50.24 4.427 ;
      RECT 50.22 4.253 50.235 4.432 ;
      RECT 50.215 4.258 50.22 4.436 ;
      RECT 50.195 4.265 50.215 4.441 ;
      RECT 50.125 4.29 50.195 4.458 ;
      RECT 50.085 4.318 50.125 4.478 ;
      RECT 50.08 4.328 50.085 4.486 ;
      RECT 50.06 4.335 50.08 4.488 ;
      RECT 50.055 4.342 50.06 4.491 ;
      RECT 50.025 4.35 50.055 4.494 ;
      RECT 50.02 4.355 50.025 4.498 ;
      RECT 49.946 4.359 50.02 4.506 ;
      RECT 49.86 4.368 49.946 4.522 ;
      RECT 49.856 4.373 49.86 4.531 ;
      RECT 49.77 4.378 49.856 4.541 ;
      RECT 49.73 4.386 49.77 4.553 ;
      RECT 49.68 4.392 49.73 4.56 ;
      RECT 49.595 4.401 49.68 4.575 ;
      RECT 49.52 4.412 49.595 4.593 ;
      RECT 49.485 4.419 49.52 4.603 ;
      RECT 49.41 4.427 49.485 4.608 ;
      RECT 49.355 4.436 49.41 4.608 ;
      RECT 49.33 4.441 49.355 4.606 ;
      RECT 49.32 4.444 49.33 4.604 ;
      RECT 49.285 4.446 49.32 4.602 ;
      RECT 49.255 4.448 49.285 4.598 ;
      RECT 49.21 4.447 49.255 4.594 ;
      RECT 49.19 4.442 49.21 4.591 ;
      RECT 49.14 4.427 49.19 4.588 ;
      RECT 49.13 4.412 49.14 4.583 ;
      RECT 49.08 4.397 49.13 4.573 ;
      RECT 49.03 4.372 49.08 4.553 ;
      RECT 49.02 4.357 49.03 4.535 ;
      RECT 49.015 4.355 49.02 4.529 ;
      RECT 48.995 4.35 49.015 4.524 ;
      RECT 48.99 4.342 48.995 4.518 ;
      RECT 48.975 4.336 48.99 4.511 ;
      RECT 48.97 4.331 48.975 4.503 ;
      RECT 48.95 4.326 48.97 4.495 ;
      RECT 48.935 4.319 48.95 4.488 ;
      RECT 48.92 4.313 48.935 4.479 ;
      RECT 48.915 4.307 48.92 4.472 ;
      RECT 48.87 4.282 48.915 4.458 ;
      RECT 48.855 4.252 48.87 4.44 ;
      RECT 48.84 4.235 48.855 4.431 ;
      RECT 48.815 4.215 48.84 4.419 ;
      RECT 48.775 4.185 48.815 4.399 ;
      RECT 48.765 4.155 48.775 4.384 ;
      RECT 48.75 4.145 48.765 4.377 ;
      RECT 48.695 4.11 48.75 4.356 ;
      RECT 48.68 4.073 48.695 4.335 ;
      RECT 48.67 4.06 48.68 4.327 ;
      RECT 48.62 4.03 48.67 4.309 ;
      RECT 48.605 3.96 48.62 4.29 ;
      RECT 48.56 3.96 48.605 4.273 ;
      RECT 48.535 3.96 48.56 4.255 ;
      RECT 48.525 3.96 48.535 4.248 ;
      RECT 48.446 3.96 48.525 4.241 ;
      RECT 48.36 3.96 48.446 4.233 ;
      RECT 48.345 3.992 48.36 4.228 ;
      RECT 48.27 4.002 48.345 4.224 ;
      RECT 48.25 4.012 48.27 4.219 ;
      RECT 48.225 4.012 48.25 4.216 ;
      RECT 48.215 4.002 48.225 4.215 ;
      RECT 48.205 3.975 48.215 4.214 ;
      RECT 48.165 3.97 48.205 4.212 ;
      RECT 48.12 3.97 48.165 4.208 ;
      RECT 48.095 3.97 48.12 4.203 ;
      RECT 48.045 3.97 48.095 4.19 ;
      RECT 48.005 3.975 48.015 4.175 ;
      RECT 48.015 3.97 48.045 4.18 ;
      RECT 50 3.75 50.26 4.01 ;
      RECT 49.995 3.772 50.26 3.968 ;
      RECT 49.235 3.6 49.455 3.965 ;
      RECT 49.217 3.687 49.455 3.964 ;
      RECT 49.2 3.692 49.455 3.961 ;
      RECT 49.2 3.692 49.475 3.96 ;
      RECT 49.17 3.702 49.475 3.958 ;
      RECT 49.165 3.717 49.475 3.954 ;
      RECT 49.165 3.717 49.48 3.953 ;
      RECT 49.16 3.775 49.48 3.951 ;
      RECT 49.16 3.775 49.49 3.948 ;
      RECT 49.155 3.84 49.49 3.943 ;
      RECT 49.235 3.6 49.495 3.86 ;
      RECT 47.98 3.43 48.24 3.69 ;
      RECT 47.98 3.473 48.326 3.664 ;
      RECT 47.98 3.473 48.37 3.663 ;
      RECT 47.98 3.473 48.39 3.661 ;
      RECT 47.98 3.473 48.49 3.66 ;
      RECT 47.98 3.473 48.51 3.658 ;
      RECT 47.98 3.473 48.52 3.653 ;
      RECT 48.39 3.44 48.58 3.65 ;
      RECT 48.39 3.442 48.585 3.648 ;
      RECT 48.38 3.447 48.59 3.64 ;
      RECT 48.326 3.471 48.59 3.64 ;
      RECT 48.37 3.465 48.38 3.662 ;
      RECT 48.38 3.445 48.585 3.648 ;
      RECT 47.335 4.505 47.54 4.735 ;
      RECT 47.275 4.455 47.33 4.715 ;
      RECT 47.335 4.455 47.535 4.735 ;
      RECT 48.305 4.77 48.31 4.797 ;
      RECT 48.295 4.68 48.305 4.802 ;
      RECT 48.29 4.602 48.295 4.808 ;
      RECT 48.28 4.592 48.29 4.815 ;
      RECT 48.275 4.582 48.28 4.821 ;
      RECT 48.265 4.577 48.275 4.823 ;
      RECT 48.25 4.569 48.265 4.831 ;
      RECT 48.235 4.56 48.25 4.843 ;
      RECT 48.225 4.552 48.235 4.853 ;
      RECT 48.19 4.47 48.225 4.871 ;
      RECT 48.155 4.47 48.19 4.89 ;
      RECT 48.14 4.47 48.155 4.898 ;
      RECT 48.085 4.47 48.14 4.898 ;
      RECT 48.051 4.47 48.085 4.889 ;
      RECT 47.965 4.47 48.051 4.865 ;
      RECT 47.955 4.53 47.965 4.847 ;
      RECT 47.915 4.532 47.955 4.838 ;
      RECT 47.91 4.534 47.915 4.828 ;
      RECT 47.89 4.536 47.91 4.823 ;
      RECT 47.88 4.539 47.89 4.818 ;
      RECT 47.87 4.54 47.88 4.813 ;
      RECT 47.846 4.541 47.87 4.805 ;
      RECT 47.76 4.546 47.846 4.783 ;
      RECT 47.705 4.545 47.76 4.756 ;
      RECT 47.69 4.538 47.705 4.743 ;
      RECT 47.655 4.533 47.69 4.739 ;
      RECT 47.6 4.525 47.655 4.738 ;
      RECT 47.54 4.512 47.6 4.736 ;
      RECT 47.33 4.455 47.335 4.723 ;
      RECT 47.405 3.825 47.59 4.035 ;
      RECT 47.395 3.83 47.605 4.028 ;
      RECT 47.435 3.735 47.695 3.995 ;
      RECT 47.39 3.892 47.695 3.918 ;
      RECT 46.735 3.685 46.74 4.485 ;
      RECT 46.68 3.735 46.71 4.485 ;
      RECT 46.67 3.735 46.675 4.045 ;
      RECT 46.655 3.735 46.66 4.04 ;
      RECT 46.2 3.78 46.215 3.995 ;
      RECT 46.13 3.78 46.215 3.99 ;
      RECT 47.395 3.36 47.465 3.57 ;
      RECT 47.465 3.367 47.475 3.565 ;
      RECT 47.361 3.36 47.395 3.577 ;
      RECT 47.275 3.36 47.361 3.601 ;
      RECT 47.265 3.365 47.275 3.62 ;
      RECT 47.26 3.377 47.265 3.623 ;
      RECT 47.245 3.392 47.26 3.627 ;
      RECT 47.24 3.41 47.245 3.631 ;
      RECT 47.2 3.42 47.24 3.64 ;
      RECT 47.185 3.427 47.2 3.652 ;
      RECT 47.17 3.432 47.185 3.657 ;
      RECT 47.155 3.435 47.17 3.662 ;
      RECT 47.145 3.437 47.155 3.666 ;
      RECT 47.11 3.444 47.145 3.674 ;
      RECT 47.075 3.452 47.11 3.688 ;
      RECT 47.065 3.458 47.075 3.697 ;
      RECT 47.06 3.46 47.065 3.699 ;
      RECT 47.04 3.463 47.06 3.705 ;
      RECT 47.01 3.47 47.04 3.716 ;
      RECT 47 3.476 47.01 3.723 ;
      RECT 46.975 3.479 47 3.73 ;
      RECT 46.965 3.483 46.975 3.738 ;
      RECT 46.96 3.484 46.965 3.76 ;
      RECT 46.955 3.485 46.96 3.775 ;
      RECT 46.95 3.486 46.955 3.79 ;
      RECT 46.945 3.487 46.95 3.805 ;
      RECT 46.94 3.488 46.945 3.835 ;
      RECT 46.93 3.49 46.94 3.868 ;
      RECT 46.915 3.494 46.93 3.915 ;
      RECT 46.905 3.497 46.915 3.96 ;
      RECT 46.9 3.5 46.905 3.988 ;
      RECT 46.89 3.502 46.9 4.015 ;
      RECT 46.885 3.505 46.89 4.05 ;
      RECT 46.855 3.51 46.885 4.108 ;
      RECT 46.85 3.515 46.855 4.193 ;
      RECT 46.845 3.517 46.85 4.228 ;
      RECT 46.84 3.519 46.845 4.31 ;
      RECT 46.835 3.521 46.84 4.398 ;
      RECT 46.825 3.523 46.835 4.48 ;
      RECT 46.81 3.537 46.825 4.485 ;
      RECT 46.775 3.582 46.81 4.485 ;
      RECT 46.765 3.622 46.775 4.485 ;
      RECT 46.75 3.65 46.765 4.485 ;
      RECT 46.745 3.667 46.75 4.485 ;
      RECT 46.74 3.675 46.745 4.485 ;
      RECT 46.73 3.69 46.735 4.485 ;
      RECT 46.725 3.697 46.73 4.485 ;
      RECT 46.715 3.717 46.725 4.485 ;
      RECT 46.71 3.73 46.715 4.485 ;
      RECT 46.675 3.735 46.68 4.07 ;
      RECT 46.66 4.125 46.68 4.485 ;
      RECT 46.66 3.735 46.67 4.043 ;
      RECT 46.655 4.165 46.66 4.485 ;
      RECT 46.605 3.735 46.655 4.038 ;
      RECT 46.65 4.202 46.655 4.485 ;
      RECT 46.64 4.225 46.65 4.485 ;
      RECT 46.635 4.27 46.64 4.485 ;
      RECT 46.625 4.28 46.635 4.478 ;
      RECT 46.551 3.735 46.605 4.032 ;
      RECT 46.465 3.735 46.551 4.025 ;
      RECT 46.416 3.782 46.465 4.018 ;
      RECT 46.33 3.79 46.416 4.011 ;
      RECT 46.315 3.787 46.33 4.006 ;
      RECT 46.301 3.78 46.315 4.005 ;
      RECT 46.215 3.78 46.301 4 ;
      RECT 46.12 3.785 46.13 3.985 ;
      RECT 45.71 3.215 45.725 3.615 ;
      RECT 45.905 3.215 45.91 3.475 ;
      RECT 45.65 3.215 45.695 3.475 ;
      RECT 46.105 4.52 46.11 4.725 ;
      RECT 46.1 4.51 46.105 4.73 ;
      RECT 46.095 4.497 46.1 4.735 ;
      RECT 46.09 4.477 46.095 4.735 ;
      RECT 46.065 4.43 46.09 4.735 ;
      RECT 46.03 4.345 46.065 4.735 ;
      RECT 46.025 4.282 46.03 4.735 ;
      RECT 46.02 4.267 46.025 4.735 ;
      RECT 46.005 4.227 46.02 4.735 ;
      RECT 46 4.202 46.005 4.735 ;
      RECT 45.99 4.185 46 4.735 ;
      RECT 45.955 4.107 45.99 4.735 ;
      RECT 45.95 4.05 45.955 4.735 ;
      RECT 45.945 4.037 45.95 4.735 ;
      RECT 45.935 4.015 45.945 4.735 ;
      RECT 45.925 3.98 45.935 4.735 ;
      RECT 45.915 3.95 45.925 4.735 ;
      RECT 45.905 3.865 45.915 4.378 ;
      RECT 45.912 4.51 45.915 4.735 ;
      RECT 45.91 4.52 45.912 4.735 ;
      RECT 45.9 4.53 45.91 4.73 ;
      RECT 45.895 3.215 45.905 3.61 ;
      RECT 45.9 3.742 45.905 4.353 ;
      RECT 45.895 3.64 45.9 4.336 ;
      RECT 45.885 3.215 45.895 4.312 ;
      RECT 45.88 3.215 45.885 4.283 ;
      RECT 45.875 3.215 45.88 4.273 ;
      RECT 45.855 3.215 45.875 4.235 ;
      RECT 45.85 3.215 45.855 4.193 ;
      RECT 45.845 3.215 45.85 4.173 ;
      RECT 45.815 3.215 45.845 4.123 ;
      RECT 45.805 3.215 45.815 4.07 ;
      RECT 45.8 3.215 45.805 4.043 ;
      RECT 45.795 3.215 45.8 4.028 ;
      RECT 45.785 3.215 45.795 4.005 ;
      RECT 45.775 3.215 45.785 3.98 ;
      RECT 45.77 3.215 45.775 3.92 ;
      RECT 45.76 3.215 45.77 3.858 ;
      RECT 45.755 3.215 45.76 3.778 ;
      RECT 45.75 3.215 45.755 3.743 ;
      RECT 45.745 3.215 45.75 3.718 ;
      RECT 45.74 3.215 45.745 3.703 ;
      RECT 45.735 3.215 45.74 3.673 ;
      RECT 45.73 3.215 45.735 3.65 ;
      RECT 45.725 3.215 45.73 3.623 ;
      RECT 45.695 3.215 45.71 3.61 ;
      RECT 44.85 4.75 45.035 4.96 ;
      RECT 44.84 4.755 45.05 4.953 ;
      RECT 44.84 4.755 45.07 4.925 ;
      RECT 44.84 4.755 45.085 4.904 ;
      RECT 44.84 4.755 45.1 4.902 ;
      RECT 44.84 4.755 45.11 4.901 ;
      RECT 44.84 4.755 45.14 4.898 ;
      RECT 45.49 4.6 45.75 4.86 ;
      RECT 45.45 4.647 45.75 4.843 ;
      RECT 45.441 4.655 45.45 4.846 ;
      RECT 45.035 4.748 45.75 4.843 ;
      RECT 45.355 4.673 45.441 4.853 ;
      RECT 45.05 4.745 45.75 4.843 ;
      RECT 45.296 4.695 45.355 4.865 ;
      RECT 45.07 4.741 45.75 4.843 ;
      RECT 45.21 4.707 45.296 4.876 ;
      RECT 45.085 4.737 45.75 4.843 ;
      RECT 45.155 4.72 45.21 4.888 ;
      RECT 45.1 4.735 45.75 4.843 ;
      RECT 45.14 4.726 45.155 4.894 ;
      RECT 45.11 4.731 45.75 4.843 ;
      RECT 45.255 4.255 45.515 4.515 ;
      RECT 45.255 4.275 45.625 4.485 ;
      RECT 45.255 4.28 45.635 4.48 ;
      RECT 45.446 3.694 45.525 3.925 ;
      RECT 45.36 3.697 45.575 3.92 ;
      RECT 45.355 3.697 45.575 3.915 ;
      RECT 45.355 3.702 45.585 3.913 ;
      RECT 45.33 3.702 45.585 3.91 ;
      RECT 45.33 3.71 45.595 3.908 ;
      RECT 45.21 3.645 45.47 3.905 ;
      RECT 45.21 3.692 45.52 3.905 ;
      RECT 44.465 4.265 44.47 4.525 ;
      RECT 44.295 4.035 44.3 4.525 ;
      RECT 44.18 4.275 44.185 4.5 ;
      RECT 44.89 3.37 44.895 3.58 ;
      RECT 44.895 3.375 44.91 3.575 ;
      RECT 44.83 3.37 44.89 3.588 ;
      RECT 44.815 3.37 44.83 3.598 ;
      RECT 44.765 3.37 44.815 3.615 ;
      RECT 44.745 3.37 44.765 3.638 ;
      RECT 44.73 3.37 44.745 3.65 ;
      RECT 44.71 3.37 44.73 3.66 ;
      RECT 44.7 3.375 44.71 3.669 ;
      RECT 44.695 3.385 44.7 3.674 ;
      RECT 44.69 3.397 44.695 3.678 ;
      RECT 44.68 3.42 44.69 3.683 ;
      RECT 44.675 3.435 44.68 3.687 ;
      RECT 44.67 3.452 44.675 3.69 ;
      RECT 44.665 3.46 44.67 3.693 ;
      RECT 44.655 3.465 44.665 3.697 ;
      RECT 44.65 3.472 44.655 3.702 ;
      RECT 44.64 3.477 44.65 3.706 ;
      RECT 44.615 3.489 44.64 3.717 ;
      RECT 44.595 3.506 44.615 3.733 ;
      RECT 44.57 3.523 44.595 3.755 ;
      RECT 44.535 3.546 44.57 3.813 ;
      RECT 44.515 3.568 44.535 3.875 ;
      RECT 44.51 3.578 44.515 3.91 ;
      RECT 44.5 3.585 44.51 3.948 ;
      RECT 44.495 3.592 44.5 3.968 ;
      RECT 44.49 3.603 44.495 4.005 ;
      RECT 44.485 3.611 44.49 4.07 ;
      RECT 44.475 3.622 44.485 4.123 ;
      RECT 44.47 3.64 44.475 4.193 ;
      RECT 44.465 3.65 44.47 4.23 ;
      RECT 44.46 3.66 44.465 4.525 ;
      RECT 44.455 3.672 44.46 4.525 ;
      RECT 44.45 3.682 44.455 4.525 ;
      RECT 44.44 3.692 44.45 4.525 ;
      RECT 44.43 3.715 44.44 4.525 ;
      RECT 44.415 3.75 44.43 4.525 ;
      RECT 44.375 3.812 44.415 4.525 ;
      RECT 44.37 3.865 44.375 4.525 ;
      RECT 44.345 3.9 44.37 4.525 ;
      RECT 44.33 3.945 44.345 4.525 ;
      RECT 44.325 3.967 44.33 4.525 ;
      RECT 44.315 3.98 44.325 4.525 ;
      RECT 44.305 4.005 44.315 4.525 ;
      RECT 44.3 4.027 44.305 4.525 ;
      RECT 44.275 4.065 44.295 4.525 ;
      RECT 44.235 4.122 44.275 4.525 ;
      RECT 44.23 4.172 44.235 4.525 ;
      RECT 44.225 4.19 44.23 4.525 ;
      RECT 44.22 4.202 44.225 4.525 ;
      RECT 44.21 4.22 44.22 4.525 ;
      RECT 44.2 4.24 44.21 4.5 ;
      RECT 44.195 4.257 44.2 4.5 ;
      RECT 44.185 4.27 44.195 4.5 ;
      RECT 44.155 4.28 44.18 4.5 ;
      RECT 44.145 4.287 44.155 4.5 ;
      RECT 44.13 4.297 44.145 4.495 ;
      RECT 43.23 10.055 43.52 10.285 ;
      RECT 43.29 8.575 43.46 10.285 ;
      RECT 43.28 8.945 43.635 9.3 ;
      RECT 43.23 8.575 43.52 8.805 ;
      RECT 42.825 3.69 42.93 4.26 ;
      RECT 42.825 4.025 43.15 4.255 ;
      RECT 42.825 4.055 43.32 4.225 ;
      RECT 42.825 3.69 43.015 4.255 ;
      RECT 42.24 3.655 42.53 3.885 ;
      RECT 42.24 3.69 43.015 3.86 ;
      RECT 42.3 2.175 42.47 3.885 ;
      RECT 42.24 2.175 42.53 2.405 ;
      RECT 42.24 10.055 42.53 10.285 ;
      RECT 42.3 8.575 42.47 10.285 ;
      RECT 42.24 8.575 42.53 8.805 ;
      RECT 42.24 8.61 43.09 8.77 ;
      RECT 42.925 8.205 43.09 8.77 ;
      RECT 42.24 8.605 42.635 8.77 ;
      RECT 42.86 8.205 43.15 8.435 ;
      RECT 42.86 8.235 43.32 8.405 ;
      RECT 41.87 4.025 42.16 4.255 ;
      RECT 41.87 4.055 42.33 4.225 ;
      RECT 41.935 2.95 42.1 4.255 ;
      RECT 40.45 2.92 40.74 3.15 ;
      RECT 40.45 2.95 42.1 3.12 ;
      RECT 40.51 2.18 40.68 3.15 ;
      RECT 40.45 2.18 40.74 2.41 ;
      RECT 40.45 10.05 40.74 10.28 ;
      RECT 40.51 9.31 40.68 10.28 ;
      RECT 40.51 9.405 42.1 9.575 ;
      RECT 41.93 8.205 42.1 9.575 ;
      RECT 40.45 9.31 40.74 9.54 ;
      RECT 41.87 8.205 42.16 8.435 ;
      RECT 41.87 8.235 42.33 8.405 ;
      RECT 40.88 3.26 41.23 3.61 ;
      RECT 38.545 3.32 41.23 3.49 ;
      RECT 38.545 2.635 38.715 3.49 ;
      RECT 38.445 2.635 38.795 2.985 ;
      RECT 40.905 8.94 41.23 9.265 ;
      RECT 36.33 8.895 36.68 9.245 ;
      RECT 40.88 8.94 41.23 9.17 ;
      RECT 36.1 8.94 36.68 9.17 ;
      RECT 35.93 8.97 41.23 9.14 ;
      RECT 40.105 3.66 40.425 3.98 ;
      RECT 40.075 3.66 40.425 3.89 ;
      RECT 39.905 3.69 40.425 3.86 ;
      RECT 40.105 8.54 40.425 8.83 ;
      RECT 40.075 8.57 40.425 8.8 ;
      RECT 39.905 8.6 40.425 8.77 ;
      RECT 36.74 3.76 36.925 3.97 ;
      RECT 36.73 3.765 36.94 3.963 ;
      RECT 36.73 3.765 37.026 3.94 ;
      RECT 36.73 3.765 37.085 3.915 ;
      RECT 36.73 3.765 37.14 3.895 ;
      RECT 36.73 3.765 37.15 3.883 ;
      RECT 36.73 3.765 37.345 3.822 ;
      RECT 36.73 3.765 37.375 3.805 ;
      RECT 36.73 3.765 37.395 3.795 ;
      RECT 37.275 3.53 37.535 3.79 ;
      RECT 37.26 3.62 37.275 3.837 ;
      RECT 36.795 3.752 37.535 3.79 ;
      RECT 37.246 3.631 37.26 3.843 ;
      RECT 36.835 3.745 37.535 3.79 ;
      RECT 37.16 3.671 37.246 3.862 ;
      RECT 37.085 3.732 37.535 3.79 ;
      RECT 37.155 3.707 37.16 3.879 ;
      RECT 37.14 3.717 37.535 3.79 ;
      RECT 37.15 3.712 37.155 3.881 ;
      RECT 37.445 4.217 37.45 4.309 ;
      RECT 37.44 4.195 37.445 4.326 ;
      RECT 37.435 4.185 37.44 4.338 ;
      RECT 37.425 4.176 37.435 4.348 ;
      RECT 37.42 4.171 37.425 4.356 ;
      RECT 37.415 4.03 37.42 4.359 ;
      RECT 37.381 4.03 37.415 4.37 ;
      RECT 37.295 4.03 37.381 4.405 ;
      RECT 37.215 4.03 37.295 4.453 ;
      RECT 37.186 4.03 37.215 4.477 ;
      RECT 37.1 4.03 37.186 4.483 ;
      RECT 37.095 4.214 37.1 4.488 ;
      RECT 37.06 4.225 37.095 4.491 ;
      RECT 37.035 4.24 37.06 4.495 ;
      RECT 37.021 4.249 37.035 4.497 ;
      RECT 36.935 4.276 37.021 4.503 ;
      RECT 36.87 4.317 36.935 4.512 ;
      RECT 36.855 4.337 36.87 4.517 ;
      RECT 36.825 4.347 36.855 4.52 ;
      RECT 36.82 4.357 36.825 4.523 ;
      RECT 36.79 4.362 36.82 4.525 ;
      RECT 36.77 4.367 36.79 4.529 ;
      RECT 36.685 4.37 36.77 4.536 ;
      RECT 36.67 4.367 36.685 4.542 ;
      RECT 36.66 4.364 36.67 4.544 ;
      RECT 36.64 4.361 36.66 4.546 ;
      RECT 36.62 4.357 36.64 4.547 ;
      RECT 36.605 4.353 36.62 4.549 ;
      RECT 36.595 4.35 36.605 4.55 ;
      RECT 36.555 4.344 36.595 4.548 ;
      RECT 36.545 4.339 36.555 4.546 ;
      RECT 36.53 4.336 36.545 4.542 ;
      RECT 36.505 4.331 36.53 4.535 ;
      RECT 36.455 4.322 36.505 4.523 ;
      RECT 36.385 4.308 36.455 4.505 ;
      RECT 36.327 4.293 36.385 4.487 ;
      RECT 36.241 4.276 36.327 4.467 ;
      RECT 36.155 4.255 36.241 4.442 ;
      RECT 36.105 4.24 36.155 4.423 ;
      RECT 36.101 4.234 36.105 4.415 ;
      RECT 36.015 4.224 36.101 4.402 ;
      RECT 35.98 4.209 36.015 4.385 ;
      RECT 35.965 4.202 35.98 4.378 ;
      RECT 35.905 4.19 35.965 4.366 ;
      RECT 35.885 4.177 35.905 4.354 ;
      RECT 35.845 4.168 35.885 4.346 ;
      RECT 35.84 4.16 35.845 4.339 ;
      RECT 35.76 4.15 35.84 4.325 ;
      RECT 35.745 4.137 35.76 4.31 ;
      RECT 35.74 4.135 35.745 4.308 ;
      RECT 35.661 4.123 35.74 4.295 ;
      RECT 35.575 4.098 35.661 4.27 ;
      RECT 35.56 4.067 35.575 4.255 ;
      RECT 35.545 4.042 35.56 4.251 ;
      RECT 35.53 4.035 35.545 4.247 ;
      RECT 35.355 4.04 35.36 4.243 ;
      RECT 35.35 4.045 35.355 4.238 ;
      RECT 35.36 4.035 35.53 4.245 ;
      RECT 36.075 3.795 36.18 4.055 ;
      RECT 36.89 3.32 36.895 3.545 ;
      RECT 37.02 3.32 37.075 3.53 ;
      RECT 37.075 3.325 37.085 3.523 ;
      RECT 36.981 3.32 37.02 3.533 ;
      RECT 36.895 3.32 36.981 3.54 ;
      RECT 36.875 3.325 36.89 3.546 ;
      RECT 36.865 3.365 36.875 3.548 ;
      RECT 36.835 3.375 36.865 3.55 ;
      RECT 36.83 3.38 36.835 3.552 ;
      RECT 36.805 3.385 36.83 3.554 ;
      RECT 36.79 3.39 36.805 3.556 ;
      RECT 36.775 3.392 36.79 3.558 ;
      RECT 36.77 3.397 36.775 3.56 ;
      RECT 36.72 3.405 36.77 3.563 ;
      RECT 36.695 3.414 36.72 3.568 ;
      RECT 36.685 3.421 36.695 3.573 ;
      RECT 36.68 3.424 36.685 3.577 ;
      RECT 36.66 3.427 36.68 3.586 ;
      RECT 36.63 3.435 36.66 3.606 ;
      RECT 36.601 3.448 36.63 3.628 ;
      RECT 36.515 3.482 36.601 3.672 ;
      RECT 36.51 3.508 36.515 3.71 ;
      RECT 36.505 3.512 36.51 3.719 ;
      RECT 36.47 3.525 36.505 3.752 ;
      RECT 36.46 3.539 36.47 3.79 ;
      RECT 36.455 3.543 36.46 3.803 ;
      RECT 36.45 3.547 36.455 3.808 ;
      RECT 36.44 3.555 36.45 3.82 ;
      RECT 36.435 3.562 36.44 3.835 ;
      RECT 36.41 3.575 36.435 3.86 ;
      RECT 36.37 3.604 36.41 3.915 ;
      RECT 36.355 3.629 36.37 3.97 ;
      RECT 36.345 3.64 36.355 3.993 ;
      RECT 36.34 3.647 36.345 4.005 ;
      RECT 36.335 3.651 36.34 4.013 ;
      RECT 36.28 3.679 36.335 4.055 ;
      RECT 36.26 3.715 36.28 4.055 ;
      RECT 36.245 3.73 36.26 4.055 ;
      RECT 36.19 3.762 36.245 4.055 ;
      RECT 36.18 3.792 36.19 4.055 ;
      RECT 35.79 3.407 35.975 3.645 ;
      RECT 35.775 3.409 35.985 3.64 ;
      RECT 35.66 3.355 35.92 3.615 ;
      RECT 35.655 3.392 35.92 3.569 ;
      RECT 35.65 3.402 35.92 3.566 ;
      RECT 35.645 3.442 35.985 3.56 ;
      RECT 35.64 3.475 35.985 3.55 ;
      RECT 35.65 3.417 36 3.488 ;
      RECT 35.947 4.515 35.96 5.045 ;
      RECT 35.861 4.515 35.96 5.044 ;
      RECT 35.861 4.515 35.965 5.043 ;
      RECT 35.775 4.515 35.965 5.041 ;
      RECT 35.77 4.515 35.965 5.038 ;
      RECT 35.77 4.515 35.975 5.036 ;
      RECT 35.765 4.807 35.975 5.033 ;
      RECT 35.765 4.817 35.98 5.03 ;
      RECT 35.765 4.885 35.985 5.026 ;
      RECT 35.755 4.89 35.985 5.025 ;
      RECT 35.755 4.982 35.99 5.022 ;
      RECT 35.74 4.515 36 4.775 ;
      RECT 35.67 10.05 35.96 10.28 ;
      RECT 35.73 9.31 35.9 10.28 ;
      RECT 35.645 9.34 35.985 9.685 ;
      RECT 35.67 9.31 35.96 9.685 ;
      RECT 34.97 3.505 35.015 5.04 ;
      RECT 35.17 3.505 35.2 3.72 ;
      RECT 33.545 3.245 33.665 3.455 ;
      RECT 33.205 3.195 33.465 3.455 ;
      RECT 33.205 3.24 33.5 3.445 ;
      RECT 35.21 3.521 35.215 3.575 ;
      RECT 35.205 3.514 35.21 3.708 ;
      RECT 35.2 3.508 35.205 3.715 ;
      RECT 35.155 3.505 35.17 3.728 ;
      RECT 35.15 3.505 35.155 3.75 ;
      RECT 35.145 3.505 35.15 3.798 ;
      RECT 35.14 3.505 35.145 3.818 ;
      RECT 35.13 3.505 35.14 3.925 ;
      RECT 35.125 3.505 35.13 3.988 ;
      RECT 35.12 3.505 35.125 4.045 ;
      RECT 35.115 3.505 35.12 4.053 ;
      RECT 35.1 3.505 35.115 4.16 ;
      RECT 35.09 3.505 35.1 4.295 ;
      RECT 35.08 3.505 35.09 4.405 ;
      RECT 35.07 3.505 35.08 4.462 ;
      RECT 35.065 3.505 35.07 4.502 ;
      RECT 35.06 3.505 35.065 4.538 ;
      RECT 35.05 3.505 35.06 4.578 ;
      RECT 35.045 3.505 35.05 4.62 ;
      RECT 35.025 3.505 35.045 4.685 ;
      RECT 35.03 4.83 35.035 5.01 ;
      RECT 35.025 4.812 35.03 5.018 ;
      RECT 35.02 3.505 35.025 4.748 ;
      RECT 35.02 4.792 35.025 5.025 ;
      RECT 35.015 3.505 35.02 5.035 ;
      RECT 34.96 3.505 34.97 3.805 ;
      RECT 34.965 4.052 34.97 5.04 ;
      RECT 34.96 4.117 34.965 5.04 ;
      RECT 34.955 3.506 34.96 3.795 ;
      RECT 34.95 4.182 34.96 5.04 ;
      RECT 34.945 3.507 34.955 3.785 ;
      RECT 34.935 4.295 34.95 5.04 ;
      RECT 34.94 3.508 34.945 3.775 ;
      RECT 34.92 3.509 34.94 3.753 ;
      RECT 34.925 4.392 34.935 5.04 ;
      RECT 34.92 4.467 34.925 5.04 ;
      RECT 34.91 3.508 34.92 3.73 ;
      RECT 34.915 4.51 34.92 5.04 ;
      RECT 34.91 4.537 34.915 5.04 ;
      RECT 34.9 3.506 34.91 3.718 ;
      RECT 34.905 4.58 34.91 5.04 ;
      RECT 34.9 4.607 34.905 5.04 ;
      RECT 34.89 3.505 34.9 3.705 ;
      RECT 34.895 4.622 34.9 5.04 ;
      RECT 34.855 4.68 34.895 5.04 ;
      RECT 34.885 3.504 34.89 3.69 ;
      RECT 34.88 3.502 34.885 3.683 ;
      RECT 34.87 3.499 34.88 3.673 ;
      RECT 34.865 3.496 34.87 3.658 ;
      RECT 34.85 3.492 34.865 3.651 ;
      RECT 34.845 4.735 34.855 5.04 ;
      RECT 34.845 3.489 34.85 3.646 ;
      RECT 34.83 3.485 34.845 3.64 ;
      RECT 34.84 4.752 34.845 5.04 ;
      RECT 34.83 4.815 34.84 5.04 ;
      RECT 34.75 3.47 34.83 3.62 ;
      RECT 34.825 4.822 34.83 5.035 ;
      RECT 34.82 4.83 34.825 5.025 ;
      RECT 34.74 3.456 34.75 3.604 ;
      RECT 34.725 3.452 34.74 3.602 ;
      RECT 34.715 3.447 34.725 3.598 ;
      RECT 34.69 3.44 34.715 3.59 ;
      RECT 34.685 3.435 34.69 3.585 ;
      RECT 34.675 3.435 34.685 3.583 ;
      RECT 34.665 3.433 34.675 3.581 ;
      RECT 34.635 3.425 34.665 3.575 ;
      RECT 34.62 3.417 34.635 3.568 ;
      RECT 34.6 3.412 34.62 3.561 ;
      RECT 34.595 3.408 34.6 3.556 ;
      RECT 34.565 3.401 34.595 3.55 ;
      RECT 34.54 3.392 34.565 3.54 ;
      RECT 34.51 3.385 34.54 3.532 ;
      RECT 34.485 3.375 34.51 3.523 ;
      RECT 34.47 3.367 34.485 3.517 ;
      RECT 34.445 3.362 34.47 3.512 ;
      RECT 34.435 3.358 34.445 3.507 ;
      RECT 34.415 3.353 34.435 3.502 ;
      RECT 34.38 3.348 34.415 3.495 ;
      RECT 34.32 3.343 34.38 3.488 ;
      RECT 34.307 3.339 34.32 3.486 ;
      RECT 34.221 3.334 34.307 3.483 ;
      RECT 34.135 3.324 34.221 3.479 ;
      RECT 34.094 3.317 34.135 3.476 ;
      RECT 34.008 3.31 34.094 3.473 ;
      RECT 33.922 3.3 34.008 3.469 ;
      RECT 33.836 3.29 33.922 3.464 ;
      RECT 33.75 3.28 33.836 3.46 ;
      RECT 33.74 3.265 33.75 3.458 ;
      RECT 33.73 3.25 33.74 3.458 ;
      RECT 33.665 3.245 33.73 3.457 ;
      RECT 33.5 3.242 33.545 3.45 ;
      RECT 34.745 4.147 34.75 4.338 ;
      RECT 34.74 4.142 34.745 4.345 ;
      RECT 34.726 4.14 34.74 4.351 ;
      RECT 34.64 4.14 34.726 4.353 ;
      RECT 34.636 4.14 34.64 4.356 ;
      RECT 34.55 4.14 34.636 4.374 ;
      RECT 34.54 4.145 34.55 4.393 ;
      RECT 34.53 4.2 34.54 4.397 ;
      RECT 34.505 4.215 34.53 4.404 ;
      RECT 34.465 4.235 34.505 4.417 ;
      RECT 34.46 4.247 34.465 4.427 ;
      RECT 34.445 4.253 34.46 4.432 ;
      RECT 34.44 4.258 34.445 4.436 ;
      RECT 34.42 4.265 34.44 4.441 ;
      RECT 34.35 4.29 34.42 4.458 ;
      RECT 34.31 4.318 34.35 4.478 ;
      RECT 34.305 4.328 34.31 4.486 ;
      RECT 34.285 4.335 34.305 4.488 ;
      RECT 34.28 4.342 34.285 4.491 ;
      RECT 34.25 4.35 34.28 4.494 ;
      RECT 34.245 4.355 34.25 4.498 ;
      RECT 34.171 4.359 34.245 4.506 ;
      RECT 34.085 4.368 34.171 4.522 ;
      RECT 34.081 4.373 34.085 4.531 ;
      RECT 33.995 4.378 34.081 4.541 ;
      RECT 33.955 4.386 33.995 4.553 ;
      RECT 33.905 4.392 33.955 4.56 ;
      RECT 33.82 4.401 33.905 4.575 ;
      RECT 33.745 4.412 33.82 4.593 ;
      RECT 33.71 4.419 33.745 4.603 ;
      RECT 33.635 4.427 33.71 4.608 ;
      RECT 33.58 4.436 33.635 4.608 ;
      RECT 33.555 4.441 33.58 4.606 ;
      RECT 33.545 4.444 33.555 4.604 ;
      RECT 33.51 4.446 33.545 4.602 ;
      RECT 33.48 4.448 33.51 4.598 ;
      RECT 33.435 4.447 33.48 4.594 ;
      RECT 33.415 4.442 33.435 4.591 ;
      RECT 33.365 4.427 33.415 4.588 ;
      RECT 33.355 4.412 33.365 4.583 ;
      RECT 33.305 4.397 33.355 4.573 ;
      RECT 33.255 4.372 33.305 4.553 ;
      RECT 33.245 4.357 33.255 4.535 ;
      RECT 33.24 4.355 33.245 4.529 ;
      RECT 33.22 4.35 33.24 4.524 ;
      RECT 33.215 4.342 33.22 4.518 ;
      RECT 33.2 4.336 33.215 4.511 ;
      RECT 33.195 4.331 33.2 4.503 ;
      RECT 33.175 4.326 33.195 4.495 ;
      RECT 33.16 4.319 33.175 4.488 ;
      RECT 33.145 4.313 33.16 4.479 ;
      RECT 33.14 4.307 33.145 4.472 ;
      RECT 33.095 4.282 33.14 4.458 ;
      RECT 33.08 4.252 33.095 4.44 ;
      RECT 33.065 4.235 33.08 4.431 ;
      RECT 33.04 4.215 33.065 4.419 ;
      RECT 33 4.185 33.04 4.399 ;
      RECT 32.99 4.155 33 4.384 ;
      RECT 32.975 4.145 32.99 4.377 ;
      RECT 32.92 4.11 32.975 4.356 ;
      RECT 32.905 4.073 32.92 4.335 ;
      RECT 32.895 4.06 32.905 4.327 ;
      RECT 32.845 4.03 32.895 4.309 ;
      RECT 32.83 3.96 32.845 4.29 ;
      RECT 32.785 3.96 32.83 4.273 ;
      RECT 32.76 3.96 32.785 4.255 ;
      RECT 32.75 3.96 32.76 4.248 ;
      RECT 32.671 3.96 32.75 4.241 ;
      RECT 32.585 3.96 32.671 4.233 ;
      RECT 32.57 3.992 32.585 4.228 ;
      RECT 32.495 4.002 32.57 4.224 ;
      RECT 32.475 4.012 32.495 4.219 ;
      RECT 32.45 4.012 32.475 4.216 ;
      RECT 32.44 4.002 32.45 4.215 ;
      RECT 32.43 3.975 32.44 4.214 ;
      RECT 32.39 3.97 32.43 4.212 ;
      RECT 32.345 3.97 32.39 4.208 ;
      RECT 32.32 3.97 32.345 4.203 ;
      RECT 32.27 3.97 32.32 4.19 ;
      RECT 32.23 3.975 32.24 4.175 ;
      RECT 32.24 3.97 32.27 4.18 ;
      RECT 34.225 3.75 34.485 4.01 ;
      RECT 34.22 3.772 34.485 3.968 ;
      RECT 33.46 3.6 33.68 3.965 ;
      RECT 33.442 3.687 33.68 3.964 ;
      RECT 33.425 3.692 33.68 3.961 ;
      RECT 33.425 3.692 33.7 3.96 ;
      RECT 33.395 3.702 33.7 3.958 ;
      RECT 33.39 3.717 33.7 3.954 ;
      RECT 33.39 3.717 33.705 3.953 ;
      RECT 33.385 3.775 33.705 3.951 ;
      RECT 33.385 3.775 33.715 3.948 ;
      RECT 33.38 3.84 33.715 3.943 ;
      RECT 33.46 3.6 33.72 3.86 ;
      RECT 32.205 3.43 32.465 3.69 ;
      RECT 32.205 3.473 32.551 3.664 ;
      RECT 32.205 3.473 32.595 3.663 ;
      RECT 32.205 3.473 32.615 3.661 ;
      RECT 32.205 3.473 32.715 3.66 ;
      RECT 32.205 3.473 32.735 3.658 ;
      RECT 32.205 3.473 32.745 3.653 ;
      RECT 32.615 3.44 32.805 3.65 ;
      RECT 32.615 3.442 32.81 3.648 ;
      RECT 32.605 3.447 32.815 3.64 ;
      RECT 32.551 3.471 32.815 3.64 ;
      RECT 32.595 3.465 32.605 3.662 ;
      RECT 32.605 3.445 32.81 3.648 ;
      RECT 31.56 4.505 31.765 4.735 ;
      RECT 31.5 4.455 31.555 4.715 ;
      RECT 31.56 4.455 31.76 4.735 ;
      RECT 32.53 4.77 32.535 4.797 ;
      RECT 32.52 4.68 32.53 4.802 ;
      RECT 32.515 4.602 32.52 4.808 ;
      RECT 32.505 4.592 32.515 4.815 ;
      RECT 32.5 4.582 32.505 4.821 ;
      RECT 32.49 4.577 32.5 4.823 ;
      RECT 32.475 4.569 32.49 4.831 ;
      RECT 32.46 4.56 32.475 4.843 ;
      RECT 32.45 4.552 32.46 4.853 ;
      RECT 32.415 4.47 32.45 4.871 ;
      RECT 32.38 4.47 32.415 4.89 ;
      RECT 32.365 4.47 32.38 4.898 ;
      RECT 32.31 4.47 32.365 4.898 ;
      RECT 32.276 4.47 32.31 4.889 ;
      RECT 32.19 4.47 32.276 4.865 ;
      RECT 32.18 4.53 32.19 4.847 ;
      RECT 32.14 4.532 32.18 4.838 ;
      RECT 32.135 4.534 32.14 4.828 ;
      RECT 32.115 4.536 32.135 4.823 ;
      RECT 32.105 4.539 32.115 4.818 ;
      RECT 32.095 4.54 32.105 4.813 ;
      RECT 32.071 4.541 32.095 4.805 ;
      RECT 31.985 4.546 32.071 4.783 ;
      RECT 31.93 4.545 31.985 4.756 ;
      RECT 31.915 4.538 31.93 4.743 ;
      RECT 31.88 4.533 31.915 4.739 ;
      RECT 31.825 4.525 31.88 4.738 ;
      RECT 31.765 4.512 31.825 4.736 ;
      RECT 31.555 4.455 31.56 4.723 ;
      RECT 31.63 3.825 31.815 4.035 ;
      RECT 31.62 3.83 31.83 4.028 ;
      RECT 31.66 3.735 31.92 3.995 ;
      RECT 31.615 3.892 31.92 3.918 ;
      RECT 30.96 3.685 30.965 4.485 ;
      RECT 30.905 3.735 30.935 4.485 ;
      RECT 30.895 3.735 30.9 4.045 ;
      RECT 30.88 3.735 30.885 4.04 ;
      RECT 30.425 3.78 30.44 3.995 ;
      RECT 30.355 3.78 30.44 3.99 ;
      RECT 31.62 3.36 31.69 3.57 ;
      RECT 31.69 3.367 31.7 3.565 ;
      RECT 31.586 3.36 31.62 3.577 ;
      RECT 31.5 3.36 31.586 3.601 ;
      RECT 31.49 3.365 31.5 3.62 ;
      RECT 31.485 3.377 31.49 3.623 ;
      RECT 31.47 3.392 31.485 3.627 ;
      RECT 31.465 3.41 31.47 3.631 ;
      RECT 31.425 3.42 31.465 3.64 ;
      RECT 31.41 3.427 31.425 3.652 ;
      RECT 31.395 3.432 31.41 3.657 ;
      RECT 31.38 3.435 31.395 3.662 ;
      RECT 31.37 3.437 31.38 3.666 ;
      RECT 31.335 3.444 31.37 3.674 ;
      RECT 31.3 3.452 31.335 3.688 ;
      RECT 31.29 3.458 31.3 3.697 ;
      RECT 31.285 3.46 31.29 3.699 ;
      RECT 31.265 3.463 31.285 3.705 ;
      RECT 31.235 3.47 31.265 3.716 ;
      RECT 31.225 3.476 31.235 3.723 ;
      RECT 31.2 3.479 31.225 3.73 ;
      RECT 31.19 3.483 31.2 3.738 ;
      RECT 31.185 3.484 31.19 3.76 ;
      RECT 31.18 3.485 31.185 3.775 ;
      RECT 31.175 3.486 31.18 3.79 ;
      RECT 31.17 3.487 31.175 3.805 ;
      RECT 31.165 3.488 31.17 3.835 ;
      RECT 31.155 3.49 31.165 3.868 ;
      RECT 31.14 3.494 31.155 3.915 ;
      RECT 31.13 3.497 31.14 3.96 ;
      RECT 31.125 3.5 31.13 3.988 ;
      RECT 31.115 3.502 31.125 4.015 ;
      RECT 31.11 3.505 31.115 4.05 ;
      RECT 31.08 3.51 31.11 4.108 ;
      RECT 31.075 3.515 31.08 4.193 ;
      RECT 31.07 3.517 31.075 4.228 ;
      RECT 31.065 3.519 31.07 4.31 ;
      RECT 31.06 3.521 31.065 4.398 ;
      RECT 31.05 3.523 31.06 4.48 ;
      RECT 31.035 3.537 31.05 4.485 ;
      RECT 31 3.582 31.035 4.485 ;
      RECT 30.99 3.622 31 4.485 ;
      RECT 30.975 3.65 30.99 4.485 ;
      RECT 30.97 3.667 30.975 4.485 ;
      RECT 30.965 3.675 30.97 4.485 ;
      RECT 30.955 3.69 30.96 4.485 ;
      RECT 30.95 3.697 30.955 4.485 ;
      RECT 30.94 3.717 30.95 4.485 ;
      RECT 30.935 3.73 30.94 4.485 ;
      RECT 30.9 3.735 30.905 4.07 ;
      RECT 30.885 4.125 30.905 4.485 ;
      RECT 30.885 3.735 30.895 4.043 ;
      RECT 30.88 4.165 30.885 4.485 ;
      RECT 30.83 3.735 30.88 4.038 ;
      RECT 30.875 4.202 30.88 4.485 ;
      RECT 30.865 4.225 30.875 4.485 ;
      RECT 30.86 4.27 30.865 4.485 ;
      RECT 30.85 4.28 30.86 4.478 ;
      RECT 30.776 3.735 30.83 4.032 ;
      RECT 30.69 3.735 30.776 4.025 ;
      RECT 30.641 3.782 30.69 4.018 ;
      RECT 30.555 3.79 30.641 4.011 ;
      RECT 30.54 3.787 30.555 4.006 ;
      RECT 30.526 3.78 30.54 4.005 ;
      RECT 30.44 3.78 30.526 4 ;
      RECT 30.345 3.785 30.355 3.985 ;
      RECT 29.935 3.215 29.95 3.615 ;
      RECT 30.13 3.215 30.135 3.475 ;
      RECT 29.875 3.215 29.92 3.475 ;
      RECT 30.33 4.52 30.335 4.725 ;
      RECT 30.325 4.51 30.33 4.73 ;
      RECT 30.32 4.497 30.325 4.735 ;
      RECT 30.315 4.477 30.32 4.735 ;
      RECT 30.29 4.43 30.315 4.735 ;
      RECT 30.255 4.345 30.29 4.735 ;
      RECT 30.25 4.282 30.255 4.735 ;
      RECT 30.245 4.267 30.25 4.735 ;
      RECT 30.23 4.227 30.245 4.735 ;
      RECT 30.225 4.202 30.23 4.735 ;
      RECT 30.215 4.185 30.225 4.735 ;
      RECT 30.18 4.107 30.215 4.735 ;
      RECT 30.175 4.05 30.18 4.735 ;
      RECT 30.17 4.037 30.175 4.735 ;
      RECT 30.16 4.015 30.17 4.735 ;
      RECT 30.15 3.98 30.16 4.735 ;
      RECT 30.14 3.95 30.15 4.735 ;
      RECT 30.13 3.865 30.14 4.378 ;
      RECT 30.137 4.51 30.14 4.735 ;
      RECT 30.135 4.52 30.137 4.735 ;
      RECT 30.125 4.53 30.135 4.73 ;
      RECT 30.12 3.215 30.13 3.61 ;
      RECT 30.125 3.742 30.13 4.353 ;
      RECT 30.12 3.64 30.125 4.336 ;
      RECT 30.11 3.215 30.12 4.312 ;
      RECT 30.105 3.215 30.11 4.283 ;
      RECT 30.1 3.215 30.105 4.273 ;
      RECT 30.08 3.215 30.1 4.235 ;
      RECT 30.075 3.215 30.08 4.193 ;
      RECT 30.07 3.215 30.075 4.173 ;
      RECT 30.04 3.215 30.07 4.123 ;
      RECT 30.03 3.215 30.04 4.07 ;
      RECT 30.025 3.215 30.03 4.043 ;
      RECT 30.02 3.215 30.025 4.028 ;
      RECT 30.01 3.215 30.02 4.005 ;
      RECT 30 3.215 30.01 3.98 ;
      RECT 29.995 3.215 30 3.92 ;
      RECT 29.985 3.215 29.995 3.858 ;
      RECT 29.98 3.215 29.985 3.778 ;
      RECT 29.975 3.215 29.98 3.743 ;
      RECT 29.97 3.215 29.975 3.718 ;
      RECT 29.965 3.215 29.97 3.703 ;
      RECT 29.96 3.215 29.965 3.673 ;
      RECT 29.955 3.215 29.96 3.65 ;
      RECT 29.95 3.215 29.955 3.623 ;
      RECT 29.92 3.215 29.935 3.61 ;
      RECT 29.075 4.75 29.26 4.96 ;
      RECT 29.065 4.755 29.275 4.953 ;
      RECT 29.065 4.755 29.295 4.925 ;
      RECT 29.065 4.755 29.31 4.904 ;
      RECT 29.065 4.755 29.325 4.902 ;
      RECT 29.065 4.755 29.335 4.901 ;
      RECT 29.065 4.755 29.365 4.898 ;
      RECT 29.715 4.6 29.975 4.86 ;
      RECT 29.675 4.647 29.975 4.843 ;
      RECT 29.666 4.655 29.675 4.846 ;
      RECT 29.26 4.748 29.975 4.843 ;
      RECT 29.58 4.673 29.666 4.853 ;
      RECT 29.275 4.745 29.975 4.843 ;
      RECT 29.521 4.695 29.58 4.865 ;
      RECT 29.295 4.741 29.975 4.843 ;
      RECT 29.435 4.707 29.521 4.876 ;
      RECT 29.31 4.737 29.975 4.843 ;
      RECT 29.38 4.72 29.435 4.888 ;
      RECT 29.325 4.735 29.975 4.843 ;
      RECT 29.365 4.726 29.38 4.894 ;
      RECT 29.335 4.731 29.975 4.843 ;
      RECT 29.48 4.255 29.74 4.515 ;
      RECT 29.48 4.275 29.85 4.485 ;
      RECT 29.48 4.28 29.86 4.48 ;
      RECT 29.671 3.694 29.75 3.925 ;
      RECT 29.585 3.697 29.8 3.92 ;
      RECT 29.58 3.697 29.8 3.915 ;
      RECT 29.58 3.702 29.81 3.913 ;
      RECT 29.555 3.702 29.81 3.91 ;
      RECT 29.555 3.71 29.82 3.908 ;
      RECT 29.435 3.645 29.695 3.905 ;
      RECT 29.435 3.692 29.745 3.905 ;
      RECT 28.69 4.265 28.695 4.525 ;
      RECT 28.52 4.035 28.525 4.525 ;
      RECT 28.405 4.275 28.41 4.5 ;
      RECT 29.115 3.37 29.12 3.58 ;
      RECT 29.12 3.375 29.135 3.575 ;
      RECT 29.055 3.37 29.115 3.588 ;
      RECT 29.04 3.37 29.055 3.598 ;
      RECT 28.99 3.37 29.04 3.615 ;
      RECT 28.97 3.37 28.99 3.638 ;
      RECT 28.955 3.37 28.97 3.65 ;
      RECT 28.935 3.37 28.955 3.66 ;
      RECT 28.925 3.375 28.935 3.669 ;
      RECT 28.92 3.385 28.925 3.674 ;
      RECT 28.915 3.397 28.92 3.678 ;
      RECT 28.905 3.42 28.915 3.683 ;
      RECT 28.9 3.435 28.905 3.687 ;
      RECT 28.895 3.452 28.9 3.69 ;
      RECT 28.89 3.46 28.895 3.693 ;
      RECT 28.88 3.465 28.89 3.697 ;
      RECT 28.875 3.472 28.88 3.702 ;
      RECT 28.865 3.477 28.875 3.706 ;
      RECT 28.84 3.489 28.865 3.717 ;
      RECT 28.82 3.506 28.84 3.733 ;
      RECT 28.795 3.523 28.82 3.755 ;
      RECT 28.76 3.546 28.795 3.813 ;
      RECT 28.74 3.568 28.76 3.875 ;
      RECT 28.735 3.578 28.74 3.91 ;
      RECT 28.725 3.585 28.735 3.948 ;
      RECT 28.72 3.592 28.725 3.968 ;
      RECT 28.715 3.603 28.72 4.005 ;
      RECT 28.71 3.611 28.715 4.07 ;
      RECT 28.7 3.622 28.71 4.123 ;
      RECT 28.695 3.64 28.7 4.193 ;
      RECT 28.69 3.65 28.695 4.23 ;
      RECT 28.685 3.66 28.69 4.525 ;
      RECT 28.68 3.672 28.685 4.525 ;
      RECT 28.675 3.682 28.68 4.525 ;
      RECT 28.665 3.692 28.675 4.525 ;
      RECT 28.655 3.715 28.665 4.525 ;
      RECT 28.64 3.75 28.655 4.525 ;
      RECT 28.6 3.812 28.64 4.525 ;
      RECT 28.595 3.865 28.6 4.525 ;
      RECT 28.57 3.9 28.595 4.525 ;
      RECT 28.555 3.945 28.57 4.525 ;
      RECT 28.55 3.967 28.555 4.525 ;
      RECT 28.54 3.98 28.55 4.525 ;
      RECT 28.53 4.005 28.54 4.525 ;
      RECT 28.525 4.027 28.53 4.525 ;
      RECT 28.5 4.065 28.52 4.525 ;
      RECT 28.46 4.122 28.5 4.525 ;
      RECT 28.455 4.172 28.46 4.525 ;
      RECT 28.45 4.19 28.455 4.525 ;
      RECT 28.445 4.202 28.45 4.525 ;
      RECT 28.435 4.22 28.445 4.525 ;
      RECT 28.425 4.24 28.435 4.5 ;
      RECT 28.42 4.257 28.425 4.5 ;
      RECT 28.41 4.27 28.42 4.5 ;
      RECT 28.38 4.28 28.405 4.5 ;
      RECT 28.37 4.287 28.38 4.5 ;
      RECT 28.355 4.297 28.37 4.495 ;
      RECT 27.45 10.055 27.74 10.285 ;
      RECT 27.51 8.575 27.68 10.285 ;
      RECT 27.505 8.94 27.855 9.29 ;
      RECT 27.45 8.575 27.74 8.805 ;
      RECT 27.045 3.69 27.15 4.26 ;
      RECT 27.045 4.025 27.37 4.255 ;
      RECT 27.045 4.055 27.54 4.225 ;
      RECT 27.045 3.69 27.235 4.255 ;
      RECT 26.46 3.655 26.75 3.885 ;
      RECT 26.46 3.69 27.235 3.86 ;
      RECT 26.52 2.175 26.69 3.885 ;
      RECT 26.46 2.175 26.75 2.405 ;
      RECT 26.46 10.055 26.75 10.285 ;
      RECT 26.52 8.575 26.69 10.285 ;
      RECT 26.46 8.575 26.75 8.805 ;
      RECT 26.46 8.61 27.31 8.77 ;
      RECT 27.145 8.205 27.31 8.77 ;
      RECT 26.46 8.605 26.855 8.77 ;
      RECT 27.08 8.205 27.37 8.435 ;
      RECT 27.08 8.235 27.54 8.405 ;
      RECT 26.09 4.025 26.38 4.255 ;
      RECT 26.09 4.055 26.55 4.225 ;
      RECT 26.155 2.95 26.32 4.255 ;
      RECT 24.67 2.92 24.96 3.15 ;
      RECT 24.67 2.95 26.32 3.12 ;
      RECT 24.73 2.18 24.9 3.15 ;
      RECT 24.67 2.18 24.96 2.41 ;
      RECT 24.67 10.05 24.96 10.28 ;
      RECT 24.73 9.31 24.9 10.28 ;
      RECT 24.73 9.405 26.32 9.575 ;
      RECT 26.15 8.205 26.32 9.575 ;
      RECT 24.67 9.31 24.96 9.54 ;
      RECT 26.09 8.205 26.38 8.435 ;
      RECT 26.09 8.235 26.55 8.405 ;
      RECT 25.1 3.26 25.45 3.61 ;
      RECT 22.765 3.32 25.45 3.49 ;
      RECT 22.765 2.635 22.935 3.49 ;
      RECT 22.665 2.635 23.015 2.985 ;
      RECT 25.125 8.94 25.45 9.265 ;
      RECT 20.52 8.89 20.87 9.24 ;
      RECT 25.1 8.94 25.45 9.17 ;
      RECT 20.32 8.94 20.87 9.17 ;
      RECT 20.15 8.97 25.45 9.14 ;
      RECT 24.325 3.66 24.645 3.98 ;
      RECT 24.295 3.66 24.645 3.89 ;
      RECT 24.125 3.69 24.645 3.86 ;
      RECT 24.325 8.54 24.645 8.83 ;
      RECT 24.295 8.57 24.645 8.8 ;
      RECT 24.125 8.6 24.645 8.77 ;
      RECT 20.96 3.76 21.145 3.97 ;
      RECT 20.95 3.765 21.16 3.963 ;
      RECT 20.95 3.765 21.246 3.94 ;
      RECT 20.95 3.765 21.305 3.915 ;
      RECT 20.95 3.765 21.36 3.895 ;
      RECT 20.95 3.765 21.37 3.883 ;
      RECT 20.95 3.765 21.565 3.822 ;
      RECT 20.95 3.765 21.595 3.805 ;
      RECT 20.95 3.765 21.615 3.795 ;
      RECT 21.495 3.53 21.755 3.79 ;
      RECT 21.48 3.62 21.495 3.837 ;
      RECT 21.015 3.752 21.755 3.79 ;
      RECT 21.466 3.631 21.48 3.843 ;
      RECT 21.055 3.745 21.755 3.79 ;
      RECT 21.38 3.671 21.466 3.862 ;
      RECT 21.305 3.732 21.755 3.79 ;
      RECT 21.375 3.707 21.38 3.879 ;
      RECT 21.36 3.717 21.755 3.79 ;
      RECT 21.37 3.712 21.375 3.881 ;
      RECT 21.665 4.217 21.67 4.309 ;
      RECT 21.66 4.195 21.665 4.326 ;
      RECT 21.655 4.185 21.66 4.338 ;
      RECT 21.645 4.176 21.655 4.348 ;
      RECT 21.64 4.171 21.645 4.356 ;
      RECT 21.635 4.03 21.64 4.359 ;
      RECT 21.601 4.03 21.635 4.37 ;
      RECT 21.515 4.03 21.601 4.405 ;
      RECT 21.435 4.03 21.515 4.453 ;
      RECT 21.406 4.03 21.435 4.477 ;
      RECT 21.32 4.03 21.406 4.483 ;
      RECT 21.315 4.214 21.32 4.488 ;
      RECT 21.28 4.225 21.315 4.491 ;
      RECT 21.255 4.24 21.28 4.495 ;
      RECT 21.241 4.249 21.255 4.497 ;
      RECT 21.155 4.276 21.241 4.503 ;
      RECT 21.09 4.317 21.155 4.512 ;
      RECT 21.075 4.337 21.09 4.517 ;
      RECT 21.045 4.347 21.075 4.52 ;
      RECT 21.04 4.357 21.045 4.523 ;
      RECT 21.01 4.362 21.04 4.525 ;
      RECT 20.99 4.367 21.01 4.529 ;
      RECT 20.905 4.37 20.99 4.536 ;
      RECT 20.89 4.367 20.905 4.542 ;
      RECT 20.88 4.364 20.89 4.544 ;
      RECT 20.86 4.361 20.88 4.546 ;
      RECT 20.84 4.357 20.86 4.547 ;
      RECT 20.825 4.353 20.84 4.549 ;
      RECT 20.815 4.35 20.825 4.55 ;
      RECT 20.775 4.344 20.815 4.548 ;
      RECT 20.765 4.339 20.775 4.546 ;
      RECT 20.75 4.336 20.765 4.542 ;
      RECT 20.725 4.331 20.75 4.535 ;
      RECT 20.675 4.322 20.725 4.523 ;
      RECT 20.605 4.308 20.675 4.505 ;
      RECT 20.547 4.293 20.605 4.487 ;
      RECT 20.461 4.276 20.547 4.467 ;
      RECT 20.375 4.255 20.461 4.442 ;
      RECT 20.325 4.24 20.375 4.423 ;
      RECT 20.321 4.234 20.325 4.415 ;
      RECT 20.235 4.224 20.321 4.402 ;
      RECT 20.2 4.209 20.235 4.385 ;
      RECT 20.185 4.202 20.2 4.378 ;
      RECT 20.125 4.19 20.185 4.366 ;
      RECT 20.105 4.177 20.125 4.354 ;
      RECT 20.065 4.168 20.105 4.346 ;
      RECT 20.06 4.16 20.065 4.339 ;
      RECT 19.98 4.15 20.06 4.325 ;
      RECT 19.965 4.137 19.98 4.31 ;
      RECT 19.96 4.135 19.965 4.308 ;
      RECT 19.881 4.123 19.96 4.295 ;
      RECT 19.795 4.098 19.881 4.27 ;
      RECT 19.78 4.067 19.795 4.255 ;
      RECT 19.765 4.042 19.78 4.251 ;
      RECT 19.75 4.035 19.765 4.247 ;
      RECT 19.575 4.04 19.58 4.243 ;
      RECT 19.57 4.045 19.575 4.238 ;
      RECT 19.58 4.035 19.75 4.245 ;
      RECT 20.295 3.795 20.4 4.055 ;
      RECT 21.11 3.32 21.115 3.545 ;
      RECT 21.24 3.32 21.295 3.53 ;
      RECT 21.295 3.325 21.305 3.523 ;
      RECT 21.201 3.32 21.24 3.533 ;
      RECT 21.115 3.32 21.201 3.54 ;
      RECT 21.095 3.325 21.11 3.546 ;
      RECT 21.085 3.365 21.095 3.548 ;
      RECT 21.055 3.375 21.085 3.55 ;
      RECT 21.05 3.38 21.055 3.552 ;
      RECT 21.025 3.385 21.05 3.554 ;
      RECT 21.01 3.39 21.025 3.556 ;
      RECT 20.995 3.392 21.01 3.558 ;
      RECT 20.99 3.397 20.995 3.56 ;
      RECT 20.94 3.405 20.99 3.563 ;
      RECT 20.915 3.414 20.94 3.568 ;
      RECT 20.905 3.421 20.915 3.573 ;
      RECT 20.9 3.424 20.905 3.577 ;
      RECT 20.88 3.427 20.9 3.586 ;
      RECT 20.85 3.435 20.88 3.606 ;
      RECT 20.821 3.448 20.85 3.628 ;
      RECT 20.735 3.482 20.821 3.672 ;
      RECT 20.73 3.508 20.735 3.71 ;
      RECT 20.725 3.512 20.73 3.719 ;
      RECT 20.69 3.525 20.725 3.752 ;
      RECT 20.68 3.539 20.69 3.79 ;
      RECT 20.675 3.543 20.68 3.803 ;
      RECT 20.67 3.547 20.675 3.808 ;
      RECT 20.66 3.555 20.67 3.82 ;
      RECT 20.655 3.562 20.66 3.835 ;
      RECT 20.63 3.575 20.655 3.86 ;
      RECT 20.59 3.604 20.63 3.915 ;
      RECT 20.575 3.629 20.59 3.97 ;
      RECT 20.565 3.64 20.575 3.993 ;
      RECT 20.56 3.647 20.565 4.005 ;
      RECT 20.555 3.651 20.56 4.013 ;
      RECT 20.5 3.679 20.555 4.055 ;
      RECT 20.48 3.715 20.5 4.055 ;
      RECT 20.465 3.73 20.48 4.055 ;
      RECT 20.41 3.762 20.465 4.055 ;
      RECT 20.4 3.792 20.41 4.055 ;
      RECT 20.01 3.407 20.195 3.645 ;
      RECT 19.995 3.409 20.205 3.64 ;
      RECT 19.88 3.355 20.14 3.615 ;
      RECT 19.875 3.392 20.14 3.569 ;
      RECT 19.87 3.402 20.14 3.566 ;
      RECT 19.865 3.442 20.205 3.56 ;
      RECT 19.86 3.475 20.205 3.55 ;
      RECT 19.87 3.417 20.22 3.488 ;
      RECT 20.167 4.515 20.18 5.045 ;
      RECT 20.081 4.515 20.18 5.044 ;
      RECT 20.081 4.515 20.185 5.043 ;
      RECT 19.995 4.515 20.185 5.041 ;
      RECT 19.99 4.515 20.185 5.038 ;
      RECT 19.99 4.515 20.195 5.036 ;
      RECT 19.985 4.807 20.195 5.033 ;
      RECT 19.985 4.817 20.2 5.03 ;
      RECT 19.985 4.885 20.205 5.026 ;
      RECT 19.975 4.89 20.205 5.025 ;
      RECT 19.975 4.982 20.21 5.022 ;
      RECT 19.96 4.515 20.22 4.775 ;
      RECT 19.89 10.05 20.18 10.28 ;
      RECT 19.95 9.31 20.12 10.28 ;
      RECT 19.865 9.34 20.205 9.685 ;
      RECT 19.89 9.31 20.18 9.685 ;
      RECT 19.19 3.505 19.235 5.04 ;
      RECT 19.39 3.505 19.42 3.72 ;
      RECT 17.765 3.245 17.885 3.455 ;
      RECT 17.425 3.195 17.685 3.455 ;
      RECT 17.425 3.24 17.72 3.445 ;
      RECT 19.43 3.521 19.435 3.575 ;
      RECT 19.425 3.514 19.43 3.708 ;
      RECT 19.42 3.508 19.425 3.715 ;
      RECT 19.375 3.505 19.39 3.728 ;
      RECT 19.37 3.505 19.375 3.75 ;
      RECT 19.365 3.505 19.37 3.798 ;
      RECT 19.36 3.505 19.365 3.818 ;
      RECT 19.35 3.505 19.36 3.925 ;
      RECT 19.345 3.505 19.35 3.988 ;
      RECT 19.34 3.505 19.345 4.045 ;
      RECT 19.335 3.505 19.34 4.053 ;
      RECT 19.32 3.505 19.335 4.16 ;
      RECT 19.31 3.505 19.32 4.295 ;
      RECT 19.3 3.505 19.31 4.405 ;
      RECT 19.29 3.505 19.3 4.462 ;
      RECT 19.285 3.505 19.29 4.502 ;
      RECT 19.28 3.505 19.285 4.538 ;
      RECT 19.27 3.505 19.28 4.578 ;
      RECT 19.265 3.505 19.27 4.62 ;
      RECT 19.245 3.505 19.265 4.685 ;
      RECT 19.25 4.83 19.255 5.01 ;
      RECT 19.245 4.812 19.25 5.018 ;
      RECT 19.24 3.505 19.245 4.748 ;
      RECT 19.24 4.792 19.245 5.025 ;
      RECT 19.235 3.505 19.24 5.035 ;
      RECT 19.18 3.505 19.19 3.805 ;
      RECT 19.185 4.052 19.19 5.04 ;
      RECT 19.18 4.117 19.185 5.04 ;
      RECT 19.175 3.506 19.18 3.795 ;
      RECT 19.17 4.182 19.18 5.04 ;
      RECT 19.165 3.507 19.175 3.785 ;
      RECT 19.155 4.295 19.17 5.04 ;
      RECT 19.16 3.508 19.165 3.775 ;
      RECT 19.14 3.509 19.16 3.753 ;
      RECT 19.145 4.392 19.155 5.04 ;
      RECT 19.14 4.467 19.145 5.04 ;
      RECT 19.13 3.508 19.14 3.73 ;
      RECT 19.135 4.51 19.14 5.04 ;
      RECT 19.13 4.537 19.135 5.04 ;
      RECT 19.12 3.506 19.13 3.718 ;
      RECT 19.125 4.58 19.13 5.04 ;
      RECT 19.12 4.607 19.125 5.04 ;
      RECT 19.11 3.505 19.12 3.705 ;
      RECT 19.115 4.622 19.12 5.04 ;
      RECT 19.075 4.68 19.115 5.04 ;
      RECT 19.105 3.504 19.11 3.69 ;
      RECT 19.1 3.502 19.105 3.683 ;
      RECT 19.09 3.499 19.1 3.673 ;
      RECT 19.085 3.496 19.09 3.658 ;
      RECT 19.07 3.492 19.085 3.651 ;
      RECT 19.065 4.735 19.075 5.04 ;
      RECT 19.065 3.489 19.07 3.646 ;
      RECT 19.05 3.485 19.065 3.64 ;
      RECT 19.06 4.752 19.065 5.04 ;
      RECT 19.05 4.815 19.06 5.04 ;
      RECT 18.97 3.47 19.05 3.62 ;
      RECT 19.045 4.822 19.05 5.035 ;
      RECT 19.04 4.83 19.045 5.025 ;
      RECT 18.96 3.456 18.97 3.604 ;
      RECT 18.945 3.452 18.96 3.602 ;
      RECT 18.935 3.447 18.945 3.598 ;
      RECT 18.91 3.44 18.935 3.59 ;
      RECT 18.905 3.435 18.91 3.585 ;
      RECT 18.895 3.435 18.905 3.583 ;
      RECT 18.885 3.433 18.895 3.581 ;
      RECT 18.855 3.425 18.885 3.575 ;
      RECT 18.84 3.417 18.855 3.568 ;
      RECT 18.82 3.412 18.84 3.561 ;
      RECT 18.815 3.408 18.82 3.556 ;
      RECT 18.785 3.401 18.815 3.55 ;
      RECT 18.76 3.392 18.785 3.54 ;
      RECT 18.73 3.385 18.76 3.532 ;
      RECT 18.705 3.375 18.73 3.523 ;
      RECT 18.69 3.367 18.705 3.517 ;
      RECT 18.665 3.362 18.69 3.512 ;
      RECT 18.655 3.358 18.665 3.507 ;
      RECT 18.635 3.353 18.655 3.502 ;
      RECT 18.6 3.348 18.635 3.495 ;
      RECT 18.54 3.343 18.6 3.488 ;
      RECT 18.527 3.339 18.54 3.486 ;
      RECT 18.441 3.334 18.527 3.483 ;
      RECT 18.355 3.324 18.441 3.479 ;
      RECT 18.314 3.317 18.355 3.476 ;
      RECT 18.228 3.31 18.314 3.473 ;
      RECT 18.142 3.3 18.228 3.469 ;
      RECT 18.056 3.29 18.142 3.464 ;
      RECT 17.97 3.28 18.056 3.46 ;
      RECT 17.96 3.265 17.97 3.458 ;
      RECT 17.95 3.25 17.96 3.458 ;
      RECT 17.885 3.245 17.95 3.457 ;
      RECT 17.72 3.242 17.765 3.45 ;
      RECT 18.965 4.147 18.97 4.338 ;
      RECT 18.96 4.142 18.965 4.345 ;
      RECT 18.946 4.14 18.96 4.351 ;
      RECT 18.86 4.14 18.946 4.353 ;
      RECT 18.856 4.14 18.86 4.356 ;
      RECT 18.77 4.14 18.856 4.374 ;
      RECT 18.76 4.145 18.77 4.393 ;
      RECT 18.75 4.2 18.76 4.397 ;
      RECT 18.725 4.215 18.75 4.404 ;
      RECT 18.685 4.235 18.725 4.417 ;
      RECT 18.68 4.247 18.685 4.427 ;
      RECT 18.665 4.253 18.68 4.432 ;
      RECT 18.66 4.258 18.665 4.436 ;
      RECT 18.64 4.265 18.66 4.441 ;
      RECT 18.57 4.29 18.64 4.458 ;
      RECT 18.53 4.318 18.57 4.478 ;
      RECT 18.525 4.328 18.53 4.486 ;
      RECT 18.505 4.335 18.525 4.488 ;
      RECT 18.5 4.342 18.505 4.491 ;
      RECT 18.47 4.35 18.5 4.494 ;
      RECT 18.465 4.355 18.47 4.498 ;
      RECT 18.391 4.359 18.465 4.506 ;
      RECT 18.305 4.368 18.391 4.522 ;
      RECT 18.301 4.373 18.305 4.531 ;
      RECT 18.215 4.378 18.301 4.541 ;
      RECT 18.175 4.386 18.215 4.553 ;
      RECT 18.125 4.392 18.175 4.56 ;
      RECT 18.04 4.401 18.125 4.575 ;
      RECT 17.965 4.412 18.04 4.593 ;
      RECT 17.93 4.419 17.965 4.603 ;
      RECT 17.855 4.427 17.93 4.608 ;
      RECT 17.8 4.436 17.855 4.608 ;
      RECT 17.775 4.441 17.8 4.606 ;
      RECT 17.765 4.444 17.775 4.604 ;
      RECT 17.73 4.446 17.765 4.602 ;
      RECT 17.7 4.448 17.73 4.598 ;
      RECT 17.655 4.447 17.7 4.594 ;
      RECT 17.635 4.442 17.655 4.591 ;
      RECT 17.585 4.427 17.635 4.588 ;
      RECT 17.575 4.412 17.585 4.583 ;
      RECT 17.525 4.397 17.575 4.573 ;
      RECT 17.475 4.372 17.525 4.553 ;
      RECT 17.465 4.357 17.475 4.535 ;
      RECT 17.46 4.355 17.465 4.529 ;
      RECT 17.44 4.35 17.46 4.524 ;
      RECT 17.435 4.342 17.44 4.518 ;
      RECT 17.42 4.336 17.435 4.511 ;
      RECT 17.415 4.331 17.42 4.503 ;
      RECT 17.395 4.326 17.415 4.495 ;
      RECT 17.38 4.319 17.395 4.488 ;
      RECT 17.365 4.313 17.38 4.479 ;
      RECT 17.36 4.307 17.365 4.472 ;
      RECT 17.315 4.282 17.36 4.458 ;
      RECT 17.3 4.252 17.315 4.44 ;
      RECT 17.285 4.235 17.3 4.431 ;
      RECT 17.26 4.215 17.285 4.419 ;
      RECT 17.22 4.185 17.26 4.399 ;
      RECT 17.21 4.155 17.22 4.384 ;
      RECT 17.195 4.145 17.21 4.377 ;
      RECT 17.14 4.11 17.195 4.356 ;
      RECT 17.125 4.073 17.14 4.335 ;
      RECT 17.115 4.06 17.125 4.327 ;
      RECT 17.065 4.03 17.115 4.309 ;
      RECT 17.05 3.96 17.065 4.29 ;
      RECT 17.005 3.96 17.05 4.273 ;
      RECT 16.98 3.96 17.005 4.255 ;
      RECT 16.97 3.96 16.98 4.248 ;
      RECT 16.891 3.96 16.97 4.241 ;
      RECT 16.805 3.96 16.891 4.233 ;
      RECT 16.79 3.992 16.805 4.228 ;
      RECT 16.715 4.002 16.79 4.224 ;
      RECT 16.695 4.012 16.715 4.219 ;
      RECT 16.67 4.012 16.695 4.216 ;
      RECT 16.66 4.002 16.67 4.215 ;
      RECT 16.65 3.975 16.66 4.214 ;
      RECT 16.61 3.97 16.65 4.212 ;
      RECT 16.565 3.97 16.61 4.208 ;
      RECT 16.54 3.97 16.565 4.203 ;
      RECT 16.49 3.97 16.54 4.19 ;
      RECT 16.45 3.975 16.46 4.175 ;
      RECT 16.46 3.97 16.49 4.18 ;
      RECT 18.445 3.75 18.705 4.01 ;
      RECT 18.44 3.772 18.705 3.968 ;
      RECT 17.68 3.6 17.9 3.965 ;
      RECT 17.662 3.687 17.9 3.964 ;
      RECT 17.645 3.692 17.9 3.961 ;
      RECT 17.645 3.692 17.92 3.96 ;
      RECT 17.615 3.702 17.92 3.958 ;
      RECT 17.61 3.717 17.92 3.954 ;
      RECT 17.61 3.717 17.925 3.953 ;
      RECT 17.605 3.775 17.925 3.951 ;
      RECT 17.605 3.775 17.935 3.948 ;
      RECT 17.6 3.84 17.935 3.943 ;
      RECT 17.68 3.6 17.94 3.86 ;
      RECT 16.425 3.43 16.685 3.69 ;
      RECT 16.425 3.473 16.771 3.664 ;
      RECT 16.425 3.473 16.815 3.663 ;
      RECT 16.425 3.473 16.835 3.661 ;
      RECT 16.425 3.473 16.935 3.66 ;
      RECT 16.425 3.473 16.955 3.658 ;
      RECT 16.425 3.473 16.965 3.653 ;
      RECT 16.835 3.44 17.025 3.65 ;
      RECT 16.835 3.442 17.03 3.648 ;
      RECT 16.825 3.447 17.035 3.64 ;
      RECT 16.771 3.471 17.035 3.64 ;
      RECT 16.815 3.465 16.825 3.662 ;
      RECT 16.825 3.445 17.03 3.648 ;
      RECT 15.78 4.505 15.985 4.735 ;
      RECT 15.72 4.455 15.775 4.715 ;
      RECT 15.78 4.455 15.98 4.735 ;
      RECT 16.75 4.77 16.755 4.797 ;
      RECT 16.74 4.68 16.75 4.802 ;
      RECT 16.735 4.602 16.74 4.808 ;
      RECT 16.725 4.592 16.735 4.815 ;
      RECT 16.72 4.582 16.725 4.821 ;
      RECT 16.71 4.577 16.72 4.823 ;
      RECT 16.695 4.569 16.71 4.831 ;
      RECT 16.68 4.56 16.695 4.843 ;
      RECT 16.67 4.552 16.68 4.853 ;
      RECT 16.635 4.47 16.67 4.871 ;
      RECT 16.6 4.47 16.635 4.89 ;
      RECT 16.585 4.47 16.6 4.898 ;
      RECT 16.53 4.47 16.585 4.898 ;
      RECT 16.496 4.47 16.53 4.889 ;
      RECT 16.41 4.47 16.496 4.865 ;
      RECT 16.4 4.53 16.41 4.847 ;
      RECT 16.36 4.532 16.4 4.838 ;
      RECT 16.355 4.534 16.36 4.828 ;
      RECT 16.335 4.536 16.355 4.823 ;
      RECT 16.325 4.539 16.335 4.818 ;
      RECT 16.315 4.54 16.325 4.813 ;
      RECT 16.291 4.541 16.315 4.805 ;
      RECT 16.205 4.546 16.291 4.783 ;
      RECT 16.15 4.545 16.205 4.756 ;
      RECT 16.135 4.538 16.15 4.743 ;
      RECT 16.1 4.533 16.135 4.739 ;
      RECT 16.045 4.525 16.1 4.738 ;
      RECT 15.985 4.512 16.045 4.736 ;
      RECT 15.775 4.455 15.78 4.723 ;
      RECT 15.85 3.825 16.035 4.035 ;
      RECT 15.84 3.83 16.05 4.028 ;
      RECT 15.88 3.735 16.14 3.995 ;
      RECT 15.835 3.892 16.14 3.918 ;
      RECT 15.18 3.685 15.185 4.485 ;
      RECT 15.125 3.735 15.155 4.485 ;
      RECT 15.115 3.735 15.12 4.045 ;
      RECT 15.1 3.735 15.105 4.04 ;
      RECT 14.645 3.78 14.66 3.995 ;
      RECT 14.575 3.78 14.66 3.99 ;
      RECT 15.84 3.36 15.91 3.57 ;
      RECT 15.91 3.367 15.92 3.565 ;
      RECT 15.806 3.36 15.84 3.577 ;
      RECT 15.72 3.36 15.806 3.601 ;
      RECT 15.71 3.365 15.72 3.62 ;
      RECT 15.705 3.377 15.71 3.623 ;
      RECT 15.69 3.392 15.705 3.627 ;
      RECT 15.685 3.41 15.69 3.631 ;
      RECT 15.645 3.42 15.685 3.64 ;
      RECT 15.63 3.427 15.645 3.652 ;
      RECT 15.615 3.432 15.63 3.657 ;
      RECT 15.6 3.435 15.615 3.662 ;
      RECT 15.59 3.437 15.6 3.666 ;
      RECT 15.555 3.444 15.59 3.674 ;
      RECT 15.52 3.452 15.555 3.688 ;
      RECT 15.51 3.458 15.52 3.697 ;
      RECT 15.505 3.46 15.51 3.699 ;
      RECT 15.485 3.463 15.505 3.705 ;
      RECT 15.455 3.47 15.485 3.716 ;
      RECT 15.445 3.476 15.455 3.723 ;
      RECT 15.42 3.479 15.445 3.73 ;
      RECT 15.41 3.483 15.42 3.738 ;
      RECT 15.405 3.484 15.41 3.76 ;
      RECT 15.4 3.485 15.405 3.775 ;
      RECT 15.395 3.486 15.4 3.79 ;
      RECT 15.39 3.487 15.395 3.805 ;
      RECT 15.385 3.488 15.39 3.835 ;
      RECT 15.375 3.49 15.385 3.868 ;
      RECT 15.36 3.494 15.375 3.915 ;
      RECT 15.35 3.497 15.36 3.96 ;
      RECT 15.345 3.5 15.35 3.988 ;
      RECT 15.335 3.502 15.345 4.015 ;
      RECT 15.33 3.505 15.335 4.05 ;
      RECT 15.3 3.51 15.33 4.108 ;
      RECT 15.295 3.515 15.3 4.193 ;
      RECT 15.29 3.517 15.295 4.228 ;
      RECT 15.285 3.519 15.29 4.31 ;
      RECT 15.28 3.521 15.285 4.398 ;
      RECT 15.27 3.523 15.28 4.48 ;
      RECT 15.255 3.537 15.27 4.485 ;
      RECT 15.22 3.582 15.255 4.485 ;
      RECT 15.21 3.622 15.22 4.485 ;
      RECT 15.195 3.65 15.21 4.485 ;
      RECT 15.19 3.667 15.195 4.485 ;
      RECT 15.185 3.675 15.19 4.485 ;
      RECT 15.175 3.69 15.18 4.485 ;
      RECT 15.17 3.697 15.175 4.485 ;
      RECT 15.16 3.717 15.17 4.485 ;
      RECT 15.155 3.73 15.16 4.485 ;
      RECT 15.12 3.735 15.125 4.07 ;
      RECT 15.105 4.125 15.125 4.485 ;
      RECT 15.105 3.735 15.115 4.043 ;
      RECT 15.1 4.165 15.105 4.485 ;
      RECT 15.05 3.735 15.1 4.038 ;
      RECT 15.095 4.202 15.1 4.485 ;
      RECT 15.085 4.225 15.095 4.485 ;
      RECT 15.08 4.27 15.085 4.485 ;
      RECT 15.07 4.28 15.08 4.478 ;
      RECT 14.996 3.735 15.05 4.032 ;
      RECT 14.91 3.735 14.996 4.025 ;
      RECT 14.861 3.782 14.91 4.018 ;
      RECT 14.775 3.79 14.861 4.011 ;
      RECT 14.76 3.787 14.775 4.006 ;
      RECT 14.746 3.78 14.76 4.005 ;
      RECT 14.66 3.78 14.746 4 ;
      RECT 14.565 3.785 14.575 3.985 ;
      RECT 14.155 3.215 14.17 3.615 ;
      RECT 14.35 3.215 14.355 3.475 ;
      RECT 14.095 3.215 14.14 3.475 ;
      RECT 14.55 4.52 14.555 4.725 ;
      RECT 14.545 4.51 14.55 4.73 ;
      RECT 14.54 4.497 14.545 4.735 ;
      RECT 14.535 4.477 14.54 4.735 ;
      RECT 14.51 4.43 14.535 4.735 ;
      RECT 14.475 4.345 14.51 4.735 ;
      RECT 14.47 4.282 14.475 4.735 ;
      RECT 14.465 4.267 14.47 4.735 ;
      RECT 14.45 4.227 14.465 4.735 ;
      RECT 14.445 4.202 14.45 4.735 ;
      RECT 14.435 4.185 14.445 4.735 ;
      RECT 14.4 4.107 14.435 4.735 ;
      RECT 14.395 4.05 14.4 4.735 ;
      RECT 14.39 4.037 14.395 4.735 ;
      RECT 14.38 4.015 14.39 4.735 ;
      RECT 14.37 3.98 14.38 4.735 ;
      RECT 14.36 3.95 14.37 4.735 ;
      RECT 14.35 3.865 14.36 4.378 ;
      RECT 14.357 4.51 14.36 4.735 ;
      RECT 14.355 4.52 14.357 4.735 ;
      RECT 14.345 4.53 14.355 4.73 ;
      RECT 14.34 3.215 14.35 3.61 ;
      RECT 14.345 3.742 14.35 4.353 ;
      RECT 14.34 3.64 14.345 4.336 ;
      RECT 14.33 3.215 14.34 4.312 ;
      RECT 14.325 3.215 14.33 4.283 ;
      RECT 14.32 3.215 14.325 4.273 ;
      RECT 14.3 3.215 14.32 4.235 ;
      RECT 14.295 3.215 14.3 4.193 ;
      RECT 14.29 3.215 14.295 4.173 ;
      RECT 14.26 3.215 14.29 4.123 ;
      RECT 14.25 3.215 14.26 4.07 ;
      RECT 14.245 3.215 14.25 4.043 ;
      RECT 14.24 3.215 14.245 4.028 ;
      RECT 14.23 3.215 14.24 4.005 ;
      RECT 14.22 3.215 14.23 3.98 ;
      RECT 14.215 3.215 14.22 3.92 ;
      RECT 14.205 3.215 14.215 3.858 ;
      RECT 14.2 3.215 14.205 3.778 ;
      RECT 14.195 3.215 14.2 3.743 ;
      RECT 14.19 3.215 14.195 3.718 ;
      RECT 14.185 3.215 14.19 3.703 ;
      RECT 14.18 3.215 14.185 3.673 ;
      RECT 14.175 3.215 14.18 3.65 ;
      RECT 14.17 3.215 14.175 3.623 ;
      RECT 14.14 3.215 14.155 3.61 ;
      RECT 13.295 4.75 13.48 4.96 ;
      RECT 13.285 4.755 13.495 4.953 ;
      RECT 13.285 4.755 13.515 4.925 ;
      RECT 13.285 4.755 13.53 4.904 ;
      RECT 13.285 4.755 13.545 4.902 ;
      RECT 13.285 4.755 13.555 4.901 ;
      RECT 13.285 4.755 13.585 4.898 ;
      RECT 13.935 4.6 14.195 4.86 ;
      RECT 13.895 4.647 14.195 4.843 ;
      RECT 13.886 4.655 13.895 4.846 ;
      RECT 13.48 4.748 14.195 4.843 ;
      RECT 13.8 4.673 13.886 4.853 ;
      RECT 13.495 4.745 14.195 4.843 ;
      RECT 13.741 4.695 13.8 4.865 ;
      RECT 13.515 4.741 14.195 4.843 ;
      RECT 13.655 4.707 13.741 4.876 ;
      RECT 13.53 4.737 14.195 4.843 ;
      RECT 13.6 4.72 13.655 4.888 ;
      RECT 13.545 4.735 14.195 4.843 ;
      RECT 13.585 4.726 13.6 4.894 ;
      RECT 13.555 4.731 14.195 4.843 ;
      RECT 13.7 4.255 13.96 4.515 ;
      RECT 13.7 4.275 14.07 4.485 ;
      RECT 13.7 4.28 14.08 4.48 ;
      RECT 13.891 3.694 13.97 3.925 ;
      RECT 13.805 3.697 14.02 3.92 ;
      RECT 13.8 3.697 14.02 3.915 ;
      RECT 13.8 3.702 14.03 3.913 ;
      RECT 13.775 3.702 14.03 3.91 ;
      RECT 13.775 3.71 14.04 3.908 ;
      RECT 13.655 3.645 13.915 3.905 ;
      RECT 13.655 3.692 13.965 3.905 ;
      RECT 12.91 4.265 12.915 4.525 ;
      RECT 12.74 4.035 12.745 4.525 ;
      RECT 12.625 4.275 12.63 4.5 ;
      RECT 13.335 3.37 13.34 3.58 ;
      RECT 13.34 3.375 13.355 3.575 ;
      RECT 13.275 3.37 13.335 3.588 ;
      RECT 13.26 3.37 13.275 3.598 ;
      RECT 13.21 3.37 13.26 3.615 ;
      RECT 13.19 3.37 13.21 3.638 ;
      RECT 13.175 3.37 13.19 3.65 ;
      RECT 13.155 3.37 13.175 3.66 ;
      RECT 13.145 3.375 13.155 3.669 ;
      RECT 13.14 3.385 13.145 3.674 ;
      RECT 13.135 3.397 13.14 3.678 ;
      RECT 13.125 3.42 13.135 3.683 ;
      RECT 13.12 3.435 13.125 3.687 ;
      RECT 13.115 3.452 13.12 3.69 ;
      RECT 13.11 3.46 13.115 3.693 ;
      RECT 13.1 3.465 13.11 3.697 ;
      RECT 13.095 3.472 13.1 3.702 ;
      RECT 13.085 3.477 13.095 3.706 ;
      RECT 13.06 3.489 13.085 3.717 ;
      RECT 13.04 3.506 13.06 3.733 ;
      RECT 13.015 3.523 13.04 3.755 ;
      RECT 12.98 3.546 13.015 3.813 ;
      RECT 12.96 3.568 12.98 3.875 ;
      RECT 12.955 3.578 12.96 3.91 ;
      RECT 12.945 3.585 12.955 3.948 ;
      RECT 12.94 3.592 12.945 3.968 ;
      RECT 12.935 3.603 12.94 4.005 ;
      RECT 12.93 3.611 12.935 4.07 ;
      RECT 12.92 3.622 12.93 4.123 ;
      RECT 12.915 3.64 12.92 4.193 ;
      RECT 12.91 3.65 12.915 4.23 ;
      RECT 12.905 3.66 12.91 4.525 ;
      RECT 12.9 3.672 12.905 4.525 ;
      RECT 12.895 3.682 12.9 4.525 ;
      RECT 12.885 3.692 12.895 4.525 ;
      RECT 12.875 3.715 12.885 4.525 ;
      RECT 12.86 3.75 12.875 4.525 ;
      RECT 12.82 3.812 12.86 4.525 ;
      RECT 12.815 3.865 12.82 4.525 ;
      RECT 12.79 3.9 12.815 4.525 ;
      RECT 12.775 3.945 12.79 4.525 ;
      RECT 12.77 3.967 12.775 4.525 ;
      RECT 12.76 3.98 12.77 4.525 ;
      RECT 12.75 4.005 12.76 4.525 ;
      RECT 12.745 4.027 12.75 4.525 ;
      RECT 12.72 4.065 12.74 4.525 ;
      RECT 12.68 4.122 12.72 4.525 ;
      RECT 12.675 4.172 12.68 4.525 ;
      RECT 12.67 4.19 12.675 4.525 ;
      RECT 12.665 4.202 12.67 4.525 ;
      RECT 12.655 4.22 12.665 4.525 ;
      RECT 12.645 4.24 12.655 4.5 ;
      RECT 12.64 4.257 12.645 4.5 ;
      RECT 12.63 4.27 12.64 4.5 ;
      RECT 12.6 4.28 12.625 4.5 ;
      RECT 12.59 4.287 12.6 4.5 ;
      RECT 12.575 4.297 12.59 4.495 ;
      RECT 11.445 8.94 11.735 9.17 ;
      RECT 11.275 8.97 11.735 9.14 ;
      RECT 11.015 10.05 11.305 10.28 ;
      RECT 11.075 9.31 11.245 10.28 ;
      RECT 10.925 9.31 11.275 9.6 ;
      RECT 10.925 9.31 11.305 9.54 ;
      RECT 10.55 8.57 10.9 8.86 ;
      RECT 10.55 8.57 10.93 8.8 ;
      RECT 10.47 8.6 10.93 8.77 ;
      RECT 85.465 4.145 85.835 4.515 ;
      RECT 69.68 4.145 70.05 4.515 ;
      RECT 53.895 4.145 54.265 4.515 ;
      RECT 38.12 4.145 38.49 4.515 ;
      RECT 22.34 4.145 22.71 4.515 ;
    LAYER mcon ;
      RECT 90.635 8.605 90.805 8.775 ;
      RECT 90.635 10.085 90.805 10.255 ;
      RECT 90.285 1.395 90.455 1.565 ;
      RECT 90.285 5.455 90.455 5.625 ;
      RECT 90.285 6.835 90.455 7.005 ;
      RECT 90.285 10.895 90.455 11.065 ;
      RECT 90.265 4.055 90.435 4.225 ;
      RECT 90.265 8.235 90.435 8.405 ;
      RECT 89.645 2.205 89.815 2.375 ;
      RECT 89.645 3.685 89.815 3.855 ;
      RECT 89.645 8.605 89.815 8.775 ;
      RECT 89.645 10.085 89.815 10.255 ;
      RECT 89.295 1.395 89.465 1.565 ;
      RECT 89.295 5.455 89.465 5.625 ;
      RECT 89.295 6.835 89.465 7.005 ;
      RECT 89.295 10.895 89.465 11.065 ;
      RECT 89.275 4.055 89.445 4.225 ;
      RECT 89.275 8.235 89.445 8.405 ;
      RECT 88.595 1.4 88.765 1.57 ;
      RECT 88.595 5.46 88.765 5.63 ;
      RECT 88.595 6.83 88.765 7 ;
      RECT 88.595 10.89 88.765 11.06 ;
      RECT 88.285 3.32 88.455 3.49 ;
      RECT 88.285 8.97 88.455 9.14 ;
      RECT 87.915 1.4 88.085 1.57 ;
      RECT 87.915 10.89 88.085 11.06 ;
      RECT 87.855 2.21 88.025 2.38 ;
      RECT 87.855 2.95 88.025 3.12 ;
      RECT 87.855 9.34 88.025 9.51 ;
      RECT 87.855 10.08 88.025 10.25 ;
      RECT 87.48 3.69 87.65 3.86 ;
      RECT 87.48 8.6 87.65 8.77 ;
      RECT 87.235 1.4 87.405 1.57 ;
      RECT 87.235 10.89 87.405 11.06 ;
      RECT 86.555 1.4 86.725 1.57 ;
      RECT 86.555 10.89 86.725 11.06 ;
      RECT 84.93 2.71 85.1 2.88 ;
      RECT 84.93 5.43 85.1 5.6 ;
      RECT 84.56 4.17 84.73 4.34 ;
      RECT 84.47 2.71 84.64 2.88 ;
      RECT 84.47 5.43 84.64 5.6 ;
      RECT 84.24 3.34 84.41 3.51 ;
      RECT 84.095 3.78 84.265 3.95 ;
      RECT 84.01 2.71 84.18 2.88 ;
      RECT 84.01 5.43 84.18 5.6 ;
      RECT 83.815 6.83 83.985 7 ;
      RECT 83.815 10.89 83.985 11.06 ;
      RECT 83.55 2.71 83.72 2.88 ;
      RECT 83.55 5.43 83.72 5.6 ;
      RECT 83.505 8.97 83.675 9.14 ;
      RECT 83.485 3.82 83.655 3.99 ;
      RECT 83.14 3.455 83.31 3.625 ;
      RECT 83.135 10.89 83.305 11.06 ;
      RECT 83.13 4.815 83.3 4.985 ;
      RECT 83.09 2.71 83.26 2.88 ;
      RECT 83.09 5.43 83.26 5.6 ;
      RECT 83.075 9.34 83.245 9.51 ;
      RECT 83.075 10.08 83.245 10.25 ;
      RECT 82.715 4.055 82.885 4.225 ;
      RECT 82.7 8.6 82.87 8.77 ;
      RECT 82.63 2.71 82.8 2.88 ;
      RECT 82.63 5.43 82.8 5.6 ;
      RECT 82.455 10.89 82.625 11.06 ;
      RECT 82.365 3.53 82.535 3.7 ;
      RECT 82.185 4.845 82.355 5.015 ;
      RECT 82.17 2.71 82.34 2.88 ;
      RECT 82.17 5.43 82.34 5.6 ;
      RECT 81.905 4.16 82.075 4.33 ;
      RECT 81.775 10.89 81.945 11.06 ;
      RECT 81.71 2.71 81.88 2.88 ;
      RECT 81.71 5.43 81.88 5.6 ;
      RECT 81.585 3.785 81.755 3.955 ;
      RECT 81.25 2.71 81.42 2.88 ;
      RECT 81.25 5.43 81.42 5.6 ;
      RECT 80.895 3.265 81.065 3.435 ;
      RECT 80.82 3.735 80.99 3.905 ;
      RECT 80.79 2.71 80.96 2.88 ;
      RECT 80.79 5.43 80.96 5.6 ;
      RECT 80.33 2.71 80.5 2.88 ;
      RECT 80.33 5.43 80.5 5.6 ;
      RECT 79.97 3.46 80.14 3.63 ;
      RECT 79.87 2.71 80.04 2.88 ;
      RECT 79.87 5.43 80.04 5.6 ;
      RECT 79.63 4.655 79.8 4.825 ;
      RECT 79.595 3.99 79.765 4.16 ;
      RECT 79.41 2.71 79.58 2.88 ;
      RECT 79.41 5.43 79.58 5.6 ;
      RECT 78.985 3.845 79.155 4.015 ;
      RECT 78.95 2.71 79.12 2.88 ;
      RECT 78.95 5.43 79.12 5.6 ;
      RECT 78.915 4.545 79.085 4.715 ;
      RECT 78.855 3.38 79.025 3.55 ;
      RECT 78.49 2.71 78.66 2.88 ;
      RECT 78.49 5.43 78.66 5.6 ;
      RECT 78.215 4.295 78.385 4.465 ;
      RECT 78.03 2.71 78.2 2.88 ;
      RECT 78.03 5.43 78.2 5.6 ;
      RECT 77.71 3.8 77.88 3.97 ;
      RECT 77.57 2.71 77.74 2.88 ;
      RECT 77.57 5.43 77.74 5.6 ;
      RECT 77.49 4.545 77.66 4.715 ;
      RECT 77.285 3.425 77.455 3.595 ;
      RECT 77.11 2.71 77.28 2.88 ;
      RECT 77.11 5.43 77.28 5.6 ;
      RECT 77.015 4.295 77.185 4.465 ;
      RECT 76.975 3.725 77.145 3.895 ;
      RECT 76.65 2.71 76.82 2.88 ;
      RECT 76.65 5.43 76.82 5.6 ;
      RECT 76.43 4.77 76.6 4.94 ;
      RECT 76.29 3.39 76.46 3.56 ;
      RECT 76.19 2.71 76.36 2.88 ;
      RECT 76.19 5.43 76.36 5.6 ;
      RECT 75.73 2.71 75.9 2.88 ;
      RECT 75.73 5.43 75.9 5.6 ;
      RECT 75.72 4.31 75.89 4.48 ;
      RECT 74.85 8.605 75.02 8.775 ;
      RECT 74.85 10.085 75.02 10.255 ;
      RECT 74.5 1.395 74.67 1.565 ;
      RECT 74.5 5.455 74.67 5.625 ;
      RECT 74.5 6.835 74.67 7.005 ;
      RECT 74.5 10.895 74.67 11.065 ;
      RECT 74.48 4.055 74.65 4.225 ;
      RECT 74.48 8.235 74.65 8.405 ;
      RECT 73.86 2.205 74.03 2.375 ;
      RECT 73.86 3.685 74.03 3.855 ;
      RECT 73.86 8.605 74.03 8.775 ;
      RECT 73.86 10.085 74.03 10.255 ;
      RECT 73.51 1.395 73.68 1.565 ;
      RECT 73.51 5.455 73.68 5.625 ;
      RECT 73.51 6.835 73.68 7.005 ;
      RECT 73.51 10.895 73.68 11.065 ;
      RECT 73.49 4.055 73.66 4.225 ;
      RECT 73.49 8.235 73.66 8.405 ;
      RECT 72.81 1.4 72.98 1.57 ;
      RECT 72.81 5.46 72.98 5.63 ;
      RECT 72.81 6.83 72.98 7 ;
      RECT 72.81 10.89 72.98 11.06 ;
      RECT 72.5 3.32 72.67 3.49 ;
      RECT 72.5 8.97 72.67 9.14 ;
      RECT 72.13 1.4 72.3 1.57 ;
      RECT 72.13 10.89 72.3 11.06 ;
      RECT 72.07 2.21 72.24 2.38 ;
      RECT 72.07 2.95 72.24 3.12 ;
      RECT 72.07 9.34 72.24 9.51 ;
      RECT 72.07 10.08 72.24 10.25 ;
      RECT 71.695 3.69 71.865 3.86 ;
      RECT 71.695 8.6 71.865 8.77 ;
      RECT 71.45 1.4 71.62 1.57 ;
      RECT 71.45 10.89 71.62 11.06 ;
      RECT 70.77 1.4 70.94 1.57 ;
      RECT 70.77 10.89 70.94 11.06 ;
      RECT 69.145 2.71 69.315 2.88 ;
      RECT 69.145 5.43 69.315 5.6 ;
      RECT 68.775 4.17 68.945 4.34 ;
      RECT 68.685 2.71 68.855 2.88 ;
      RECT 68.685 5.43 68.855 5.6 ;
      RECT 68.455 3.34 68.625 3.51 ;
      RECT 68.31 3.78 68.48 3.95 ;
      RECT 68.225 2.71 68.395 2.88 ;
      RECT 68.225 5.43 68.395 5.6 ;
      RECT 68.03 6.83 68.2 7 ;
      RECT 68.03 10.89 68.2 11.06 ;
      RECT 67.765 2.71 67.935 2.88 ;
      RECT 67.765 5.43 67.935 5.6 ;
      RECT 67.72 8.97 67.89 9.14 ;
      RECT 67.7 3.82 67.87 3.99 ;
      RECT 67.355 3.455 67.525 3.625 ;
      RECT 67.35 10.89 67.52 11.06 ;
      RECT 67.345 4.815 67.515 4.985 ;
      RECT 67.305 2.71 67.475 2.88 ;
      RECT 67.305 5.43 67.475 5.6 ;
      RECT 67.29 9.34 67.46 9.51 ;
      RECT 67.29 10.08 67.46 10.25 ;
      RECT 66.93 4.055 67.1 4.225 ;
      RECT 66.915 8.6 67.085 8.77 ;
      RECT 66.845 2.71 67.015 2.88 ;
      RECT 66.845 5.43 67.015 5.6 ;
      RECT 66.67 10.89 66.84 11.06 ;
      RECT 66.58 3.53 66.75 3.7 ;
      RECT 66.4 4.845 66.57 5.015 ;
      RECT 66.385 2.71 66.555 2.88 ;
      RECT 66.385 5.43 66.555 5.6 ;
      RECT 66.12 4.16 66.29 4.33 ;
      RECT 65.99 10.89 66.16 11.06 ;
      RECT 65.925 2.71 66.095 2.88 ;
      RECT 65.925 5.43 66.095 5.6 ;
      RECT 65.8 3.785 65.97 3.955 ;
      RECT 65.465 2.71 65.635 2.88 ;
      RECT 65.465 5.43 65.635 5.6 ;
      RECT 65.11 3.265 65.28 3.435 ;
      RECT 65.035 3.735 65.205 3.905 ;
      RECT 65.005 2.71 65.175 2.88 ;
      RECT 65.005 5.43 65.175 5.6 ;
      RECT 64.545 2.71 64.715 2.88 ;
      RECT 64.545 5.43 64.715 5.6 ;
      RECT 64.185 3.46 64.355 3.63 ;
      RECT 64.085 2.71 64.255 2.88 ;
      RECT 64.085 5.43 64.255 5.6 ;
      RECT 63.845 4.655 64.015 4.825 ;
      RECT 63.81 3.99 63.98 4.16 ;
      RECT 63.625 2.71 63.795 2.88 ;
      RECT 63.625 5.43 63.795 5.6 ;
      RECT 63.2 3.845 63.37 4.015 ;
      RECT 63.165 2.71 63.335 2.88 ;
      RECT 63.165 5.43 63.335 5.6 ;
      RECT 63.13 4.545 63.3 4.715 ;
      RECT 63.07 3.38 63.24 3.55 ;
      RECT 62.705 2.71 62.875 2.88 ;
      RECT 62.705 5.43 62.875 5.6 ;
      RECT 62.43 4.295 62.6 4.465 ;
      RECT 62.245 2.71 62.415 2.88 ;
      RECT 62.245 5.43 62.415 5.6 ;
      RECT 61.925 3.8 62.095 3.97 ;
      RECT 61.785 2.71 61.955 2.88 ;
      RECT 61.785 5.43 61.955 5.6 ;
      RECT 61.705 4.545 61.875 4.715 ;
      RECT 61.5 3.425 61.67 3.595 ;
      RECT 61.325 2.71 61.495 2.88 ;
      RECT 61.325 5.43 61.495 5.6 ;
      RECT 61.23 4.295 61.4 4.465 ;
      RECT 61.19 3.725 61.36 3.895 ;
      RECT 60.865 2.71 61.035 2.88 ;
      RECT 60.865 5.43 61.035 5.6 ;
      RECT 60.645 4.77 60.815 4.94 ;
      RECT 60.505 3.39 60.675 3.56 ;
      RECT 60.405 2.71 60.575 2.88 ;
      RECT 60.405 5.43 60.575 5.6 ;
      RECT 59.945 2.71 60.115 2.88 ;
      RECT 59.945 5.43 60.115 5.6 ;
      RECT 59.935 4.31 60.105 4.48 ;
      RECT 59.065 8.605 59.235 8.775 ;
      RECT 59.065 10.085 59.235 10.255 ;
      RECT 58.715 1.395 58.885 1.565 ;
      RECT 58.715 5.455 58.885 5.625 ;
      RECT 58.715 6.835 58.885 7.005 ;
      RECT 58.715 10.895 58.885 11.065 ;
      RECT 58.695 4.055 58.865 4.225 ;
      RECT 58.695 8.235 58.865 8.405 ;
      RECT 58.075 2.205 58.245 2.375 ;
      RECT 58.075 3.685 58.245 3.855 ;
      RECT 58.075 8.605 58.245 8.775 ;
      RECT 58.075 10.085 58.245 10.255 ;
      RECT 57.725 1.395 57.895 1.565 ;
      RECT 57.725 5.455 57.895 5.625 ;
      RECT 57.725 6.835 57.895 7.005 ;
      RECT 57.725 10.895 57.895 11.065 ;
      RECT 57.705 4.055 57.875 4.225 ;
      RECT 57.705 8.235 57.875 8.405 ;
      RECT 57.025 1.4 57.195 1.57 ;
      RECT 57.025 5.46 57.195 5.63 ;
      RECT 57.025 6.83 57.195 7 ;
      RECT 57.025 10.89 57.195 11.06 ;
      RECT 56.715 3.32 56.885 3.49 ;
      RECT 56.715 8.97 56.885 9.14 ;
      RECT 56.345 1.4 56.515 1.57 ;
      RECT 56.345 10.89 56.515 11.06 ;
      RECT 56.285 2.21 56.455 2.38 ;
      RECT 56.285 2.95 56.455 3.12 ;
      RECT 56.285 9.34 56.455 9.51 ;
      RECT 56.285 10.08 56.455 10.25 ;
      RECT 55.91 3.69 56.08 3.86 ;
      RECT 55.91 8.6 56.08 8.77 ;
      RECT 55.665 1.4 55.835 1.57 ;
      RECT 55.665 10.89 55.835 11.06 ;
      RECT 54.985 1.4 55.155 1.57 ;
      RECT 54.985 10.89 55.155 11.06 ;
      RECT 53.36 2.71 53.53 2.88 ;
      RECT 53.36 5.43 53.53 5.6 ;
      RECT 52.99 4.17 53.16 4.34 ;
      RECT 52.9 2.71 53.07 2.88 ;
      RECT 52.9 5.43 53.07 5.6 ;
      RECT 52.67 3.34 52.84 3.51 ;
      RECT 52.525 3.78 52.695 3.95 ;
      RECT 52.44 2.71 52.61 2.88 ;
      RECT 52.44 5.43 52.61 5.6 ;
      RECT 52.245 6.83 52.415 7 ;
      RECT 52.245 10.89 52.415 11.06 ;
      RECT 51.98 2.71 52.15 2.88 ;
      RECT 51.98 5.43 52.15 5.6 ;
      RECT 51.935 8.97 52.105 9.14 ;
      RECT 51.915 3.82 52.085 3.99 ;
      RECT 51.57 3.455 51.74 3.625 ;
      RECT 51.565 10.89 51.735 11.06 ;
      RECT 51.56 4.815 51.73 4.985 ;
      RECT 51.52 2.71 51.69 2.88 ;
      RECT 51.52 5.43 51.69 5.6 ;
      RECT 51.505 9.34 51.675 9.51 ;
      RECT 51.505 10.08 51.675 10.25 ;
      RECT 51.145 4.055 51.315 4.225 ;
      RECT 51.13 8.6 51.3 8.77 ;
      RECT 51.06 2.71 51.23 2.88 ;
      RECT 51.06 5.43 51.23 5.6 ;
      RECT 50.885 10.89 51.055 11.06 ;
      RECT 50.795 3.53 50.965 3.7 ;
      RECT 50.615 4.845 50.785 5.015 ;
      RECT 50.6 2.71 50.77 2.88 ;
      RECT 50.6 5.43 50.77 5.6 ;
      RECT 50.335 4.16 50.505 4.33 ;
      RECT 50.205 10.89 50.375 11.06 ;
      RECT 50.14 2.71 50.31 2.88 ;
      RECT 50.14 5.43 50.31 5.6 ;
      RECT 50.015 3.785 50.185 3.955 ;
      RECT 49.68 2.71 49.85 2.88 ;
      RECT 49.68 5.43 49.85 5.6 ;
      RECT 49.325 3.265 49.495 3.435 ;
      RECT 49.25 3.735 49.42 3.905 ;
      RECT 49.22 2.71 49.39 2.88 ;
      RECT 49.22 5.43 49.39 5.6 ;
      RECT 48.76 2.71 48.93 2.88 ;
      RECT 48.76 5.43 48.93 5.6 ;
      RECT 48.4 3.46 48.57 3.63 ;
      RECT 48.3 2.71 48.47 2.88 ;
      RECT 48.3 5.43 48.47 5.6 ;
      RECT 48.06 4.655 48.23 4.825 ;
      RECT 48.025 3.99 48.195 4.16 ;
      RECT 47.84 2.71 48.01 2.88 ;
      RECT 47.84 5.43 48.01 5.6 ;
      RECT 47.415 3.845 47.585 4.015 ;
      RECT 47.38 2.71 47.55 2.88 ;
      RECT 47.38 5.43 47.55 5.6 ;
      RECT 47.345 4.545 47.515 4.715 ;
      RECT 47.285 3.38 47.455 3.55 ;
      RECT 46.92 2.71 47.09 2.88 ;
      RECT 46.92 5.43 47.09 5.6 ;
      RECT 46.645 4.295 46.815 4.465 ;
      RECT 46.46 2.71 46.63 2.88 ;
      RECT 46.46 5.43 46.63 5.6 ;
      RECT 46.14 3.8 46.31 3.97 ;
      RECT 46 2.71 46.17 2.88 ;
      RECT 46 5.43 46.17 5.6 ;
      RECT 45.92 4.545 46.09 4.715 ;
      RECT 45.715 3.425 45.885 3.595 ;
      RECT 45.54 2.71 45.71 2.88 ;
      RECT 45.54 5.43 45.71 5.6 ;
      RECT 45.445 4.295 45.615 4.465 ;
      RECT 45.405 3.725 45.575 3.895 ;
      RECT 45.08 2.71 45.25 2.88 ;
      RECT 45.08 5.43 45.25 5.6 ;
      RECT 44.86 4.77 45.03 4.94 ;
      RECT 44.72 3.39 44.89 3.56 ;
      RECT 44.62 2.71 44.79 2.88 ;
      RECT 44.62 5.43 44.79 5.6 ;
      RECT 44.16 2.71 44.33 2.88 ;
      RECT 44.16 5.43 44.33 5.6 ;
      RECT 44.15 4.31 44.32 4.48 ;
      RECT 43.29 8.605 43.46 8.775 ;
      RECT 43.29 10.085 43.46 10.255 ;
      RECT 42.94 1.395 43.11 1.565 ;
      RECT 42.94 5.455 43.11 5.625 ;
      RECT 42.94 6.835 43.11 7.005 ;
      RECT 42.94 10.895 43.11 11.065 ;
      RECT 42.92 4.055 43.09 4.225 ;
      RECT 42.92 8.235 43.09 8.405 ;
      RECT 42.3 2.205 42.47 2.375 ;
      RECT 42.3 3.685 42.47 3.855 ;
      RECT 42.3 8.605 42.47 8.775 ;
      RECT 42.3 10.085 42.47 10.255 ;
      RECT 41.95 1.395 42.12 1.565 ;
      RECT 41.95 5.455 42.12 5.625 ;
      RECT 41.95 6.835 42.12 7.005 ;
      RECT 41.95 10.895 42.12 11.065 ;
      RECT 41.93 4.055 42.1 4.225 ;
      RECT 41.93 8.235 42.1 8.405 ;
      RECT 41.25 1.4 41.42 1.57 ;
      RECT 41.25 5.46 41.42 5.63 ;
      RECT 41.25 6.83 41.42 7 ;
      RECT 41.25 10.89 41.42 11.06 ;
      RECT 40.94 3.32 41.11 3.49 ;
      RECT 40.94 8.97 41.11 9.14 ;
      RECT 40.57 1.4 40.74 1.57 ;
      RECT 40.57 10.89 40.74 11.06 ;
      RECT 40.51 2.21 40.68 2.38 ;
      RECT 40.51 2.95 40.68 3.12 ;
      RECT 40.51 9.34 40.68 9.51 ;
      RECT 40.51 10.08 40.68 10.25 ;
      RECT 40.135 3.69 40.305 3.86 ;
      RECT 40.135 8.6 40.305 8.77 ;
      RECT 39.89 1.4 40.06 1.57 ;
      RECT 39.89 10.89 40.06 11.06 ;
      RECT 39.21 1.4 39.38 1.57 ;
      RECT 39.21 10.89 39.38 11.06 ;
      RECT 37.585 2.71 37.755 2.88 ;
      RECT 37.585 5.43 37.755 5.6 ;
      RECT 37.215 4.17 37.385 4.34 ;
      RECT 37.125 2.71 37.295 2.88 ;
      RECT 37.125 5.43 37.295 5.6 ;
      RECT 36.895 3.34 37.065 3.51 ;
      RECT 36.75 3.78 36.92 3.95 ;
      RECT 36.665 2.71 36.835 2.88 ;
      RECT 36.665 5.43 36.835 5.6 ;
      RECT 36.47 6.83 36.64 7 ;
      RECT 36.47 10.89 36.64 11.06 ;
      RECT 36.205 2.71 36.375 2.88 ;
      RECT 36.205 5.43 36.375 5.6 ;
      RECT 36.16 8.97 36.33 9.14 ;
      RECT 36.14 3.82 36.31 3.99 ;
      RECT 35.795 3.455 35.965 3.625 ;
      RECT 35.79 10.89 35.96 11.06 ;
      RECT 35.785 4.815 35.955 4.985 ;
      RECT 35.745 2.71 35.915 2.88 ;
      RECT 35.745 5.43 35.915 5.6 ;
      RECT 35.73 9.34 35.9 9.51 ;
      RECT 35.73 10.08 35.9 10.25 ;
      RECT 35.37 4.055 35.54 4.225 ;
      RECT 35.355 8.6 35.525 8.77 ;
      RECT 35.285 2.71 35.455 2.88 ;
      RECT 35.285 5.43 35.455 5.6 ;
      RECT 35.11 10.89 35.28 11.06 ;
      RECT 35.02 3.53 35.19 3.7 ;
      RECT 34.84 4.845 35.01 5.015 ;
      RECT 34.825 2.71 34.995 2.88 ;
      RECT 34.825 5.43 34.995 5.6 ;
      RECT 34.56 4.16 34.73 4.33 ;
      RECT 34.43 10.89 34.6 11.06 ;
      RECT 34.365 2.71 34.535 2.88 ;
      RECT 34.365 5.43 34.535 5.6 ;
      RECT 34.24 3.785 34.41 3.955 ;
      RECT 33.905 2.71 34.075 2.88 ;
      RECT 33.905 5.43 34.075 5.6 ;
      RECT 33.55 3.265 33.72 3.435 ;
      RECT 33.475 3.735 33.645 3.905 ;
      RECT 33.445 2.71 33.615 2.88 ;
      RECT 33.445 5.43 33.615 5.6 ;
      RECT 32.985 2.71 33.155 2.88 ;
      RECT 32.985 5.43 33.155 5.6 ;
      RECT 32.625 3.46 32.795 3.63 ;
      RECT 32.525 2.71 32.695 2.88 ;
      RECT 32.525 5.43 32.695 5.6 ;
      RECT 32.285 4.655 32.455 4.825 ;
      RECT 32.25 3.99 32.42 4.16 ;
      RECT 32.065 2.71 32.235 2.88 ;
      RECT 32.065 5.43 32.235 5.6 ;
      RECT 31.64 3.845 31.81 4.015 ;
      RECT 31.605 2.71 31.775 2.88 ;
      RECT 31.605 5.43 31.775 5.6 ;
      RECT 31.57 4.545 31.74 4.715 ;
      RECT 31.51 3.38 31.68 3.55 ;
      RECT 31.145 2.71 31.315 2.88 ;
      RECT 31.145 5.43 31.315 5.6 ;
      RECT 30.87 4.295 31.04 4.465 ;
      RECT 30.685 2.71 30.855 2.88 ;
      RECT 30.685 5.43 30.855 5.6 ;
      RECT 30.365 3.8 30.535 3.97 ;
      RECT 30.225 2.71 30.395 2.88 ;
      RECT 30.225 5.43 30.395 5.6 ;
      RECT 30.145 4.545 30.315 4.715 ;
      RECT 29.94 3.425 30.11 3.595 ;
      RECT 29.765 2.71 29.935 2.88 ;
      RECT 29.765 5.43 29.935 5.6 ;
      RECT 29.67 4.295 29.84 4.465 ;
      RECT 29.63 3.725 29.8 3.895 ;
      RECT 29.305 2.71 29.475 2.88 ;
      RECT 29.305 5.43 29.475 5.6 ;
      RECT 29.085 4.77 29.255 4.94 ;
      RECT 28.945 3.39 29.115 3.56 ;
      RECT 28.845 2.71 29.015 2.88 ;
      RECT 28.845 5.43 29.015 5.6 ;
      RECT 28.385 2.71 28.555 2.88 ;
      RECT 28.385 5.43 28.555 5.6 ;
      RECT 28.375 4.31 28.545 4.48 ;
      RECT 27.51 8.605 27.68 8.775 ;
      RECT 27.51 10.085 27.68 10.255 ;
      RECT 27.16 1.395 27.33 1.565 ;
      RECT 27.16 5.455 27.33 5.625 ;
      RECT 27.16 6.835 27.33 7.005 ;
      RECT 27.16 10.895 27.33 11.065 ;
      RECT 27.14 4.055 27.31 4.225 ;
      RECT 27.14 8.235 27.31 8.405 ;
      RECT 26.52 2.205 26.69 2.375 ;
      RECT 26.52 3.685 26.69 3.855 ;
      RECT 26.52 8.605 26.69 8.775 ;
      RECT 26.52 10.085 26.69 10.255 ;
      RECT 26.17 1.395 26.34 1.565 ;
      RECT 26.17 5.455 26.34 5.625 ;
      RECT 26.17 6.835 26.34 7.005 ;
      RECT 26.17 10.895 26.34 11.065 ;
      RECT 26.15 4.055 26.32 4.225 ;
      RECT 26.15 8.235 26.32 8.405 ;
      RECT 25.47 1.4 25.64 1.57 ;
      RECT 25.47 5.46 25.64 5.63 ;
      RECT 25.47 6.83 25.64 7 ;
      RECT 25.47 10.89 25.64 11.06 ;
      RECT 25.16 3.32 25.33 3.49 ;
      RECT 25.16 8.97 25.33 9.14 ;
      RECT 24.79 1.4 24.96 1.57 ;
      RECT 24.79 10.89 24.96 11.06 ;
      RECT 24.73 2.21 24.9 2.38 ;
      RECT 24.73 2.95 24.9 3.12 ;
      RECT 24.73 9.34 24.9 9.51 ;
      RECT 24.73 10.08 24.9 10.25 ;
      RECT 24.355 3.69 24.525 3.86 ;
      RECT 24.355 8.6 24.525 8.77 ;
      RECT 24.11 1.4 24.28 1.57 ;
      RECT 24.11 10.89 24.28 11.06 ;
      RECT 23.43 1.4 23.6 1.57 ;
      RECT 23.43 10.89 23.6 11.06 ;
      RECT 21.805 2.71 21.975 2.88 ;
      RECT 21.805 5.43 21.975 5.6 ;
      RECT 21.435 4.17 21.605 4.34 ;
      RECT 21.345 2.71 21.515 2.88 ;
      RECT 21.345 5.43 21.515 5.6 ;
      RECT 21.115 3.34 21.285 3.51 ;
      RECT 20.97 3.78 21.14 3.95 ;
      RECT 20.885 2.71 21.055 2.88 ;
      RECT 20.885 5.43 21.055 5.6 ;
      RECT 20.69 6.83 20.86 7 ;
      RECT 20.69 10.89 20.86 11.06 ;
      RECT 20.425 2.71 20.595 2.88 ;
      RECT 20.425 5.43 20.595 5.6 ;
      RECT 20.38 8.97 20.55 9.14 ;
      RECT 20.36 3.82 20.53 3.99 ;
      RECT 20.015 3.455 20.185 3.625 ;
      RECT 20.01 10.89 20.18 11.06 ;
      RECT 20.005 4.815 20.175 4.985 ;
      RECT 19.965 2.71 20.135 2.88 ;
      RECT 19.965 5.43 20.135 5.6 ;
      RECT 19.95 9.34 20.12 9.51 ;
      RECT 19.95 10.08 20.12 10.25 ;
      RECT 19.59 4.055 19.76 4.225 ;
      RECT 19.575 8.6 19.745 8.77 ;
      RECT 19.505 2.71 19.675 2.88 ;
      RECT 19.505 5.43 19.675 5.6 ;
      RECT 19.33 10.89 19.5 11.06 ;
      RECT 19.24 3.53 19.41 3.7 ;
      RECT 19.06 4.845 19.23 5.015 ;
      RECT 19.045 2.71 19.215 2.88 ;
      RECT 19.045 5.43 19.215 5.6 ;
      RECT 18.78 4.16 18.95 4.33 ;
      RECT 18.65 10.89 18.82 11.06 ;
      RECT 18.585 2.71 18.755 2.88 ;
      RECT 18.585 5.43 18.755 5.6 ;
      RECT 18.46 3.785 18.63 3.955 ;
      RECT 18.125 2.71 18.295 2.88 ;
      RECT 18.125 5.43 18.295 5.6 ;
      RECT 17.77 3.265 17.94 3.435 ;
      RECT 17.695 3.735 17.865 3.905 ;
      RECT 17.665 2.71 17.835 2.88 ;
      RECT 17.665 5.43 17.835 5.6 ;
      RECT 17.205 2.71 17.375 2.88 ;
      RECT 17.205 5.43 17.375 5.6 ;
      RECT 16.845 3.46 17.015 3.63 ;
      RECT 16.745 2.71 16.915 2.88 ;
      RECT 16.745 5.43 16.915 5.6 ;
      RECT 16.505 4.655 16.675 4.825 ;
      RECT 16.47 3.99 16.64 4.16 ;
      RECT 16.285 2.71 16.455 2.88 ;
      RECT 16.285 5.43 16.455 5.6 ;
      RECT 15.86 3.845 16.03 4.015 ;
      RECT 15.825 2.71 15.995 2.88 ;
      RECT 15.825 5.43 15.995 5.6 ;
      RECT 15.79 4.545 15.96 4.715 ;
      RECT 15.73 3.38 15.9 3.55 ;
      RECT 15.365 2.71 15.535 2.88 ;
      RECT 15.365 5.43 15.535 5.6 ;
      RECT 15.09 4.295 15.26 4.465 ;
      RECT 14.905 2.71 15.075 2.88 ;
      RECT 14.905 5.43 15.075 5.6 ;
      RECT 14.585 3.8 14.755 3.97 ;
      RECT 14.445 2.71 14.615 2.88 ;
      RECT 14.445 5.43 14.615 5.6 ;
      RECT 14.365 4.545 14.535 4.715 ;
      RECT 14.16 3.425 14.33 3.595 ;
      RECT 13.985 2.71 14.155 2.88 ;
      RECT 13.985 5.43 14.155 5.6 ;
      RECT 13.89 4.295 14.06 4.465 ;
      RECT 13.85 3.725 14.02 3.895 ;
      RECT 13.525 2.71 13.695 2.88 ;
      RECT 13.525 5.43 13.695 5.6 ;
      RECT 13.305 4.77 13.475 4.94 ;
      RECT 13.165 3.39 13.335 3.56 ;
      RECT 13.065 2.71 13.235 2.88 ;
      RECT 13.065 5.43 13.235 5.6 ;
      RECT 12.605 2.71 12.775 2.88 ;
      RECT 12.605 5.43 12.775 5.6 ;
      RECT 12.595 4.31 12.765 4.48 ;
      RECT 11.815 6.83 11.985 7 ;
      RECT 11.815 10.89 11.985 11.06 ;
      RECT 11.505 8.97 11.675 9.14 ;
      RECT 11.135 10.89 11.305 11.06 ;
      RECT 11.075 9.34 11.245 9.51 ;
      RECT 11.075 10.08 11.245 10.25 ;
      RECT 10.7 8.6 10.87 8.77 ;
      RECT 10.455 10.89 10.625 11.06 ;
      RECT 9.775 10.89 9.945 11.06 ;
    LAYER li1 ;
      RECT 83.715 0 83.885 3.38 ;
      RECT 81.755 0 81.925 3.38 ;
      RECT 79.315 0 79.485 3.38 ;
      RECT 78.355 0 78.525 3.38 ;
      RECT 77.835 0 78.005 3.38 ;
      RECT 76.875 0 77.045 3.38 ;
      RECT 75.915 0 76.085 3.38 ;
      RECT 67.93 0 68.1 3.38 ;
      RECT 65.97 0 66.14 3.38 ;
      RECT 63.53 0 63.7 3.38 ;
      RECT 62.57 0 62.74 3.38 ;
      RECT 62.05 0 62.22 3.38 ;
      RECT 61.09 0 61.26 3.38 ;
      RECT 60.13 0 60.3 3.38 ;
      RECT 52.145 0 52.315 3.38 ;
      RECT 50.185 0 50.355 3.38 ;
      RECT 47.745 0 47.915 3.38 ;
      RECT 46.785 0 46.955 3.38 ;
      RECT 46.265 0 46.435 3.38 ;
      RECT 45.305 0 45.475 3.38 ;
      RECT 44.345 0 44.515 3.38 ;
      RECT 36.37 0 36.54 3.38 ;
      RECT 34.41 0 34.58 3.38 ;
      RECT 31.97 0 32.14 3.38 ;
      RECT 31.01 0 31.18 3.38 ;
      RECT 30.49 0 30.66 3.38 ;
      RECT 29.53 0 29.7 3.38 ;
      RECT 28.57 0 28.74 3.38 ;
      RECT 20.59 0 20.76 3.38 ;
      RECT 18.63 0 18.8 3.38 ;
      RECT 16.19 0 16.36 3.38 ;
      RECT 15.23 0 15.4 3.38 ;
      RECT 14.71 0 14.88 3.38 ;
      RECT 13.75 0 13.92 3.38 ;
      RECT 12.79 0 12.96 3.38 ;
      RECT 75.7 0 85.3 2.885 ;
      RECT 59.915 0 69.515 2.885 ;
      RECT 44.13 0 53.73 2.885 ;
      RECT 28.355 0 37.955 2.885 ;
      RECT 12.575 0 22.175 2.885 ;
      RECT 75.585 2.71 85.415 2.88 ;
      RECT 75.7 0 85.415 2.88 ;
      RECT 59.8 2.71 69.63 2.88 ;
      RECT 59.915 0 69.63 2.88 ;
      RECT 44.015 2.71 53.845 2.88 ;
      RECT 44.13 0 53.845 2.88 ;
      RECT 28.24 2.71 38.07 2.88 ;
      RECT 28.355 0 38.07 2.88 ;
      RECT 12.46 2.71 22.29 2.88 ;
      RECT 12.575 0 22.29 2.88 ;
      RECT 86.475 0 86.645 2.23 ;
      RECT 70.69 0 70.86 2.23 ;
      RECT 54.905 0 55.075 2.23 ;
      RECT 39.13 0 39.3 2.23 ;
      RECT 23.35 0 23.52 2.23 ;
      RECT 90.205 0 90.375 2.225 ;
      RECT 89.215 0 89.385 2.225 ;
      RECT 74.42 0 74.59 2.225 ;
      RECT 73.43 0 73.6 2.225 ;
      RECT 58.635 0 58.805 2.225 ;
      RECT 57.645 0 57.815 2.225 ;
      RECT 42.86 0 43.03 2.225 ;
      RECT 41.87 0 42.04 2.225 ;
      RECT 27.08 0 27.25 2.225 ;
      RECT 26.09 0 26.26 2.225 ;
      RECT 9.415 0 91.185 1.6 ;
      RECT 9.41 10.86 91.185 12.46 ;
      RECT 90.205 10.235 90.375 12.46 ;
      RECT 89.215 10.235 89.385 12.46 ;
      RECT 86.475 10.23 86.645 12.46 ;
      RECT 81.695 10.23 81.865 12.46 ;
      RECT 74.42 10.235 74.59 12.46 ;
      RECT 73.43 10.235 73.6 12.46 ;
      RECT 70.69 10.23 70.86 12.46 ;
      RECT 65.91 10.23 66.08 12.46 ;
      RECT 58.635 10.235 58.805 12.46 ;
      RECT 57.645 10.235 57.815 12.46 ;
      RECT 54.905 10.23 55.075 12.46 ;
      RECT 50.125 10.23 50.295 12.46 ;
      RECT 42.86 10.235 43.03 12.46 ;
      RECT 41.87 10.235 42.04 12.46 ;
      RECT 39.13 10.23 39.3 12.46 ;
      RECT 34.35 10.23 34.52 12.46 ;
      RECT 27.08 10.235 27.25 12.46 ;
      RECT 26.09 10.235 26.26 12.46 ;
      RECT 23.35 10.23 23.52 12.46 ;
      RECT 18.57 10.23 18.74 12.46 ;
      RECT 9.41 10.85 10.22 12.46 ;
      RECT 9.695 10.83 9.88 12.46 ;
      RECT 9.695 10.23 9.865 12.46 ;
      RECT 11.505 5.43 11.675 10.59 ;
      RECT 90.205 4.695 90.375 7.765 ;
      RECT 89.215 4.695 89.385 7.765 ;
      RECT 74.42 4.695 74.59 7.765 ;
      RECT 73.43 4.695 73.6 7.765 ;
      RECT 58.635 4.695 58.805 7.765 ;
      RECT 57.645 4.695 57.815 7.765 ;
      RECT 42.86 4.695 43.03 7.765 ;
      RECT 41.87 4.695 42.04 7.765 ;
      RECT 27.08 4.695 27.25 7.765 ;
      RECT 26.09 4.695 26.26 7.765 ;
      RECT 86.475 4.7 86.645 7.76 ;
      RECT 81.695 5.43 81.865 7.76 ;
      RECT 70.69 4.7 70.86 7.76 ;
      RECT 65.91 5.43 66.08 7.76 ;
      RECT 54.905 4.7 55.075 7.76 ;
      RECT 50.125 5.43 50.295 7.76 ;
      RECT 39.13 4.7 39.3 7.76 ;
      RECT 34.35 5.43 34.52 7.76 ;
      RECT 23.35 4.7 23.52 7.76 ;
      RECT 18.57 5.43 18.74 7.76 ;
      RECT 9.695 5.43 9.865 7.76 ;
      RECT 89.045 5.425 91.025 7.035 ;
      RECT 73.26 5.425 75.24 7.035 ;
      RECT 57.475 5.425 59.455 7.035 ;
      RECT 41.7 5.425 43.68 7.035 ;
      RECT 25.92 5.425 27.9 7.035 ;
      RECT 9.415 5.43 91.18 7.03 ;
      RECT 84.675 4.93 84.845 7.03 ;
      RECT 83.715 4.93 83.885 7.03 ;
      RECT 81.275 4.93 81.445 7.03 ;
      RECT 80.275 4.93 80.445 7.03 ;
      RECT 79.315 4.93 79.485 7.03 ;
      RECT 76.875 4.93 77.045 7.03 ;
      RECT 68.89 4.93 69.06 7.03 ;
      RECT 67.93 4.93 68.1 7.03 ;
      RECT 65.49 4.93 65.66 7.03 ;
      RECT 64.49 4.93 64.66 7.03 ;
      RECT 63.53 4.93 63.7 7.03 ;
      RECT 61.09 4.93 61.26 7.03 ;
      RECT 53.105 4.93 53.275 7.03 ;
      RECT 52.145 4.93 52.315 7.03 ;
      RECT 49.705 4.93 49.875 7.03 ;
      RECT 48.705 4.93 48.875 7.03 ;
      RECT 47.745 4.93 47.915 7.03 ;
      RECT 45.305 4.93 45.475 7.03 ;
      RECT 37.33 4.93 37.5 7.03 ;
      RECT 36.37 4.93 36.54 7.03 ;
      RECT 33.93 4.93 34.1 7.03 ;
      RECT 32.93 4.93 33.1 7.03 ;
      RECT 31.97 4.93 32.14 7.03 ;
      RECT 29.53 4.93 29.7 7.03 ;
      RECT 21.55 4.93 21.72 7.03 ;
      RECT 20.59 4.93 20.76 7.03 ;
      RECT 18.15 4.93 18.32 7.03 ;
      RECT 17.15 4.93 17.32 7.03 ;
      RECT 16.19 4.93 16.36 7.03 ;
      RECT 13.75 4.93 13.92 7.03 ;
      RECT 90.265 3.035 90.435 4.225 ;
      RECT 90.265 3.035 90.735 3.205 ;
      RECT 90.265 9.255 90.735 9.425 ;
      RECT 90.265 8.235 90.435 9.425 ;
      RECT 89.275 3.035 89.445 4.225 ;
      RECT 89.275 3.035 89.745 3.205 ;
      RECT 89.275 9.255 89.745 9.425 ;
      RECT 89.275 8.235 89.445 9.425 ;
      RECT 87.425 3.93 87.595 5.16 ;
      RECT 87.48 2.15 87.65 4.1 ;
      RECT 87.425 1.87 87.595 2.32 ;
      RECT 87.425 10.14 87.595 10.59 ;
      RECT 87.48 8.36 87.65 10.31 ;
      RECT 87.425 7.3 87.595 8.53 ;
      RECT 86.905 1.87 87.075 5.16 ;
      RECT 86.905 3.37 87.31 3.7 ;
      RECT 86.905 2.53 87.31 2.86 ;
      RECT 86.905 7.3 87.075 10.59 ;
      RECT 86.905 9.6 87.31 9.93 ;
      RECT 86.905 8.76 87.31 9.09 ;
      RECT 84.24 3.27 84.97 3.51 ;
      RECT 84.782 3.065 84.97 3.51 ;
      RECT 84.61 3.077 84.985 3.504 ;
      RECT 84.525 3.092 85.005 3.489 ;
      RECT 84.525 3.107 85.01 3.479 ;
      RECT 84.48 3.127 85.025 3.471 ;
      RECT 84.457 3.162 85.04 3.425 ;
      RECT 84.371 3.185 85.045 3.385 ;
      RECT 84.371 3.203 85.055 3.355 ;
      RECT 84.24 3.272 85.06 3.318 ;
      RECT 84.285 3.215 85.055 3.355 ;
      RECT 84.371 3.167 85.04 3.425 ;
      RECT 84.457 3.136 85.025 3.471 ;
      RECT 84.48 3.117 85.01 3.479 ;
      RECT 84.525 3.09 84.985 3.504 ;
      RECT 84.61 3.072 84.97 3.51 ;
      RECT 84.696 3.066 84.97 3.51 ;
      RECT 84.782 3.061 84.915 3.51 ;
      RECT 84.868 3.056 84.915 3.51 ;
      RECT 84.56 3.954 84.73 4.34 ;
      RECT 84.555 3.954 84.73 4.335 ;
      RECT 84.53 3.954 84.73 4.3 ;
      RECT 84.53 3.982 84.74 4.29 ;
      RECT 84.51 3.982 84.74 4.25 ;
      RECT 84.505 3.982 84.74 4.223 ;
      RECT 84.505 4 84.745 4.215 ;
      RECT 84.45 4 84.745 4.15 ;
      RECT 84.45 4.017 84.755 4.133 ;
      RECT 84.44 4.017 84.755 4.073 ;
      RECT 84.44 4.034 84.76 4.07 ;
      RECT 84.435 3.87 84.605 4.048 ;
      RECT 84.435 3.904 84.691 4.048 ;
      RECT 84.43 4.67 84.435 4.683 ;
      RECT 84.425 4.565 84.43 4.688 ;
      RECT 84.4 4.425 84.425 4.703 ;
      RECT 84.365 4.376 84.4 4.735 ;
      RECT 84.36 4.344 84.365 4.755 ;
      RECT 84.355 4.335 84.36 4.755 ;
      RECT 84.275 4.3 84.355 4.755 ;
      RECT 84.212 4.27 84.275 4.755 ;
      RECT 84.126 4.258 84.212 4.755 ;
      RECT 84.04 4.244 84.126 4.755 ;
      RECT 83.96 4.231 84.04 4.741 ;
      RECT 83.925 4.223 83.96 4.721 ;
      RECT 83.915 4.22 83.925 4.712 ;
      RECT 83.885 4.215 83.915 4.699 ;
      RECT 83.835 4.19 83.885 4.675 ;
      RECT 83.821 4.164 83.835 4.657 ;
      RECT 83.735 4.124 83.821 4.633 ;
      RECT 83.69 4.072 83.735 4.602 ;
      RECT 83.68 4.047 83.69 4.589 ;
      RECT 83.675 3.828 83.68 3.85 ;
      RECT 83.67 4.03 83.68 4.585 ;
      RECT 83.67 3.826 83.675 3.94 ;
      RECT 83.66 3.822 83.67 4.581 ;
      RECT 83.616 3.82 83.66 4.569 ;
      RECT 83.53 3.82 83.616 4.54 ;
      RECT 83.5 3.82 83.53 4.513 ;
      RECT 83.485 3.82 83.5 4.501 ;
      RECT 83.445 3.832 83.485 4.486 ;
      RECT 83.425 3.851 83.445 4.465 ;
      RECT 83.415 3.861 83.425 4.449 ;
      RECT 83.405 3.867 83.415 4.438 ;
      RECT 83.385 3.877 83.405 4.421 ;
      RECT 83.38 3.886 83.385 4.408 ;
      RECT 83.375 3.89 83.38 4.358 ;
      RECT 83.365 3.896 83.375 4.275 ;
      RECT 83.36 3.9 83.365 4.189 ;
      RECT 83.355 3.92 83.36 4.126 ;
      RECT 83.35 3.943 83.355 4.073 ;
      RECT 83.345 3.961 83.35 4.018 ;
      RECT 83.955 3.78 84.125 4.04 ;
      RECT 84.125 3.745 84.17 4.026 ;
      RECT 84.086 3.747 84.175 4.009 ;
      RECT 83.975 3.764 84.261 3.98 ;
      RECT 83.975 3.779 84.265 3.952 ;
      RECT 83.975 3.76 84.175 4.009 ;
      RECT 84 3.748 84.125 4.04 ;
      RECT 84.086 3.746 84.17 4.026 ;
      RECT 83.14 3.135 83.31 3.625 ;
      RECT 83.14 3.135 83.345 3.605 ;
      RECT 83.275 3.055 83.385 3.565 ;
      RECT 83.256 3.059 83.405 3.535 ;
      RECT 83.17 3.067 83.425 3.518 ;
      RECT 83.17 3.073 83.43 3.508 ;
      RECT 83.17 3.082 83.45 3.496 ;
      RECT 83.145 3.107 83.48 3.474 ;
      RECT 83.145 3.127 83.485 3.454 ;
      RECT 83.14 3.14 83.495 3.434 ;
      RECT 83.14 3.207 83.5 3.415 ;
      RECT 83.14 3.34 83.505 3.402 ;
      RECT 83.135 3.145 83.495 3.235 ;
      RECT 83.145 3.102 83.45 3.496 ;
      RECT 83.256 3.057 83.385 3.565 ;
      RECT 83.13 4.81 83.43 5.065 ;
      RECT 83.215 4.776 83.43 5.065 ;
      RECT 83.215 4.779 83.435 4.925 ;
      RECT 83.15 4.8 83.435 4.925 ;
      RECT 83.185 4.79 83.43 5.065 ;
      RECT 83.18 4.795 83.435 4.925 ;
      RECT 83.215 4.774 83.416 5.065 ;
      RECT 83.301 4.765 83.416 5.065 ;
      RECT 83.301 4.759 83.33 5.065 ;
      RECT 82.79 4.4 82.8 4.89 ;
      RECT 82.45 4.335 82.46 4.635 ;
      RECT 82.965 4.507 82.97 4.726 ;
      RECT 82.955 4.487 82.965 4.743 ;
      RECT 82.945 4.467 82.955 4.773 ;
      RECT 82.94 4.457 82.945 4.788 ;
      RECT 82.935 4.453 82.94 4.793 ;
      RECT 82.92 4.445 82.935 4.8 ;
      RECT 82.88 4.425 82.92 4.825 ;
      RECT 82.855 4.407 82.88 4.858 ;
      RECT 82.85 4.405 82.855 4.871 ;
      RECT 82.83 4.402 82.85 4.875 ;
      RECT 82.8 4.4 82.83 4.885 ;
      RECT 82.73 4.402 82.79 4.886 ;
      RECT 82.71 4.402 82.73 4.88 ;
      RECT 82.685 4.4 82.71 4.877 ;
      RECT 82.65 4.395 82.685 4.873 ;
      RECT 82.63 4.389 82.65 4.86 ;
      RECT 82.62 4.386 82.63 4.848 ;
      RECT 82.6 4.383 82.62 4.833 ;
      RECT 82.58 4.379 82.6 4.815 ;
      RECT 82.575 4.376 82.58 4.805 ;
      RECT 82.57 4.375 82.575 4.803 ;
      RECT 82.56 4.372 82.57 4.795 ;
      RECT 82.55 4.366 82.56 4.778 ;
      RECT 82.54 4.36 82.55 4.76 ;
      RECT 82.53 4.354 82.54 4.748 ;
      RECT 82.52 4.348 82.53 4.728 ;
      RECT 82.515 4.344 82.52 4.713 ;
      RECT 82.51 4.342 82.515 4.705 ;
      RECT 82.505 4.34 82.51 4.698 ;
      RECT 82.5 4.338 82.505 4.688 ;
      RECT 82.495 4.336 82.5 4.682 ;
      RECT 82.485 4.335 82.495 4.672 ;
      RECT 82.475 4.335 82.485 4.663 ;
      RECT 82.46 4.335 82.475 4.648 ;
      RECT 82.42 4.335 82.45 4.632 ;
      RECT 82.4 4.337 82.42 4.627 ;
      RECT 82.395 4.342 82.4 4.625 ;
      RECT 82.365 4.35 82.395 4.623 ;
      RECT 82.335 4.365 82.365 4.622 ;
      RECT 82.29 4.387 82.335 4.627 ;
      RECT 82.285 4.402 82.29 4.631 ;
      RECT 82.27 4.407 82.285 4.633 ;
      RECT 82.265 4.411 82.27 4.635 ;
      RECT 82.205 4.434 82.265 4.644 ;
      RECT 82.185 4.46 82.205 4.657 ;
      RECT 82.175 4.467 82.185 4.661 ;
      RECT 82.16 4.474 82.175 4.664 ;
      RECT 82.14 4.484 82.16 4.667 ;
      RECT 82.135 4.492 82.14 4.67 ;
      RECT 82.09 4.497 82.135 4.677 ;
      RECT 82.08 4.5 82.09 4.684 ;
      RECT 82.07 4.5 82.08 4.688 ;
      RECT 82.035 4.502 82.07 4.7 ;
      RECT 82.015 4.505 82.035 4.713 ;
      RECT 81.975 4.508 82.015 4.724 ;
      RECT 81.96 4.51 81.975 4.737 ;
      RECT 81.95 4.51 81.96 4.742 ;
      RECT 81.925 4.511 81.95 4.75 ;
      RECT 81.915 4.513 81.925 4.755 ;
      RECT 81.91 4.514 81.915 4.758 ;
      RECT 81.885 4.512 81.91 4.761 ;
      RECT 81.87 4.51 81.885 4.762 ;
      RECT 81.85 4.507 81.87 4.764 ;
      RECT 81.83 4.502 81.85 4.764 ;
      RECT 81.77 4.497 81.83 4.761 ;
      RECT 81.735 4.472 81.77 4.757 ;
      RECT 81.725 4.449 81.735 4.755 ;
      RECT 81.695 4.426 81.725 4.755 ;
      RECT 81.685 4.405 81.695 4.755 ;
      RECT 81.66 4.387 81.685 4.753 ;
      RECT 81.645 4.365 81.66 4.75 ;
      RECT 81.63 4.347 81.645 4.748 ;
      RECT 81.61 4.337 81.63 4.746 ;
      RECT 81.595 4.332 81.61 4.745 ;
      RECT 81.58 4.33 81.595 4.744 ;
      RECT 81.55 4.331 81.58 4.742 ;
      RECT 81.53 4.334 81.55 4.74 ;
      RECT 81.473 4.338 81.53 4.74 ;
      RECT 81.387 4.347 81.473 4.74 ;
      RECT 81.301 4.358 81.387 4.74 ;
      RECT 81.215 4.369 81.301 4.74 ;
      RECT 81.195 4.376 81.215 4.748 ;
      RECT 81.185 4.379 81.195 4.755 ;
      RECT 81.12 4.384 81.185 4.773 ;
      RECT 81.09 4.391 81.12 4.798 ;
      RECT 81.08 4.394 81.09 4.805 ;
      RECT 81.035 4.398 81.08 4.81 ;
      RECT 81.005 4.403 81.035 4.815 ;
      RECT 81.004 4.405 81.005 4.815 ;
      RECT 80.918 4.411 81.004 4.815 ;
      RECT 80.832 4.422 80.918 4.815 ;
      RECT 80.746 4.434 80.832 4.815 ;
      RECT 80.66 4.445 80.746 4.815 ;
      RECT 80.645 4.452 80.66 4.81 ;
      RECT 80.64 4.454 80.645 4.804 ;
      RECT 80.62 4.465 80.64 4.799 ;
      RECT 80.61 4.483 80.62 4.793 ;
      RECT 80.605 4.495 80.61 4.593 ;
      RECT 82.9 3.248 82.92 3.335 ;
      RECT 82.895 3.183 82.9 3.367 ;
      RECT 82.885 3.15 82.895 3.372 ;
      RECT 82.88 3.13 82.885 3.378 ;
      RECT 82.85 3.13 82.88 3.395 ;
      RECT 82.801 3.13 82.85 3.431 ;
      RECT 82.715 3.13 82.801 3.489 ;
      RECT 82.686 3.14 82.715 3.538 ;
      RECT 82.6 3.182 82.686 3.591 ;
      RECT 82.58 3.22 82.6 3.638 ;
      RECT 82.555 3.237 82.58 3.658 ;
      RECT 82.545 3.251 82.555 3.678 ;
      RECT 82.54 3.257 82.545 3.688 ;
      RECT 82.535 3.261 82.54 3.695 ;
      RECT 82.485 3.281 82.535 3.7 ;
      RECT 82.42 3.325 82.485 3.7 ;
      RECT 82.395 3.375 82.42 3.7 ;
      RECT 82.385 3.405 82.395 3.7 ;
      RECT 82.38 3.432 82.385 3.7 ;
      RECT 82.375 3.45 82.38 3.7 ;
      RECT 82.365 3.492 82.375 3.7 ;
      RECT 82.715 4.05 82.885 4.225 ;
      RECT 82.655 3.878 82.715 4.213 ;
      RECT 82.645 3.871 82.655 4.196 ;
      RECT 82.6 4.05 82.885 4.176 ;
      RECT 82.581 4.05 82.885 4.154 ;
      RECT 82.495 4.05 82.885 4.119 ;
      RECT 82.475 3.87 82.645 4.075 ;
      RECT 82.475 4.017 82.88 4.075 ;
      RECT 82.475 3.965 82.855 4.075 ;
      RECT 82.475 3.92 82.82 4.075 ;
      RECT 82.475 3.902 82.785 4.075 ;
      RECT 82.475 3.892 82.78 4.075 ;
      RECT 82.645 10.14 82.815 10.59 ;
      RECT 82.7 8.36 82.87 10.31 ;
      RECT 82.645 7.3 82.815 8.53 ;
      RECT 82.125 7.3 82.295 10.59 ;
      RECT 82.125 9.6 82.53 9.93 ;
      RECT 82.125 8.76 82.53 9.09 ;
      RECT 82.195 4.85 82.385 5.075 ;
      RECT 82.185 4.851 82.39 5.07 ;
      RECT 82.185 4.853 82.4 5.05 ;
      RECT 82.185 4.857 82.405 5.035 ;
      RECT 82.185 4.844 82.355 5.07 ;
      RECT 82.185 4.847 82.38 5.07 ;
      RECT 82.195 4.843 82.355 5.075 ;
      RECT 82.281 4.841 82.355 5.075 ;
      RECT 81.905 4.092 82.075 4.33 ;
      RECT 81.905 4.092 82.161 4.244 ;
      RECT 81.905 4.092 82.165 4.154 ;
      RECT 81.955 3.865 82.175 4.133 ;
      RECT 81.95 3.882 82.18 4.106 ;
      RECT 81.915 4.04 82.18 4.106 ;
      RECT 81.935 3.89 82.075 4.33 ;
      RECT 81.925 3.972 82.185 4.089 ;
      RECT 81.92 4.02 82.185 4.089 ;
      RECT 81.925 3.93 82.18 4.106 ;
      RECT 81.95 3.867 82.175 4.133 ;
      RECT 81.515 3.842 81.685 4.04 ;
      RECT 81.515 3.842 81.73 4.015 ;
      RECT 81.585 3.785 81.755 3.973 ;
      RECT 81.56 3.8 81.755 3.973 ;
      RECT 81.175 3.846 81.205 4.04 ;
      RECT 81.17 3.818 81.175 4.04 ;
      RECT 81.14 3.792 81.17 4.042 ;
      RECT 81.115 3.75 81.14 4.045 ;
      RECT 81.105 3.722 81.115 4.047 ;
      RECT 81.07 3.702 81.105 4.049 ;
      RECT 81.005 3.687 81.07 4.055 ;
      RECT 80.955 3.685 81.005 4.061 ;
      RECT 80.932 3.687 80.955 4.066 ;
      RECT 80.846 3.698 80.932 4.072 ;
      RECT 80.76 3.716 80.846 4.082 ;
      RECT 80.745 3.727 80.76 4.088 ;
      RECT 80.675 3.75 80.745 4.094 ;
      RECT 80.62 3.782 80.675 4.102 ;
      RECT 80.58 3.805 80.62 4.108 ;
      RECT 80.566 3.818 80.58 4.111 ;
      RECT 80.48 3.84 80.566 4.117 ;
      RECT 80.465 3.865 80.48 4.123 ;
      RECT 80.425 3.88 80.465 4.127 ;
      RECT 80.375 3.895 80.425 4.132 ;
      RECT 80.35 3.902 80.375 4.136 ;
      RECT 80.29 3.897 80.35 4.14 ;
      RECT 80.275 3.888 80.29 4.144 ;
      RECT 80.205 3.878 80.275 4.14 ;
      RECT 80.18 3.87 80.2 4.13 ;
      RECT 80.121 3.87 80.18 4.108 ;
      RECT 80.035 3.87 80.121 4.065 ;
      RECT 80.2 3.87 80.205 4.135 ;
      RECT 80.895 3.101 81.065 3.435 ;
      RECT 80.865 3.101 81.065 3.43 ;
      RECT 80.805 3.068 80.865 3.418 ;
      RECT 80.805 3.124 81.075 3.413 ;
      RECT 80.78 3.124 81.075 3.407 ;
      RECT 80.775 3.065 80.805 3.404 ;
      RECT 80.76 3.071 80.895 3.402 ;
      RECT 80.755 3.079 80.98 3.39 ;
      RECT 80.755 3.131 81.09 3.343 ;
      RECT 80.74 3.087 80.98 3.338 ;
      RECT 80.74 3.157 81.1 3.279 ;
      RECT 80.71 3.107 81.065 3.24 ;
      RECT 80.71 3.197 81.11 3.236 ;
      RECT 80.76 3.076 80.98 3.402 ;
      RECT 80.1 3.406 80.155 3.67 ;
      RECT 80.1 3.406 80.22 3.669 ;
      RECT 80.1 3.406 80.245 3.668 ;
      RECT 80.1 3.406 80.31 3.667 ;
      RECT 80.245 3.372 80.325 3.666 ;
      RECT 80.06 3.416 80.47 3.665 ;
      RECT 80.1 3.413 80.47 3.665 ;
      RECT 80.06 3.421 80.475 3.658 ;
      RECT 80.045 3.423 80.475 3.657 ;
      RECT 80.045 3.43 80.48 3.653 ;
      RECT 80.025 3.429 80.475 3.649 ;
      RECT 80.025 3.437 80.485 3.648 ;
      RECT 80.02 3.434 80.48 3.644 ;
      RECT 80.02 3.447 80.495 3.643 ;
      RECT 80.005 3.437 80.485 3.642 ;
      RECT 79.97 3.45 80.495 3.635 ;
      RECT 80.155 3.405 80.465 3.665 ;
      RECT 80.155 3.39 80.415 3.665 ;
      RECT 80.22 3.377 80.35 3.665 ;
      RECT 79.765 4.466 79.78 4.859 ;
      RECT 79.73 4.471 79.78 4.858 ;
      RECT 79.765 4.47 79.825 4.857 ;
      RECT 79.71 4.481 79.825 4.856 ;
      RECT 79.725 4.477 79.825 4.856 ;
      RECT 79.69 4.487 79.9 4.853 ;
      RECT 79.69 4.506 79.945 4.851 ;
      RECT 79.69 4.513 79.95 4.848 ;
      RECT 79.675 4.49 79.9 4.845 ;
      RECT 79.655 4.495 79.9 4.838 ;
      RECT 79.65 4.499 79.9 4.834 ;
      RECT 79.65 4.516 79.96 4.833 ;
      RECT 79.63 4.51 79.945 4.829 ;
      RECT 79.63 4.519 79.965 4.823 ;
      RECT 79.625 4.525 79.965 4.595 ;
      RECT 79.69 4.485 79.825 4.853 ;
      RECT 79.565 3.848 79.765 4.16 ;
      RECT 79.64 3.826 79.765 4.16 ;
      RECT 79.58 3.845 79.77 4.145 ;
      RECT 79.55 3.856 79.77 4.143 ;
      RECT 79.565 3.851 79.775 4.109 ;
      RECT 79.55 3.955 79.78 4.076 ;
      RECT 79.58 3.827 79.765 4.16 ;
      RECT 79.64 3.805 79.74 4.16 ;
      RECT 79.665 3.802 79.74 4.16 ;
      RECT 79.665 3.797 79.685 4.16 ;
      RECT 79.07 3.865 79.245 4.04 ;
      RECT 79.065 3.865 79.245 4.038 ;
      RECT 79.04 3.865 79.245 4.033 ;
      RECT 78.985 3.845 79.155 4.023 ;
      RECT 78.985 3.852 79.22 4.023 ;
      RECT 79.07 4.532 79.085 4.715 ;
      RECT 79.06 4.51 79.07 4.715 ;
      RECT 79.045 4.49 79.06 4.715 ;
      RECT 79.035 4.465 79.045 4.715 ;
      RECT 79.005 4.43 79.035 4.715 ;
      RECT 78.97 4.37 79.005 4.715 ;
      RECT 78.965 4.332 78.97 4.715 ;
      RECT 78.915 4.283 78.965 4.715 ;
      RECT 78.905 4.233 78.915 4.703 ;
      RECT 78.89 4.212 78.905 4.663 ;
      RECT 78.87 4.18 78.89 4.613 ;
      RECT 78.845 4.136 78.87 4.553 ;
      RECT 78.84 4.108 78.845 4.508 ;
      RECT 78.835 4.099 78.84 4.494 ;
      RECT 78.83 4.092 78.835 4.481 ;
      RECT 78.825 4.087 78.83 4.47 ;
      RECT 78.82 4.072 78.825 4.46 ;
      RECT 78.815 4.05 78.82 4.447 ;
      RECT 78.805 4.01 78.815 4.422 ;
      RECT 78.78 3.94 78.805 4.378 ;
      RECT 78.775 3.88 78.78 4.343 ;
      RECT 78.76 3.86 78.775 4.31 ;
      RECT 78.755 3.86 78.76 4.285 ;
      RECT 78.725 3.86 78.755 4.24 ;
      RECT 78.68 3.86 78.725 4.18 ;
      RECT 78.605 3.86 78.68 4.128 ;
      RECT 78.6 3.86 78.605 4.093 ;
      RECT 78.595 3.86 78.6 4.083 ;
      RECT 78.59 3.86 78.595 4.063 ;
      RECT 78.855 3.08 79.025 3.55 ;
      RECT 78.8 3.073 78.995 3.534 ;
      RECT 78.8 3.087 79.03 3.533 ;
      RECT 78.785 3.088 79.03 3.514 ;
      RECT 78.78 3.106 79.03 3.5 ;
      RECT 78.785 3.089 79.035 3.498 ;
      RECT 78.77 3.12 79.035 3.483 ;
      RECT 78.785 3.095 79.04 3.468 ;
      RECT 78.765 3.135 79.04 3.465 ;
      RECT 78.78 3.107 79.045 3.45 ;
      RECT 78.78 3.119 79.05 3.43 ;
      RECT 78.765 3.135 79.055 3.413 ;
      RECT 78.765 3.145 79.06 3.268 ;
      RECT 78.76 3.145 79.06 3.225 ;
      RECT 78.76 3.16 79.065 3.203 ;
      RECT 78.855 3.07 78.995 3.55 ;
      RECT 78.855 3.068 78.965 3.55 ;
      RECT 78.941 3.065 78.965 3.55 ;
      RECT 78.6 4.732 78.605 4.778 ;
      RECT 78.59 4.58 78.6 4.802 ;
      RECT 78.585 4.425 78.59 4.827 ;
      RECT 78.57 4.387 78.585 4.838 ;
      RECT 78.565 4.37 78.57 4.845 ;
      RECT 78.555 4.358 78.565 4.852 ;
      RECT 78.55 4.349 78.555 4.854 ;
      RECT 78.545 4.347 78.55 4.858 ;
      RECT 78.5 4.338 78.545 4.873 ;
      RECT 78.495 4.33 78.5 4.887 ;
      RECT 78.49 4.327 78.495 4.891 ;
      RECT 78.475 4.322 78.49 4.899 ;
      RECT 78.42 4.312 78.475 4.91 ;
      RECT 78.385 4.3 78.42 4.911 ;
      RECT 78.376 4.295 78.385 4.905 ;
      RECT 78.29 4.295 78.376 4.895 ;
      RECT 78.26 4.295 78.29 4.873 ;
      RECT 78.25 4.295 78.255 4.853 ;
      RECT 78.245 4.295 78.25 4.815 ;
      RECT 78.24 4.295 78.245 4.773 ;
      RECT 78.235 4.295 78.24 4.733 ;
      RECT 78.23 4.295 78.235 4.663 ;
      RECT 78.22 4.295 78.23 4.585 ;
      RECT 78.215 4.295 78.22 4.485 ;
      RECT 78.255 4.295 78.26 4.855 ;
      RECT 77.75 4.377 77.84 4.855 ;
      RECT 77.735 4.38 77.855 4.853 ;
      RECT 77.75 4.379 77.855 4.853 ;
      RECT 77.715 4.386 77.88 4.843 ;
      RECT 77.735 4.38 77.88 4.843 ;
      RECT 77.7 4.392 77.88 4.831 ;
      RECT 77.735 4.383 77.93 4.824 ;
      RECT 77.686 4.4 77.93 4.822 ;
      RECT 77.715 4.39 77.94 4.81 ;
      RECT 77.686 4.411 77.97 4.801 ;
      RECT 77.6 4.435 77.97 4.795 ;
      RECT 77.6 4.448 78.01 4.778 ;
      RECT 77.595 4.47 78.01 4.771 ;
      RECT 77.565 4.485 78.01 4.761 ;
      RECT 77.56 4.496 78.01 4.751 ;
      RECT 77.53 4.509 78.01 4.742 ;
      RECT 77.515 4.527 78.01 4.731 ;
      RECT 77.49 4.54 78.01 4.721 ;
      RECT 77.75 4.376 77.76 4.855 ;
      RECT 77.796 3.8 77.835 4.045 ;
      RECT 77.71 3.8 77.845 4.043 ;
      RECT 77.595 3.825 77.845 4.04 ;
      RECT 77.595 3.825 77.85 4.038 ;
      RECT 77.595 3.825 77.865 4.033 ;
      RECT 77.701 3.8 77.88 4.013 ;
      RECT 77.615 3.808 77.88 4.013 ;
      RECT 77.285 3.16 77.455 3.595 ;
      RECT 77.275 3.194 77.455 3.578 ;
      RECT 77.355 3.13 77.525 3.565 ;
      RECT 77.26 3.205 77.525 3.543 ;
      RECT 77.355 3.14 77.53 3.533 ;
      RECT 77.285 3.192 77.56 3.518 ;
      RECT 77.245 3.218 77.56 3.503 ;
      RECT 77.245 3.26 77.57 3.483 ;
      RECT 77.24 3.285 77.575 3.465 ;
      RECT 77.24 3.295 77.58 3.45 ;
      RECT 77.235 3.232 77.56 3.448 ;
      RECT 77.235 3.305 77.585 3.433 ;
      RECT 77.23 3.242 77.56 3.43 ;
      RECT 77.225 3.326 77.59 3.413 ;
      RECT 77.225 3.358 77.595 3.393 ;
      RECT 77.22 3.272 77.57 3.385 ;
      RECT 77.225 3.257 77.56 3.413 ;
      RECT 77.24 3.227 77.56 3.465 ;
      RECT 77.085 3.814 77.31 4.07 ;
      RECT 77.085 3.847 77.33 4.06 ;
      RECT 77.05 3.847 77.33 4.058 ;
      RECT 77.05 3.86 77.335 4.048 ;
      RECT 77.05 3.88 77.345 4.04 ;
      RECT 77.05 3.977 77.35 4.033 ;
      RECT 77.03 3.725 77.16 4.023 ;
      RECT 76.985 3.88 77.345 3.965 ;
      RECT 76.975 3.725 77.16 3.91 ;
      RECT 76.975 3.757 77.246 3.91 ;
      RECT 76.94 4.287 76.96 4.465 ;
      RECT 76.905 4.24 76.94 4.465 ;
      RECT 76.89 4.18 76.905 4.465 ;
      RECT 76.865 4.127 76.89 4.465 ;
      RECT 76.85 4.08 76.865 4.465 ;
      RECT 76.83 4.057 76.85 4.465 ;
      RECT 76.805 4.022 76.83 4.465 ;
      RECT 76.795 3.868 76.805 4.465 ;
      RECT 76.765 3.863 76.795 4.456 ;
      RECT 76.76 3.86 76.765 4.446 ;
      RECT 76.745 3.86 76.76 4.42 ;
      RECT 76.74 3.86 76.745 4.383 ;
      RECT 76.715 3.86 76.74 4.335 ;
      RECT 76.695 3.86 76.715 4.26 ;
      RECT 76.685 3.86 76.695 4.22 ;
      RECT 76.68 3.86 76.685 4.195 ;
      RECT 76.675 3.86 76.68 4.178 ;
      RECT 76.67 3.86 76.675 4.16 ;
      RECT 76.665 3.861 76.67 4.15 ;
      RECT 76.655 3.863 76.665 4.118 ;
      RECT 76.645 3.865 76.655 4.085 ;
      RECT 76.635 3.868 76.645 4.058 ;
      RECT 76.96 4.295 77.185 4.465 ;
      RECT 76.29 3.107 76.46 3.56 ;
      RECT 76.29 3.107 76.55 3.526 ;
      RECT 76.29 3.107 76.58 3.51 ;
      RECT 76.29 3.107 76.61 3.483 ;
      RECT 76.546 3.085 76.625 3.465 ;
      RECT 76.325 3.092 76.63 3.45 ;
      RECT 76.325 3.1 76.64 3.413 ;
      RECT 76.285 3.127 76.64 3.385 ;
      RECT 76.27 3.14 76.64 3.35 ;
      RECT 76.29 3.115 76.66 3.34 ;
      RECT 76.265 3.18 76.66 3.31 ;
      RECT 76.265 3.21 76.665 3.293 ;
      RECT 76.26 3.24 76.665 3.28 ;
      RECT 76.325 3.089 76.625 3.465 ;
      RECT 76.46 3.086 76.546 3.544 ;
      RECT 76.411 3.087 76.625 3.465 ;
      RECT 76.555 4.747 76.6 4.94 ;
      RECT 76.545 4.717 76.555 4.94 ;
      RECT 76.54 4.702 76.545 4.94 ;
      RECT 76.5 4.612 76.54 4.94 ;
      RECT 76.495 4.525 76.5 4.94 ;
      RECT 76.485 4.495 76.495 4.94 ;
      RECT 76.48 4.455 76.485 4.94 ;
      RECT 76.47 4.417 76.48 4.94 ;
      RECT 76.465 4.382 76.47 4.94 ;
      RECT 76.445 4.335 76.465 4.94 ;
      RECT 76.43 4.26 76.445 4.94 ;
      RECT 76.425 4.215 76.43 4.935 ;
      RECT 76.42 4.195 76.425 4.908 ;
      RECT 76.415 4.175 76.42 4.893 ;
      RECT 76.41 4.15 76.415 4.873 ;
      RECT 76.405 4.128 76.41 4.858 ;
      RECT 76.4 4.106 76.405 4.84 ;
      RECT 76.395 4.085 76.4 4.83 ;
      RECT 76.385 4.057 76.395 4.8 ;
      RECT 76.375 4.02 76.385 4.768 ;
      RECT 76.365 3.98 76.375 4.735 ;
      RECT 76.355 3.958 76.365 4.705 ;
      RECT 76.325 3.91 76.355 4.637 ;
      RECT 76.31 3.87 76.325 4.564 ;
      RECT 76.3 3.87 76.31 4.53 ;
      RECT 76.295 3.87 76.3 4.505 ;
      RECT 76.29 3.87 76.295 4.49 ;
      RECT 76.285 3.87 76.29 4.468 ;
      RECT 76.28 3.87 76.285 4.455 ;
      RECT 76.265 3.87 76.28 4.42 ;
      RECT 76.245 3.87 76.265 4.36 ;
      RECT 76.235 3.87 76.245 4.31 ;
      RECT 76.215 3.87 76.235 4.258 ;
      RECT 76.195 3.87 76.215 4.215 ;
      RECT 76.185 3.87 76.195 4.203 ;
      RECT 76.155 3.87 76.185 4.19 ;
      RECT 76.125 3.891 76.155 4.17 ;
      RECT 76.115 3.919 76.125 4.15 ;
      RECT 76.1 3.936 76.115 4.118 ;
      RECT 76.095 3.95 76.1 4.085 ;
      RECT 76.09 3.958 76.095 4.058 ;
      RECT 76.085 3.966 76.09 4.02 ;
      RECT 76.09 4.49 76.095 4.825 ;
      RECT 76.055 4.477 76.09 4.824 ;
      RECT 75.985 4.417 76.055 4.823 ;
      RECT 75.905 4.36 75.985 4.822 ;
      RECT 75.77 4.32 75.905 4.821 ;
      RECT 75.77 4.507 76.105 4.81 ;
      RECT 75.73 4.507 76.105 4.8 ;
      RECT 75.73 4.525 76.11 4.795 ;
      RECT 75.73 4.615 76.115 4.785 ;
      RECT 75.725 4.31 75.89 4.765 ;
      RECT 75.72 4.31 75.89 4.508 ;
      RECT 75.72 4.467 76.085 4.508 ;
      RECT 75.72 4.455 76.08 4.508 ;
      RECT 74.48 3.035 74.65 4.225 ;
      RECT 74.48 3.035 74.95 3.205 ;
      RECT 74.48 9.255 74.95 9.425 ;
      RECT 74.48 8.235 74.65 9.425 ;
      RECT 73.49 3.035 73.66 4.225 ;
      RECT 73.49 3.035 73.96 3.205 ;
      RECT 73.49 9.255 73.96 9.425 ;
      RECT 73.49 8.235 73.66 9.425 ;
      RECT 71.64 3.93 71.81 5.16 ;
      RECT 71.695 2.15 71.865 4.1 ;
      RECT 71.64 1.87 71.81 2.32 ;
      RECT 71.64 10.14 71.81 10.59 ;
      RECT 71.695 8.36 71.865 10.31 ;
      RECT 71.64 7.3 71.81 8.53 ;
      RECT 71.12 1.87 71.29 5.16 ;
      RECT 71.12 3.37 71.525 3.7 ;
      RECT 71.12 2.53 71.525 2.86 ;
      RECT 71.12 7.3 71.29 10.59 ;
      RECT 71.12 9.6 71.525 9.93 ;
      RECT 71.12 8.76 71.525 9.09 ;
      RECT 68.455 3.27 69.185 3.51 ;
      RECT 68.997 3.065 69.185 3.51 ;
      RECT 68.825 3.077 69.2 3.504 ;
      RECT 68.74 3.092 69.22 3.489 ;
      RECT 68.74 3.107 69.225 3.479 ;
      RECT 68.695 3.127 69.24 3.471 ;
      RECT 68.672 3.162 69.255 3.425 ;
      RECT 68.586 3.185 69.26 3.385 ;
      RECT 68.586 3.203 69.27 3.355 ;
      RECT 68.455 3.272 69.275 3.318 ;
      RECT 68.5 3.215 69.27 3.355 ;
      RECT 68.586 3.167 69.255 3.425 ;
      RECT 68.672 3.136 69.24 3.471 ;
      RECT 68.695 3.117 69.225 3.479 ;
      RECT 68.74 3.09 69.2 3.504 ;
      RECT 68.825 3.072 69.185 3.51 ;
      RECT 68.911 3.066 69.185 3.51 ;
      RECT 68.997 3.061 69.13 3.51 ;
      RECT 69.083 3.056 69.13 3.51 ;
      RECT 68.775 3.954 68.945 4.34 ;
      RECT 68.77 3.954 68.945 4.335 ;
      RECT 68.745 3.954 68.945 4.3 ;
      RECT 68.745 3.982 68.955 4.29 ;
      RECT 68.725 3.982 68.955 4.25 ;
      RECT 68.72 3.982 68.955 4.223 ;
      RECT 68.72 4 68.96 4.215 ;
      RECT 68.665 4 68.96 4.15 ;
      RECT 68.665 4.017 68.97 4.133 ;
      RECT 68.655 4.017 68.97 4.073 ;
      RECT 68.655 4.034 68.975 4.07 ;
      RECT 68.65 3.87 68.82 4.048 ;
      RECT 68.65 3.904 68.906 4.048 ;
      RECT 68.645 4.67 68.65 4.683 ;
      RECT 68.64 4.565 68.645 4.688 ;
      RECT 68.615 4.425 68.64 4.703 ;
      RECT 68.58 4.376 68.615 4.735 ;
      RECT 68.575 4.344 68.58 4.755 ;
      RECT 68.57 4.335 68.575 4.755 ;
      RECT 68.49 4.3 68.57 4.755 ;
      RECT 68.427 4.27 68.49 4.755 ;
      RECT 68.341 4.258 68.427 4.755 ;
      RECT 68.255 4.244 68.341 4.755 ;
      RECT 68.175 4.231 68.255 4.741 ;
      RECT 68.14 4.223 68.175 4.721 ;
      RECT 68.13 4.22 68.14 4.712 ;
      RECT 68.1 4.215 68.13 4.699 ;
      RECT 68.05 4.19 68.1 4.675 ;
      RECT 68.036 4.164 68.05 4.657 ;
      RECT 67.95 4.124 68.036 4.633 ;
      RECT 67.905 4.072 67.95 4.602 ;
      RECT 67.895 4.047 67.905 4.589 ;
      RECT 67.89 3.828 67.895 3.85 ;
      RECT 67.885 4.03 67.895 4.585 ;
      RECT 67.885 3.826 67.89 3.94 ;
      RECT 67.875 3.822 67.885 4.581 ;
      RECT 67.831 3.82 67.875 4.569 ;
      RECT 67.745 3.82 67.831 4.54 ;
      RECT 67.715 3.82 67.745 4.513 ;
      RECT 67.7 3.82 67.715 4.501 ;
      RECT 67.66 3.832 67.7 4.486 ;
      RECT 67.64 3.851 67.66 4.465 ;
      RECT 67.63 3.861 67.64 4.449 ;
      RECT 67.62 3.867 67.63 4.438 ;
      RECT 67.6 3.877 67.62 4.421 ;
      RECT 67.595 3.886 67.6 4.408 ;
      RECT 67.59 3.89 67.595 4.358 ;
      RECT 67.58 3.896 67.59 4.275 ;
      RECT 67.575 3.9 67.58 4.189 ;
      RECT 67.57 3.92 67.575 4.126 ;
      RECT 67.565 3.943 67.57 4.073 ;
      RECT 67.56 3.961 67.565 4.018 ;
      RECT 68.17 3.78 68.34 4.04 ;
      RECT 68.34 3.745 68.385 4.026 ;
      RECT 68.301 3.747 68.39 4.009 ;
      RECT 68.19 3.764 68.476 3.98 ;
      RECT 68.19 3.779 68.48 3.952 ;
      RECT 68.19 3.76 68.39 4.009 ;
      RECT 68.215 3.748 68.34 4.04 ;
      RECT 68.301 3.746 68.385 4.026 ;
      RECT 67.355 3.135 67.525 3.625 ;
      RECT 67.355 3.135 67.56 3.605 ;
      RECT 67.49 3.055 67.6 3.565 ;
      RECT 67.471 3.059 67.62 3.535 ;
      RECT 67.385 3.067 67.64 3.518 ;
      RECT 67.385 3.073 67.645 3.508 ;
      RECT 67.385 3.082 67.665 3.496 ;
      RECT 67.36 3.107 67.695 3.474 ;
      RECT 67.36 3.127 67.7 3.454 ;
      RECT 67.355 3.14 67.71 3.434 ;
      RECT 67.355 3.207 67.715 3.415 ;
      RECT 67.355 3.34 67.72 3.402 ;
      RECT 67.35 3.145 67.71 3.235 ;
      RECT 67.36 3.102 67.665 3.496 ;
      RECT 67.471 3.057 67.6 3.565 ;
      RECT 67.345 4.81 67.645 5.065 ;
      RECT 67.43 4.776 67.645 5.065 ;
      RECT 67.43 4.779 67.65 4.925 ;
      RECT 67.365 4.8 67.65 4.925 ;
      RECT 67.4 4.79 67.645 5.065 ;
      RECT 67.395 4.795 67.65 4.925 ;
      RECT 67.43 4.774 67.631 5.065 ;
      RECT 67.516 4.765 67.631 5.065 ;
      RECT 67.516 4.759 67.545 5.065 ;
      RECT 67.005 4.4 67.015 4.89 ;
      RECT 66.665 4.335 66.675 4.635 ;
      RECT 67.18 4.507 67.185 4.726 ;
      RECT 67.17 4.487 67.18 4.743 ;
      RECT 67.16 4.467 67.17 4.773 ;
      RECT 67.155 4.457 67.16 4.788 ;
      RECT 67.15 4.453 67.155 4.793 ;
      RECT 67.135 4.445 67.15 4.8 ;
      RECT 67.095 4.425 67.135 4.825 ;
      RECT 67.07 4.407 67.095 4.858 ;
      RECT 67.065 4.405 67.07 4.871 ;
      RECT 67.045 4.402 67.065 4.875 ;
      RECT 67.015 4.4 67.045 4.885 ;
      RECT 66.945 4.402 67.005 4.886 ;
      RECT 66.925 4.402 66.945 4.88 ;
      RECT 66.9 4.4 66.925 4.877 ;
      RECT 66.865 4.395 66.9 4.873 ;
      RECT 66.845 4.389 66.865 4.86 ;
      RECT 66.835 4.386 66.845 4.848 ;
      RECT 66.815 4.383 66.835 4.833 ;
      RECT 66.795 4.379 66.815 4.815 ;
      RECT 66.79 4.376 66.795 4.805 ;
      RECT 66.785 4.375 66.79 4.803 ;
      RECT 66.775 4.372 66.785 4.795 ;
      RECT 66.765 4.366 66.775 4.778 ;
      RECT 66.755 4.36 66.765 4.76 ;
      RECT 66.745 4.354 66.755 4.748 ;
      RECT 66.735 4.348 66.745 4.728 ;
      RECT 66.73 4.344 66.735 4.713 ;
      RECT 66.725 4.342 66.73 4.705 ;
      RECT 66.72 4.34 66.725 4.698 ;
      RECT 66.715 4.338 66.72 4.688 ;
      RECT 66.71 4.336 66.715 4.682 ;
      RECT 66.7 4.335 66.71 4.672 ;
      RECT 66.69 4.335 66.7 4.663 ;
      RECT 66.675 4.335 66.69 4.648 ;
      RECT 66.635 4.335 66.665 4.632 ;
      RECT 66.615 4.337 66.635 4.627 ;
      RECT 66.61 4.342 66.615 4.625 ;
      RECT 66.58 4.35 66.61 4.623 ;
      RECT 66.55 4.365 66.58 4.622 ;
      RECT 66.505 4.387 66.55 4.627 ;
      RECT 66.5 4.402 66.505 4.631 ;
      RECT 66.485 4.407 66.5 4.633 ;
      RECT 66.48 4.411 66.485 4.635 ;
      RECT 66.42 4.434 66.48 4.644 ;
      RECT 66.4 4.46 66.42 4.657 ;
      RECT 66.39 4.467 66.4 4.661 ;
      RECT 66.375 4.474 66.39 4.664 ;
      RECT 66.355 4.484 66.375 4.667 ;
      RECT 66.35 4.492 66.355 4.67 ;
      RECT 66.305 4.497 66.35 4.677 ;
      RECT 66.295 4.5 66.305 4.684 ;
      RECT 66.285 4.5 66.295 4.688 ;
      RECT 66.25 4.502 66.285 4.7 ;
      RECT 66.23 4.505 66.25 4.713 ;
      RECT 66.19 4.508 66.23 4.724 ;
      RECT 66.175 4.51 66.19 4.737 ;
      RECT 66.165 4.51 66.175 4.742 ;
      RECT 66.14 4.511 66.165 4.75 ;
      RECT 66.13 4.513 66.14 4.755 ;
      RECT 66.125 4.514 66.13 4.758 ;
      RECT 66.1 4.512 66.125 4.761 ;
      RECT 66.085 4.51 66.1 4.762 ;
      RECT 66.065 4.507 66.085 4.764 ;
      RECT 66.045 4.502 66.065 4.764 ;
      RECT 65.985 4.497 66.045 4.761 ;
      RECT 65.95 4.472 65.985 4.757 ;
      RECT 65.94 4.449 65.95 4.755 ;
      RECT 65.91 4.426 65.94 4.755 ;
      RECT 65.9 4.405 65.91 4.755 ;
      RECT 65.875 4.387 65.9 4.753 ;
      RECT 65.86 4.365 65.875 4.75 ;
      RECT 65.845 4.347 65.86 4.748 ;
      RECT 65.825 4.337 65.845 4.746 ;
      RECT 65.81 4.332 65.825 4.745 ;
      RECT 65.795 4.33 65.81 4.744 ;
      RECT 65.765 4.331 65.795 4.742 ;
      RECT 65.745 4.334 65.765 4.74 ;
      RECT 65.688 4.338 65.745 4.74 ;
      RECT 65.602 4.347 65.688 4.74 ;
      RECT 65.516 4.358 65.602 4.74 ;
      RECT 65.43 4.369 65.516 4.74 ;
      RECT 65.41 4.376 65.43 4.748 ;
      RECT 65.4 4.379 65.41 4.755 ;
      RECT 65.335 4.384 65.4 4.773 ;
      RECT 65.305 4.391 65.335 4.798 ;
      RECT 65.295 4.394 65.305 4.805 ;
      RECT 65.25 4.398 65.295 4.81 ;
      RECT 65.22 4.403 65.25 4.815 ;
      RECT 65.219 4.405 65.22 4.815 ;
      RECT 65.133 4.411 65.219 4.815 ;
      RECT 65.047 4.422 65.133 4.815 ;
      RECT 64.961 4.434 65.047 4.815 ;
      RECT 64.875 4.445 64.961 4.815 ;
      RECT 64.86 4.452 64.875 4.81 ;
      RECT 64.855 4.454 64.86 4.804 ;
      RECT 64.835 4.465 64.855 4.799 ;
      RECT 64.825 4.483 64.835 4.793 ;
      RECT 64.82 4.495 64.825 4.593 ;
      RECT 67.115 3.248 67.135 3.335 ;
      RECT 67.11 3.183 67.115 3.367 ;
      RECT 67.1 3.15 67.11 3.372 ;
      RECT 67.095 3.13 67.1 3.378 ;
      RECT 67.065 3.13 67.095 3.395 ;
      RECT 67.016 3.13 67.065 3.431 ;
      RECT 66.93 3.13 67.016 3.489 ;
      RECT 66.901 3.14 66.93 3.538 ;
      RECT 66.815 3.182 66.901 3.591 ;
      RECT 66.795 3.22 66.815 3.638 ;
      RECT 66.77 3.237 66.795 3.658 ;
      RECT 66.76 3.251 66.77 3.678 ;
      RECT 66.755 3.257 66.76 3.688 ;
      RECT 66.75 3.261 66.755 3.695 ;
      RECT 66.7 3.281 66.75 3.7 ;
      RECT 66.635 3.325 66.7 3.7 ;
      RECT 66.61 3.375 66.635 3.7 ;
      RECT 66.6 3.405 66.61 3.7 ;
      RECT 66.595 3.432 66.6 3.7 ;
      RECT 66.59 3.45 66.595 3.7 ;
      RECT 66.58 3.492 66.59 3.7 ;
      RECT 66.93 4.05 67.1 4.225 ;
      RECT 66.87 3.878 66.93 4.213 ;
      RECT 66.86 3.871 66.87 4.196 ;
      RECT 66.815 4.05 67.1 4.176 ;
      RECT 66.796 4.05 67.1 4.154 ;
      RECT 66.71 4.05 67.1 4.119 ;
      RECT 66.69 3.87 66.86 4.075 ;
      RECT 66.69 4.017 67.095 4.075 ;
      RECT 66.69 3.965 67.07 4.075 ;
      RECT 66.69 3.92 67.035 4.075 ;
      RECT 66.69 3.902 67 4.075 ;
      RECT 66.69 3.892 66.995 4.075 ;
      RECT 66.86 10.14 67.03 10.59 ;
      RECT 66.915 8.36 67.085 10.31 ;
      RECT 66.86 7.3 67.03 8.53 ;
      RECT 66.34 7.3 66.51 10.59 ;
      RECT 66.34 9.6 66.745 9.93 ;
      RECT 66.34 8.76 66.745 9.09 ;
      RECT 66.41 4.85 66.6 5.075 ;
      RECT 66.4 4.851 66.605 5.07 ;
      RECT 66.4 4.853 66.615 5.05 ;
      RECT 66.4 4.857 66.62 5.035 ;
      RECT 66.4 4.844 66.57 5.07 ;
      RECT 66.4 4.847 66.595 5.07 ;
      RECT 66.41 4.843 66.57 5.075 ;
      RECT 66.496 4.841 66.57 5.075 ;
      RECT 66.12 4.092 66.29 4.33 ;
      RECT 66.12 4.092 66.376 4.244 ;
      RECT 66.12 4.092 66.38 4.154 ;
      RECT 66.17 3.865 66.39 4.133 ;
      RECT 66.165 3.882 66.395 4.106 ;
      RECT 66.13 4.04 66.395 4.106 ;
      RECT 66.15 3.89 66.29 4.33 ;
      RECT 66.14 3.972 66.4 4.089 ;
      RECT 66.135 4.02 66.4 4.089 ;
      RECT 66.14 3.93 66.395 4.106 ;
      RECT 66.165 3.867 66.39 4.133 ;
      RECT 65.73 3.842 65.9 4.04 ;
      RECT 65.73 3.842 65.945 4.015 ;
      RECT 65.8 3.785 65.97 3.973 ;
      RECT 65.775 3.8 65.97 3.973 ;
      RECT 65.39 3.846 65.42 4.04 ;
      RECT 65.385 3.818 65.39 4.04 ;
      RECT 65.355 3.792 65.385 4.042 ;
      RECT 65.33 3.75 65.355 4.045 ;
      RECT 65.32 3.722 65.33 4.047 ;
      RECT 65.285 3.702 65.32 4.049 ;
      RECT 65.22 3.687 65.285 4.055 ;
      RECT 65.17 3.685 65.22 4.061 ;
      RECT 65.147 3.687 65.17 4.066 ;
      RECT 65.061 3.698 65.147 4.072 ;
      RECT 64.975 3.716 65.061 4.082 ;
      RECT 64.96 3.727 64.975 4.088 ;
      RECT 64.89 3.75 64.96 4.094 ;
      RECT 64.835 3.782 64.89 4.102 ;
      RECT 64.795 3.805 64.835 4.108 ;
      RECT 64.781 3.818 64.795 4.111 ;
      RECT 64.695 3.84 64.781 4.117 ;
      RECT 64.68 3.865 64.695 4.123 ;
      RECT 64.64 3.88 64.68 4.127 ;
      RECT 64.59 3.895 64.64 4.132 ;
      RECT 64.565 3.902 64.59 4.136 ;
      RECT 64.505 3.897 64.565 4.14 ;
      RECT 64.49 3.888 64.505 4.144 ;
      RECT 64.42 3.878 64.49 4.14 ;
      RECT 64.395 3.87 64.415 4.13 ;
      RECT 64.336 3.87 64.395 4.108 ;
      RECT 64.25 3.87 64.336 4.065 ;
      RECT 64.415 3.87 64.42 4.135 ;
      RECT 65.11 3.101 65.28 3.435 ;
      RECT 65.08 3.101 65.28 3.43 ;
      RECT 65.02 3.068 65.08 3.418 ;
      RECT 65.02 3.124 65.29 3.413 ;
      RECT 64.995 3.124 65.29 3.407 ;
      RECT 64.99 3.065 65.02 3.404 ;
      RECT 64.975 3.071 65.11 3.402 ;
      RECT 64.97 3.079 65.195 3.39 ;
      RECT 64.97 3.131 65.305 3.343 ;
      RECT 64.955 3.087 65.195 3.338 ;
      RECT 64.955 3.157 65.315 3.279 ;
      RECT 64.925 3.107 65.28 3.24 ;
      RECT 64.925 3.197 65.325 3.236 ;
      RECT 64.975 3.076 65.195 3.402 ;
      RECT 64.315 3.406 64.37 3.67 ;
      RECT 64.315 3.406 64.435 3.669 ;
      RECT 64.315 3.406 64.46 3.668 ;
      RECT 64.315 3.406 64.525 3.667 ;
      RECT 64.46 3.372 64.54 3.666 ;
      RECT 64.275 3.416 64.685 3.665 ;
      RECT 64.315 3.413 64.685 3.665 ;
      RECT 64.275 3.421 64.69 3.658 ;
      RECT 64.26 3.423 64.69 3.657 ;
      RECT 64.26 3.43 64.695 3.653 ;
      RECT 64.24 3.429 64.69 3.649 ;
      RECT 64.24 3.437 64.7 3.648 ;
      RECT 64.235 3.434 64.695 3.644 ;
      RECT 64.235 3.447 64.71 3.643 ;
      RECT 64.22 3.437 64.7 3.642 ;
      RECT 64.185 3.45 64.71 3.635 ;
      RECT 64.37 3.405 64.68 3.665 ;
      RECT 64.37 3.39 64.63 3.665 ;
      RECT 64.435 3.377 64.565 3.665 ;
      RECT 63.98 4.466 63.995 4.859 ;
      RECT 63.945 4.471 63.995 4.858 ;
      RECT 63.98 4.47 64.04 4.857 ;
      RECT 63.925 4.481 64.04 4.856 ;
      RECT 63.94 4.477 64.04 4.856 ;
      RECT 63.905 4.487 64.115 4.853 ;
      RECT 63.905 4.506 64.16 4.851 ;
      RECT 63.905 4.513 64.165 4.848 ;
      RECT 63.89 4.49 64.115 4.845 ;
      RECT 63.87 4.495 64.115 4.838 ;
      RECT 63.865 4.499 64.115 4.834 ;
      RECT 63.865 4.516 64.175 4.833 ;
      RECT 63.845 4.51 64.16 4.829 ;
      RECT 63.845 4.519 64.18 4.823 ;
      RECT 63.84 4.525 64.18 4.595 ;
      RECT 63.905 4.485 64.04 4.853 ;
      RECT 63.78 3.848 63.98 4.16 ;
      RECT 63.855 3.826 63.98 4.16 ;
      RECT 63.795 3.845 63.985 4.145 ;
      RECT 63.765 3.856 63.985 4.143 ;
      RECT 63.78 3.851 63.99 4.109 ;
      RECT 63.765 3.955 63.995 4.076 ;
      RECT 63.795 3.827 63.98 4.16 ;
      RECT 63.855 3.805 63.955 4.16 ;
      RECT 63.88 3.802 63.955 4.16 ;
      RECT 63.88 3.797 63.9 4.16 ;
      RECT 63.285 3.865 63.46 4.04 ;
      RECT 63.28 3.865 63.46 4.038 ;
      RECT 63.255 3.865 63.46 4.033 ;
      RECT 63.2 3.845 63.37 4.023 ;
      RECT 63.2 3.852 63.435 4.023 ;
      RECT 63.285 4.532 63.3 4.715 ;
      RECT 63.275 4.51 63.285 4.715 ;
      RECT 63.26 4.49 63.275 4.715 ;
      RECT 63.25 4.465 63.26 4.715 ;
      RECT 63.22 4.43 63.25 4.715 ;
      RECT 63.185 4.37 63.22 4.715 ;
      RECT 63.18 4.332 63.185 4.715 ;
      RECT 63.13 4.283 63.18 4.715 ;
      RECT 63.12 4.233 63.13 4.703 ;
      RECT 63.105 4.212 63.12 4.663 ;
      RECT 63.085 4.18 63.105 4.613 ;
      RECT 63.06 4.136 63.085 4.553 ;
      RECT 63.055 4.108 63.06 4.508 ;
      RECT 63.05 4.099 63.055 4.494 ;
      RECT 63.045 4.092 63.05 4.481 ;
      RECT 63.04 4.087 63.045 4.47 ;
      RECT 63.035 4.072 63.04 4.46 ;
      RECT 63.03 4.05 63.035 4.447 ;
      RECT 63.02 4.01 63.03 4.422 ;
      RECT 62.995 3.94 63.02 4.378 ;
      RECT 62.99 3.88 62.995 4.343 ;
      RECT 62.975 3.86 62.99 4.31 ;
      RECT 62.97 3.86 62.975 4.285 ;
      RECT 62.94 3.86 62.97 4.24 ;
      RECT 62.895 3.86 62.94 4.18 ;
      RECT 62.82 3.86 62.895 4.128 ;
      RECT 62.815 3.86 62.82 4.093 ;
      RECT 62.81 3.86 62.815 4.083 ;
      RECT 62.805 3.86 62.81 4.063 ;
      RECT 63.07 3.08 63.24 3.55 ;
      RECT 63.015 3.073 63.21 3.534 ;
      RECT 63.015 3.087 63.245 3.533 ;
      RECT 63 3.088 63.245 3.514 ;
      RECT 62.995 3.106 63.245 3.5 ;
      RECT 63 3.089 63.25 3.498 ;
      RECT 62.985 3.12 63.25 3.483 ;
      RECT 63 3.095 63.255 3.468 ;
      RECT 62.98 3.135 63.255 3.465 ;
      RECT 62.995 3.107 63.26 3.45 ;
      RECT 62.995 3.119 63.265 3.43 ;
      RECT 62.98 3.135 63.27 3.413 ;
      RECT 62.98 3.145 63.275 3.268 ;
      RECT 62.975 3.145 63.275 3.225 ;
      RECT 62.975 3.16 63.28 3.203 ;
      RECT 63.07 3.07 63.21 3.55 ;
      RECT 63.07 3.068 63.18 3.55 ;
      RECT 63.156 3.065 63.18 3.55 ;
      RECT 62.815 4.732 62.82 4.778 ;
      RECT 62.805 4.58 62.815 4.802 ;
      RECT 62.8 4.425 62.805 4.827 ;
      RECT 62.785 4.387 62.8 4.838 ;
      RECT 62.78 4.37 62.785 4.845 ;
      RECT 62.77 4.358 62.78 4.852 ;
      RECT 62.765 4.349 62.77 4.854 ;
      RECT 62.76 4.347 62.765 4.858 ;
      RECT 62.715 4.338 62.76 4.873 ;
      RECT 62.71 4.33 62.715 4.887 ;
      RECT 62.705 4.327 62.71 4.891 ;
      RECT 62.69 4.322 62.705 4.899 ;
      RECT 62.635 4.312 62.69 4.91 ;
      RECT 62.6 4.3 62.635 4.911 ;
      RECT 62.591 4.295 62.6 4.905 ;
      RECT 62.505 4.295 62.591 4.895 ;
      RECT 62.475 4.295 62.505 4.873 ;
      RECT 62.465 4.295 62.47 4.853 ;
      RECT 62.46 4.295 62.465 4.815 ;
      RECT 62.455 4.295 62.46 4.773 ;
      RECT 62.45 4.295 62.455 4.733 ;
      RECT 62.445 4.295 62.45 4.663 ;
      RECT 62.435 4.295 62.445 4.585 ;
      RECT 62.43 4.295 62.435 4.485 ;
      RECT 62.47 4.295 62.475 4.855 ;
      RECT 61.965 4.377 62.055 4.855 ;
      RECT 61.95 4.38 62.07 4.853 ;
      RECT 61.965 4.379 62.07 4.853 ;
      RECT 61.93 4.386 62.095 4.843 ;
      RECT 61.95 4.38 62.095 4.843 ;
      RECT 61.915 4.392 62.095 4.831 ;
      RECT 61.95 4.383 62.145 4.824 ;
      RECT 61.901 4.4 62.145 4.822 ;
      RECT 61.93 4.39 62.155 4.81 ;
      RECT 61.901 4.411 62.185 4.801 ;
      RECT 61.815 4.435 62.185 4.795 ;
      RECT 61.815 4.448 62.225 4.778 ;
      RECT 61.81 4.47 62.225 4.771 ;
      RECT 61.78 4.485 62.225 4.761 ;
      RECT 61.775 4.496 62.225 4.751 ;
      RECT 61.745 4.509 62.225 4.742 ;
      RECT 61.73 4.527 62.225 4.731 ;
      RECT 61.705 4.54 62.225 4.721 ;
      RECT 61.965 4.376 61.975 4.855 ;
      RECT 62.011 3.8 62.05 4.045 ;
      RECT 61.925 3.8 62.06 4.043 ;
      RECT 61.81 3.825 62.06 4.04 ;
      RECT 61.81 3.825 62.065 4.038 ;
      RECT 61.81 3.825 62.08 4.033 ;
      RECT 61.916 3.8 62.095 4.013 ;
      RECT 61.83 3.808 62.095 4.013 ;
      RECT 61.5 3.16 61.67 3.595 ;
      RECT 61.49 3.194 61.67 3.578 ;
      RECT 61.57 3.13 61.74 3.565 ;
      RECT 61.475 3.205 61.74 3.543 ;
      RECT 61.57 3.14 61.745 3.533 ;
      RECT 61.5 3.192 61.775 3.518 ;
      RECT 61.46 3.218 61.775 3.503 ;
      RECT 61.46 3.26 61.785 3.483 ;
      RECT 61.455 3.285 61.79 3.465 ;
      RECT 61.455 3.295 61.795 3.45 ;
      RECT 61.45 3.232 61.775 3.448 ;
      RECT 61.45 3.305 61.8 3.433 ;
      RECT 61.445 3.242 61.775 3.43 ;
      RECT 61.44 3.326 61.805 3.413 ;
      RECT 61.44 3.358 61.81 3.393 ;
      RECT 61.435 3.272 61.785 3.385 ;
      RECT 61.44 3.257 61.775 3.413 ;
      RECT 61.455 3.227 61.775 3.465 ;
      RECT 61.3 3.814 61.525 4.07 ;
      RECT 61.3 3.847 61.545 4.06 ;
      RECT 61.265 3.847 61.545 4.058 ;
      RECT 61.265 3.86 61.55 4.048 ;
      RECT 61.265 3.88 61.56 4.04 ;
      RECT 61.265 3.977 61.565 4.033 ;
      RECT 61.245 3.725 61.375 4.023 ;
      RECT 61.2 3.88 61.56 3.965 ;
      RECT 61.19 3.725 61.375 3.91 ;
      RECT 61.19 3.757 61.461 3.91 ;
      RECT 61.155 4.287 61.175 4.465 ;
      RECT 61.12 4.24 61.155 4.465 ;
      RECT 61.105 4.18 61.12 4.465 ;
      RECT 61.08 4.127 61.105 4.465 ;
      RECT 61.065 4.08 61.08 4.465 ;
      RECT 61.045 4.057 61.065 4.465 ;
      RECT 61.02 4.022 61.045 4.465 ;
      RECT 61.01 3.868 61.02 4.465 ;
      RECT 60.98 3.863 61.01 4.456 ;
      RECT 60.975 3.86 60.98 4.446 ;
      RECT 60.96 3.86 60.975 4.42 ;
      RECT 60.955 3.86 60.96 4.383 ;
      RECT 60.93 3.86 60.955 4.335 ;
      RECT 60.91 3.86 60.93 4.26 ;
      RECT 60.9 3.86 60.91 4.22 ;
      RECT 60.895 3.86 60.9 4.195 ;
      RECT 60.89 3.86 60.895 4.178 ;
      RECT 60.885 3.86 60.89 4.16 ;
      RECT 60.88 3.861 60.885 4.15 ;
      RECT 60.87 3.863 60.88 4.118 ;
      RECT 60.86 3.865 60.87 4.085 ;
      RECT 60.85 3.868 60.86 4.058 ;
      RECT 61.175 4.295 61.4 4.465 ;
      RECT 60.505 3.107 60.675 3.56 ;
      RECT 60.505 3.107 60.765 3.526 ;
      RECT 60.505 3.107 60.795 3.51 ;
      RECT 60.505 3.107 60.825 3.483 ;
      RECT 60.761 3.085 60.84 3.465 ;
      RECT 60.54 3.092 60.845 3.45 ;
      RECT 60.54 3.1 60.855 3.413 ;
      RECT 60.5 3.127 60.855 3.385 ;
      RECT 60.485 3.14 60.855 3.35 ;
      RECT 60.505 3.115 60.875 3.34 ;
      RECT 60.48 3.18 60.875 3.31 ;
      RECT 60.48 3.21 60.88 3.293 ;
      RECT 60.475 3.24 60.88 3.28 ;
      RECT 60.54 3.089 60.84 3.465 ;
      RECT 60.675 3.086 60.761 3.544 ;
      RECT 60.626 3.087 60.84 3.465 ;
      RECT 60.77 4.747 60.815 4.94 ;
      RECT 60.76 4.717 60.77 4.94 ;
      RECT 60.755 4.702 60.76 4.94 ;
      RECT 60.715 4.612 60.755 4.94 ;
      RECT 60.71 4.525 60.715 4.94 ;
      RECT 60.7 4.495 60.71 4.94 ;
      RECT 60.695 4.455 60.7 4.94 ;
      RECT 60.685 4.417 60.695 4.94 ;
      RECT 60.68 4.382 60.685 4.94 ;
      RECT 60.66 4.335 60.68 4.94 ;
      RECT 60.645 4.26 60.66 4.94 ;
      RECT 60.64 4.215 60.645 4.935 ;
      RECT 60.635 4.195 60.64 4.908 ;
      RECT 60.63 4.175 60.635 4.893 ;
      RECT 60.625 4.15 60.63 4.873 ;
      RECT 60.62 4.128 60.625 4.858 ;
      RECT 60.615 4.106 60.62 4.84 ;
      RECT 60.61 4.085 60.615 4.83 ;
      RECT 60.6 4.057 60.61 4.8 ;
      RECT 60.59 4.02 60.6 4.768 ;
      RECT 60.58 3.98 60.59 4.735 ;
      RECT 60.57 3.958 60.58 4.705 ;
      RECT 60.54 3.91 60.57 4.637 ;
      RECT 60.525 3.87 60.54 4.564 ;
      RECT 60.515 3.87 60.525 4.53 ;
      RECT 60.51 3.87 60.515 4.505 ;
      RECT 60.505 3.87 60.51 4.49 ;
      RECT 60.5 3.87 60.505 4.468 ;
      RECT 60.495 3.87 60.5 4.455 ;
      RECT 60.48 3.87 60.495 4.42 ;
      RECT 60.46 3.87 60.48 4.36 ;
      RECT 60.45 3.87 60.46 4.31 ;
      RECT 60.43 3.87 60.45 4.258 ;
      RECT 60.41 3.87 60.43 4.215 ;
      RECT 60.4 3.87 60.41 4.203 ;
      RECT 60.37 3.87 60.4 4.19 ;
      RECT 60.34 3.891 60.37 4.17 ;
      RECT 60.33 3.919 60.34 4.15 ;
      RECT 60.315 3.936 60.33 4.118 ;
      RECT 60.31 3.95 60.315 4.085 ;
      RECT 60.305 3.958 60.31 4.058 ;
      RECT 60.3 3.966 60.305 4.02 ;
      RECT 60.305 4.49 60.31 4.825 ;
      RECT 60.27 4.477 60.305 4.824 ;
      RECT 60.2 4.417 60.27 4.823 ;
      RECT 60.12 4.36 60.2 4.822 ;
      RECT 59.985 4.32 60.12 4.821 ;
      RECT 59.985 4.507 60.32 4.81 ;
      RECT 59.945 4.507 60.32 4.8 ;
      RECT 59.945 4.525 60.325 4.795 ;
      RECT 59.945 4.615 60.33 4.785 ;
      RECT 59.94 4.31 60.105 4.765 ;
      RECT 59.935 4.31 60.105 4.508 ;
      RECT 59.935 4.467 60.3 4.508 ;
      RECT 59.935 4.455 60.295 4.508 ;
      RECT 58.695 3.035 58.865 4.225 ;
      RECT 58.695 3.035 59.165 3.205 ;
      RECT 58.695 9.255 59.165 9.425 ;
      RECT 58.695 8.235 58.865 9.425 ;
      RECT 57.705 3.035 57.875 4.225 ;
      RECT 57.705 3.035 58.175 3.205 ;
      RECT 57.705 9.255 58.175 9.425 ;
      RECT 57.705 8.235 57.875 9.425 ;
      RECT 55.855 3.93 56.025 5.16 ;
      RECT 55.91 2.15 56.08 4.1 ;
      RECT 55.855 1.87 56.025 2.32 ;
      RECT 55.855 10.14 56.025 10.59 ;
      RECT 55.91 8.36 56.08 10.31 ;
      RECT 55.855 7.3 56.025 8.53 ;
      RECT 55.335 1.87 55.505 5.16 ;
      RECT 55.335 3.37 55.74 3.7 ;
      RECT 55.335 2.53 55.74 2.86 ;
      RECT 55.335 7.3 55.505 10.59 ;
      RECT 55.335 9.6 55.74 9.93 ;
      RECT 55.335 8.76 55.74 9.09 ;
      RECT 52.67 3.27 53.4 3.51 ;
      RECT 53.212 3.065 53.4 3.51 ;
      RECT 53.04 3.077 53.415 3.504 ;
      RECT 52.955 3.092 53.435 3.489 ;
      RECT 52.955 3.107 53.44 3.479 ;
      RECT 52.91 3.127 53.455 3.471 ;
      RECT 52.887 3.162 53.47 3.425 ;
      RECT 52.801 3.185 53.475 3.385 ;
      RECT 52.801 3.203 53.485 3.355 ;
      RECT 52.67 3.272 53.49 3.318 ;
      RECT 52.715 3.215 53.485 3.355 ;
      RECT 52.801 3.167 53.47 3.425 ;
      RECT 52.887 3.136 53.455 3.471 ;
      RECT 52.91 3.117 53.44 3.479 ;
      RECT 52.955 3.09 53.415 3.504 ;
      RECT 53.04 3.072 53.4 3.51 ;
      RECT 53.126 3.066 53.4 3.51 ;
      RECT 53.212 3.061 53.345 3.51 ;
      RECT 53.298 3.056 53.345 3.51 ;
      RECT 52.99 3.954 53.16 4.34 ;
      RECT 52.985 3.954 53.16 4.335 ;
      RECT 52.96 3.954 53.16 4.3 ;
      RECT 52.96 3.982 53.17 4.29 ;
      RECT 52.94 3.982 53.17 4.25 ;
      RECT 52.935 3.982 53.17 4.223 ;
      RECT 52.935 4 53.175 4.215 ;
      RECT 52.88 4 53.175 4.15 ;
      RECT 52.88 4.017 53.185 4.133 ;
      RECT 52.87 4.017 53.185 4.073 ;
      RECT 52.87 4.034 53.19 4.07 ;
      RECT 52.865 3.87 53.035 4.048 ;
      RECT 52.865 3.904 53.121 4.048 ;
      RECT 52.86 4.67 52.865 4.683 ;
      RECT 52.855 4.565 52.86 4.688 ;
      RECT 52.83 4.425 52.855 4.703 ;
      RECT 52.795 4.376 52.83 4.735 ;
      RECT 52.79 4.344 52.795 4.755 ;
      RECT 52.785 4.335 52.79 4.755 ;
      RECT 52.705 4.3 52.785 4.755 ;
      RECT 52.642 4.27 52.705 4.755 ;
      RECT 52.556 4.258 52.642 4.755 ;
      RECT 52.47 4.244 52.556 4.755 ;
      RECT 52.39 4.231 52.47 4.741 ;
      RECT 52.355 4.223 52.39 4.721 ;
      RECT 52.345 4.22 52.355 4.712 ;
      RECT 52.315 4.215 52.345 4.699 ;
      RECT 52.265 4.19 52.315 4.675 ;
      RECT 52.251 4.164 52.265 4.657 ;
      RECT 52.165 4.124 52.251 4.633 ;
      RECT 52.12 4.072 52.165 4.602 ;
      RECT 52.11 4.047 52.12 4.589 ;
      RECT 52.105 3.828 52.11 3.85 ;
      RECT 52.1 4.03 52.11 4.585 ;
      RECT 52.1 3.826 52.105 3.94 ;
      RECT 52.09 3.822 52.1 4.581 ;
      RECT 52.046 3.82 52.09 4.569 ;
      RECT 51.96 3.82 52.046 4.54 ;
      RECT 51.93 3.82 51.96 4.513 ;
      RECT 51.915 3.82 51.93 4.501 ;
      RECT 51.875 3.832 51.915 4.486 ;
      RECT 51.855 3.851 51.875 4.465 ;
      RECT 51.845 3.861 51.855 4.449 ;
      RECT 51.835 3.867 51.845 4.438 ;
      RECT 51.815 3.877 51.835 4.421 ;
      RECT 51.81 3.886 51.815 4.408 ;
      RECT 51.805 3.89 51.81 4.358 ;
      RECT 51.795 3.896 51.805 4.275 ;
      RECT 51.79 3.9 51.795 4.189 ;
      RECT 51.785 3.92 51.79 4.126 ;
      RECT 51.78 3.943 51.785 4.073 ;
      RECT 51.775 3.961 51.78 4.018 ;
      RECT 52.385 3.78 52.555 4.04 ;
      RECT 52.555 3.745 52.6 4.026 ;
      RECT 52.516 3.747 52.605 4.009 ;
      RECT 52.405 3.764 52.691 3.98 ;
      RECT 52.405 3.779 52.695 3.952 ;
      RECT 52.405 3.76 52.605 4.009 ;
      RECT 52.43 3.748 52.555 4.04 ;
      RECT 52.516 3.746 52.6 4.026 ;
      RECT 51.57 3.135 51.74 3.625 ;
      RECT 51.57 3.135 51.775 3.605 ;
      RECT 51.705 3.055 51.815 3.565 ;
      RECT 51.686 3.059 51.835 3.535 ;
      RECT 51.6 3.067 51.855 3.518 ;
      RECT 51.6 3.073 51.86 3.508 ;
      RECT 51.6 3.082 51.88 3.496 ;
      RECT 51.575 3.107 51.91 3.474 ;
      RECT 51.575 3.127 51.915 3.454 ;
      RECT 51.57 3.14 51.925 3.434 ;
      RECT 51.57 3.207 51.93 3.415 ;
      RECT 51.57 3.34 51.935 3.402 ;
      RECT 51.565 3.145 51.925 3.235 ;
      RECT 51.575 3.102 51.88 3.496 ;
      RECT 51.686 3.057 51.815 3.565 ;
      RECT 51.56 4.81 51.86 5.065 ;
      RECT 51.645 4.776 51.86 5.065 ;
      RECT 51.645 4.779 51.865 4.925 ;
      RECT 51.58 4.8 51.865 4.925 ;
      RECT 51.615 4.79 51.86 5.065 ;
      RECT 51.61 4.795 51.865 4.925 ;
      RECT 51.645 4.774 51.846 5.065 ;
      RECT 51.731 4.765 51.846 5.065 ;
      RECT 51.731 4.759 51.76 5.065 ;
      RECT 51.22 4.4 51.23 4.89 ;
      RECT 50.88 4.335 50.89 4.635 ;
      RECT 51.395 4.507 51.4 4.726 ;
      RECT 51.385 4.487 51.395 4.743 ;
      RECT 51.375 4.467 51.385 4.773 ;
      RECT 51.37 4.457 51.375 4.788 ;
      RECT 51.365 4.453 51.37 4.793 ;
      RECT 51.35 4.445 51.365 4.8 ;
      RECT 51.31 4.425 51.35 4.825 ;
      RECT 51.285 4.407 51.31 4.858 ;
      RECT 51.28 4.405 51.285 4.871 ;
      RECT 51.26 4.402 51.28 4.875 ;
      RECT 51.23 4.4 51.26 4.885 ;
      RECT 51.16 4.402 51.22 4.886 ;
      RECT 51.14 4.402 51.16 4.88 ;
      RECT 51.115 4.4 51.14 4.877 ;
      RECT 51.08 4.395 51.115 4.873 ;
      RECT 51.06 4.389 51.08 4.86 ;
      RECT 51.05 4.386 51.06 4.848 ;
      RECT 51.03 4.383 51.05 4.833 ;
      RECT 51.01 4.379 51.03 4.815 ;
      RECT 51.005 4.376 51.01 4.805 ;
      RECT 51 4.375 51.005 4.803 ;
      RECT 50.99 4.372 51 4.795 ;
      RECT 50.98 4.366 50.99 4.778 ;
      RECT 50.97 4.36 50.98 4.76 ;
      RECT 50.96 4.354 50.97 4.748 ;
      RECT 50.95 4.348 50.96 4.728 ;
      RECT 50.945 4.344 50.95 4.713 ;
      RECT 50.94 4.342 50.945 4.705 ;
      RECT 50.935 4.34 50.94 4.698 ;
      RECT 50.93 4.338 50.935 4.688 ;
      RECT 50.925 4.336 50.93 4.682 ;
      RECT 50.915 4.335 50.925 4.672 ;
      RECT 50.905 4.335 50.915 4.663 ;
      RECT 50.89 4.335 50.905 4.648 ;
      RECT 50.85 4.335 50.88 4.632 ;
      RECT 50.83 4.337 50.85 4.627 ;
      RECT 50.825 4.342 50.83 4.625 ;
      RECT 50.795 4.35 50.825 4.623 ;
      RECT 50.765 4.365 50.795 4.622 ;
      RECT 50.72 4.387 50.765 4.627 ;
      RECT 50.715 4.402 50.72 4.631 ;
      RECT 50.7 4.407 50.715 4.633 ;
      RECT 50.695 4.411 50.7 4.635 ;
      RECT 50.635 4.434 50.695 4.644 ;
      RECT 50.615 4.46 50.635 4.657 ;
      RECT 50.605 4.467 50.615 4.661 ;
      RECT 50.59 4.474 50.605 4.664 ;
      RECT 50.57 4.484 50.59 4.667 ;
      RECT 50.565 4.492 50.57 4.67 ;
      RECT 50.52 4.497 50.565 4.677 ;
      RECT 50.51 4.5 50.52 4.684 ;
      RECT 50.5 4.5 50.51 4.688 ;
      RECT 50.465 4.502 50.5 4.7 ;
      RECT 50.445 4.505 50.465 4.713 ;
      RECT 50.405 4.508 50.445 4.724 ;
      RECT 50.39 4.51 50.405 4.737 ;
      RECT 50.38 4.51 50.39 4.742 ;
      RECT 50.355 4.511 50.38 4.75 ;
      RECT 50.345 4.513 50.355 4.755 ;
      RECT 50.34 4.514 50.345 4.758 ;
      RECT 50.315 4.512 50.34 4.761 ;
      RECT 50.3 4.51 50.315 4.762 ;
      RECT 50.28 4.507 50.3 4.764 ;
      RECT 50.26 4.502 50.28 4.764 ;
      RECT 50.2 4.497 50.26 4.761 ;
      RECT 50.165 4.472 50.2 4.757 ;
      RECT 50.155 4.449 50.165 4.755 ;
      RECT 50.125 4.426 50.155 4.755 ;
      RECT 50.115 4.405 50.125 4.755 ;
      RECT 50.09 4.387 50.115 4.753 ;
      RECT 50.075 4.365 50.09 4.75 ;
      RECT 50.06 4.347 50.075 4.748 ;
      RECT 50.04 4.337 50.06 4.746 ;
      RECT 50.025 4.332 50.04 4.745 ;
      RECT 50.01 4.33 50.025 4.744 ;
      RECT 49.98 4.331 50.01 4.742 ;
      RECT 49.96 4.334 49.98 4.74 ;
      RECT 49.903 4.338 49.96 4.74 ;
      RECT 49.817 4.347 49.903 4.74 ;
      RECT 49.731 4.358 49.817 4.74 ;
      RECT 49.645 4.369 49.731 4.74 ;
      RECT 49.625 4.376 49.645 4.748 ;
      RECT 49.615 4.379 49.625 4.755 ;
      RECT 49.55 4.384 49.615 4.773 ;
      RECT 49.52 4.391 49.55 4.798 ;
      RECT 49.51 4.394 49.52 4.805 ;
      RECT 49.465 4.398 49.51 4.81 ;
      RECT 49.435 4.403 49.465 4.815 ;
      RECT 49.434 4.405 49.435 4.815 ;
      RECT 49.348 4.411 49.434 4.815 ;
      RECT 49.262 4.422 49.348 4.815 ;
      RECT 49.176 4.434 49.262 4.815 ;
      RECT 49.09 4.445 49.176 4.815 ;
      RECT 49.075 4.452 49.09 4.81 ;
      RECT 49.07 4.454 49.075 4.804 ;
      RECT 49.05 4.465 49.07 4.799 ;
      RECT 49.04 4.483 49.05 4.793 ;
      RECT 49.035 4.495 49.04 4.593 ;
      RECT 51.33 3.248 51.35 3.335 ;
      RECT 51.325 3.183 51.33 3.367 ;
      RECT 51.315 3.15 51.325 3.372 ;
      RECT 51.31 3.13 51.315 3.378 ;
      RECT 51.28 3.13 51.31 3.395 ;
      RECT 51.231 3.13 51.28 3.431 ;
      RECT 51.145 3.13 51.231 3.489 ;
      RECT 51.116 3.14 51.145 3.538 ;
      RECT 51.03 3.182 51.116 3.591 ;
      RECT 51.01 3.22 51.03 3.638 ;
      RECT 50.985 3.237 51.01 3.658 ;
      RECT 50.975 3.251 50.985 3.678 ;
      RECT 50.97 3.257 50.975 3.688 ;
      RECT 50.965 3.261 50.97 3.695 ;
      RECT 50.915 3.281 50.965 3.7 ;
      RECT 50.85 3.325 50.915 3.7 ;
      RECT 50.825 3.375 50.85 3.7 ;
      RECT 50.815 3.405 50.825 3.7 ;
      RECT 50.81 3.432 50.815 3.7 ;
      RECT 50.805 3.45 50.81 3.7 ;
      RECT 50.795 3.492 50.805 3.7 ;
      RECT 51.145 4.05 51.315 4.225 ;
      RECT 51.085 3.878 51.145 4.213 ;
      RECT 51.075 3.871 51.085 4.196 ;
      RECT 51.03 4.05 51.315 4.176 ;
      RECT 51.011 4.05 51.315 4.154 ;
      RECT 50.925 4.05 51.315 4.119 ;
      RECT 50.905 3.87 51.075 4.075 ;
      RECT 50.905 4.017 51.31 4.075 ;
      RECT 50.905 3.965 51.285 4.075 ;
      RECT 50.905 3.92 51.25 4.075 ;
      RECT 50.905 3.902 51.215 4.075 ;
      RECT 50.905 3.892 51.21 4.075 ;
      RECT 51.075 10.14 51.245 10.59 ;
      RECT 51.13 8.36 51.3 10.31 ;
      RECT 51.075 7.3 51.245 8.53 ;
      RECT 50.555 7.3 50.725 10.59 ;
      RECT 50.555 9.6 50.96 9.93 ;
      RECT 50.555 8.76 50.96 9.09 ;
      RECT 50.625 4.85 50.815 5.075 ;
      RECT 50.615 4.851 50.82 5.07 ;
      RECT 50.615 4.853 50.83 5.05 ;
      RECT 50.615 4.857 50.835 5.035 ;
      RECT 50.615 4.844 50.785 5.07 ;
      RECT 50.615 4.847 50.81 5.07 ;
      RECT 50.625 4.843 50.785 5.075 ;
      RECT 50.711 4.841 50.785 5.075 ;
      RECT 50.335 4.092 50.505 4.33 ;
      RECT 50.335 4.092 50.591 4.244 ;
      RECT 50.335 4.092 50.595 4.154 ;
      RECT 50.385 3.865 50.605 4.133 ;
      RECT 50.38 3.882 50.61 4.106 ;
      RECT 50.345 4.04 50.61 4.106 ;
      RECT 50.365 3.89 50.505 4.33 ;
      RECT 50.355 3.972 50.615 4.089 ;
      RECT 50.35 4.02 50.615 4.089 ;
      RECT 50.355 3.93 50.61 4.106 ;
      RECT 50.38 3.867 50.605 4.133 ;
      RECT 49.945 3.842 50.115 4.04 ;
      RECT 49.945 3.842 50.16 4.015 ;
      RECT 50.015 3.785 50.185 3.973 ;
      RECT 49.99 3.8 50.185 3.973 ;
      RECT 49.605 3.846 49.635 4.04 ;
      RECT 49.6 3.818 49.605 4.04 ;
      RECT 49.57 3.792 49.6 4.042 ;
      RECT 49.545 3.75 49.57 4.045 ;
      RECT 49.535 3.722 49.545 4.047 ;
      RECT 49.5 3.702 49.535 4.049 ;
      RECT 49.435 3.687 49.5 4.055 ;
      RECT 49.385 3.685 49.435 4.061 ;
      RECT 49.362 3.687 49.385 4.066 ;
      RECT 49.276 3.698 49.362 4.072 ;
      RECT 49.19 3.716 49.276 4.082 ;
      RECT 49.175 3.727 49.19 4.088 ;
      RECT 49.105 3.75 49.175 4.094 ;
      RECT 49.05 3.782 49.105 4.102 ;
      RECT 49.01 3.805 49.05 4.108 ;
      RECT 48.996 3.818 49.01 4.111 ;
      RECT 48.91 3.84 48.996 4.117 ;
      RECT 48.895 3.865 48.91 4.123 ;
      RECT 48.855 3.88 48.895 4.127 ;
      RECT 48.805 3.895 48.855 4.132 ;
      RECT 48.78 3.902 48.805 4.136 ;
      RECT 48.72 3.897 48.78 4.14 ;
      RECT 48.705 3.888 48.72 4.144 ;
      RECT 48.635 3.878 48.705 4.14 ;
      RECT 48.61 3.87 48.63 4.13 ;
      RECT 48.551 3.87 48.61 4.108 ;
      RECT 48.465 3.87 48.551 4.065 ;
      RECT 48.63 3.87 48.635 4.135 ;
      RECT 49.325 3.101 49.495 3.435 ;
      RECT 49.295 3.101 49.495 3.43 ;
      RECT 49.235 3.068 49.295 3.418 ;
      RECT 49.235 3.124 49.505 3.413 ;
      RECT 49.21 3.124 49.505 3.407 ;
      RECT 49.205 3.065 49.235 3.404 ;
      RECT 49.19 3.071 49.325 3.402 ;
      RECT 49.185 3.079 49.41 3.39 ;
      RECT 49.185 3.131 49.52 3.343 ;
      RECT 49.17 3.087 49.41 3.338 ;
      RECT 49.17 3.157 49.53 3.279 ;
      RECT 49.14 3.107 49.495 3.24 ;
      RECT 49.14 3.197 49.54 3.236 ;
      RECT 49.19 3.076 49.41 3.402 ;
      RECT 48.53 3.406 48.585 3.67 ;
      RECT 48.53 3.406 48.65 3.669 ;
      RECT 48.53 3.406 48.675 3.668 ;
      RECT 48.53 3.406 48.74 3.667 ;
      RECT 48.675 3.372 48.755 3.666 ;
      RECT 48.49 3.416 48.9 3.665 ;
      RECT 48.53 3.413 48.9 3.665 ;
      RECT 48.49 3.421 48.905 3.658 ;
      RECT 48.475 3.423 48.905 3.657 ;
      RECT 48.475 3.43 48.91 3.653 ;
      RECT 48.455 3.429 48.905 3.649 ;
      RECT 48.455 3.437 48.915 3.648 ;
      RECT 48.45 3.434 48.91 3.644 ;
      RECT 48.45 3.447 48.925 3.643 ;
      RECT 48.435 3.437 48.915 3.642 ;
      RECT 48.4 3.45 48.925 3.635 ;
      RECT 48.585 3.405 48.895 3.665 ;
      RECT 48.585 3.39 48.845 3.665 ;
      RECT 48.65 3.377 48.78 3.665 ;
      RECT 48.195 4.466 48.21 4.859 ;
      RECT 48.16 4.471 48.21 4.858 ;
      RECT 48.195 4.47 48.255 4.857 ;
      RECT 48.14 4.481 48.255 4.856 ;
      RECT 48.155 4.477 48.255 4.856 ;
      RECT 48.12 4.487 48.33 4.853 ;
      RECT 48.12 4.506 48.375 4.851 ;
      RECT 48.12 4.513 48.38 4.848 ;
      RECT 48.105 4.49 48.33 4.845 ;
      RECT 48.085 4.495 48.33 4.838 ;
      RECT 48.08 4.499 48.33 4.834 ;
      RECT 48.08 4.516 48.39 4.833 ;
      RECT 48.06 4.51 48.375 4.829 ;
      RECT 48.06 4.519 48.395 4.823 ;
      RECT 48.055 4.525 48.395 4.595 ;
      RECT 48.12 4.485 48.255 4.853 ;
      RECT 47.995 3.848 48.195 4.16 ;
      RECT 48.07 3.826 48.195 4.16 ;
      RECT 48.01 3.845 48.2 4.145 ;
      RECT 47.98 3.856 48.2 4.143 ;
      RECT 47.995 3.851 48.205 4.109 ;
      RECT 47.98 3.955 48.21 4.076 ;
      RECT 48.01 3.827 48.195 4.16 ;
      RECT 48.07 3.805 48.17 4.16 ;
      RECT 48.095 3.802 48.17 4.16 ;
      RECT 48.095 3.797 48.115 4.16 ;
      RECT 47.5 3.865 47.675 4.04 ;
      RECT 47.495 3.865 47.675 4.038 ;
      RECT 47.47 3.865 47.675 4.033 ;
      RECT 47.415 3.845 47.585 4.023 ;
      RECT 47.415 3.852 47.65 4.023 ;
      RECT 47.5 4.532 47.515 4.715 ;
      RECT 47.49 4.51 47.5 4.715 ;
      RECT 47.475 4.49 47.49 4.715 ;
      RECT 47.465 4.465 47.475 4.715 ;
      RECT 47.435 4.43 47.465 4.715 ;
      RECT 47.4 4.37 47.435 4.715 ;
      RECT 47.395 4.332 47.4 4.715 ;
      RECT 47.345 4.283 47.395 4.715 ;
      RECT 47.335 4.233 47.345 4.703 ;
      RECT 47.32 4.212 47.335 4.663 ;
      RECT 47.3 4.18 47.32 4.613 ;
      RECT 47.275 4.136 47.3 4.553 ;
      RECT 47.27 4.108 47.275 4.508 ;
      RECT 47.265 4.099 47.27 4.494 ;
      RECT 47.26 4.092 47.265 4.481 ;
      RECT 47.255 4.087 47.26 4.47 ;
      RECT 47.25 4.072 47.255 4.46 ;
      RECT 47.245 4.05 47.25 4.447 ;
      RECT 47.235 4.01 47.245 4.422 ;
      RECT 47.21 3.94 47.235 4.378 ;
      RECT 47.205 3.88 47.21 4.343 ;
      RECT 47.19 3.86 47.205 4.31 ;
      RECT 47.185 3.86 47.19 4.285 ;
      RECT 47.155 3.86 47.185 4.24 ;
      RECT 47.11 3.86 47.155 4.18 ;
      RECT 47.035 3.86 47.11 4.128 ;
      RECT 47.03 3.86 47.035 4.093 ;
      RECT 47.025 3.86 47.03 4.083 ;
      RECT 47.02 3.86 47.025 4.063 ;
      RECT 47.285 3.08 47.455 3.55 ;
      RECT 47.23 3.073 47.425 3.534 ;
      RECT 47.23 3.087 47.46 3.533 ;
      RECT 47.215 3.088 47.46 3.514 ;
      RECT 47.21 3.106 47.46 3.5 ;
      RECT 47.215 3.089 47.465 3.498 ;
      RECT 47.2 3.12 47.465 3.483 ;
      RECT 47.215 3.095 47.47 3.468 ;
      RECT 47.195 3.135 47.47 3.465 ;
      RECT 47.21 3.107 47.475 3.45 ;
      RECT 47.21 3.119 47.48 3.43 ;
      RECT 47.195 3.135 47.485 3.413 ;
      RECT 47.195 3.145 47.49 3.268 ;
      RECT 47.19 3.145 47.49 3.225 ;
      RECT 47.19 3.16 47.495 3.203 ;
      RECT 47.285 3.07 47.425 3.55 ;
      RECT 47.285 3.068 47.395 3.55 ;
      RECT 47.371 3.065 47.395 3.55 ;
      RECT 47.03 4.732 47.035 4.778 ;
      RECT 47.02 4.58 47.03 4.802 ;
      RECT 47.015 4.425 47.02 4.827 ;
      RECT 47 4.387 47.015 4.838 ;
      RECT 46.995 4.37 47 4.845 ;
      RECT 46.985 4.358 46.995 4.852 ;
      RECT 46.98 4.349 46.985 4.854 ;
      RECT 46.975 4.347 46.98 4.858 ;
      RECT 46.93 4.338 46.975 4.873 ;
      RECT 46.925 4.33 46.93 4.887 ;
      RECT 46.92 4.327 46.925 4.891 ;
      RECT 46.905 4.322 46.92 4.899 ;
      RECT 46.85 4.312 46.905 4.91 ;
      RECT 46.815 4.3 46.85 4.911 ;
      RECT 46.806 4.295 46.815 4.905 ;
      RECT 46.72 4.295 46.806 4.895 ;
      RECT 46.69 4.295 46.72 4.873 ;
      RECT 46.68 4.295 46.685 4.853 ;
      RECT 46.675 4.295 46.68 4.815 ;
      RECT 46.67 4.295 46.675 4.773 ;
      RECT 46.665 4.295 46.67 4.733 ;
      RECT 46.66 4.295 46.665 4.663 ;
      RECT 46.65 4.295 46.66 4.585 ;
      RECT 46.645 4.295 46.65 4.485 ;
      RECT 46.685 4.295 46.69 4.855 ;
      RECT 46.18 4.377 46.27 4.855 ;
      RECT 46.165 4.38 46.285 4.853 ;
      RECT 46.18 4.379 46.285 4.853 ;
      RECT 46.145 4.386 46.31 4.843 ;
      RECT 46.165 4.38 46.31 4.843 ;
      RECT 46.13 4.392 46.31 4.831 ;
      RECT 46.165 4.383 46.36 4.824 ;
      RECT 46.116 4.4 46.36 4.822 ;
      RECT 46.145 4.39 46.37 4.81 ;
      RECT 46.116 4.411 46.4 4.801 ;
      RECT 46.03 4.435 46.4 4.795 ;
      RECT 46.03 4.448 46.44 4.778 ;
      RECT 46.025 4.47 46.44 4.771 ;
      RECT 45.995 4.485 46.44 4.761 ;
      RECT 45.99 4.496 46.44 4.751 ;
      RECT 45.96 4.509 46.44 4.742 ;
      RECT 45.945 4.527 46.44 4.731 ;
      RECT 45.92 4.54 46.44 4.721 ;
      RECT 46.18 4.376 46.19 4.855 ;
      RECT 46.226 3.8 46.265 4.045 ;
      RECT 46.14 3.8 46.275 4.043 ;
      RECT 46.025 3.825 46.275 4.04 ;
      RECT 46.025 3.825 46.28 4.038 ;
      RECT 46.025 3.825 46.295 4.033 ;
      RECT 46.131 3.8 46.31 4.013 ;
      RECT 46.045 3.808 46.31 4.013 ;
      RECT 45.715 3.16 45.885 3.595 ;
      RECT 45.705 3.194 45.885 3.578 ;
      RECT 45.785 3.13 45.955 3.565 ;
      RECT 45.69 3.205 45.955 3.543 ;
      RECT 45.785 3.14 45.96 3.533 ;
      RECT 45.715 3.192 45.99 3.518 ;
      RECT 45.675 3.218 45.99 3.503 ;
      RECT 45.675 3.26 46 3.483 ;
      RECT 45.67 3.285 46.005 3.465 ;
      RECT 45.67 3.295 46.01 3.45 ;
      RECT 45.665 3.232 45.99 3.448 ;
      RECT 45.665 3.305 46.015 3.433 ;
      RECT 45.66 3.242 45.99 3.43 ;
      RECT 45.655 3.326 46.02 3.413 ;
      RECT 45.655 3.358 46.025 3.393 ;
      RECT 45.65 3.272 46 3.385 ;
      RECT 45.655 3.257 45.99 3.413 ;
      RECT 45.67 3.227 45.99 3.465 ;
      RECT 45.515 3.814 45.74 4.07 ;
      RECT 45.515 3.847 45.76 4.06 ;
      RECT 45.48 3.847 45.76 4.058 ;
      RECT 45.48 3.86 45.765 4.048 ;
      RECT 45.48 3.88 45.775 4.04 ;
      RECT 45.48 3.977 45.78 4.033 ;
      RECT 45.46 3.725 45.59 4.023 ;
      RECT 45.415 3.88 45.775 3.965 ;
      RECT 45.405 3.725 45.59 3.91 ;
      RECT 45.405 3.757 45.676 3.91 ;
      RECT 45.37 4.287 45.39 4.465 ;
      RECT 45.335 4.24 45.37 4.465 ;
      RECT 45.32 4.18 45.335 4.465 ;
      RECT 45.295 4.127 45.32 4.465 ;
      RECT 45.28 4.08 45.295 4.465 ;
      RECT 45.26 4.057 45.28 4.465 ;
      RECT 45.235 4.022 45.26 4.465 ;
      RECT 45.225 3.868 45.235 4.465 ;
      RECT 45.195 3.863 45.225 4.456 ;
      RECT 45.19 3.86 45.195 4.446 ;
      RECT 45.175 3.86 45.19 4.42 ;
      RECT 45.17 3.86 45.175 4.383 ;
      RECT 45.145 3.86 45.17 4.335 ;
      RECT 45.125 3.86 45.145 4.26 ;
      RECT 45.115 3.86 45.125 4.22 ;
      RECT 45.11 3.86 45.115 4.195 ;
      RECT 45.105 3.86 45.11 4.178 ;
      RECT 45.1 3.86 45.105 4.16 ;
      RECT 45.095 3.861 45.1 4.15 ;
      RECT 45.085 3.863 45.095 4.118 ;
      RECT 45.075 3.865 45.085 4.085 ;
      RECT 45.065 3.868 45.075 4.058 ;
      RECT 45.39 4.295 45.615 4.465 ;
      RECT 44.72 3.107 44.89 3.56 ;
      RECT 44.72 3.107 44.98 3.526 ;
      RECT 44.72 3.107 45.01 3.51 ;
      RECT 44.72 3.107 45.04 3.483 ;
      RECT 44.976 3.085 45.055 3.465 ;
      RECT 44.755 3.092 45.06 3.45 ;
      RECT 44.755 3.1 45.07 3.413 ;
      RECT 44.715 3.127 45.07 3.385 ;
      RECT 44.7 3.14 45.07 3.35 ;
      RECT 44.72 3.115 45.09 3.34 ;
      RECT 44.695 3.18 45.09 3.31 ;
      RECT 44.695 3.21 45.095 3.293 ;
      RECT 44.69 3.24 45.095 3.28 ;
      RECT 44.755 3.089 45.055 3.465 ;
      RECT 44.89 3.086 44.976 3.544 ;
      RECT 44.841 3.087 45.055 3.465 ;
      RECT 44.985 4.747 45.03 4.94 ;
      RECT 44.975 4.717 44.985 4.94 ;
      RECT 44.97 4.702 44.975 4.94 ;
      RECT 44.93 4.612 44.97 4.94 ;
      RECT 44.925 4.525 44.93 4.94 ;
      RECT 44.915 4.495 44.925 4.94 ;
      RECT 44.91 4.455 44.915 4.94 ;
      RECT 44.9 4.417 44.91 4.94 ;
      RECT 44.895 4.382 44.9 4.94 ;
      RECT 44.875 4.335 44.895 4.94 ;
      RECT 44.86 4.26 44.875 4.94 ;
      RECT 44.855 4.215 44.86 4.935 ;
      RECT 44.85 4.195 44.855 4.908 ;
      RECT 44.845 4.175 44.85 4.893 ;
      RECT 44.84 4.15 44.845 4.873 ;
      RECT 44.835 4.128 44.84 4.858 ;
      RECT 44.83 4.106 44.835 4.84 ;
      RECT 44.825 4.085 44.83 4.83 ;
      RECT 44.815 4.057 44.825 4.8 ;
      RECT 44.805 4.02 44.815 4.768 ;
      RECT 44.795 3.98 44.805 4.735 ;
      RECT 44.785 3.958 44.795 4.705 ;
      RECT 44.755 3.91 44.785 4.637 ;
      RECT 44.74 3.87 44.755 4.564 ;
      RECT 44.73 3.87 44.74 4.53 ;
      RECT 44.725 3.87 44.73 4.505 ;
      RECT 44.72 3.87 44.725 4.49 ;
      RECT 44.715 3.87 44.72 4.468 ;
      RECT 44.71 3.87 44.715 4.455 ;
      RECT 44.695 3.87 44.71 4.42 ;
      RECT 44.675 3.87 44.695 4.36 ;
      RECT 44.665 3.87 44.675 4.31 ;
      RECT 44.645 3.87 44.665 4.258 ;
      RECT 44.625 3.87 44.645 4.215 ;
      RECT 44.615 3.87 44.625 4.203 ;
      RECT 44.585 3.87 44.615 4.19 ;
      RECT 44.555 3.891 44.585 4.17 ;
      RECT 44.545 3.919 44.555 4.15 ;
      RECT 44.53 3.936 44.545 4.118 ;
      RECT 44.525 3.95 44.53 4.085 ;
      RECT 44.52 3.958 44.525 4.058 ;
      RECT 44.515 3.966 44.52 4.02 ;
      RECT 44.52 4.49 44.525 4.825 ;
      RECT 44.485 4.477 44.52 4.824 ;
      RECT 44.415 4.417 44.485 4.823 ;
      RECT 44.335 4.36 44.415 4.822 ;
      RECT 44.2 4.32 44.335 4.821 ;
      RECT 44.2 4.507 44.535 4.81 ;
      RECT 44.16 4.507 44.535 4.8 ;
      RECT 44.16 4.525 44.54 4.795 ;
      RECT 44.16 4.615 44.545 4.785 ;
      RECT 44.155 4.31 44.32 4.765 ;
      RECT 44.15 4.31 44.32 4.508 ;
      RECT 44.15 4.467 44.515 4.508 ;
      RECT 44.15 4.455 44.51 4.508 ;
      RECT 42.92 3.035 43.09 4.225 ;
      RECT 42.92 3.035 43.39 3.205 ;
      RECT 42.92 9.255 43.39 9.425 ;
      RECT 42.92 8.235 43.09 9.425 ;
      RECT 41.93 3.035 42.1 4.225 ;
      RECT 41.93 3.035 42.4 3.205 ;
      RECT 41.93 9.255 42.4 9.425 ;
      RECT 41.93 8.235 42.1 9.425 ;
      RECT 40.08 3.93 40.25 5.16 ;
      RECT 40.135 2.15 40.305 4.1 ;
      RECT 40.08 1.87 40.25 2.32 ;
      RECT 40.08 10.14 40.25 10.59 ;
      RECT 40.135 8.36 40.305 10.31 ;
      RECT 40.08 7.3 40.25 8.53 ;
      RECT 39.56 1.87 39.73 5.16 ;
      RECT 39.56 3.37 39.965 3.7 ;
      RECT 39.56 2.53 39.965 2.86 ;
      RECT 39.56 7.3 39.73 10.59 ;
      RECT 39.56 9.6 39.965 9.93 ;
      RECT 39.56 8.76 39.965 9.09 ;
      RECT 36.895 3.27 37.625 3.51 ;
      RECT 37.437 3.065 37.625 3.51 ;
      RECT 37.265 3.077 37.64 3.504 ;
      RECT 37.18 3.092 37.66 3.489 ;
      RECT 37.18 3.107 37.665 3.479 ;
      RECT 37.135 3.127 37.68 3.471 ;
      RECT 37.112 3.162 37.695 3.425 ;
      RECT 37.026 3.185 37.7 3.385 ;
      RECT 37.026 3.203 37.71 3.355 ;
      RECT 36.895 3.272 37.715 3.318 ;
      RECT 36.94 3.215 37.71 3.355 ;
      RECT 37.026 3.167 37.695 3.425 ;
      RECT 37.112 3.136 37.68 3.471 ;
      RECT 37.135 3.117 37.665 3.479 ;
      RECT 37.18 3.09 37.64 3.504 ;
      RECT 37.265 3.072 37.625 3.51 ;
      RECT 37.351 3.066 37.625 3.51 ;
      RECT 37.437 3.061 37.57 3.51 ;
      RECT 37.523 3.056 37.57 3.51 ;
      RECT 37.215 3.954 37.385 4.34 ;
      RECT 37.21 3.954 37.385 4.335 ;
      RECT 37.185 3.954 37.385 4.3 ;
      RECT 37.185 3.982 37.395 4.29 ;
      RECT 37.165 3.982 37.395 4.25 ;
      RECT 37.16 3.982 37.395 4.223 ;
      RECT 37.16 4 37.4 4.215 ;
      RECT 37.105 4 37.4 4.15 ;
      RECT 37.105 4.017 37.41 4.133 ;
      RECT 37.095 4.017 37.41 4.073 ;
      RECT 37.095 4.034 37.415 4.07 ;
      RECT 37.09 3.87 37.26 4.048 ;
      RECT 37.09 3.904 37.346 4.048 ;
      RECT 37.085 4.67 37.09 4.683 ;
      RECT 37.08 4.565 37.085 4.688 ;
      RECT 37.055 4.425 37.08 4.703 ;
      RECT 37.02 4.376 37.055 4.735 ;
      RECT 37.015 4.344 37.02 4.755 ;
      RECT 37.01 4.335 37.015 4.755 ;
      RECT 36.93 4.3 37.01 4.755 ;
      RECT 36.867 4.27 36.93 4.755 ;
      RECT 36.781 4.258 36.867 4.755 ;
      RECT 36.695 4.244 36.781 4.755 ;
      RECT 36.615 4.231 36.695 4.741 ;
      RECT 36.58 4.223 36.615 4.721 ;
      RECT 36.57 4.22 36.58 4.712 ;
      RECT 36.54 4.215 36.57 4.699 ;
      RECT 36.49 4.19 36.54 4.675 ;
      RECT 36.476 4.164 36.49 4.657 ;
      RECT 36.39 4.124 36.476 4.633 ;
      RECT 36.345 4.072 36.39 4.602 ;
      RECT 36.335 4.047 36.345 4.589 ;
      RECT 36.33 3.828 36.335 3.85 ;
      RECT 36.325 4.03 36.335 4.585 ;
      RECT 36.325 3.826 36.33 3.94 ;
      RECT 36.315 3.822 36.325 4.581 ;
      RECT 36.271 3.82 36.315 4.569 ;
      RECT 36.185 3.82 36.271 4.54 ;
      RECT 36.155 3.82 36.185 4.513 ;
      RECT 36.14 3.82 36.155 4.501 ;
      RECT 36.1 3.832 36.14 4.486 ;
      RECT 36.08 3.851 36.1 4.465 ;
      RECT 36.07 3.861 36.08 4.449 ;
      RECT 36.06 3.867 36.07 4.438 ;
      RECT 36.04 3.877 36.06 4.421 ;
      RECT 36.035 3.886 36.04 4.408 ;
      RECT 36.03 3.89 36.035 4.358 ;
      RECT 36.02 3.896 36.03 4.275 ;
      RECT 36.015 3.9 36.02 4.189 ;
      RECT 36.01 3.92 36.015 4.126 ;
      RECT 36.005 3.943 36.01 4.073 ;
      RECT 36 3.961 36.005 4.018 ;
      RECT 36.61 3.78 36.78 4.04 ;
      RECT 36.78 3.745 36.825 4.026 ;
      RECT 36.741 3.747 36.83 4.009 ;
      RECT 36.63 3.764 36.916 3.98 ;
      RECT 36.63 3.779 36.92 3.952 ;
      RECT 36.63 3.76 36.83 4.009 ;
      RECT 36.655 3.748 36.78 4.04 ;
      RECT 36.741 3.746 36.825 4.026 ;
      RECT 35.795 3.135 35.965 3.625 ;
      RECT 35.795 3.135 36 3.605 ;
      RECT 35.93 3.055 36.04 3.565 ;
      RECT 35.911 3.059 36.06 3.535 ;
      RECT 35.825 3.067 36.08 3.518 ;
      RECT 35.825 3.073 36.085 3.508 ;
      RECT 35.825 3.082 36.105 3.496 ;
      RECT 35.8 3.107 36.135 3.474 ;
      RECT 35.8 3.127 36.14 3.454 ;
      RECT 35.795 3.14 36.15 3.434 ;
      RECT 35.795 3.207 36.155 3.415 ;
      RECT 35.795 3.34 36.16 3.402 ;
      RECT 35.79 3.145 36.15 3.235 ;
      RECT 35.8 3.102 36.105 3.496 ;
      RECT 35.911 3.057 36.04 3.565 ;
      RECT 35.785 4.81 36.085 5.065 ;
      RECT 35.87 4.776 36.085 5.065 ;
      RECT 35.87 4.779 36.09 4.925 ;
      RECT 35.805 4.8 36.09 4.925 ;
      RECT 35.84 4.79 36.085 5.065 ;
      RECT 35.835 4.795 36.09 4.925 ;
      RECT 35.87 4.774 36.071 5.065 ;
      RECT 35.956 4.765 36.071 5.065 ;
      RECT 35.956 4.759 35.985 5.065 ;
      RECT 35.445 4.4 35.455 4.89 ;
      RECT 35.105 4.335 35.115 4.635 ;
      RECT 35.62 4.507 35.625 4.726 ;
      RECT 35.61 4.487 35.62 4.743 ;
      RECT 35.6 4.467 35.61 4.773 ;
      RECT 35.595 4.457 35.6 4.788 ;
      RECT 35.59 4.453 35.595 4.793 ;
      RECT 35.575 4.445 35.59 4.8 ;
      RECT 35.535 4.425 35.575 4.825 ;
      RECT 35.51 4.407 35.535 4.858 ;
      RECT 35.505 4.405 35.51 4.871 ;
      RECT 35.485 4.402 35.505 4.875 ;
      RECT 35.455 4.4 35.485 4.885 ;
      RECT 35.385 4.402 35.445 4.886 ;
      RECT 35.365 4.402 35.385 4.88 ;
      RECT 35.34 4.4 35.365 4.877 ;
      RECT 35.305 4.395 35.34 4.873 ;
      RECT 35.285 4.389 35.305 4.86 ;
      RECT 35.275 4.386 35.285 4.848 ;
      RECT 35.255 4.383 35.275 4.833 ;
      RECT 35.235 4.379 35.255 4.815 ;
      RECT 35.23 4.376 35.235 4.805 ;
      RECT 35.225 4.375 35.23 4.803 ;
      RECT 35.215 4.372 35.225 4.795 ;
      RECT 35.205 4.366 35.215 4.778 ;
      RECT 35.195 4.36 35.205 4.76 ;
      RECT 35.185 4.354 35.195 4.748 ;
      RECT 35.175 4.348 35.185 4.728 ;
      RECT 35.17 4.344 35.175 4.713 ;
      RECT 35.165 4.342 35.17 4.705 ;
      RECT 35.16 4.34 35.165 4.698 ;
      RECT 35.155 4.338 35.16 4.688 ;
      RECT 35.15 4.336 35.155 4.682 ;
      RECT 35.14 4.335 35.15 4.672 ;
      RECT 35.13 4.335 35.14 4.663 ;
      RECT 35.115 4.335 35.13 4.648 ;
      RECT 35.075 4.335 35.105 4.632 ;
      RECT 35.055 4.337 35.075 4.627 ;
      RECT 35.05 4.342 35.055 4.625 ;
      RECT 35.02 4.35 35.05 4.623 ;
      RECT 34.99 4.365 35.02 4.622 ;
      RECT 34.945 4.387 34.99 4.627 ;
      RECT 34.94 4.402 34.945 4.631 ;
      RECT 34.925 4.407 34.94 4.633 ;
      RECT 34.92 4.411 34.925 4.635 ;
      RECT 34.86 4.434 34.92 4.644 ;
      RECT 34.84 4.46 34.86 4.657 ;
      RECT 34.83 4.467 34.84 4.661 ;
      RECT 34.815 4.474 34.83 4.664 ;
      RECT 34.795 4.484 34.815 4.667 ;
      RECT 34.79 4.492 34.795 4.67 ;
      RECT 34.745 4.497 34.79 4.677 ;
      RECT 34.735 4.5 34.745 4.684 ;
      RECT 34.725 4.5 34.735 4.688 ;
      RECT 34.69 4.502 34.725 4.7 ;
      RECT 34.67 4.505 34.69 4.713 ;
      RECT 34.63 4.508 34.67 4.724 ;
      RECT 34.615 4.51 34.63 4.737 ;
      RECT 34.605 4.51 34.615 4.742 ;
      RECT 34.58 4.511 34.605 4.75 ;
      RECT 34.57 4.513 34.58 4.755 ;
      RECT 34.565 4.514 34.57 4.758 ;
      RECT 34.54 4.512 34.565 4.761 ;
      RECT 34.525 4.51 34.54 4.762 ;
      RECT 34.505 4.507 34.525 4.764 ;
      RECT 34.485 4.502 34.505 4.764 ;
      RECT 34.425 4.497 34.485 4.761 ;
      RECT 34.39 4.472 34.425 4.757 ;
      RECT 34.38 4.449 34.39 4.755 ;
      RECT 34.35 4.426 34.38 4.755 ;
      RECT 34.34 4.405 34.35 4.755 ;
      RECT 34.315 4.387 34.34 4.753 ;
      RECT 34.3 4.365 34.315 4.75 ;
      RECT 34.285 4.347 34.3 4.748 ;
      RECT 34.265 4.337 34.285 4.746 ;
      RECT 34.25 4.332 34.265 4.745 ;
      RECT 34.235 4.33 34.25 4.744 ;
      RECT 34.205 4.331 34.235 4.742 ;
      RECT 34.185 4.334 34.205 4.74 ;
      RECT 34.128 4.338 34.185 4.74 ;
      RECT 34.042 4.347 34.128 4.74 ;
      RECT 33.956 4.358 34.042 4.74 ;
      RECT 33.87 4.369 33.956 4.74 ;
      RECT 33.85 4.376 33.87 4.748 ;
      RECT 33.84 4.379 33.85 4.755 ;
      RECT 33.775 4.384 33.84 4.773 ;
      RECT 33.745 4.391 33.775 4.798 ;
      RECT 33.735 4.394 33.745 4.805 ;
      RECT 33.69 4.398 33.735 4.81 ;
      RECT 33.66 4.403 33.69 4.815 ;
      RECT 33.659 4.405 33.66 4.815 ;
      RECT 33.573 4.411 33.659 4.815 ;
      RECT 33.487 4.422 33.573 4.815 ;
      RECT 33.401 4.434 33.487 4.815 ;
      RECT 33.315 4.445 33.401 4.815 ;
      RECT 33.3 4.452 33.315 4.81 ;
      RECT 33.295 4.454 33.3 4.804 ;
      RECT 33.275 4.465 33.295 4.799 ;
      RECT 33.265 4.483 33.275 4.793 ;
      RECT 33.26 4.495 33.265 4.593 ;
      RECT 35.555 3.248 35.575 3.335 ;
      RECT 35.55 3.183 35.555 3.367 ;
      RECT 35.54 3.15 35.55 3.372 ;
      RECT 35.535 3.13 35.54 3.378 ;
      RECT 35.505 3.13 35.535 3.395 ;
      RECT 35.456 3.13 35.505 3.431 ;
      RECT 35.37 3.13 35.456 3.489 ;
      RECT 35.341 3.14 35.37 3.538 ;
      RECT 35.255 3.182 35.341 3.591 ;
      RECT 35.235 3.22 35.255 3.638 ;
      RECT 35.21 3.237 35.235 3.658 ;
      RECT 35.2 3.251 35.21 3.678 ;
      RECT 35.195 3.257 35.2 3.688 ;
      RECT 35.19 3.261 35.195 3.695 ;
      RECT 35.14 3.281 35.19 3.7 ;
      RECT 35.075 3.325 35.14 3.7 ;
      RECT 35.05 3.375 35.075 3.7 ;
      RECT 35.04 3.405 35.05 3.7 ;
      RECT 35.035 3.432 35.04 3.7 ;
      RECT 35.03 3.45 35.035 3.7 ;
      RECT 35.02 3.492 35.03 3.7 ;
      RECT 35.37 4.05 35.54 4.225 ;
      RECT 35.31 3.878 35.37 4.213 ;
      RECT 35.3 3.871 35.31 4.196 ;
      RECT 35.255 4.05 35.54 4.176 ;
      RECT 35.236 4.05 35.54 4.154 ;
      RECT 35.15 4.05 35.54 4.119 ;
      RECT 35.13 3.87 35.3 4.075 ;
      RECT 35.13 4.017 35.535 4.075 ;
      RECT 35.13 3.965 35.51 4.075 ;
      RECT 35.13 3.92 35.475 4.075 ;
      RECT 35.13 3.902 35.44 4.075 ;
      RECT 35.13 3.892 35.435 4.075 ;
      RECT 35.3 10.14 35.47 10.59 ;
      RECT 35.355 8.36 35.525 10.31 ;
      RECT 35.3 7.3 35.47 8.53 ;
      RECT 34.78 7.3 34.95 10.59 ;
      RECT 34.78 9.6 35.185 9.93 ;
      RECT 34.78 8.76 35.185 9.09 ;
      RECT 34.85 4.85 35.04 5.075 ;
      RECT 34.84 4.851 35.045 5.07 ;
      RECT 34.84 4.853 35.055 5.05 ;
      RECT 34.84 4.857 35.06 5.035 ;
      RECT 34.84 4.844 35.01 5.07 ;
      RECT 34.84 4.847 35.035 5.07 ;
      RECT 34.85 4.843 35.01 5.075 ;
      RECT 34.936 4.841 35.01 5.075 ;
      RECT 34.56 4.092 34.73 4.33 ;
      RECT 34.56 4.092 34.816 4.244 ;
      RECT 34.56 4.092 34.82 4.154 ;
      RECT 34.61 3.865 34.83 4.133 ;
      RECT 34.605 3.882 34.835 4.106 ;
      RECT 34.57 4.04 34.835 4.106 ;
      RECT 34.59 3.89 34.73 4.33 ;
      RECT 34.58 3.972 34.84 4.089 ;
      RECT 34.575 4.02 34.84 4.089 ;
      RECT 34.58 3.93 34.835 4.106 ;
      RECT 34.605 3.867 34.83 4.133 ;
      RECT 34.17 3.842 34.34 4.04 ;
      RECT 34.17 3.842 34.385 4.015 ;
      RECT 34.24 3.785 34.41 3.973 ;
      RECT 34.215 3.8 34.41 3.973 ;
      RECT 33.83 3.846 33.86 4.04 ;
      RECT 33.825 3.818 33.83 4.04 ;
      RECT 33.795 3.792 33.825 4.042 ;
      RECT 33.77 3.75 33.795 4.045 ;
      RECT 33.76 3.722 33.77 4.047 ;
      RECT 33.725 3.702 33.76 4.049 ;
      RECT 33.66 3.687 33.725 4.055 ;
      RECT 33.61 3.685 33.66 4.061 ;
      RECT 33.587 3.687 33.61 4.066 ;
      RECT 33.501 3.698 33.587 4.072 ;
      RECT 33.415 3.716 33.501 4.082 ;
      RECT 33.4 3.727 33.415 4.088 ;
      RECT 33.33 3.75 33.4 4.094 ;
      RECT 33.275 3.782 33.33 4.102 ;
      RECT 33.235 3.805 33.275 4.108 ;
      RECT 33.221 3.818 33.235 4.111 ;
      RECT 33.135 3.84 33.221 4.117 ;
      RECT 33.12 3.865 33.135 4.123 ;
      RECT 33.08 3.88 33.12 4.127 ;
      RECT 33.03 3.895 33.08 4.132 ;
      RECT 33.005 3.902 33.03 4.136 ;
      RECT 32.945 3.897 33.005 4.14 ;
      RECT 32.93 3.888 32.945 4.144 ;
      RECT 32.86 3.878 32.93 4.14 ;
      RECT 32.835 3.87 32.855 4.13 ;
      RECT 32.776 3.87 32.835 4.108 ;
      RECT 32.69 3.87 32.776 4.065 ;
      RECT 32.855 3.87 32.86 4.135 ;
      RECT 33.55 3.101 33.72 3.435 ;
      RECT 33.52 3.101 33.72 3.43 ;
      RECT 33.46 3.068 33.52 3.418 ;
      RECT 33.46 3.124 33.73 3.413 ;
      RECT 33.435 3.124 33.73 3.407 ;
      RECT 33.43 3.065 33.46 3.404 ;
      RECT 33.415 3.071 33.55 3.402 ;
      RECT 33.41 3.079 33.635 3.39 ;
      RECT 33.41 3.131 33.745 3.343 ;
      RECT 33.395 3.087 33.635 3.338 ;
      RECT 33.395 3.157 33.755 3.279 ;
      RECT 33.365 3.107 33.72 3.24 ;
      RECT 33.365 3.197 33.765 3.236 ;
      RECT 33.415 3.076 33.635 3.402 ;
      RECT 32.755 3.406 32.81 3.67 ;
      RECT 32.755 3.406 32.875 3.669 ;
      RECT 32.755 3.406 32.9 3.668 ;
      RECT 32.755 3.406 32.965 3.667 ;
      RECT 32.9 3.372 32.98 3.666 ;
      RECT 32.715 3.416 33.125 3.665 ;
      RECT 32.755 3.413 33.125 3.665 ;
      RECT 32.715 3.421 33.13 3.658 ;
      RECT 32.7 3.423 33.13 3.657 ;
      RECT 32.7 3.43 33.135 3.653 ;
      RECT 32.68 3.429 33.13 3.649 ;
      RECT 32.68 3.437 33.14 3.648 ;
      RECT 32.675 3.434 33.135 3.644 ;
      RECT 32.675 3.447 33.15 3.643 ;
      RECT 32.66 3.437 33.14 3.642 ;
      RECT 32.625 3.45 33.15 3.635 ;
      RECT 32.81 3.405 33.12 3.665 ;
      RECT 32.81 3.39 33.07 3.665 ;
      RECT 32.875 3.377 33.005 3.665 ;
      RECT 32.42 4.466 32.435 4.859 ;
      RECT 32.385 4.471 32.435 4.858 ;
      RECT 32.42 4.47 32.48 4.857 ;
      RECT 32.365 4.481 32.48 4.856 ;
      RECT 32.38 4.477 32.48 4.856 ;
      RECT 32.345 4.487 32.555 4.853 ;
      RECT 32.345 4.506 32.6 4.851 ;
      RECT 32.345 4.513 32.605 4.848 ;
      RECT 32.33 4.49 32.555 4.845 ;
      RECT 32.31 4.495 32.555 4.838 ;
      RECT 32.305 4.499 32.555 4.834 ;
      RECT 32.305 4.516 32.615 4.833 ;
      RECT 32.285 4.51 32.6 4.829 ;
      RECT 32.285 4.519 32.62 4.823 ;
      RECT 32.28 4.525 32.62 4.595 ;
      RECT 32.345 4.485 32.48 4.853 ;
      RECT 32.22 3.848 32.42 4.16 ;
      RECT 32.295 3.826 32.42 4.16 ;
      RECT 32.235 3.845 32.425 4.145 ;
      RECT 32.205 3.856 32.425 4.143 ;
      RECT 32.22 3.851 32.43 4.109 ;
      RECT 32.205 3.955 32.435 4.076 ;
      RECT 32.235 3.827 32.42 4.16 ;
      RECT 32.295 3.805 32.395 4.16 ;
      RECT 32.32 3.802 32.395 4.16 ;
      RECT 32.32 3.797 32.34 4.16 ;
      RECT 31.725 3.865 31.9 4.04 ;
      RECT 31.72 3.865 31.9 4.038 ;
      RECT 31.695 3.865 31.9 4.033 ;
      RECT 31.64 3.845 31.81 4.023 ;
      RECT 31.64 3.852 31.875 4.023 ;
      RECT 31.725 4.532 31.74 4.715 ;
      RECT 31.715 4.51 31.725 4.715 ;
      RECT 31.7 4.49 31.715 4.715 ;
      RECT 31.69 4.465 31.7 4.715 ;
      RECT 31.66 4.43 31.69 4.715 ;
      RECT 31.625 4.37 31.66 4.715 ;
      RECT 31.62 4.332 31.625 4.715 ;
      RECT 31.57 4.283 31.62 4.715 ;
      RECT 31.56 4.233 31.57 4.703 ;
      RECT 31.545 4.212 31.56 4.663 ;
      RECT 31.525 4.18 31.545 4.613 ;
      RECT 31.5 4.136 31.525 4.553 ;
      RECT 31.495 4.108 31.5 4.508 ;
      RECT 31.49 4.099 31.495 4.494 ;
      RECT 31.485 4.092 31.49 4.481 ;
      RECT 31.48 4.087 31.485 4.47 ;
      RECT 31.475 4.072 31.48 4.46 ;
      RECT 31.47 4.05 31.475 4.447 ;
      RECT 31.46 4.01 31.47 4.422 ;
      RECT 31.435 3.94 31.46 4.378 ;
      RECT 31.43 3.88 31.435 4.343 ;
      RECT 31.415 3.86 31.43 4.31 ;
      RECT 31.41 3.86 31.415 4.285 ;
      RECT 31.38 3.86 31.41 4.24 ;
      RECT 31.335 3.86 31.38 4.18 ;
      RECT 31.26 3.86 31.335 4.128 ;
      RECT 31.255 3.86 31.26 4.093 ;
      RECT 31.25 3.86 31.255 4.083 ;
      RECT 31.245 3.86 31.25 4.063 ;
      RECT 31.51 3.08 31.68 3.55 ;
      RECT 31.455 3.073 31.65 3.534 ;
      RECT 31.455 3.087 31.685 3.533 ;
      RECT 31.44 3.088 31.685 3.514 ;
      RECT 31.435 3.106 31.685 3.5 ;
      RECT 31.44 3.089 31.69 3.498 ;
      RECT 31.425 3.12 31.69 3.483 ;
      RECT 31.44 3.095 31.695 3.468 ;
      RECT 31.42 3.135 31.695 3.465 ;
      RECT 31.435 3.107 31.7 3.45 ;
      RECT 31.435 3.119 31.705 3.43 ;
      RECT 31.42 3.135 31.71 3.413 ;
      RECT 31.42 3.145 31.715 3.268 ;
      RECT 31.415 3.145 31.715 3.225 ;
      RECT 31.415 3.16 31.72 3.203 ;
      RECT 31.51 3.07 31.65 3.55 ;
      RECT 31.51 3.068 31.62 3.55 ;
      RECT 31.596 3.065 31.62 3.55 ;
      RECT 31.255 4.732 31.26 4.778 ;
      RECT 31.245 4.58 31.255 4.802 ;
      RECT 31.24 4.425 31.245 4.827 ;
      RECT 31.225 4.387 31.24 4.838 ;
      RECT 31.22 4.37 31.225 4.845 ;
      RECT 31.21 4.358 31.22 4.852 ;
      RECT 31.205 4.349 31.21 4.854 ;
      RECT 31.2 4.347 31.205 4.858 ;
      RECT 31.155 4.338 31.2 4.873 ;
      RECT 31.15 4.33 31.155 4.887 ;
      RECT 31.145 4.327 31.15 4.891 ;
      RECT 31.13 4.322 31.145 4.899 ;
      RECT 31.075 4.312 31.13 4.91 ;
      RECT 31.04 4.3 31.075 4.911 ;
      RECT 31.031 4.295 31.04 4.905 ;
      RECT 30.945 4.295 31.031 4.895 ;
      RECT 30.915 4.295 30.945 4.873 ;
      RECT 30.905 4.295 30.91 4.853 ;
      RECT 30.9 4.295 30.905 4.815 ;
      RECT 30.895 4.295 30.9 4.773 ;
      RECT 30.89 4.295 30.895 4.733 ;
      RECT 30.885 4.295 30.89 4.663 ;
      RECT 30.875 4.295 30.885 4.585 ;
      RECT 30.87 4.295 30.875 4.485 ;
      RECT 30.91 4.295 30.915 4.855 ;
      RECT 30.405 4.377 30.495 4.855 ;
      RECT 30.39 4.38 30.51 4.853 ;
      RECT 30.405 4.379 30.51 4.853 ;
      RECT 30.37 4.386 30.535 4.843 ;
      RECT 30.39 4.38 30.535 4.843 ;
      RECT 30.355 4.392 30.535 4.831 ;
      RECT 30.39 4.383 30.585 4.824 ;
      RECT 30.341 4.4 30.585 4.822 ;
      RECT 30.37 4.39 30.595 4.81 ;
      RECT 30.341 4.411 30.625 4.801 ;
      RECT 30.255 4.435 30.625 4.795 ;
      RECT 30.255 4.448 30.665 4.778 ;
      RECT 30.25 4.47 30.665 4.771 ;
      RECT 30.22 4.485 30.665 4.761 ;
      RECT 30.215 4.496 30.665 4.751 ;
      RECT 30.185 4.509 30.665 4.742 ;
      RECT 30.17 4.527 30.665 4.731 ;
      RECT 30.145 4.54 30.665 4.721 ;
      RECT 30.405 4.376 30.415 4.855 ;
      RECT 30.451 3.8 30.49 4.045 ;
      RECT 30.365 3.8 30.5 4.043 ;
      RECT 30.25 3.825 30.5 4.04 ;
      RECT 30.25 3.825 30.505 4.038 ;
      RECT 30.25 3.825 30.52 4.033 ;
      RECT 30.356 3.8 30.535 4.013 ;
      RECT 30.27 3.808 30.535 4.013 ;
      RECT 29.94 3.16 30.11 3.595 ;
      RECT 29.93 3.194 30.11 3.578 ;
      RECT 30.01 3.13 30.18 3.565 ;
      RECT 29.915 3.205 30.18 3.543 ;
      RECT 30.01 3.14 30.185 3.533 ;
      RECT 29.94 3.192 30.215 3.518 ;
      RECT 29.9 3.218 30.215 3.503 ;
      RECT 29.9 3.26 30.225 3.483 ;
      RECT 29.895 3.285 30.23 3.465 ;
      RECT 29.895 3.295 30.235 3.45 ;
      RECT 29.89 3.232 30.215 3.448 ;
      RECT 29.89 3.305 30.24 3.433 ;
      RECT 29.885 3.242 30.215 3.43 ;
      RECT 29.88 3.326 30.245 3.413 ;
      RECT 29.88 3.358 30.25 3.393 ;
      RECT 29.875 3.272 30.225 3.385 ;
      RECT 29.88 3.257 30.215 3.413 ;
      RECT 29.895 3.227 30.215 3.465 ;
      RECT 29.74 3.814 29.965 4.07 ;
      RECT 29.74 3.847 29.985 4.06 ;
      RECT 29.705 3.847 29.985 4.058 ;
      RECT 29.705 3.86 29.99 4.048 ;
      RECT 29.705 3.88 30 4.04 ;
      RECT 29.705 3.977 30.005 4.033 ;
      RECT 29.685 3.725 29.815 4.023 ;
      RECT 29.64 3.88 30 3.965 ;
      RECT 29.63 3.725 29.815 3.91 ;
      RECT 29.63 3.757 29.901 3.91 ;
      RECT 29.595 4.287 29.615 4.465 ;
      RECT 29.56 4.24 29.595 4.465 ;
      RECT 29.545 4.18 29.56 4.465 ;
      RECT 29.52 4.127 29.545 4.465 ;
      RECT 29.505 4.08 29.52 4.465 ;
      RECT 29.485 4.057 29.505 4.465 ;
      RECT 29.46 4.022 29.485 4.465 ;
      RECT 29.45 3.868 29.46 4.465 ;
      RECT 29.42 3.863 29.45 4.456 ;
      RECT 29.415 3.86 29.42 4.446 ;
      RECT 29.4 3.86 29.415 4.42 ;
      RECT 29.395 3.86 29.4 4.383 ;
      RECT 29.37 3.86 29.395 4.335 ;
      RECT 29.35 3.86 29.37 4.26 ;
      RECT 29.34 3.86 29.35 4.22 ;
      RECT 29.335 3.86 29.34 4.195 ;
      RECT 29.33 3.86 29.335 4.178 ;
      RECT 29.325 3.86 29.33 4.16 ;
      RECT 29.32 3.861 29.325 4.15 ;
      RECT 29.31 3.863 29.32 4.118 ;
      RECT 29.3 3.865 29.31 4.085 ;
      RECT 29.29 3.868 29.3 4.058 ;
      RECT 29.615 4.295 29.84 4.465 ;
      RECT 28.945 3.107 29.115 3.56 ;
      RECT 28.945 3.107 29.205 3.526 ;
      RECT 28.945 3.107 29.235 3.51 ;
      RECT 28.945 3.107 29.265 3.483 ;
      RECT 29.201 3.085 29.28 3.465 ;
      RECT 28.98 3.092 29.285 3.45 ;
      RECT 28.98 3.1 29.295 3.413 ;
      RECT 28.94 3.127 29.295 3.385 ;
      RECT 28.925 3.14 29.295 3.35 ;
      RECT 28.945 3.115 29.315 3.34 ;
      RECT 28.92 3.18 29.315 3.31 ;
      RECT 28.92 3.21 29.32 3.293 ;
      RECT 28.915 3.24 29.32 3.28 ;
      RECT 28.98 3.089 29.28 3.465 ;
      RECT 29.115 3.086 29.201 3.544 ;
      RECT 29.066 3.087 29.28 3.465 ;
      RECT 29.21 4.747 29.255 4.94 ;
      RECT 29.2 4.717 29.21 4.94 ;
      RECT 29.195 4.702 29.2 4.94 ;
      RECT 29.155 4.612 29.195 4.94 ;
      RECT 29.15 4.525 29.155 4.94 ;
      RECT 29.14 4.495 29.15 4.94 ;
      RECT 29.135 4.455 29.14 4.94 ;
      RECT 29.125 4.417 29.135 4.94 ;
      RECT 29.12 4.382 29.125 4.94 ;
      RECT 29.1 4.335 29.12 4.94 ;
      RECT 29.085 4.26 29.1 4.94 ;
      RECT 29.08 4.215 29.085 4.935 ;
      RECT 29.075 4.195 29.08 4.908 ;
      RECT 29.07 4.175 29.075 4.893 ;
      RECT 29.065 4.15 29.07 4.873 ;
      RECT 29.06 4.128 29.065 4.858 ;
      RECT 29.055 4.106 29.06 4.84 ;
      RECT 29.05 4.085 29.055 4.83 ;
      RECT 29.04 4.057 29.05 4.8 ;
      RECT 29.03 4.02 29.04 4.768 ;
      RECT 29.02 3.98 29.03 4.735 ;
      RECT 29.01 3.958 29.02 4.705 ;
      RECT 28.98 3.91 29.01 4.637 ;
      RECT 28.965 3.87 28.98 4.564 ;
      RECT 28.955 3.87 28.965 4.53 ;
      RECT 28.95 3.87 28.955 4.505 ;
      RECT 28.945 3.87 28.95 4.49 ;
      RECT 28.94 3.87 28.945 4.468 ;
      RECT 28.935 3.87 28.94 4.455 ;
      RECT 28.92 3.87 28.935 4.42 ;
      RECT 28.9 3.87 28.92 4.36 ;
      RECT 28.89 3.87 28.9 4.31 ;
      RECT 28.87 3.87 28.89 4.258 ;
      RECT 28.85 3.87 28.87 4.215 ;
      RECT 28.84 3.87 28.85 4.203 ;
      RECT 28.81 3.87 28.84 4.19 ;
      RECT 28.78 3.891 28.81 4.17 ;
      RECT 28.77 3.919 28.78 4.15 ;
      RECT 28.755 3.936 28.77 4.118 ;
      RECT 28.75 3.95 28.755 4.085 ;
      RECT 28.745 3.958 28.75 4.058 ;
      RECT 28.74 3.966 28.745 4.02 ;
      RECT 28.745 4.49 28.75 4.825 ;
      RECT 28.71 4.477 28.745 4.824 ;
      RECT 28.64 4.417 28.71 4.823 ;
      RECT 28.56 4.36 28.64 4.822 ;
      RECT 28.425 4.32 28.56 4.821 ;
      RECT 28.425 4.507 28.76 4.81 ;
      RECT 28.385 4.507 28.76 4.8 ;
      RECT 28.385 4.525 28.765 4.795 ;
      RECT 28.385 4.615 28.77 4.785 ;
      RECT 28.38 4.31 28.545 4.765 ;
      RECT 28.375 4.31 28.545 4.508 ;
      RECT 28.375 4.467 28.74 4.508 ;
      RECT 28.375 4.455 28.735 4.508 ;
      RECT 27.14 3.035 27.31 4.225 ;
      RECT 27.14 3.035 27.61 3.205 ;
      RECT 27.14 9.255 27.61 9.425 ;
      RECT 27.14 8.235 27.31 9.425 ;
      RECT 26.15 3.035 26.32 4.225 ;
      RECT 26.15 3.035 26.62 3.205 ;
      RECT 26.15 9.255 26.62 9.425 ;
      RECT 26.15 8.235 26.32 9.425 ;
      RECT 24.3 3.93 24.47 5.16 ;
      RECT 24.355 2.15 24.525 4.1 ;
      RECT 24.3 1.87 24.47 2.32 ;
      RECT 24.3 10.14 24.47 10.59 ;
      RECT 24.355 8.36 24.525 10.31 ;
      RECT 24.3 7.3 24.47 8.53 ;
      RECT 23.78 1.87 23.95 5.16 ;
      RECT 23.78 3.37 24.185 3.7 ;
      RECT 23.78 2.53 24.185 2.86 ;
      RECT 23.78 7.3 23.95 10.59 ;
      RECT 23.78 9.6 24.185 9.93 ;
      RECT 23.78 8.76 24.185 9.09 ;
      RECT 21.115 3.27 21.845 3.51 ;
      RECT 21.657 3.065 21.845 3.51 ;
      RECT 21.485 3.077 21.86 3.504 ;
      RECT 21.4 3.092 21.88 3.489 ;
      RECT 21.4 3.107 21.885 3.479 ;
      RECT 21.355 3.127 21.9 3.471 ;
      RECT 21.332 3.162 21.915 3.425 ;
      RECT 21.246 3.185 21.92 3.385 ;
      RECT 21.246 3.203 21.93 3.355 ;
      RECT 21.115 3.272 21.935 3.318 ;
      RECT 21.16 3.215 21.93 3.355 ;
      RECT 21.246 3.167 21.915 3.425 ;
      RECT 21.332 3.136 21.9 3.471 ;
      RECT 21.355 3.117 21.885 3.479 ;
      RECT 21.4 3.09 21.86 3.504 ;
      RECT 21.485 3.072 21.845 3.51 ;
      RECT 21.571 3.066 21.845 3.51 ;
      RECT 21.657 3.061 21.79 3.51 ;
      RECT 21.743 3.056 21.79 3.51 ;
      RECT 21.435 3.954 21.605 4.34 ;
      RECT 21.43 3.954 21.605 4.335 ;
      RECT 21.405 3.954 21.605 4.3 ;
      RECT 21.405 3.982 21.615 4.29 ;
      RECT 21.385 3.982 21.615 4.25 ;
      RECT 21.38 3.982 21.615 4.223 ;
      RECT 21.38 4 21.62 4.215 ;
      RECT 21.325 4 21.62 4.15 ;
      RECT 21.325 4.017 21.63 4.133 ;
      RECT 21.315 4.017 21.63 4.073 ;
      RECT 21.315 4.034 21.635 4.07 ;
      RECT 21.31 3.87 21.48 4.048 ;
      RECT 21.31 3.904 21.566 4.048 ;
      RECT 21.305 4.67 21.31 4.683 ;
      RECT 21.3 4.565 21.305 4.688 ;
      RECT 21.275 4.425 21.3 4.703 ;
      RECT 21.24 4.376 21.275 4.735 ;
      RECT 21.235 4.344 21.24 4.755 ;
      RECT 21.23 4.335 21.235 4.755 ;
      RECT 21.15 4.3 21.23 4.755 ;
      RECT 21.087 4.27 21.15 4.755 ;
      RECT 21.001 4.258 21.087 4.755 ;
      RECT 20.915 4.244 21.001 4.755 ;
      RECT 20.835 4.231 20.915 4.741 ;
      RECT 20.8 4.223 20.835 4.721 ;
      RECT 20.79 4.22 20.8 4.712 ;
      RECT 20.76 4.215 20.79 4.699 ;
      RECT 20.71 4.19 20.76 4.675 ;
      RECT 20.696 4.164 20.71 4.657 ;
      RECT 20.61 4.124 20.696 4.633 ;
      RECT 20.565 4.072 20.61 4.602 ;
      RECT 20.555 4.047 20.565 4.589 ;
      RECT 20.55 3.828 20.555 3.85 ;
      RECT 20.545 4.03 20.555 4.585 ;
      RECT 20.545 3.826 20.55 3.94 ;
      RECT 20.535 3.822 20.545 4.581 ;
      RECT 20.491 3.82 20.535 4.569 ;
      RECT 20.405 3.82 20.491 4.54 ;
      RECT 20.375 3.82 20.405 4.513 ;
      RECT 20.36 3.82 20.375 4.501 ;
      RECT 20.32 3.832 20.36 4.486 ;
      RECT 20.3 3.851 20.32 4.465 ;
      RECT 20.29 3.861 20.3 4.449 ;
      RECT 20.28 3.867 20.29 4.438 ;
      RECT 20.26 3.877 20.28 4.421 ;
      RECT 20.255 3.886 20.26 4.408 ;
      RECT 20.25 3.89 20.255 4.358 ;
      RECT 20.24 3.896 20.25 4.275 ;
      RECT 20.235 3.9 20.24 4.189 ;
      RECT 20.23 3.92 20.235 4.126 ;
      RECT 20.225 3.943 20.23 4.073 ;
      RECT 20.22 3.961 20.225 4.018 ;
      RECT 20.83 3.78 21 4.04 ;
      RECT 21 3.745 21.045 4.026 ;
      RECT 20.961 3.747 21.05 4.009 ;
      RECT 20.85 3.764 21.136 3.98 ;
      RECT 20.85 3.779 21.14 3.952 ;
      RECT 20.85 3.76 21.05 4.009 ;
      RECT 20.875 3.748 21 4.04 ;
      RECT 20.961 3.746 21.045 4.026 ;
      RECT 20.015 3.135 20.185 3.625 ;
      RECT 20.015 3.135 20.22 3.605 ;
      RECT 20.15 3.055 20.26 3.565 ;
      RECT 20.131 3.059 20.28 3.535 ;
      RECT 20.045 3.067 20.3 3.518 ;
      RECT 20.045 3.073 20.305 3.508 ;
      RECT 20.045 3.082 20.325 3.496 ;
      RECT 20.02 3.107 20.355 3.474 ;
      RECT 20.02 3.127 20.36 3.454 ;
      RECT 20.015 3.14 20.37 3.434 ;
      RECT 20.015 3.207 20.375 3.415 ;
      RECT 20.015 3.34 20.38 3.402 ;
      RECT 20.01 3.145 20.37 3.235 ;
      RECT 20.02 3.102 20.325 3.496 ;
      RECT 20.131 3.057 20.26 3.565 ;
      RECT 20.005 4.81 20.305 5.065 ;
      RECT 20.09 4.776 20.305 5.065 ;
      RECT 20.09 4.779 20.31 4.925 ;
      RECT 20.025 4.8 20.31 4.925 ;
      RECT 20.06 4.79 20.305 5.065 ;
      RECT 20.055 4.795 20.31 4.925 ;
      RECT 20.09 4.774 20.291 5.065 ;
      RECT 20.176 4.765 20.291 5.065 ;
      RECT 20.176 4.759 20.205 5.065 ;
      RECT 19.665 4.4 19.675 4.89 ;
      RECT 19.325 4.335 19.335 4.635 ;
      RECT 19.84 4.507 19.845 4.726 ;
      RECT 19.83 4.487 19.84 4.743 ;
      RECT 19.82 4.467 19.83 4.773 ;
      RECT 19.815 4.457 19.82 4.788 ;
      RECT 19.81 4.453 19.815 4.793 ;
      RECT 19.795 4.445 19.81 4.8 ;
      RECT 19.755 4.425 19.795 4.825 ;
      RECT 19.73 4.407 19.755 4.858 ;
      RECT 19.725 4.405 19.73 4.871 ;
      RECT 19.705 4.402 19.725 4.875 ;
      RECT 19.675 4.4 19.705 4.885 ;
      RECT 19.605 4.402 19.665 4.886 ;
      RECT 19.585 4.402 19.605 4.88 ;
      RECT 19.56 4.4 19.585 4.877 ;
      RECT 19.525 4.395 19.56 4.873 ;
      RECT 19.505 4.389 19.525 4.86 ;
      RECT 19.495 4.386 19.505 4.848 ;
      RECT 19.475 4.383 19.495 4.833 ;
      RECT 19.455 4.379 19.475 4.815 ;
      RECT 19.45 4.376 19.455 4.805 ;
      RECT 19.445 4.375 19.45 4.803 ;
      RECT 19.435 4.372 19.445 4.795 ;
      RECT 19.425 4.366 19.435 4.778 ;
      RECT 19.415 4.36 19.425 4.76 ;
      RECT 19.405 4.354 19.415 4.748 ;
      RECT 19.395 4.348 19.405 4.728 ;
      RECT 19.39 4.344 19.395 4.713 ;
      RECT 19.385 4.342 19.39 4.705 ;
      RECT 19.38 4.34 19.385 4.698 ;
      RECT 19.375 4.338 19.38 4.688 ;
      RECT 19.37 4.336 19.375 4.682 ;
      RECT 19.36 4.335 19.37 4.672 ;
      RECT 19.35 4.335 19.36 4.663 ;
      RECT 19.335 4.335 19.35 4.648 ;
      RECT 19.295 4.335 19.325 4.632 ;
      RECT 19.275 4.337 19.295 4.627 ;
      RECT 19.27 4.342 19.275 4.625 ;
      RECT 19.24 4.35 19.27 4.623 ;
      RECT 19.21 4.365 19.24 4.622 ;
      RECT 19.165 4.387 19.21 4.627 ;
      RECT 19.16 4.402 19.165 4.631 ;
      RECT 19.145 4.407 19.16 4.633 ;
      RECT 19.14 4.411 19.145 4.635 ;
      RECT 19.08 4.434 19.14 4.644 ;
      RECT 19.06 4.46 19.08 4.657 ;
      RECT 19.05 4.467 19.06 4.661 ;
      RECT 19.035 4.474 19.05 4.664 ;
      RECT 19.015 4.484 19.035 4.667 ;
      RECT 19.01 4.492 19.015 4.67 ;
      RECT 18.965 4.497 19.01 4.677 ;
      RECT 18.955 4.5 18.965 4.684 ;
      RECT 18.945 4.5 18.955 4.688 ;
      RECT 18.91 4.502 18.945 4.7 ;
      RECT 18.89 4.505 18.91 4.713 ;
      RECT 18.85 4.508 18.89 4.724 ;
      RECT 18.835 4.51 18.85 4.737 ;
      RECT 18.825 4.51 18.835 4.742 ;
      RECT 18.8 4.511 18.825 4.75 ;
      RECT 18.79 4.513 18.8 4.755 ;
      RECT 18.785 4.514 18.79 4.758 ;
      RECT 18.76 4.512 18.785 4.761 ;
      RECT 18.745 4.51 18.76 4.762 ;
      RECT 18.725 4.507 18.745 4.764 ;
      RECT 18.705 4.502 18.725 4.764 ;
      RECT 18.645 4.497 18.705 4.761 ;
      RECT 18.61 4.472 18.645 4.757 ;
      RECT 18.6 4.449 18.61 4.755 ;
      RECT 18.57 4.426 18.6 4.755 ;
      RECT 18.56 4.405 18.57 4.755 ;
      RECT 18.535 4.387 18.56 4.753 ;
      RECT 18.52 4.365 18.535 4.75 ;
      RECT 18.505 4.347 18.52 4.748 ;
      RECT 18.485 4.337 18.505 4.746 ;
      RECT 18.47 4.332 18.485 4.745 ;
      RECT 18.455 4.33 18.47 4.744 ;
      RECT 18.425 4.331 18.455 4.742 ;
      RECT 18.405 4.334 18.425 4.74 ;
      RECT 18.348 4.338 18.405 4.74 ;
      RECT 18.262 4.347 18.348 4.74 ;
      RECT 18.176 4.358 18.262 4.74 ;
      RECT 18.09 4.369 18.176 4.74 ;
      RECT 18.07 4.376 18.09 4.748 ;
      RECT 18.06 4.379 18.07 4.755 ;
      RECT 17.995 4.384 18.06 4.773 ;
      RECT 17.965 4.391 17.995 4.798 ;
      RECT 17.955 4.394 17.965 4.805 ;
      RECT 17.91 4.398 17.955 4.81 ;
      RECT 17.88 4.403 17.91 4.815 ;
      RECT 17.879 4.405 17.88 4.815 ;
      RECT 17.793 4.411 17.879 4.815 ;
      RECT 17.707 4.422 17.793 4.815 ;
      RECT 17.621 4.434 17.707 4.815 ;
      RECT 17.535 4.445 17.621 4.815 ;
      RECT 17.52 4.452 17.535 4.81 ;
      RECT 17.515 4.454 17.52 4.804 ;
      RECT 17.495 4.465 17.515 4.799 ;
      RECT 17.485 4.483 17.495 4.793 ;
      RECT 17.48 4.495 17.485 4.593 ;
      RECT 19.775 3.248 19.795 3.335 ;
      RECT 19.77 3.183 19.775 3.367 ;
      RECT 19.76 3.15 19.77 3.372 ;
      RECT 19.755 3.13 19.76 3.378 ;
      RECT 19.725 3.13 19.755 3.395 ;
      RECT 19.676 3.13 19.725 3.431 ;
      RECT 19.59 3.13 19.676 3.489 ;
      RECT 19.561 3.14 19.59 3.538 ;
      RECT 19.475 3.182 19.561 3.591 ;
      RECT 19.455 3.22 19.475 3.638 ;
      RECT 19.43 3.237 19.455 3.658 ;
      RECT 19.42 3.251 19.43 3.678 ;
      RECT 19.415 3.257 19.42 3.688 ;
      RECT 19.41 3.261 19.415 3.695 ;
      RECT 19.36 3.281 19.41 3.7 ;
      RECT 19.295 3.325 19.36 3.7 ;
      RECT 19.27 3.375 19.295 3.7 ;
      RECT 19.26 3.405 19.27 3.7 ;
      RECT 19.255 3.432 19.26 3.7 ;
      RECT 19.25 3.45 19.255 3.7 ;
      RECT 19.24 3.492 19.25 3.7 ;
      RECT 19.59 4.05 19.76 4.225 ;
      RECT 19.53 3.878 19.59 4.213 ;
      RECT 19.52 3.871 19.53 4.196 ;
      RECT 19.475 4.05 19.76 4.176 ;
      RECT 19.456 4.05 19.76 4.154 ;
      RECT 19.37 4.05 19.76 4.119 ;
      RECT 19.35 3.87 19.52 4.075 ;
      RECT 19.35 4.017 19.755 4.075 ;
      RECT 19.35 3.965 19.73 4.075 ;
      RECT 19.35 3.92 19.695 4.075 ;
      RECT 19.35 3.902 19.66 4.075 ;
      RECT 19.35 3.892 19.655 4.075 ;
      RECT 19.52 10.14 19.69 10.59 ;
      RECT 19.575 8.36 19.745 10.31 ;
      RECT 19.52 7.3 19.69 8.53 ;
      RECT 19 7.3 19.17 10.59 ;
      RECT 19 9.6 19.405 9.93 ;
      RECT 19 8.76 19.405 9.09 ;
      RECT 19.07 4.85 19.26 5.075 ;
      RECT 19.06 4.851 19.265 5.07 ;
      RECT 19.06 4.853 19.275 5.05 ;
      RECT 19.06 4.857 19.28 5.035 ;
      RECT 19.06 4.844 19.23 5.07 ;
      RECT 19.06 4.847 19.255 5.07 ;
      RECT 19.07 4.843 19.23 5.075 ;
      RECT 19.156 4.841 19.23 5.075 ;
      RECT 18.78 4.092 18.95 4.33 ;
      RECT 18.78 4.092 19.036 4.244 ;
      RECT 18.78 4.092 19.04 4.154 ;
      RECT 18.83 3.865 19.05 4.133 ;
      RECT 18.825 3.882 19.055 4.106 ;
      RECT 18.79 4.04 19.055 4.106 ;
      RECT 18.81 3.89 18.95 4.33 ;
      RECT 18.8 3.972 19.06 4.089 ;
      RECT 18.795 4.02 19.06 4.089 ;
      RECT 18.8 3.93 19.055 4.106 ;
      RECT 18.825 3.867 19.05 4.133 ;
      RECT 18.39 3.842 18.56 4.04 ;
      RECT 18.39 3.842 18.605 4.015 ;
      RECT 18.46 3.785 18.63 3.973 ;
      RECT 18.435 3.8 18.63 3.973 ;
      RECT 18.05 3.846 18.08 4.04 ;
      RECT 18.045 3.818 18.05 4.04 ;
      RECT 18.015 3.792 18.045 4.042 ;
      RECT 17.99 3.75 18.015 4.045 ;
      RECT 17.98 3.722 17.99 4.047 ;
      RECT 17.945 3.702 17.98 4.049 ;
      RECT 17.88 3.687 17.945 4.055 ;
      RECT 17.83 3.685 17.88 4.061 ;
      RECT 17.807 3.687 17.83 4.066 ;
      RECT 17.721 3.698 17.807 4.072 ;
      RECT 17.635 3.716 17.721 4.082 ;
      RECT 17.62 3.727 17.635 4.088 ;
      RECT 17.55 3.75 17.62 4.094 ;
      RECT 17.495 3.782 17.55 4.102 ;
      RECT 17.455 3.805 17.495 4.108 ;
      RECT 17.441 3.818 17.455 4.111 ;
      RECT 17.355 3.84 17.441 4.117 ;
      RECT 17.34 3.865 17.355 4.123 ;
      RECT 17.3 3.88 17.34 4.127 ;
      RECT 17.25 3.895 17.3 4.132 ;
      RECT 17.225 3.902 17.25 4.136 ;
      RECT 17.165 3.897 17.225 4.14 ;
      RECT 17.15 3.888 17.165 4.144 ;
      RECT 17.08 3.878 17.15 4.14 ;
      RECT 17.055 3.87 17.075 4.13 ;
      RECT 16.996 3.87 17.055 4.108 ;
      RECT 16.91 3.87 16.996 4.065 ;
      RECT 17.075 3.87 17.08 4.135 ;
      RECT 17.77 3.101 17.94 3.435 ;
      RECT 17.74 3.101 17.94 3.43 ;
      RECT 17.68 3.068 17.74 3.418 ;
      RECT 17.68 3.124 17.95 3.413 ;
      RECT 17.655 3.124 17.95 3.407 ;
      RECT 17.65 3.065 17.68 3.404 ;
      RECT 17.635 3.071 17.77 3.402 ;
      RECT 17.63 3.079 17.855 3.39 ;
      RECT 17.63 3.131 17.965 3.343 ;
      RECT 17.615 3.087 17.855 3.338 ;
      RECT 17.615 3.157 17.975 3.279 ;
      RECT 17.585 3.107 17.94 3.24 ;
      RECT 17.585 3.197 17.985 3.236 ;
      RECT 17.635 3.076 17.855 3.402 ;
      RECT 16.975 3.406 17.03 3.67 ;
      RECT 16.975 3.406 17.095 3.669 ;
      RECT 16.975 3.406 17.12 3.668 ;
      RECT 16.975 3.406 17.185 3.667 ;
      RECT 17.12 3.372 17.2 3.666 ;
      RECT 16.935 3.416 17.345 3.665 ;
      RECT 16.975 3.413 17.345 3.665 ;
      RECT 16.935 3.421 17.35 3.658 ;
      RECT 16.92 3.423 17.35 3.657 ;
      RECT 16.92 3.43 17.355 3.653 ;
      RECT 16.9 3.429 17.35 3.649 ;
      RECT 16.9 3.437 17.36 3.648 ;
      RECT 16.895 3.434 17.355 3.644 ;
      RECT 16.895 3.447 17.37 3.643 ;
      RECT 16.88 3.437 17.36 3.642 ;
      RECT 16.845 3.45 17.37 3.635 ;
      RECT 17.03 3.405 17.34 3.665 ;
      RECT 17.03 3.39 17.29 3.665 ;
      RECT 17.095 3.377 17.225 3.665 ;
      RECT 16.64 4.466 16.655 4.859 ;
      RECT 16.605 4.471 16.655 4.858 ;
      RECT 16.64 4.47 16.7 4.857 ;
      RECT 16.585 4.481 16.7 4.856 ;
      RECT 16.6 4.477 16.7 4.856 ;
      RECT 16.565 4.487 16.775 4.853 ;
      RECT 16.565 4.506 16.82 4.851 ;
      RECT 16.565 4.513 16.825 4.848 ;
      RECT 16.55 4.49 16.775 4.845 ;
      RECT 16.53 4.495 16.775 4.838 ;
      RECT 16.525 4.499 16.775 4.834 ;
      RECT 16.525 4.516 16.835 4.833 ;
      RECT 16.505 4.51 16.82 4.829 ;
      RECT 16.505 4.519 16.84 4.823 ;
      RECT 16.5 4.525 16.84 4.595 ;
      RECT 16.565 4.485 16.7 4.853 ;
      RECT 16.44 3.848 16.64 4.16 ;
      RECT 16.515 3.826 16.64 4.16 ;
      RECT 16.455 3.845 16.645 4.145 ;
      RECT 16.425 3.856 16.645 4.143 ;
      RECT 16.44 3.851 16.65 4.109 ;
      RECT 16.425 3.955 16.655 4.076 ;
      RECT 16.455 3.827 16.64 4.16 ;
      RECT 16.515 3.805 16.615 4.16 ;
      RECT 16.54 3.802 16.615 4.16 ;
      RECT 16.54 3.797 16.56 4.16 ;
      RECT 15.945 3.865 16.12 4.04 ;
      RECT 15.94 3.865 16.12 4.038 ;
      RECT 15.915 3.865 16.12 4.033 ;
      RECT 15.86 3.845 16.03 4.023 ;
      RECT 15.86 3.852 16.095 4.023 ;
      RECT 15.945 4.532 15.96 4.715 ;
      RECT 15.935 4.51 15.945 4.715 ;
      RECT 15.92 4.49 15.935 4.715 ;
      RECT 15.91 4.465 15.92 4.715 ;
      RECT 15.88 4.43 15.91 4.715 ;
      RECT 15.845 4.37 15.88 4.715 ;
      RECT 15.84 4.332 15.845 4.715 ;
      RECT 15.79 4.283 15.84 4.715 ;
      RECT 15.78 4.233 15.79 4.703 ;
      RECT 15.765 4.212 15.78 4.663 ;
      RECT 15.745 4.18 15.765 4.613 ;
      RECT 15.72 4.136 15.745 4.553 ;
      RECT 15.715 4.108 15.72 4.508 ;
      RECT 15.71 4.099 15.715 4.494 ;
      RECT 15.705 4.092 15.71 4.481 ;
      RECT 15.7 4.087 15.705 4.47 ;
      RECT 15.695 4.072 15.7 4.46 ;
      RECT 15.69 4.05 15.695 4.447 ;
      RECT 15.68 4.01 15.69 4.422 ;
      RECT 15.655 3.94 15.68 4.378 ;
      RECT 15.65 3.88 15.655 4.343 ;
      RECT 15.635 3.86 15.65 4.31 ;
      RECT 15.63 3.86 15.635 4.285 ;
      RECT 15.6 3.86 15.63 4.24 ;
      RECT 15.555 3.86 15.6 4.18 ;
      RECT 15.48 3.86 15.555 4.128 ;
      RECT 15.475 3.86 15.48 4.093 ;
      RECT 15.47 3.86 15.475 4.083 ;
      RECT 15.465 3.86 15.47 4.063 ;
      RECT 15.73 3.08 15.9 3.55 ;
      RECT 15.675 3.073 15.87 3.534 ;
      RECT 15.675 3.087 15.905 3.533 ;
      RECT 15.66 3.088 15.905 3.514 ;
      RECT 15.655 3.106 15.905 3.5 ;
      RECT 15.66 3.089 15.91 3.498 ;
      RECT 15.645 3.12 15.91 3.483 ;
      RECT 15.66 3.095 15.915 3.468 ;
      RECT 15.64 3.135 15.915 3.465 ;
      RECT 15.655 3.107 15.92 3.45 ;
      RECT 15.655 3.119 15.925 3.43 ;
      RECT 15.64 3.135 15.93 3.413 ;
      RECT 15.64 3.145 15.935 3.268 ;
      RECT 15.635 3.145 15.935 3.225 ;
      RECT 15.635 3.16 15.94 3.203 ;
      RECT 15.73 3.07 15.87 3.55 ;
      RECT 15.73 3.068 15.84 3.55 ;
      RECT 15.816 3.065 15.84 3.55 ;
      RECT 15.475 4.732 15.48 4.778 ;
      RECT 15.465 4.58 15.475 4.802 ;
      RECT 15.46 4.425 15.465 4.827 ;
      RECT 15.445 4.387 15.46 4.838 ;
      RECT 15.44 4.37 15.445 4.845 ;
      RECT 15.43 4.358 15.44 4.852 ;
      RECT 15.425 4.349 15.43 4.854 ;
      RECT 15.42 4.347 15.425 4.858 ;
      RECT 15.375 4.338 15.42 4.873 ;
      RECT 15.37 4.33 15.375 4.887 ;
      RECT 15.365 4.327 15.37 4.891 ;
      RECT 15.35 4.322 15.365 4.899 ;
      RECT 15.295 4.312 15.35 4.91 ;
      RECT 15.26 4.3 15.295 4.911 ;
      RECT 15.251 4.295 15.26 4.905 ;
      RECT 15.165 4.295 15.251 4.895 ;
      RECT 15.135 4.295 15.165 4.873 ;
      RECT 15.125 4.295 15.13 4.853 ;
      RECT 15.12 4.295 15.125 4.815 ;
      RECT 15.115 4.295 15.12 4.773 ;
      RECT 15.11 4.295 15.115 4.733 ;
      RECT 15.105 4.295 15.11 4.663 ;
      RECT 15.095 4.295 15.105 4.585 ;
      RECT 15.09 4.295 15.095 4.485 ;
      RECT 15.13 4.295 15.135 4.855 ;
      RECT 14.625 4.377 14.715 4.855 ;
      RECT 14.61 4.38 14.73 4.853 ;
      RECT 14.625 4.379 14.73 4.853 ;
      RECT 14.59 4.386 14.755 4.843 ;
      RECT 14.61 4.38 14.755 4.843 ;
      RECT 14.575 4.392 14.755 4.831 ;
      RECT 14.61 4.383 14.805 4.824 ;
      RECT 14.561 4.4 14.805 4.822 ;
      RECT 14.59 4.39 14.815 4.81 ;
      RECT 14.561 4.411 14.845 4.801 ;
      RECT 14.475 4.435 14.845 4.795 ;
      RECT 14.475 4.448 14.885 4.778 ;
      RECT 14.47 4.47 14.885 4.771 ;
      RECT 14.44 4.485 14.885 4.761 ;
      RECT 14.435 4.496 14.885 4.751 ;
      RECT 14.405 4.509 14.885 4.742 ;
      RECT 14.39 4.527 14.885 4.731 ;
      RECT 14.365 4.54 14.885 4.721 ;
      RECT 14.625 4.376 14.635 4.855 ;
      RECT 14.671 3.8 14.71 4.045 ;
      RECT 14.585 3.8 14.72 4.043 ;
      RECT 14.47 3.825 14.72 4.04 ;
      RECT 14.47 3.825 14.725 4.038 ;
      RECT 14.47 3.825 14.74 4.033 ;
      RECT 14.576 3.8 14.755 4.013 ;
      RECT 14.49 3.808 14.755 4.013 ;
      RECT 14.16 3.16 14.33 3.595 ;
      RECT 14.15 3.194 14.33 3.578 ;
      RECT 14.23 3.13 14.4 3.565 ;
      RECT 14.135 3.205 14.4 3.543 ;
      RECT 14.23 3.14 14.405 3.533 ;
      RECT 14.16 3.192 14.435 3.518 ;
      RECT 14.12 3.218 14.435 3.503 ;
      RECT 14.12 3.26 14.445 3.483 ;
      RECT 14.115 3.285 14.45 3.465 ;
      RECT 14.115 3.295 14.455 3.45 ;
      RECT 14.11 3.232 14.435 3.448 ;
      RECT 14.11 3.305 14.46 3.433 ;
      RECT 14.105 3.242 14.435 3.43 ;
      RECT 14.1 3.326 14.465 3.413 ;
      RECT 14.1 3.358 14.47 3.393 ;
      RECT 14.095 3.272 14.445 3.385 ;
      RECT 14.1 3.257 14.435 3.413 ;
      RECT 14.115 3.227 14.435 3.465 ;
      RECT 13.96 3.814 14.185 4.07 ;
      RECT 13.96 3.847 14.205 4.06 ;
      RECT 13.925 3.847 14.205 4.058 ;
      RECT 13.925 3.86 14.21 4.048 ;
      RECT 13.925 3.88 14.22 4.04 ;
      RECT 13.925 3.977 14.225 4.033 ;
      RECT 13.905 3.725 14.035 4.023 ;
      RECT 13.86 3.88 14.22 3.965 ;
      RECT 13.85 3.725 14.035 3.91 ;
      RECT 13.85 3.757 14.121 3.91 ;
      RECT 13.815 4.287 13.835 4.465 ;
      RECT 13.78 4.24 13.815 4.465 ;
      RECT 13.765 4.18 13.78 4.465 ;
      RECT 13.74 4.127 13.765 4.465 ;
      RECT 13.725 4.08 13.74 4.465 ;
      RECT 13.705 4.057 13.725 4.465 ;
      RECT 13.68 4.022 13.705 4.465 ;
      RECT 13.67 3.868 13.68 4.465 ;
      RECT 13.64 3.863 13.67 4.456 ;
      RECT 13.635 3.86 13.64 4.446 ;
      RECT 13.62 3.86 13.635 4.42 ;
      RECT 13.615 3.86 13.62 4.383 ;
      RECT 13.59 3.86 13.615 4.335 ;
      RECT 13.57 3.86 13.59 4.26 ;
      RECT 13.56 3.86 13.57 4.22 ;
      RECT 13.555 3.86 13.56 4.195 ;
      RECT 13.55 3.86 13.555 4.178 ;
      RECT 13.545 3.86 13.55 4.16 ;
      RECT 13.54 3.861 13.545 4.15 ;
      RECT 13.53 3.863 13.54 4.118 ;
      RECT 13.52 3.865 13.53 4.085 ;
      RECT 13.51 3.868 13.52 4.058 ;
      RECT 13.835 4.295 14.06 4.465 ;
      RECT 13.165 3.107 13.335 3.56 ;
      RECT 13.165 3.107 13.425 3.526 ;
      RECT 13.165 3.107 13.455 3.51 ;
      RECT 13.165 3.107 13.485 3.483 ;
      RECT 13.421 3.085 13.5 3.465 ;
      RECT 13.2 3.092 13.505 3.45 ;
      RECT 13.2 3.1 13.515 3.413 ;
      RECT 13.16 3.127 13.515 3.385 ;
      RECT 13.145 3.14 13.515 3.35 ;
      RECT 13.165 3.115 13.535 3.34 ;
      RECT 13.14 3.18 13.535 3.31 ;
      RECT 13.14 3.21 13.54 3.293 ;
      RECT 13.135 3.24 13.54 3.28 ;
      RECT 13.2 3.089 13.5 3.465 ;
      RECT 13.335 3.086 13.421 3.544 ;
      RECT 13.286 3.087 13.5 3.465 ;
      RECT 13.43 4.747 13.475 4.94 ;
      RECT 13.42 4.717 13.43 4.94 ;
      RECT 13.415 4.702 13.42 4.94 ;
      RECT 13.375 4.612 13.415 4.94 ;
      RECT 13.37 4.525 13.375 4.94 ;
      RECT 13.36 4.495 13.37 4.94 ;
      RECT 13.355 4.455 13.36 4.94 ;
      RECT 13.345 4.417 13.355 4.94 ;
      RECT 13.34 4.382 13.345 4.94 ;
      RECT 13.32 4.335 13.34 4.94 ;
      RECT 13.305 4.26 13.32 4.94 ;
      RECT 13.3 4.215 13.305 4.935 ;
      RECT 13.295 4.195 13.3 4.908 ;
      RECT 13.29 4.175 13.295 4.893 ;
      RECT 13.285 4.15 13.29 4.873 ;
      RECT 13.28 4.128 13.285 4.858 ;
      RECT 13.275 4.106 13.28 4.84 ;
      RECT 13.27 4.085 13.275 4.83 ;
      RECT 13.26 4.057 13.27 4.8 ;
      RECT 13.25 4.02 13.26 4.768 ;
      RECT 13.24 3.98 13.25 4.735 ;
      RECT 13.23 3.958 13.24 4.705 ;
      RECT 13.2 3.91 13.23 4.637 ;
      RECT 13.185 3.87 13.2 4.564 ;
      RECT 13.175 3.87 13.185 4.53 ;
      RECT 13.17 3.87 13.175 4.505 ;
      RECT 13.165 3.87 13.17 4.49 ;
      RECT 13.16 3.87 13.165 4.468 ;
      RECT 13.155 3.87 13.16 4.455 ;
      RECT 13.14 3.87 13.155 4.42 ;
      RECT 13.12 3.87 13.14 4.36 ;
      RECT 13.11 3.87 13.12 4.31 ;
      RECT 13.09 3.87 13.11 4.258 ;
      RECT 13.07 3.87 13.09 4.215 ;
      RECT 13.06 3.87 13.07 4.203 ;
      RECT 13.03 3.87 13.06 4.19 ;
      RECT 13 3.891 13.03 4.17 ;
      RECT 12.99 3.919 13 4.15 ;
      RECT 12.975 3.936 12.99 4.118 ;
      RECT 12.97 3.95 12.975 4.085 ;
      RECT 12.965 3.958 12.97 4.058 ;
      RECT 12.96 3.966 12.965 4.02 ;
      RECT 12.965 4.49 12.97 4.825 ;
      RECT 12.93 4.477 12.965 4.824 ;
      RECT 12.86 4.417 12.93 4.823 ;
      RECT 12.78 4.36 12.86 4.822 ;
      RECT 12.645 4.32 12.78 4.821 ;
      RECT 12.645 4.507 12.98 4.81 ;
      RECT 12.605 4.507 12.98 4.8 ;
      RECT 12.605 4.525 12.985 4.795 ;
      RECT 12.605 4.615 12.99 4.785 ;
      RECT 12.6 4.31 12.765 4.765 ;
      RECT 12.595 4.31 12.765 4.508 ;
      RECT 12.595 4.467 12.96 4.508 ;
      RECT 12.595 4.455 12.955 4.508 ;
      RECT 10.645 10.14 10.815 10.59 ;
      RECT 10.7 8.36 10.87 10.31 ;
      RECT 10.645 7.3 10.815 8.53 ;
      RECT 10.125 7.3 10.295 10.59 ;
      RECT 10.125 9.6 10.53 9.93 ;
      RECT 10.125 8.76 10.53 9.09 ;
      RECT 90.635 7.305 90.805 8.775 ;
      RECT 90.635 10.085 90.805 10.595 ;
      RECT 89.645 1.865 89.815 2.375 ;
      RECT 89.645 3.685 89.815 5.155 ;
      RECT 89.645 7.305 89.815 8.775 ;
      RECT 89.645 10.085 89.815 10.595 ;
      RECT 88.285 1.87 88.455 5.16 ;
      RECT 88.285 7.3 88.455 10.59 ;
      RECT 87.855 1.87 88.025 2.38 ;
      RECT 87.855 2.95 88.025 5.16 ;
      RECT 87.855 7.3 88.025 9.51 ;
      RECT 87.855 10.08 88.025 10.59 ;
      RECT 85.465 4.145 85.835 4.515 ;
      RECT 83.505 7.3 83.675 10.59 ;
      RECT 83.075 7.3 83.245 9.51 ;
      RECT 83.075 10.08 83.245 10.59 ;
      RECT 74.85 7.305 75.02 8.775 ;
      RECT 74.85 10.085 75.02 10.595 ;
      RECT 73.86 1.865 74.03 2.375 ;
      RECT 73.86 3.685 74.03 5.155 ;
      RECT 73.86 7.305 74.03 8.775 ;
      RECT 73.86 10.085 74.03 10.595 ;
      RECT 72.5 1.87 72.67 5.16 ;
      RECT 72.5 7.3 72.67 10.59 ;
      RECT 72.07 1.87 72.24 2.38 ;
      RECT 72.07 2.95 72.24 5.16 ;
      RECT 72.07 7.3 72.24 9.51 ;
      RECT 72.07 10.08 72.24 10.59 ;
      RECT 69.68 4.145 70.05 4.515 ;
      RECT 67.72 7.3 67.89 10.59 ;
      RECT 67.29 7.3 67.46 9.51 ;
      RECT 67.29 10.08 67.46 10.59 ;
      RECT 59.065 7.305 59.235 8.775 ;
      RECT 59.065 10.085 59.235 10.595 ;
      RECT 58.075 1.865 58.245 2.375 ;
      RECT 58.075 3.685 58.245 5.155 ;
      RECT 58.075 7.305 58.245 8.775 ;
      RECT 58.075 10.085 58.245 10.595 ;
      RECT 56.715 1.87 56.885 5.16 ;
      RECT 56.715 7.3 56.885 10.59 ;
      RECT 56.285 1.87 56.455 2.38 ;
      RECT 56.285 2.95 56.455 5.16 ;
      RECT 56.285 7.3 56.455 9.51 ;
      RECT 56.285 10.08 56.455 10.59 ;
      RECT 53.895 4.145 54.265 4.515 ;
      RECT 51.935 7.3 52.105 10.59 ;
      RECT 51.505 7.3 51.675 9.51 ;
      RECT 51.505 10.08 51.675 10.59 ;
      RECT 43.29 7.305 43.46 8.775 ;
      RECT 43.29 10.085 43.46 10.595 ;
      RECT 42.3 1.865 42.47 2.375 ;
      RECT 42.3 3.685 42.47 5.155 ;
      RECT 42.3 7.305 42.47 8.775 ;
      RECT 42.3 10.085 42.47 10.595 ;
      RECT 40.94 1.87 41.11 5.16 ;
      RECT 40.94 7.3 41.11 10.59 ;
      RECT 40.51 1.87 40.68 2.38 ;
      RECT 40.51 2.95 40.68 5.16 ;
      RECT 40.51 7.3 40.68 9.51 ;
      RECT 40.51 10.08 40.68 10.59 ;
      RECT 38.12 4.145 38.49 4.515 ;
      RECT 36.16 7.3 36.33 10.59 ;
      RECT 35.73 7.3 35.9 9.51 ;
      RECT 35.73 10.08 35.9 10.59 ;
      RECT 27.51 7.305 27.68 8.775 ;
      RECT 27.51 10.085 27.68 10.595 ;
      RECT 26.52 1.865 26.69 2.375 ;
      RECT 26.52 3.685 26.69 5.155 ;
      RECT 26.52 7.305 26.69 8.775 ;
      RECT 26.52 10.085 26.69 10.595 ;
      RECT 25.16 1.87 25.33 5.16 ;
      RECT 25.16 7.3 25.33 10.59 ;
      RECT 24.73 1.87 24.9 2.38 ;
      RECT 24.73 2.95 24.9 5.16 ;
      RECT 24.73 7.3 24.9 9.51 ;
      RECT 24.73 10.08 24.9 10.59 ;
      RECT 22.34 4.145 22.71 4.515 ;
      RECT 20.38 7.3 20.55 10.59 ;
      RECT 19.95 7.3 20.12 9.51 ;
      RECT 19.95 10.08 20.12 10.59 ;
      RECT 11.075 7.3 11.245 9.51 ;
      RECT 11.075 10.08 11.245 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r1
  CLASS BLOCK ;
  ORIGIN -12.955 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r1 ;
  SIZE 92.44 BY 12.61 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 33.145 1.865 33.315 2.375 ;
        RECT 33.145 3.685 33.315 5.155 ;
      LAYER met1 ;
        RECT 33.085 3.655 33.375 3.885 ;
        RECT 33.085 2.175 33.375 2.405 ;
        RECT 33.145 2.175 33.315 3.885 ;
      LAYER mcon ;
        RECT 33.145 3.685 33.315 3.855 ;
        RECT 33.145 2.205 33.315 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 51.07 1.865 51.24 2.375 ;
        RECT 51.07 3.685 51.24 5.155 ;
      LAYER met1 ;
        RECT 51.01 3.655 51.3 3.885 ;
        RECT 51.01 2.175 51.3 2.405 ;
        RECT 51.07 2.175 51.24 3.885 ;
      LAYER mcon ;
        RECT 51.07 3.685 51.24 3.855 ;
        RECT 51.07 2.205 51.24 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 68.995 1.865 69.165 2.375 ;
        RECT 68.995 3.685 69.165 5.155 ;
      LAYER met1 ;
        RECT 68.935 3.655 69.225 3.885 ;
        RECT 68.935 2.175 69.225 2.405 ;
        RECT 68.995 2.175 69.165 3.885 ;
      LAYER mcon ;
        RECT 68.995 3.685 69.165 3.855 ;
        RECT 68.995 2.205 69.165 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 86.92 1.865 87.09 2.375 ;
        RECT 86.92 3.685 87.09 5.155 ;
      LAYER met1 ;
        RECT 86.86 3.655 87.15 3.885 ;
        RECT 86.86 2.175 87.15 2.405 ;
        RECT 86.92 2.175 87.09 3.885 ;
      LAYER mcon ;
        RECT 86.92 3.685 87.09 3.855 ;
        RECT 86.92 2.205 87.09 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 104.845 1.865 105.015 2.375 ;
        RECT 104.845 3.685 105.015 5.155 ;
      LAYER met1 ;
        RECT 104.785 3.655 105.075 3.885 ;
        RECT 104.785 2.175 105.075 2.405 ;
        RECT 104.845 2.175 105.015 3.885 ;
      LAYER mcon ;
        RECT 104.845 3.685 105.015 3.855 ;
        RECT 104.845 2.205 105.015 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 28.995 2.955 29.165 4.23 ;
        RECT 28.995 8.38 29.165 9.655 ;
        RECT 24.235 8.38 24.405 9.655 ;
      LAYER met2 ;
        RECT 28.915 4 29.265 4.35 ;
        RECT 28.905 8.275 29.255 8.625 ;
        RECT 28.98 4 29.155 8.625 ;
      LAYER met1 ;
        RECT 28.915 4.06 29.395 4.23 ;
        RECT 28.915 4 29.265 4.35 ;
        RECT 24.175 8.38 29.395 8.55 ;
        RECT 28.905 8.275 29.255 8.625 ;
        RECT 24.175 8.35 24.465 8.58 ;
      LAYER via1 ;
        RECT 29.005 8.375 29.155 8.525 ;
        RECT 29.015 4.1 29.165 4.25 ;
      LAYER mcon ;
        RECT 24.235 8.38 24.405 8.55 ;
        RECT 28.995 8.38 29.165 8.55 ;
        RECT 28.995 4.06 29.165 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 46.92 2.955 47.09 4.23 ;
        RECT 46.92 8.38 47.09 9.655 ;
        RECT 42.16 8.38 42.33 9.655 ;
      LAYER met2 ;
        RECT 46.84 4 47.19 4.35 ;
        RECT 46.83 8.275 47.18 8.625 ;
        RECT 46.905 4 47.08 8.625 ;
      LAYER met1 ;
        RECT 46.84 4.06 47.32 4.23 ;
        RECT 46.84 4 47.19 4.35 ;
        RECT 42.1 8.38 47.32 8.55 ;
        RECT 46.83 8.275 47.18 8.625 ;
        RECT 42.1 8.35 42.39 8.58 ;
      LAYER via1 ;
        RECT 46.93 8.375 47.08 8.525 ;
        RECT 46.94 4.1 47.09 4.25 ;
      LAYER mcon ;
        RECT 42.16 8.38 42.33 8.55 ;
        RECT 46.92 8.38 47.09 8.55 ;
        RECT 46.92 4.06 47.09 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 64.845 2.955 65.015 4.23 ;
        RECT 64.845 8.38 65.015 9.655 ;
        RECT 60.085 8.38 60.255 9.655 ;
      LAYER met2 ;
        RECT 64.765 4 65.115 4.35 ;
        RECT 64.755 8.275 65.105 8.625 ;
        RECT 64.83 4 65.005 8.625 ;
      LAYER met1 ;
        RECT 64.765 4.06 65.245 4.23 ;
        RECT 64.765 4 65.115 4.35 ;
        RECT 60.025 8.38 65.245 8.55 ;
        RECT 64.755 8.275 65.105 8.625 ;
        RECT 60.025 8.35 60.315 8.58 ;
      LAYER via1 ;
        RECT 64.855 8.375 65.005 8.525 ;
        RECT 64.865 4.1 65.015 4.25 ;
      LAYER mcon ;
        RECT 60.085 8.38 60.255 8.55 ;
        RECT 64.845 8.38 65.015 8.55 ;
        RECT 64.845 4.06 65.015 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 82.77 2.955 82.94 4.23 ;
        RECT 82.77 8.38 82.94 9.655 ;
        RECT 78.01 8.38 78.18 9.655 ;
      LAYER met2 ;
        RECT 82.69 4 83.04 4.35 ;
        RECT 82.68 8.275 83.03 8.625 ;
        RECT 82.755 4 82.93 8.625 ;
      LAYER met1 ;
        RECT 82.69 4.06 83.17 4.23 ;
        RECT 82.69 4 83.04 4.35 ;
        RECT 77.95 8.38 83.17 8.55 ;
        RECT 82.68 8.275 83.03 8.625 ;
        RECT 77.95 8.35 78.24 8.58 ;
      LAYER via1 ;
        RECT 82.78 8.375 82.93 8.525 ;
        RECT 82.79 4.1 82.94 4.25 ;
      LAYER mcon ;
        RECT 78.01 8.38 78.18 8.55 ;
        RECT 82.77 8.38 82.94 8.55 ;
        RECT 82.77 4.06 82.94 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 100.695 2.955 100.865 4.23 ;
        RECT 100.695 8.38 100.865 9.655 ;
        RECT 95.935 8.38 96.105 9.655 ;
      LAYER met2 ;
        RECT 100.615 4 100.965 4.35 ;
        RECT 100.605 8.275 100.955 8.625 ;
        RECT 100.68 4 100.855 8.625 ;
      LAYER met1 ;
        RECT 100.615 4.06 101.095 4.23 ;
        RECT 100.615 4 100.965 4.35 ;
        RECT 95.875 8.38 101.095 8.55 ;
        RECT 100.605 8.275 100.955 8.625 ;
        RECT 95.875 8.35 96.165 8.58 ;
      LAYER via1 ;
        RECT 100.705 8.375 100.855 8.525 ;
        RECT 100.715 4.1 100.865 4.25 ;
      LAYER mcon ;
        RECT 95.935 8.38 96.105 8.55 ;
        RECT 100.695 8.38 100.865 8.55 ;
        RECT 100.695 4.06 100.865 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 13.205 8.38 13.375 9.655 ;
      LAYER met1 ;
        RECT 13.145 8.38 13.605 8.55 ;
        RECT 13.145 8.35 13.435 8.58 ;
      LAYER mcon ;
        RECT 13.205 8.38 13.375 8.55 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 12.97 5.58 105.39 7.18 ;
        RECT 99.43 5.43 105.39 7.18 ;
        RECT 103.255 5.425 105.235 7.185 ;
        RECT 104.415 4.695 104.585 7.915 ;
        RECT 103.425 4.695 103.595 7.915 ;
        RECT 100.685 4.7 100.855 7.91 ;
        RECT 97.93 5.08 98.1 7.18 ;
        RECT 95.925 5.58 96.095 7.91 ;
        RECT 95.49 5.08 95.66 7.18 ;
        RECT 93.53 5.08 93.7 7.18 ;
        RECT 92.57 5.08 92.74 7.18 ;
        RECT 90.61 5.08 90.78 7.18 ;
        RECT 89.61 5.08 89.78 7.18 ;
        RECT 88.65 5.08 88.82 7.18 ;
        RECT 81.505 5.43 87.465 7.18 ;
        RECT 85.33 5.425 87.31 7.185 ;
        RECT 86.49 4.695 86.66 7.915 ;
        RECT 85.5 4.695 85.67 7.915 ;
        RECT 82.76 4.7 82.93 7.91 ;
        RECT 80.005 5.08 80.175 7.18 ;
        RECT 78 5.58 78.17 7.91 ;
        RECT 77.565 5.08 77.735 7.18 ;
        RECT 75.605 5.08 75.775 7.18 ;
        RECT 74.645 5.08 74.815 7.18 ;
        RECT 72.685 5.08 72.855 7.18 ;
        RECT 71.685 5.08 71.855 7.18 ;
        RECT 70.725 5.08 70.895 7.18 ;
        RECT 63.58 5.43 69.54 7.18 ;
        RECT 67.405 5.425 69.385 7.185 ;
        RECT 68.565 4.695 68.735 7.915 ;
        RECT 67.575 4.695 67.745 7.915 ;
        RECT 64.835 4.7 65.005 7.91 ;
        RECT 62.08 5.08 62.25 7.18 ;
        RECT 60.075 5.58 60.245 7.91 ;
        RECT 59.64 5.08 59.81 7.18 ;
        RECT 57.68 5.08 57.85 7.18 ;
        RECT 56.72 5.08 56.89 7.18 ;
        RECT 54.76 5.08 54.93 7.18 ;
        RECT 53.76 5.08 53.93 7.18 ;
        RECT 52.8 5.08 52.97 7.18 ;
        RECT 45.655 5.43 51.615 7.18 ;
        RECT 49.48 5.425 51.46 7.185 ;
        RECT 50.64 4.695 50.81 7.915 ;
        RECT 49.65 4.695 49.82 7.915 ;
        RECT 46.91 4.7 47.08 7.91 ;
        RECT 44.155 5.08 44.325 7.18 ;
        RECT 42.15 5.58 42.32 7.91 ;
        RECT 41.715 5.08 41.885 7.18 ;
        RECT 39.755 5.08 39.925 7.18 ;
        RECT 38.795 5.08 38.965 7.18 ;
        RECT 36.835 5.08 37.005 7.18 ;
        RECT 35.835 5.08 36.005 7.18 ;
        RECT 34.875 5.08 35.045 7.18 ;
        RECT 27.73 5.43 33.69 7.18 ;
        RECT 31.555 5.425 33.535 7.185 ;
        RECT 32.715 4.695 32.885 7.915 ;
        RECT 31.725 4.695 31.895 7.915 ;
        RECT 28.985 4.7 29.155 7.91 ;
        RECT 26.23 5.08 26.4 7.18 ;
        RECT 24.225 5.58 24.395 7.91 ;
        RECT 23.79 5.08 23.96 7.18 ;
        RECT 21.83 5.08 22 7.18 ;
        RECT 20.87 5.08 21.04 7.18 ;
        RECT 18.91 5.08 19.08 7.18 ;
        RECT 17.91 5.08 18.08 7.18 ;
        RECT 16.95 5.08 17.12 7.18 ;
        RECT 15.005 5.58 15.175 10.74 ;
        RECT 13.195 5.58 13.365 7.91 ;
      LAYER met1 ;
        RECT 12.97 5.58 105.39 7.18 ;
        RECT 87.84 5.43 105.39 7.18 ;
        RECT 103.255 5.425 105.235 7.185 ;
        RECT 87.84 5.425 99.8 7.18 ;
        RECT 69.915 5.43 87.465 7.18 ;
        RECT 85.33 5.425 87.31 7.185 ;
        RECT 69.915 5.425 81.875 7.18 ;
        RECT 51.99 5.43 69.54 7.18 ;
        RECT 67.405 5.425 69.385 7.185 ;
        RECT 51.99 5.425 63.95 7.18 ;
        RECT 34.065 5.43 51.615 7.18 ;
        RECT 49.48 5.425 51.46 7.185 ;
        RECT 34.065 5.425 46.025 7.18 ;
        RECT 16.14 5.43 33.69 7.18 ;
        RECT 31.555 5.425 33.535 7.185 ;
        RECT 16.14 5.425 28.1 7.18 ;
        RECT 14.945 9.09 15.235 9.32 ;
        RECT 14.775 9.12 15.235 9.29 ;
      LAYER mcon ;
        RECT 15.005 9.12 15.175 9.29 ;
        RECT 15.315 6.98 15.485 7.15 ;
        RECT 16.285 5.58 16.455 5.75 ;
        RECT 16.745 5.58 16.915 5.75 ;
        RECT 17.205 5.58 17.375 5.75 ;
        RECT 17.665 5.58 17.835 5.75 ;
        RECT 18.125 5.58 18.295 5.75 ;
        RECT 18.585 5.58 18.755 5.75 ;
        RECT 19.045 5.58 19.215 5.75 ;
        RECT 19.505 5.58 19.675 5.75 ;
        RECT 19.965 5.58 20.135 5.75 ;
        RECT 20.425 5.58 20.595 5.75 ;
        RECT 20.885 5.58 21.055 5.75 ;
        RECT 21.345 5.58 21.515 5.75 ;
        RECT 21.805 5.58 21.975 5.75 ;
        RECT 22.265 5.58 22.435 5.75 ;
        RECT 22.725 5.58 22.895 5.75 ;
        RECT 23.185 5.58 23.355 5.75 ;
        RECT 23.645 5.58 23.815 5.75 ;
        RECT 24.105 5.58 24.275 5.75 ;
        RECT 24.565 5.58 24.735 5.75 ;
        RECT 25.025 5.58 25.195 5.75 ;
        RECT 25.485 5.58 25.655 5.75 ;
        RECT 25.945 5.58 26.115 5.75 ;
        RECT 26.345 6.98 26.515 7.15 ;
        RECT 26.405 5.58 26.575 5.75 ;
        RECT 26.865 5.58 27.035 5.75 ;
        RECT 27.325 5.58 27.495 5.75 ;
        RECT 27.785 5.58 27.955 5.75 ;
        RECT 31.105 6.98 31.275 7.15 ;
        RECT 31.105 5.46 31.275 5.63 ;
        RECT 31.805 6.985 31.975 7.155 ;
        RECT 31.805 5.455 31.975 5.625 ;
        RECT 32.795 6.985 32.965 7.155 ;
        RECT 32.795 5.455 32.965 5.625 ;
        RECT 34.21 5.58 34.38 5.75 ;
        RECT 34.67 5.58 34.84 5.75 ;
        RECT 35.13 5.58 35.3 5.75 ;
        RECT 35.59 5.58 35.76 5.75 ;
        RECT 36.05 5.58 36.22 5.75 ;
        RECT 36.51 5.58 36.68 5.75 ;
        RECT 36.97 5.58 37.14 5.75 ;
        RECT 37.43 5.58 37.6 5.75 ;
        RECT 37.89 5.58 38.06 5.75 ;
        RECT 38.35 5.58 38.52 5.75 ;
        RECT 38.81 5.58 38.98 5.75 ;
        RECT 39.27 5.58 39.44 5.75 ;
        RECT 39.73 5.58 39.9 5.75 ;
        RECT 40.19 5.58 40.36 5.75 ;
        RECT 40.65 5.58 40.82 5.75 ;
        RECT 41.11 5.58 41.28 5.75 ;
        RECT 41.57 5.58 41.74 5.75 ;
        RECT 42.03 5.58 42.2 5.75 ;
        RECT 42.49 5.58 42.66 5.75 ;
        RECT 42.95 5.58 43.12 5.75 ;
        RECT 43.41 5.58 43.58 5.75 ;
        RECT 43.87 5.58 44.04 5.75 ;
        RECT 44.27 6.98 44.44 7.15 ;
        RECT 44.33 5.58 44.5 5.75 ;
        RECT 44.79 5.58 44.96 5.75 ;
        RECT 45.25 5.58 45.42 5.75 ;
        RECT 45.71 5.58 45.88 5.75 ;
        RECT 49.03 6.98 49.2 7.15 ;
        RECT 49.03 5.46 49.2 5.63 ;
        RECT 49.73 6.985 49.9 7.155 ;
        RECT 49.73 5.455 49.9 5.625 ;
        RECT 50.72 6.985 50.89 7.155 ;
        RECT 50.72 5.455 50.89 5.625 ;
        RECT 52.135 5.58 52.305 5.75 ;
        RECT 52.595 5.58 52.765 5.75 ;
        RECT 53.055 5.58 53.225 5.75 ;
        RECT 53.515 5.58 53.685 5.75 ;
        RECT 53.975 5.58 54.145 5.75 ;
        RECT 54.435 5.58 54.605 5.75 ;
        RECT 54.895 5.58 55.065 5.75 ;
        RECT 55.355 5.58 55.525 5.75 ;
        RECT 55.815 5.58 55.985 5.75 ;
        RECT 56.275 5.58 56.445 5.75 ;
        RECT 56.735 5.58 56.905 5.75 ;
        RECT 57.195 5.58 57.365 5.75 ;
        RECT 57.655 5.58 57.825 5.75 ;
        RECT 58.115 5.58 58.285 5.75 ;
        RECT 58.575 5.58 58.745 5.75 ;
        RECT 59.035 5.58 59.205 5.75 ;
        RECT 59.495 5.58 59.665 5.75 ;
        RECT 59.955 5.58 60.125 5.75 ;
        RECT 60.415 5.58 60.585 5.75 ;
        RECT 60.875 5.58 61.045 5.75 ;
        RECT 61.335 5.58 61.505 5.75 ;
        RECT 61.795 5.58 61.965 5.75 ;
        RECT 62.195 6.98 62.365 7.15 ;
        RECT 62.255 5.58 62.425 5.75 ;
        RECT 62.715 5.58 62.885 5.75 ;
        RECT 63.175 5.58 63.345 5.75 ;
        RECT 63.635 5.58 63.805 5.75 ;
        RECT 66.955 6.98 67.125 7.15 ;
        RECT 66.955 5.46 67.125 5.63 ;
        RECT 67.655 6.985 67.825 7.155 ;
        RECT 67.655 5.455 67.825 5.625 ;
        RECT 68.645 6.985 68.815 7.155 ;
        RECT 68.645 5.455 68.815 5.625 ;
        RECT 70.06 5.58 70.23 5.75 ;
        RECT 70.52 5.58 70.69 5.75 ;
        RECT 70.98 5.58 71.15 5.75 ;
        RECT 71.44 5.58 71.61 5.75 ;
        RECT 71.9 5.58 72.07 5.75 ;
        RECT 72.36 5.58 72.53 5.75 ;
        RECT 72.82 5.58 72.99 5.75 ;
        RECT 73.28 5.58 73.45 5.75 ;
        RECT 73.74 5.58 73.91 5.75 ;
        RECT 74.2 5.58 74.37 5.75 ;
        RECT 74.66 5.58 74.83 5.75 ;
        RECT 75.12 5.58 75.29 5.75 ;
        RECT 75.58 5.58 75.75 5.75 ;
        RECT 76.04 5.58 76.21 5.75 ;
        RECT 76.5 5.58 76.67 5.75 ;
        RECT 76.96 5.58 77.13 5.75 ;
        RECT 77.42 5.58 77.59 5.75 ;
        RECT 77.88 5.58 78.05 5.75 ;
        RECT 78.34 5.58 78.51 5.75 ;
        RECT 78.8 5.58 78.97 5.75 ;
        RECT 79.26 5.58 79.43 5.75 ;
        RECT 79.72 5.58 79.89 5.75 ;
        RECT 80.12 6.98 80.29 7.15 ;
        RECT 80.18 5.58 80.35 5.75 ;
        RECT 80.64 5.58 80.81 5.75 ;
        RECT 81.1 5.58 81.27 5.75 ;
        RECT 81.56 5.58 81.73 5.75 ;
        RECT 84.88 6.98 85.05 7.15 ;
        RECT 84.88 5.46 85.05 5.63 ;
        RECT 85.58 6.985 85.75 7.155 ;
        RECT 85.58 5.455 85.75 5.625 ;
        RECT 86.57 6.985 86.74 7.155 ;
        RECT 86.57 5.455 86.74 5.625 ;
        RECT 87.985 5.58 88.155 5.75 ;
        RECT 88.445 5.58 88.615 5.75 ;
        RECT 88.905 5.58 89.075 5.75 ;
        RECT 89.365 5.58 89.535 5.75 ;
        RECT 89.825 5.58 89.995 5.75 ;
        RECT 90.285 5.58 90.455 5.75 ;
        RECT 90.745 5.58 90.915 5.75 ;
        RECT 91.205 5.58 91.375 5.75 ;
        RECT 91.665 5.58 91.835 5.75 ;
        RECT 92.125 5.58 92.295 5.75 ;
        RECT 92.585 5.58 92.755 5.75 ;
        RECT 93.045 5.58 93.215 5.75 ;
        RECT 93.505 5.58 93.675 5.75 ;
        RECT 93.965 5.58 94.135 5.75 ;
        RECT 94.425 5.58 94.595 5.75 ;
        RECT 94.885 5.58 95.055 5.75 ;
        RECT 95.345 5.58 95.515 5.75 ;
        RECT 95.805 5.58 95.975 5.75 ;
        RECT 96.265 5.58 96.435 5.75 ;
        RECT 96.725 5.58 96.895 5.75 ;
        RECT 97.185 5.58 97.355 5.75 ;
        RECT 97.645 5.58 97.815 5.75 ;
        RECT 98.045 6.98 98.215 7.15 ;
        RECT 98.105 5.58 98.275 5.75 ;
        RECT 98.565 5.58 98.735 5.75 ;
        RECT 99.025 5.58 99.195 5.75 ;
        RECT 99.485 5.58 99.655 5.75 ;
        RECT 102.805 6.98 102.975 7.15 ;
        RECT 102.805 5.46 102.975 5.63 ;
        RECT 103.505 6.985 103.675 7.155 ;
        RECT 103.505 5.455 103.675 5.625 ;
        RECT 104.495 6.985 104.665 7.155 ;
        RECT 104.495 5.455 104.665 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 12.955 11.01 105.395 12.61 ;
        RECT 104.415 10.385 104.585 12.61 ;
        RECT 103.425 10.385 103.595 12.61 ;
        RECT 100.685 10.38 100.855 12.61 ;
        RECT 95.925 10.38 96.095 12.61 ;
        RECT 86.49 10.385 86.66 12.61 ;
        RECT 85.5 10.385 85.67 12.61 ;
        RECT 82.76 10.38 82.93 12.61 ;
        RECT 78 10.38 78.17 12.61 ;
        RECT 68.565 10.385 68.735 12.61 ;
        RECT 67.575 10.385 67.745 12.61 ;
        RECT 64.835 10.38 65.005 12.61 ;
        RECT 60.075 10.38 60.245 12.61 ;
        RECT 50.64 10.385 50.81 12.61 ;
        RECT 49.65 10.385 49.82 12.61 ;
        RECT 46.91 10.38 47.08 12.61 ;
        RECT 42.15 10.38 42.32 12.61 ;
        RECT 32.715 10.385 32.885 12.61 ;
        RECT 31.725 10.385 31.895 12.61 ;
        RECT 28.985 10.38 29.155 12.61 ;
        RECT 24.225 10.38 24.395 12.61 ;
        RECT 13.195 10.38 13.365 12.61 ;
        RECT 96.93 8.51 97.1 10.46 ;
        RECT 96.875 10.29 97.045 10.74 ;
        RECT 96.875 7.45 97.045 8.68 ;
        RECT 79.005 8.51 79.175 10.46 ;
        RECT 78.95 10.29 79.12 10.74 ;
        RECT 78.95 7.45 79.12 8.68 ;
        RECT 61.08 8.51 61.25 10.46 ;
        RECT 61.025 10.29 61.195 10.74 ;
        RECT 61.025 7.45 61.195 8.68 ;
        RECT 43.155 8.51 43.325 10.46 ;
        RECT 43.1 10.29 43.27 10.74 ;
        RECT 43.1 7.45 43.27 8.68 ;
        RECT 25.23 8.51 25.4 10.46 ;
        RECT 25.175 10.29 25.345 10.74 ;
        RECT 25.175 7.45 25.345 8.68 ;
      LAYER met1 ;
        RECT 12.955 11.01 105.395 12.61 ;
        RECT 96.87 8.72 97.16 8.95 ;
        RECT 96.535 8.75 97.16 8.92 ;
        RECT 96.535 8.75 96.705 12.61 ;
        RECT 78.945 8.72 79.235 8.95 ;
        RECT 78.61 8.75 79.235 8.92 ;
        RECT 78.61 8.75 78.78 12.61 ;
        RECT 61.02 8.72 61.31 8.95 ;
        RECT 60.685 8.75 61.31 8.92 ;
        RECT 60.685 8.75 60.855 12.61 ;
        RECT 43.095 8.72 43.385 8.95 ;
        RECT 42.76 8.75 43.385 8.92 ;
        RECT 42.76 8.75 42.93 12.61 ;
        RECT 25.17 8.72 25.46 8.95 ;
        RECT 24.835 8.75 25.46 8.92 ;
        RECT 24.835 8.75 25.005 12.61 ;
      LAYER mcon ;
        RECT 13.275 11.04 13.445 11.21 ;
        RECT 13.955 11.04 14.125 11.21 ;
        RECT 14.635 11.04 14.805 11.21 ;
        RECT 15.315 11.04 15.485 11.21 ;
        RECT 24.305 11.04 24.475 11.21 ;
        RECT 24.985 11.04 25.155 11.21 ;
        RECT 25.23 8.75 25.4 8.92 ;
        RECT 25.665 11.04 25.835 11.21 ;
        RECT 26.345 11.04 26.515 11.21 ;
        RECT 29.065 11.04 29.235 11.21 ;
        RECT 29.745 11.04 29.915 11.21 ;
        RECT 30.425 11.04 30.595 11.21 ;
        RECT 31.105 11.04 31.275 11.21 ;
        RECT 31.805 11.045 31.975 11.215 ;
        RECT 32.795 11.045 32.965 11.215 ;
        RECT 42.23 11.04 42.4 11.21 ;
        RECT 42.91 11.04 43.08 11.21 ;
        RECT 43.155 8.75 43.325 8.92 ;
        RECT 43.59 11.04 43.76 11.21 ;
        RECT 44.27 11.04 44.44 11.21 ;
        RECT 46.99 11.04 47.16 11.21 ;
        RECT 47.67 11.04 47.84 11.21 ;
        RECT 48.35 11.04 48.52 11.21 ;
        RECT 49.03 11.04 49.2 11.21 ;
        RECT 49.73 11.045 49.9 11.215 ;
        RECT 50.72 11.045 50.89 11.215 ;
        RECT 60.155 11.04 60.325 11.21 ;
        RECT 60.835 11.04 61.005 11.21 ;
        RECT 61.08 8.75 61.25 8.92 ;
        RECT 61.515 11.04 61.685 11.21 ;
        RECT 62.195 11.04 62.365 11.21 ;
        RECT 64.915 11.04 65.085 11.21 ;
        RECT 65.595 11.04 65.765 11.21 ;
        RECT 66.275 11.04 66.445 11.21 ;
        RECT 66.955 11.04 67.125 11.21 ;
        RECT 67.655 11.045 67.825 11.215 ;
        RECT 68.645 11.045 68.815 11.215 ;
        RECT 78.08 11.04 78.25 11.21 ;
        RECT 78.76 11.04 78.93 11.21 ;
        RECT 79.005 8.75 79.175 8.92 ;
        RECT 79.44 11.04 79.61 11.21 ;
        RECT 80.12 11.04 80.29 11.21 ;
        RECT 82.84 11.04 83.01 11.21 ;
        RECT 83.52 11.04 83.69 11.21 ;
        RECT 84.2 11.04 84.37 11.21 ;
        RECT 84.88 11.04 85.05 11.21 ;
        RECT 85.58 11.045 85.75 11.215 ;
        RECT 86.57 11.045 86.74 11.215 ;
        RECT 96.005 11.04 96.175 11.21 ;
        RECT 96.685 11.04 96.855 11.21 ;
        RECT 96.93 8.75 97.1 8.92 ;
        RECT 97.365 11.04 97.535 11.21 ;
        RECT 98.045 11.04 98.215 11.21 ;
        RECT 100.765 11.04 100.935 11.21 ;
        RECT 101.445 11.04 101.615 11.21 ;
        RECT 102.125 11.04 102.295 11.21 ;
        RECT 102.805 11.04 102.975 11.21 ;
        RECT 103.505 11.045 103.675 11.215 ;
        RECT 104.495 11.045 104.665 11.215 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 97.195 9.49 97.57 9.86 ;
      RECT 97.23 7.36 97.54 9.86 ;
      RECT 97.23 7.36 100.325 7.67 ;
      RECT 100.015 2.42 100.325 7.67 ;
      RECT 100.015 2.435 100.39 2.805 ;
      RECT 97.145 4.98 97.7 5.31 ;
      RECT 97.145 3.315 97.445 5.31 ;
      RECT 93.21 4.42 93.765 4.75 ;
      RECT 93.465 3.315 93.765 4.75 ;
      RECT 94.26 3.18 94.41 3.83 ;
      RECT 93.465 3.315 97.445 3.615 ;
      RECT 91.98 2.255 92.28 5.205 ;
      RECT 91.97 3.86 92.7 4.19 ;
      RECT 91.935 2.255 92.31 2.625 ;
      RECT 90.53 4.42 91.26 4.75 ;
      RECT 90.545 2.255 90.845 4.75 ;
      RECT 88.42 3.86 89.15 4.19 ;
      RECT 88.575 2.225 88.875 4.19 ;
      RECT 90.5 2.255 90.875 2.625 ;
      RECT 88.53 2.225 88.905 2.595 ;
      RECT 88.53 2.265 90.875 2.565 ;
      RECT 79.27 9.49 79.645 9.86 ;
      RECT 79.305 7.36 79.615 9.86 ;
      RECT 79.305 7.36 82.4 7.67 ;
      RECT 82.09 2.42 82.4 7.67 ;
      RECT 82.09 2.435 82.465 2.805 ;
      RECT 79.22 4.98 79.775 5.31 ;
      RECT 79.22 3.315 79.52 5.31 ;
      RECT 75.285 4.42 75.84 4.75 ;
      RECT 75.54 3.315 75.84 4.75 ;
      RECT 76.335 3.18 76.485 3.83 ;
      RECT 75.54 3.315 79.52 3.615 ;
      RECT 74.055 2.255 74.355 5.205 ;
      RECT 74.045 3.86 74.775 4.19 ;
      RECT 74.01 2.255 74.385 2.625 ;
      RECT 72.605 4.42 73.335 4.75 ;
      RECT 72.62 2.255 72.92 4.75 ;
      RECT 70.495 3.86 71.225 4.19 ;
      RECT 70.65 2.225 70.95 4.19 ;
      RECT 72.575 2.255 72.95 2.625 ;
      RECT 70.605 2.225 70.98 2.595 ;
      RECT 70.605 2.265 72.95 2.565 ;
      RECT 61.345 9.49 61.72 9.86 ;
      RECT 61.38 7.36 61.69 9.86 ;
      RECT 61.38 7.36 64.475 7.67 ;
      RECT 64.165 2.42 64.475 7.67 ;
      RECT 64.165 2.435 64.54 2.805 ;
      RECT 61.295 4.98 61.85 5.31 ;
      RECT 61.295 3.315 61.595 5.31 ;
      RECT 57.36 4.42 57.915 4.75 ;
      RECT 57.615 3.315 57.915 4.75 ;
      RECT 58.41 3.18 58.56 3.83 ;
      RECT 57.615 3.315 61.595 3.615 ;
      RECT 56.13 2.255 56.43 5.205 ;
      RECT 56.12 3.86 56.85 4.19 ;
      RECT 56.085 2.255 56.46 2.625 ;
      RECT 54.68 4.42 55.41 4.75 ;
      RECT 54.695 2.255 54.995 4.75 ;
      RECT 52.57 3.86 53.3 4.19 ;
      RECT 52.725 2.225 53.025 4.19 ;
      RECT 54.65 2.255 55.025 2.625 ;
      RECT 52.68 2.225 53.055 2.595 ;
      RECT 52.68 2.265 55.025 2.565 ;
      RECT 43.42 9.49 43.795 9.86 ;
      RECT 43.455 7.36 43.765 9.86 ;
      RECT 43.455 7.36 46.55 7.67 ;
      RECT 46.24 2.42 46.55 7.67 ;
      RECT 46.24 2.435 46.615 2.805 ;
      RECT 43.37 4.98 43.925 5.31 ;
      RECT 43.37 3.315 43.67 5.31 ;
      RECT 39.435 4.42 39.99 4.75 ;
      RECT 39.69 3.315 39.99 4.75 ;
      RECT 40.485 3.18 40.635 3.83 ;
      RECT 39.69 3.315 43.67 3.615 ;
      RECT 38.205 2.255 38.505 5.205 ;
      RECT 38.195 3.86 38.925 4.19 ;
      RECT 38.16 2.255 38.535 2.625 ;
      RECT 36.755 4.42 37.485 4.75 ;
      RECT 36.77 2.255 37.07 4.75 ;
      RECT 34.645 3.86 35.375 4.19 ;
      RECT 34.8 2.225 35.1 4.19 ;
      RECT 36.725 2.255 37.1 2.625 ;
      RECT 34.755 2.225 35.13 2.595 ;
      RECT 34.755 2.265 37.1 2.565 ;
      RECT 25.495 9.49 25.87 9.86 ;
      RECT 25.53 7.36 25.84 9.86 ;
      RECT 25.53 7.36 28.625 7.67 ;
      RECT 28.315 2.42 28.625 7.67 ;
      RECT 28.315 2.435 28.69 2.805 ;
      RECT 25.445 4.98 26 5.31 ;
      RECT 25.445 3.315 25.745 5.31 ;
      RECT 21.51 4.42 22.065 4.75 ;
      RECT 21.765 3.315 22.065 4.75 ;
      RECT 22.56 3.18 22.71 3.83 ;
      RECT 21.765 3.315 25.745 3.615 ;
      RECT 20.28 2.255 20.58 5.205 ;
      RECT 20.27 3.86 21 4.19 ;
      RECT 20.235 2.255 20.61 2.625 ;
      RECT 18.83 4.42 19.56 4.75 ;
      RECT 18.845 2.255 19.145 4.75 ;
      RECT 16.72 3.86 17.45 4.19 ;
      RECT 16.875 2.225 17.175 4.19 ;
      RECT 18.8 2.255 19.175 2.625 ;
      RECT 16.83 2.225 17.205 2.595 ;
      RECT 16.83 2.265 19.175 2.565 ;
      RECT 98.33 3.3 99.06 3.63 ;
      RECT 96.11 4.98 96.84 5.31 ;
      RECT 94.41 4.98 95.14 5.31 ;
      RECT 89.455 3.86 90.185 4.19 ;
      RECT 88.09 4.98 88.82 5.31 ;
      RECT 80.405 3.3 81.135 3.63 ;
      RECT 78.185 4.98 78.915 5.31 ;
      RECT 76.485 4.98 77.215 5.31 ;
      RECT 71.53 3.86 72.26 4.19 ;
      RECT 70.165 4.98 70.895 5.31 ;
      RECT 62.48 3.3 63.21 3.63 ;
      RECT 60.26 4.98 60.99 5.31 ;
      RECT 58.56 4.98 59.29 5.31 ;
      RECT 53.605 3.86 54.335 4.19 ;
      RECT 52.24 4.98 52.97 5.31 ;
      RECT 44.555 3.3 45.285 3.63 ;
      RECT 42.335 4.98 43.065 5.31 ;
      RECT 40.635 4.98 41.365 5.31 ;
      RECT 35.68 3.86 36.41 4.19 ;
      RECT 34.315 4.98 35.045 5.31 ;
      RECT 26.63 3.3 27.36 3.63 ;
      RECT 24.41 4.98 25.14 5.31 ;
      RECT 22.71 4.98 23.44 5.31 ;
      RECT 17.755 3.86 18.485 4.19 ;
      RECT 16.39 4.98 17.12 5.31 ;
    LAYER via2 ;
      RECT 100.105 2.52 100.305 2.72 ;
      RECT 98.395 3.365 98.595 3.565 ;
      RECT 97.435 5.045 97.635 5.245 ;
      RECT 97.285 9.575 97.485 9.775 ;
      RECT 96.435 5.045 96.635 5.245 ;
      RECT 94.475 5.045 94.675 5.245 ;
      RECT 93.275 4.485 93.475 4.685 ;
      RECT 92.035 3.925 92.235 4.125 ;
      RECT 92.025 2.34 92.225 2.54 ;
      RECT 90.595 4.485 90.795 4.685 ;
      RECT 90.59 2.335 90.79 2.535 ;
      RECT 89.855 3.925 90.055 4.125 ;
      RECT 88.635 3.925 88.835 4.125 ;
      RECT 88.62 2.31 88.82 2.51 ;
      RECT 88.155 5.045 88.355 5.245 ;
      RECT 82.18 2.52 82.38 2.72 ;
      RECT 80.47 3.365 80.67 3.565 ;
      RECT 79.51 5.045 79.71 5.245 ;
      RECT 79.36 9.575 79.56 9.775 ;
      RECT 78.51 5.045 78.71 5.245 ;
      RECT 76.55 5.045 76.75 5.245 ;
      RECT 75.35 4.485 75.55 4.685 ;
      RECT 74.11 3.925 74.31 4.125 ;
      RECT 74.1 2.34 74.3 2.54 ;
      RECT 72.67 4.485 72.87 4.685 ;
      RECT 72.665 2.335 72.865 2.535 ;
      RECT 71.93 3.925 72.13 4.125 ;
      RECT 70.71 3.925 70.91 4.125 ;
      RECT 70.695 2.31 70.895 2.51 ;
      RECT 70.23 5.045 70.43 5.245 ;
      RECT 64.255 2.52 64.455 2.72 ;
      RECT 62.545 3.365 62.745 3.565 ;
      RECT 61.585 5.045 61.785 5.245 ;
      RECT 61.435 9.575 61.635 9.775 ;
      RECT 60.585 5.045 60.785 5.245 ;
      RECT 58.625 5.045 58.825 5.245 ;
      RECT 57.425 4.485 57.625 4.685 ;
      RECT 56.185 3.925 56.385 4.125 ;
      RECT 56.175 2.34 56.375 2.54 ;
      RECT 54.745 4.485 54.945 4.685 ;
      RECT 54.74 2.335 54.94 2.535 ;
      RECT 54.005 3.925 54.205 4.125 ;
      RECT 52.785 3.925 52.985 4.125 ;
      RECT 52.77 2.31 52.97 2.51 ;
      RECT 52.305 5.045 52.505 5.245 ;
      RECT 46.33 2.52 46.53 2.72 ;
      RECT 44.62 3.365 44.82 3.565 ;
      RECT 43.66 5.045 43.86 5.245 ;
      RECT 43.51 9.575 43.71 9.775 ;
      RECT 42.66 5.045 42.86 5.245 ;
      RECT 40.7 5.045 40.9 5.245 ;
      RECT 39.5 4.485 39.7 4.685 ;
      RECT 38.26 3.925 38.46 4.125 ;
      RECT 38.25 2.34 38.45 2.54 ;
      RECT 36.82 4.485 37.02 4.685 ;
      RECT 36.815 2.335 37.015 2.535 ;
      RECT 36.08 3.925 36.28 4.125 ;
      RECT 34.86 3.925 35.06 4.125 ;
      RECT 34.845 2.31 35.045 2.51 ;
      RECT 34.38 5.045 34.58 5.245 ;
      RECT 28.405 2.52 28.605 2.72 ;
      RECT 26.695 3.365 26.895 3.565 ;
      RECT 25.735 5.045 25.935 5.245 ;
      RECT 25.585 9.575 25.785 9.775 ;
      RECT 24.735 5.045 24.935 5.245 ;
      RECT 22.775 5.045 22.975 5.245 ;
      RECT 21.575 4.485 21.775 4.685 ;
      RECT 20.335 3.925 20.535 4.125 ;
      RECT 20.325 2.34 20.525 2.54 ;
      RECT 18.895 4.485 19.095 4.685 ;
      RECT 18.89 2.335 19.09 2.535 ;
      RECT 18.155 3.925 18.355 4.125 ;
      RECT 16.935 3.925 17.135 4.125 ;
      RECT 16.92 2.31 17.12 2.51 ;
      RECT 16.455 5.045 16.655 5.245 ;
    LAYER met2 ;
      RECT 14.195 10.835 105.015 11.005 ;
      RECT 104.845 9.71 105.015 11.005 ;
      RECT 14.195 8.69 14.365 11.005 ;
      RECT 104.815 9.71 105.165 10.06 ;
      RECT 14.14 8.69 14.43 9.04 ;
      RECT 101.66 8.66 101.98 8.98 ;
      RECT 101.69 8.13 101.86 8.98 ;
      RECT 101.69 8.13 101.865 8.48 ;
      RECT 101.69 8.13 102.665 8.305 ;
      RECT 102.49 3.26 102.665 8.305 ;
      RECT 102.435 3.26 102.785 3.61 ;
      RECT 102.46 9.09 102.785 9.415 ;
      RECT 101.345 9.18 102.785 9.35 ;
      RECT 101.345 3.69 101.505 9.35 ;
      RECT 101.66 3.66 101.98 3.98 ;
      RECT 101.345 3.69 101.98 3.86 ;
      RECT 100.015 2.435 100.39 2.805 ;
      RECT 91.935 2.255 92.31 2.625 ;
      RECT 90.5 2.255 90.875 2.625 ;
      RECT 90.5 2.375 100.32 2.545 ;
      RECT 96.445 5.655 100.3 5.825 ;
      RECT 100.13 4.72 100.3 5.825 ;
      RECT 96.445 4.965 96.615 5.825 ;
      RECT 96.395 5.005 96.675 5.285 ;
      RECT 96.415 4.965 96.675 5.285 ;
      RECT 96.055 4.92 96.16 5.18 ;
      RECT 100.04 4.725 100.39 5.075 ;
      RECT 95.91 3.41 96 3.67 ;
      RECT 96.45 4.475 96.455 4.515 ;
      RECT 96.445 4.465 96.45 4.6 ;
      RECT 96.44 4.455 96.445 4.693 ;
      RECT 96.43 4.435 96.44 4.749 ;
      RECT 96.35 4.363 96.43 4.829 ;
      RECT 96.385 5.007 96.395 5.232 ;
      RECT 96.38 5.004 96.385 5.227 ;
      RECT 96.365 5.001 96.38 5.22 ;
      RECT 96.33 4.995 96.365 5.202 ;
      RECT 96.345 4.298 96.35 4.903 ;
      RECT 96.325 4.249 96.345 4.918 ;
      RECT 96.315 4.982 96.33 5.185 ;
      RECT 96.32 4.191 96.325 4.933 ;
      RECT 96.315 4.169 96.32 4.943 ;
      RECT 96.28 4.079 96.315 5.18 ;
      RECT 96.265 3.957 96.28 5.18 ;
      RECT 96.26 3.91 96.265 5.18 ;
      RECT 96.235 3.835 96.26 5.18 ;
      RECT 96.22 3.75 96.235 5.18 ;
      RECT 96.215 3.697 96.22 5.18 ;
      RECT 96.21 3.677 96.215 5.18 ;
      RECT 96.205 3.652 96.21 4.414 ;
      RECT 96.19 4.612 96.21 5.18 ;
      RECT 96.2 3.63 96.205 4.391 ;
      RECT 96.19 3.582 96.2 4.356 ;
      RECT 96.185 3.545 96.19 4.322 ;
      RECT 96.185 4.692 96.19 5.18 ;
      RECT 96.17 3.522 96.185 4.277 ;
      RECT 96.165 4.79 96.185 5.18 ;
      RECT 96.115 3.41 96.17 4.119 ;
      RECT 96.16 4.912 96.165 5.18 ;
      RECT 96.1 3.41 96.115 3.958 ;
      RECT 96.095 3.41 96.1 3.91 ;
      RECT 96.09 3.41 96.095 3.898 ;
      RECT 96.045 3.41 96.09 3.835 ;
      RECT 96.02 3.41 96.045 3.753 ;
      RECT 96.005 3.41 96.02 3.705 ;
      RECT 96 3.41 96.005 3.675 ;
      RECT 98.39 3.455 98.65 3.715 ;
      RECT 98.385 3.455 98.65 3.663 ;
      RECT 98.38 3.455 98.65 3.633 ;
      RECT 98.355 3.325 98.635 3.605 ;
      RECT 86.87 9.09 87.22 9.44 ;
      RECT 98.115 9.045 98.465 9.395 ;
      RECT 86.87 9.12 98.465 9.32 ;
      RECT 97.395 5.005 97.675 5.285 ;
      RECT 97.435 4.96 97.7 5.22 ;
      RECT 97.425 4.995 97.7 5.22 ;
      RECT 97.43 4.98 97.675 5.285 ;
      RECT 97.435 4.957 97.645 5.285 ;
      RECT 97.435 4.955 97.63 5.285 ;
      RECT 97.475 4.945 97.63 5.285 ;
      RECT 97.445 4.95 97.63 5.285 ;
      RECT 97.475 4.942 97.575 5.285 ;
      RECT 97.5 4.935 97.575 5.285 ;
      RECT 97.48 4.937 97.575 5.285 ;
      RECT 96.81 4.45 97.07 4.71 ;
      RECT 96.86 4.442 97.05 4.71 ;
      RECT 96.865 4.362 97.05 4.71 ;
      RECT 96.985 3.75 97.05 4.71 ;
      RECT 96.89 4.147 97.05 4.71 ;
      RECT 96.965 3.835 97.05 4.71 ;
      RECT 97 3.46 97.136 4.188 ;
      RECT 96.945 3.957 97.136 4.188 ;
      RECT 96.96 3.897 97.05 4.71 ;
      RECT 97 3.46 97.16 3.853 ;
      RECT 97 3.46 97.17 3.75 ;
      RECT 96.99 3.46 97.25 3.72 ;
      RECT 95.325 4.86 95.37 5.12 ;
      RECT 95.23 3.395 95.375 3.655 ;
      RECT 95.735 4.017 95.745 4.108 ;
      RECT 95.72 3.955 95.735 4.164 ;
      RECT 95.715 3.902 95.72 4.21 ;
      RECT 95.665 3.849 95.715 4.336 ;
      RECT 95.66 3.804 95.665 4.483 ;
      RECT 95.65 3.792 95.66 4.525 ;
      RECT 95.615 3.756 95.65 4.63 ;
      RECT 95.61 3.724 95.615 4.736 ;
      RECT 95.595 3.706 95.61 4.781 ;
      RECT 95.59 3.689 95.595 4.015 ;
      RECT 95.585 4.07 95.595 4.838 ;
      RECT 95.58 3.675 95.59 3.988 ;
      RECT 95.575 4.125 95.585 5.12 ;
      RECT 95.57 3.661 95.58 3.973 ;
      RECT 95.57 4.175 95.575 5.12 ;
      RECT 95.555 3.638 95.57 3.953 ;
      RECT 95.535 4.297 95.57 5.12 ;
      RECT 95.55 3.62 95.555 3.935 ;
      RECT 95.545 3.612 95.55 3.925 ;
      RECT 95.515 3.58 95.545 3.889 ;
      RECT 95.525 4.425 95.535 5.12 ;
      RECT 95.52 4.452 95.525 5.12 ;
      RECT 95.515 4.502 95.52 5.12 ;
      RECT 95.505 3.546 95.515 3.854 ;
      RECT 95.465 4.57 95.515 5.12 ;
      RECT 95.49 3.523 95.505 3.83 ;
      RECT 95.465 3.395 95.49 3.793 ;
      RECT 95.46 3.395 95.465 3.765 ;
      RECT 95.43 4.67 95.465 5.12 ;
      RECT 95.455 3.395 95.46 3.758 ;
      RECT 95.45 3.395 95.455 3.748 ;
      RECT 95.435 3.395 95.45 3.733 ;
      RECT 95.42 3.395 95.435 3.705 ;
      RECT 95.385 4.775 95.43 5.12 ;
      RECT 95.405 3.395 95.42 3.678 ;
      RECT 95.375 3.395 95.405 3.663 ;
      RECT 95.37 4.847 95.385 5.12 ;
      RECT 95.295 3.93 95.335 4.19 ;
      RECT 95.07 3.877 95.075 4.135 ;
      RECT 91.025 3.355 91.285 3.615 ;
      RECT 91.025 3.38 91.3 3.595 ;
      RECT 93.415 3.205 93.42 3.35 ;
      RECT 95.285 3.925 95.295 4.19 ;
      RECT 95.265 3.917 95.285 4.19 ;
      RECT 95.247 3.913 95.265 4.19 ;
      RECT 95.161 3.902 95.247 4.19 ;
      RECT 95.075 3.885 95.161 4.19 ;
      RECT 95.02 3.872 95.07 4.12 ;
      RECT 94.986 3.864 95.02 4.095 ;
      RECT 94.9 3.853 94.986 4.06 ;
      RECT 94.865 3.83 94.9 4.025 ;
      RECT 94.855 3.792 94.865 4.011 ;
      RECT 94.85 3.765 94.855 4.007 ;
      RECT 94.845 3.752 94.85 4.004 ;
      RECT 94.835 3.732 94.845 4 ;
      RECT 94.83 3.707 94.835 3.996 ;
      RECT 94.805 3.662 94.83 3.99 ;
      RECT 94.795 3.603 94.805 3.982 ;
      RECT 94.785 3.571 94.795 3.973 ;
      RECT 94.765 3.523 94.785 3.953 ;
      RECT 94.76 3.483 94.765 3.923 ;
      RECT 94.745 3.457 94.76 3.897 ;
      RECT 94.74 3.435 94.745 3.873 ;
      RECT 94.725 3.407 94.74 3.849 ;
      RECT 94.71 3.38 94.725 3.813 ;
      RECT 94.695 3.357 94.71 3.775 ;
      RECT 94.69 3.347 94.695 3.75 ;
      RECT 94.68 3.34 94.69 3.733 ;
      RECT 94.665 3.327 94.68 3.703 ;
      RECT 94.66 3.317 94.665 3.678 ;
      RECT 94.655 3.312 94.66 3.665 ;
      RECT 94.645 3.305 94.655 3.645 ;
      RECT 94.64 3.298 94.645 3.63 ;
      RECT 94.615 3.291 94.64 3.588 ;
      RECT 94.6 3.281 94.615 3.538 ;
      RECT 94.59 3.276 94.6 3.508 ;
      RECT 94.58 3.272 94.59 3.483 ;
      RECT 94.565 3.269 94.58 3.473 ;
      RECT 94.515 3.266 94.565 3.458 ;
      RECT 94.495 3.264 94.515 3.443 ;
      RECT 94.446 3.262 94.495 3.438 ;
      RECT 94.36 3.258 94.446 3.433 ;
      RECT 94.321 3.255 94.36 3.429 ;
      RECT 94.235 3.251 94.321 3.424 ;
      RECT 94.185 3.248 94.235 3.418 ;
      RECT 94.136 3.245 94.185 3.413 ;
      RECT 94.05 3.242 94.136 3.408 ;
      RECT 94.046 3.24 94.05 3.405 ;
      RECT 93.96 3.237 94.046 3.4 ;
      RECT 93.911 3.233 93.96 3.393 ;
      RECT 93.825 3.23 93.911 3.388 ;
      RECT 93.801 3.227 93.825 3.384 ;
      RECT 93.715 3.225 93.801 3.379 ;
      RECT 93.65 3.221 93.715 3.372 ;
      RECT 93.647 3.22 93.65 3.369 ;
      RECT 93.561 3.217 93.647 3.366 ;
      RECT 93.475 3.211 93.561 3.359 ;
      RECT 93.445 3.207 93.475 3.355 ;
      RECT 93.42 3.205 93.445 3.353 ;
      RECT 93.365 3.202 93.415 3.35 ;
      RECT 93.285 3.201 93.365 3.35 ;
      RECT 93.23 3.203 93.285 3.353 ;
      RECT 93.215 3.204 93.23 3.357 ;
      RECT 93.16 3.212 93.215 3.367 ;
      RECT 93.13 3.22 93.16 3.38 ;
      RECT 93.111 3.221 93.13 3.386 ;
      RECT 93.025 3.224 93.111 3.391 ;
      RECT 92.955 3.229 93.025 3.4 ;
      RECT 92.936 3.232 92.955 3.406 ;
      RECT 92.85 3.236 92.936 3.411 ;
      RECT 92.81 3.24 92.85 3.418 ;
      RECT 92.801 3.242 92.81 3.421 ;
      RECT 92.715 3.246 92.801 3.426 ;
      RECT 92.712 3.249 92.715 3.43 ;
      RECT 92.626 3.252 92.712 3.434 ;
      RECT 92.54 3.258 92.626 3.442 ;
      RECT 92.516 3.262 92.54 3.446 ;
      RECT 92.43 3.266 92.516 3.451 ;
      RECT 92.385 3.271 92.43 3.458 ;
      RECT 92.305 3.276 92.385 3.465 ;
      RECT 92.225 3.282 92.305 3.48 ;
      RECT 92.2 3.286 92.225 3.493 ;
      RECT 92.135 3.289 92.2 3.505 ;
      RECT 92.08 3.294 92.135 3.52 ;
      RECT 92.05 3.297 92.08 3.538 ;
      RECT 92.04 3.299 92.05 3.551 ;
      RECT 91.98 3.314 92.04 3.561 ;
      RECT 91.965 3.331 91.98 3.57 ;
      RECT 91.96 3.34 91.965 3.57 ;
      RECT 91.95 3.35 91.96 3.57 ;
      RECT 91.94 3.367 91.95 3.57 ;
      RECT 91.92 3.377 91.94 3.571 ;
      RECT 91.875 3.387 91.92 3.572 ;
      RECT 91.84 3.396 91.875 3.574 ;
      RECT 91.775 3.401 91.84 3.576 ;
      RECT 91.695 3.402 91.775 3.579 ;
      RECT 91.691 3.4 91.695 3.58 ;
      RECT 91.605 3.397 91.691 3.582 ;
      RECT 91.558 3.394 91.605 3.584 ;
      RECT 91.472 3.39 91.558 3.587 ;
      RECT 91.386 3.386 91.472 3.59 ;
      RECT 91.3 3.382 91.386 3.594 ;
      RECT 94.685 5.005 94.715 5.285 ;
      RECT 94.435 4.895 94.455 5.285 ;
      RECT 94.39 4.895 94.455 5.155 ;
      RECT 94.22 3.52 94.255 3.78 ;
      RECT 93.995 3.52 94.055 3.78 ;
      RECT 94.675 4.985 94.685 5.285 ;
      RECT 94.67 4.945 94.675 5.285 ;
      RECT 94.655 4.9 94.67 5.285 ;
      RECT 94.65 4.865 94.655 5.285 ;
      RECT 94.645 4.845 94.65 5.285 ;
      RECT 94.615 4.772 94.645 5.285 ;
      RECT 94.595 4.67 94.615 5.285 ;
      RECT 94.585 4.6 94.595 5.285 ;
      RECT 94.54 4.54 94.585 5.285 ;
      RECT 94.455 4.501 94.54 5.285 ;
      RECT 94.45 4.492 94.455 4.865 ;
      RECT 94.44 4.491 94.45 4.848 ;
      RECT 94.415 4.472 94.44 4.818 ;
      RECT 94.41 4.447 94.415 4.797 ;
      RECT 94.4 4.425 94.41 4.788 ;
      RECT 94.395 4.396 94.4 4.778 ;
      RECT 94.355 4.322 94.395 4.75 ;
      RECT 94.335 4.223 94.355 4.715 ;
      RECT 94.32 4.159 94.335 4.698 ;
      RECT 94.29 4.083 94.32 4.67 ;
      RECT 94.27 3.998 94.29 4.643 ;
      RECT 94.23 3.894 94.27 4.55 ;
      RECT 94.225 3.815 94.23 4.458 ;
      RECT 94.22 3.798 94.225 4.435 ;
      RECT 94.215 3.52 94.22 4.415 ;
      RECT 94.185 3.52 94.215 4.353 ;
      RECT 94.18 3.52 94.185 4.285 ;
      RECT 94.17 3.52 94.18 4.25 ;
      RECT 94.16 3.52 94.17 4.215 ;
      RECT 94.095 3.52 94.16 4.07 ;
      RECT 94.09 3.52 94.095 3.94 ;
      RECT 94.06 3.52 94.09 3.873 ;
      RECT 94.055 3.52 94.06 3.798 ;
      RECT 93.235 4.445 93.515 4.725 ;
      RECT 93.275 4.425 93.535 4.685 ;
      RECT 93.265 4.435 93.535 4.685 ;
      RECT 93.275 4.362 93.49 4.725 ;
      RECT 93.33 4.285 93.485 4.725 ;
      RECT 93.335 4.07 93.485 4.725 ;
      RECT 93.325 3.872 93.475 4.123 ;
      RECT 93.315 3.872 93.475 3.99 ;
      RECT 93.31 3.75 93.47 3.893 ;
      RECT 93.295 3.75 93.47 3.798 ;
      RECT 93.29 3.46 93.465 3.775 ;
      RECT 93.275 3.46 93.465 3.745 ;
      RECT 93.235 3.46 93.495 3.72 ;
      RECT 93.145 4.93 93.225 5.19 ;
      RECT 92.55 3.65 92.555 3.915 ;
      RECT 92.43 3.65 92.555 3.91 ;
      RECT 93.105 4.895 93.145 5.19 ;
      RECT 93.06 4.817 93.105 5.19 ;
      RECT 93.04 4.745 93.06 5.19 ;
      RECT 93.03 4.697 93.04 5.19 ;
      RECT 92.995 4.63 93.03 5.19 ;
      RECT 92.965 4.53 92.995 5.19 ;
      RECT 92.945 4.455 92.965 4.99 ;
      RECT 92.935 4.405 92.945 4.945 ;
      RECT 92.93 4.382 92.935 4.918 ;
      RECT 92.925 4.367 92.93 4.905 ;
      RECT 92.92 4.352 92.925 4.883 ;
      RECT 92.915 4.337 92.92 4.865 ;
      RECT 92.89 4.292 92.915 4.82 ;
      RECT 92.88 4.24 92.89 4.763 ;
      RECT 92.87 4.21 92.88 4.73 ;
      RECT 92.86 4.175 92.87 4.698 ;
      RECT 92.825 4.107 92.86 4.63 ;
      RECT 92.82 4.046 92.825 4.565 ;
      RECT 92.81 4.034 92.82 4.545 ;
      RECT 92.805 4.022 92.81 4.525 ;
      RECT 92.8 4.014 92.805 4.513 ;
      RECT 92.795 4.006 92.8 4.493 ;
      RECT 92.785 3.994 92.795 4.465 ;
      RECT 92.775 3.978 92.785 4.435 ;
      RECT 92.75 3.95 92.775 4.373 ;
      RECT 92.74 3.921 92.75 4.318 ;
      RECT 92.725 3.9 92.74 4.278 ;
      RECT 92.72 3.884 92.725 4.25 ;
      RECT 92.715 3.872 92.72 4.24 ;
      RECT 92.71 3.867 92.715 4.213 ;
      RECT 92.705 3.86 92.71 4.2 ;
      RECT 92.69 3.843 92.705 4.173 ;
      RECT 92.68 3.65 92.69 4.133 ;
      RECT 92.67 3.65 92.68 4.1 ;
      RECT 92.66 3.65 92.67 4.075 ;
      RECT 92.59 3.65 92.66 4.01 ;
      RECT 92.58 3.65 92.59 3.958 ;
      RECT 92.565 3.65 92.58 3.94 ;
      RECT 92.555 3.65 92.565 3.925 ;
      RECT 92.385 4.52 92.645 4.78 ;
      RECT 90.92 4.555 90.925 4.762 ;
      RECT 90.555 4.445 90.63 4.76 ;
      RECT 90.37 4.5 90.525 4.76 ;
      RECT 90.555 4.445 90.66 4.725 ;
      RECT 92.37 4.617 92.385 4.778 ;
      RECT 92.345 4.625 92.37 4.783 ;
      RECT 92.32 4.632 92.345 4.788 ;
      RECT 92.257 4.643 92.32 4.797 ;
      RECT 92.171 4.662 92.257 4.814 ;
      RECT 92.085 4.684 92.171 4.833 ;
      RECT 92.07 4.697 92.085 4.844 ;
      RECT 92.03 4.705 92.07 4.851 ;
      RECT 92.01 4.71 92.03 4.858 ;
      RECT 91.972 4.711 92.01 4.861 ;
      RECT 91.886 4.714 91.972 4.862 ;
      RECT 91.8 4.718 91.886 4.863 ;
      RECT 91.751 4.72 91.8 4.865 ;
      RECT 91.665 4.72 91.751 4.867 ;
      RECT 91.625 4.715 91.665 4.869 ;
      RECT 91.615 4.709 91.625 4.87 ;
      RECT 91.575 4.704 91.615 4.867 ;
      RECT 91.565 4.697 91.575 4.863 ;
      RECT 91.55 4.693 91.565 4.861 ;
      RECT 91.533 4.689 91.55 4.859 ;
      RECT 91.447 4.679 91.533 4.851 ;
      RECT 91.361 4.661 91.447 4.837 ;
      RECT 91.275 4.644 91.361 4.823 ;
      RECT 91.25 4.632 91.275 4.814 ;
      RECT 91.18 4.622 91.25 4.807 ;
      RECT 91.135 4.61 91.18 4.798 ;
      RECT 91.075 4.597 91.135 4.79 ;
      RECT 91.07 4.589 91.075 4.785 ;
      RECT 91.035 4.584 91.07 4.783 ;
      RECT 90.98 4.575 91.035 4.776 ;
      RECT 90.94 4.564 90.98 4.768 ;
      RECT 90.925 4.557 90.94 4.764 ;
      RECT 90.905 4.55 90.92 4.761 ;
      RECT 90.89 4.54 90.905 4.759 ;
      RECT 90.875 4.527 90.89 4.756 ;
      RECT 90.85 4.51 90.875 4.752 ;
      RECT 90.835 4.492 90.85 4.749 ;
      RECT 90.81 4.445 90.835 4.747 ;
      RECT 90.786 4.445 90.81 4.744 ;
      RECT 90.7 4.445 90.786 4.736 ;
      RECT 90.66 4.445 90.7 4.728 ;
      RECT 90.525 4.492 90.555 4.76 ;
      RECT 92.205 4.075 92.465 4.335 ;
      RECT 92.165 4.075 92.465 4.213 ;
      RECT 92.13 4.075 92.465 4.198 ;
      RECT 92.075 4.075 92.465 4.178 ;
      RECT 91.995 3.885 92.275 4.165 ;
      RECT 91.995 4.067 92.345 4.165 ;
      RECT 91.995 4.01 92.33 4.165 ;
      RECT 91.995 3.957 92.28 4.165 ;
      RECT 89.825 3.885 90.02 4.67 ;
      RECT 89.905 2.5 90.02 4.67 ;
      RECT 89.76 4.41 89.82 4.67 ;
      RECT 91.13 3.93 91.39 4.19 ;
      RECT 89.815 3.885 90.02 4.165 ;
      RECT 91.125 3.94 91.39 4.125 ;
      RECT 90.84 3.915 90.85 4.065 ;
      RECT 90.075 2.5 90.155 2.845 ;
      RECT 89.81 2.5 90.02 2.845 ;
      RECT 91.115 3.94 91.125 4.124 ;
      RECT 91.105 3.939 91.115 4.121 ;
      RECT 91.096 3.938 91.105 4.119 ;
      RECT 91.01 3.934 91.096 4.109 ;
      RECT 90.936 3.926 91.01 4.091 ;
      RECT 90.85 3.919 90.936 4.074 ;
      RECT 90.79 3.915 90.84 4.064 ;
      RECT 90.755 3.914 90.79 4.061 ;
      RECT 90.7 3.914 90.755 4.063 ;
      RECT 90.665 3.914 90.7 4.067 ;
      RECT 90.579 3.913 90.665 4.074 ;
      RECT 90.493 3.912 90.579 4.084 ;
      RECT 90.407 3.911 90.493 4.095 ;
      RECT 90.321 3.911 90.407 4.105 ;
      RECT 90.235 3.91 90.321 4.115 ;
      RECT 90.2 3.91 90.235 4.155 ;
      RECT 90.195 3.91 90.2 4.198 ;
      RECT 90.17 3.91 90.195 4.215 ;
      RECT 90.095 3.91 90.17 4.23 ;
      RECT 90.075 3.885 90.095 4.243 ;
      RECT 90.07 2.5 90.075 4.253 ;
      RECT 90.045 2.5 90.07 4.295 ;
      RECT 90.02 2.5 90.045 4.373 ;
      RECT 89.82 4.292 89.825 4.67 ;
      RECT 89.155 4.244 89.17 4.7 ;
      RECT 89.15 4.316 89.256 4.698 ;
      RECT 89.17 3.41 89.305 4.696 ;
      RECT 89.155 4.26 89.31 4.695 ;
      RECT 89.155 4.31 89.315 4.693 ;
      RECT 89.14 4.375 89.315 4.692 ;
      RECT 89.15 4.367 89.32 4.689 ;
      RECT 89.13 4.415 89.32 4.684 ;
      RECT 89.13 4.415 89.335 4.681 ;
      RECT 89.125 4.415 89.335 4.678 ;
      RECT 89.1 4.415 89.36 4.675 ;
      RECT 89.17 3.41 89.33 4.063 ;
      RECT 89.165 3.41 89.33 4.035 ;
      RECT 89.16 3.41 89.33 3.863 ;
      RECT 89.16 3.41 89.35 3.803 ;
      RECT 89.115 3.41 89.375 3.67 ;
      RECT 88.595 3.885 88.875 4.165 ;
      RECT 88.585 3.9 88.875 4.16 ;
      RECT 88.54 3.962 88.875 4.158 ;
      RECT 88.615 3.877 88.78 4.165 ;
      RECT 88.615 3.862 88.736 4.165 ;
      RECT 88.65 3.855 88.736 4.165 ;
      RECT 88.115 5.005 88.395 5.285 ;
      RECT 88.075 4.967 88.37 5.078 ;
      RECT 88.06 4.917 88.35 4.973 ;
      RECT 88.005 4.68 88.265 4.94 ;
      RECT 88.005 4.882 88.345 4.94 ;
      RECT 88.005 4.822 88.34 4.94 ;
      RECT 88.005 4.772 88.32 4.94 ;
      RECT 88.005 4.752 88.315 4.94 ;
      RECT 88.005 4.73 88.31 4.94 ;
      RECT 88.005 4.715 88.28 4.94 ;
      RECT 83.735 8.66 84.055 8.98 ;
      RECT 83.765 8.13 83.935 8.98 ;
      RECT 83.765 8.13 83.94 8.48 ;
      RECT 83.765 8.13 84.74 8.305 ;
      RECT 84.565 3.26 84.74 8.305 ;
      RECT 84.51 3.26 84.86 3.61 ;
      RECT 84.535 9.09 84.86 9.415 ;
      RECT 83.42 9.18 84.86 9.35 ;
      RECT 83.42 3.69 83.58 9.35 ;
      RECT 83.735 3.66 84.055 3.98 ;
      RECT 83.42 3.69 84.055 3.86 ;
      RECT 82.09 2.435 82.465 2.805 ;
      RECT 74.01 2.255 74.385 2.625 ;
      RECT 72.575 2.255 72.95 2.625 ;
      RECT 72.575 2.375 82.395 2.545 ;
      RECT 78.52 5.655 82.375 5.825 ;
      RECT 82.205 4.72 82.375 5.825 ;
      RECT 78.52 4.965 78.69 5.825 ;
      RECT 78.47 5.005 78.75 5.285 ;
      RECT 78.49 4.965 78.75 5.285 ;
      RECT 78.13 4.92 78.235 5.18 ;
      RECT 82.115 4.725 82.465 5.075 ;
      RECT 77.985 3.41 78.075 3.67 ;
      RECT 78.525 4.475 78.53 4.515 ;
      RECT 78.52 4.465 78.525 4.6 ;
      RECT 78.515 4.455 78.52 4.693 ;
      RECT 78.505 4.435 78.515 4.749 ;
      RECT 78.425 4.363 78.505 4.829 ;
      RECT 78.46 5.007 78.47 5.232 ;
      RECT 78.455 5.004 78.46 5.227 ;
      RECT 78.44 5.001 78.455 5.22 ;
      RECT 78.405 4.995 78.44 5.202 ;
      RECT 78.42 4.298 78.425 4.903 ;
      RECT 78.4 4.249 78.42 4.918 ;
      RECT 78.39 4.982 78.405 5.185 ;
      RECT 78.395 4.191 78.4 4.933 ;
      RECT 78.39 4.169 78.395 4.943 ;
      RECT 78.355 4.079 78.39 5.18 ;
      RECT 78.34 3.957 78.355 5.18 ;
      RECT 78.335 3.91 78.34 5.18 ;
      RECT 78.31 3.835 78.335 5.18 ;
      RECT 78.295 3.75 78.31 5.18 ;
      RECT 78.29 3.697 78.295 5.18 ;
      RECT 78.285 3.677 78.29 5.18 ;
      RECT 78.28 3.652 78.285 4.414 ;
      RECT 78.265 4.612 78.285 5.18 ;
      RECT 78.275 3.63 78.28 4.391 ;
      RECT 78.265 3.582 78.275 4.356 ;
      RECT 78.26 3.545 78.265 4.322 ;
      RECT 78.26 4.692 78.265 5.18 ;
      RECT 78.245 3.522 78.26 4.277 ;
      RECT 78.24 4.79 78.26 5.18 ;
      RECT 78.19 3.41 78.245 4.119 ;
      RECT 78.235 4.912 78.24 5.18 ;
      RECT 78.175 3.41 78.19 3.958 ;
      RECT 78.17 3.41 78.175 3.91 ;
      RECT 78.165 3.41 78.17 3.898 ;
      RECT 78.12 3.41 78.165 3.835 ;
      RECT 78.095 3.41 78.12 3.753 ;
      RECT 78.08 3.41 78.095 3.705 ;
      RECT 78.075 3.41 78.08 3.675 ;
      RECT 80.465 3.455 80.725 3.715 ;
      RECT 80.46 3.455 80.725 3.663 ;
      RECT 80.455 3.455 80.725 3.633 ;
      RECT 80.43 3.325 80.71 3.605 ;
      RECT 68.945 9.09 69.295 9.44 ;
      RECT 79.91 9.045 80.26 9.395 ;
      RECT 68.945 9.12 80.26 9.32 ;
      RECT 79.47 5.005 79.75 5.285 ;
      RECT 79.51 4.96 79.775 5.22 ;
      RECT 79.5 4.995 79.775 5.22 ;
      RECT 79.505 4.98 79.75 5.285 ;
      RECT 79.51 4.957 79.72 5.285 ;
      RECT 79.51 4.955 79.705 5.285 ;
      RECT 79.55 4.945 79.705 5.285 ;
      RECT 79.52 4.95 79.705 5.285 ;
      RECT 79.55 4.942 79.65 5.285 ;
      RECT 79.575 4.935 79.65 5.285 ;
      RECT 79.555 4.937 79.65 5.285 ;
      RECT 78.885 4.45 79.145 4.71 ;
      RECT 78.935 4.442 79.125 4.71 ;
      RECT 78.94 4.362 79.125 4.71 ;
      RECT 79.06 3.75 79.125 4.71 ;
      RECT 78.965 4.147 79.125 4.71 ;
      RECT 79.04 3.835 79.125 4.71 ;
      RECT 79.075 3.46 79.211 4.188 ;
      RECT 79.02 3.957 79.211 4.188 ;
      RECT 79.035 3.897 79.125 4.71 ;
      RECT 79.075 3.46 79.235 3.853 ;
      RECT 79.075 3.46 79.245 3.75 ;
      RECT 79.065 3.46 79.325 3.72 ;
      RECT 77.4 4.86 77.445 5.12 ;
      RECT 77.305 3.395 77.45 3.655 ;
      RECT 77.81 4.017 77.82 4.108 ;
      RECT 77.795 3.955 77.81 4.164 ;
      RECT 77.79 3.902 77.795 4.21 ;
      RECT 77.74 3.849 77.79 4.336 ;
      RECT 77.735 3.804 77.74 4.483 ;
      RECT 77.725 3.792 77.735 4.525 ;
      RECT 77.69 3.756 77.725 4.63 ;
      RECT 77.685 3.724 77.69 4.736 ;
      RECT 77.67 3.706 77.685 4.781 ;
      RECT 77.665 3.689 77.67 4.015 ;
      RECT 77.66 4.07 77.67 4.838 ;
      RECT 77.655 3.675 77.665 3.988 ;
      RECT 77.65 4.125 77.66 5.12 ;
      RECT 77.645 3.661 77.655 3.973 ;
      RECT 77.645 4.175 77.65 5.12 ;
      RECT 77.63 3.638 77.645 3.953 ;
      RECT 77.61 4.297 77.645 5.12 ;
      RECT 77.625 3.62 77.63 3.935 ;
      RECT 77.62 3.612 77.625 3.925 ;
      RECT 77.59 3.58 77.62 3.889 ;
      RECT 77.6 4.425 77.61 5.12 ;
      RECT 77.595 4.452 77.6 5.12 ;
      RECT 77.59 4.502 77.595 5.12 ;
      RECT 77.58 3.546 77.59 3.854 ;
      RECT 77.54 4.57 77.59 5.12 ;
      RECT 77.565 3.523 77.58 3.83 ;
      RECT 77.54 3.395 77.565 3.793 ;
      RECT 77.535 3.395 77.54 3.765 ;
      RECT 77.505 4.67 77.54 5.12 ;
      RECT 77.53 3.395 77.535 3.758 ;
      RECT 77.525 3.395 77.53 3.748 ;
      RECT 77.51 3.395 77.525 3.733 ;
      RECT 77.495 3.395 77.51 3.705 ;
      RECT 77.46 4.775 77.505 5.12 ;
      RECT 77.48 3.395 77.495 3.678 ;
      RECT 77.45 3.395 77.48 3.663 ;
      RECT 77.445 4.847 77.46 5.12 ;
      RECT 77.37 3.93 77.41 4.19 ;
      RECT 77.145 3.877 77.15 4.135 ;
      RECT 73.1 3.355 73.36 3.615 ;
      RECT 73.1 3.38 73.375 3.595 ;
      RECT 75.49 3.205 75.495 3.35 ;
      RECT 77.36 3.925 77.37 4.19 ;
      RECT 77.34 3.917 77.36 4.19 ;
      RECT 77.322 3.913 77.34 4.19 ;
      RECT 77.236 3.902 77.322 4.19 ;
      RECT 77.15 3.885 77.236 4.19 ;
      RECT 77.095 3.872 77.145 4.12 ;
      RECT 77.061 3.864 77.095 4.095 ;
      RECT 76.975 3.853 77.061 4.06 ;
      RECT 76.94 3.83 76.975 4.025 ;
      RECT 76.93 3.792 76.94 4.011 ;
      RECT 76.925 3.765 76.93 4.007 ;
      RECT 76.92 3.752 76.925 4.004 ;
      RECT 76.91 3.732 76.92 4 ;
      RECT 76.905 3.707 76.91 3.996 ;
      RECT 76.88 3.662 76.905 3.99 ;
      RECT 76.87 3.603 76.88 3.982 ;
      RECT 76.86 3.571 76.87 3.973 ;
      RECT 76.84 3.523 76.86 3.953 ;
      RECT 76.835 3.483 76.84 3.923 ;
      RECT 76.82 3.457 76.835 3.897 ;
      RECT 76.815 3.435 76.82 3.873 ;
      RECT 76.8 3.407 76.815 3.849 ;
      RECT 76.785 3.38 76.8 3.813 ;
      RECT 76.77 3.357 76.785 3.775 ;
      RECT 76.765 3.347 76.77 3.75 ;
      RECT 76.755 3.34 76.765 3.733 ;
      RECT 76.74 3.327 76.755 3.703 ;
      RECT 76.735 3.317 76.74 3.678 ;
      RECT 76.73 3.312 76.735 3.665 ;
      RECT 76.72 3.305 76.73 3.645 ;
      RECT 76.715 3.298 76.72 3.63 ;
      RECT 76.69 3.291 76.715 3.588 ;
      RECT 76.675 3.281 76.69 3.538 ;
      RECT 76.665 3.276 76.675 3.508 ;
      RECT 76.655 3.272 76.665 3.483 ;
      RECT 76.64 3.269 76.655 3.473 ;
      RECT 76.59 3.266 76.64 3.458 ;
      RECT 76.57 3.264 76.59 3.443 ;
      RECT 76.521 3.262 76.57 3.438 ;
      RECT 76.435 3.258 76.521 3.433 ;
      RECT 76.396 3.255 76.435 3.429 ;
      RECT 76.31 3.251 76.396 3.424 ;
      RECT 76.26 3.248 76.31 3.418 ;
      RECT 76.211 3.245 76.26 3.413 ;
      RECT 76.125 3.242 76.211 3.408 ;
      RECT 76.121 3.24 76.125 3.405 ;
      RECT 76.035 3.237 76.121 3.4 ;
      RECT 75.986 3.233 76.035 3.393 ;
      RECT 75.9 3.23 75.986 3.388 ;
      RECT 75.876 3.227 75.9 3.384 ;
      RECT 75.79 3.225 75.876 3.379 ;
      RECT 75.725 3.221 75.79 3.372 ;
      RECT 75.722 3.22 75.725 3.369 ;
      RECT 75.636 3.217 75.722 3.366 ;
      RECT 75.55 3.211 75.636 3.359 ;
      RECT 75.52 3.207 75.55 3.355 ;
      RECT 75.495 3.205 75.52 3.353 ;
      RECT 75.44 3.202 75.49 3.35 ;
      RECT 75.36 3.201 75.44 3.35 ;
      RECT 75.305 3.203 75.36 3.353 ;
      RECT 75.29 3.204 75.305 3.357 ;
      RECT 75.235 3.212 75.29 3.367 ;
      RECT 75.205 3.22 75.235 3.38 ;
      RECT 75.186 3.221 75.205 3.386 ;
      RECT 75.1 3.224 75.186 3.391 ;
      RECT 75.03 3.229 75.1 3.4 ;
      RECT 75.011 3.232 75.03 3.406 ;
      RECT 74.925 3.236 75.011 3.411 ;
      RECT 74.885 3.24 74.925 3.418 ;
      RECT 74.876 3.242 74.885 3.421 ;
      RECT 74.79 3.246 74.876 3.426 ;
      RECT 74.787 3.249 74.79 3.43 ;
      RECT 74.701 3.252 74.787 3.434 ;
      RECT 74.615 3.258 74.701 3.442 ;
      RECT 74.591 3.262 74.615 3.446 ;
      RECT 74.505 3.266 74.591 3.451 ;
      RECT 74.46 3.271 74.505 3.458 ;
      RECT 74.38 3.276 74.46 3.465 ;
      RECT 74.3 3.282 74.38 3.48 ;
      RECT 74.275 3.286 74.3 3.493 ;
      RECT 74.21 3.289 74.275 3.505 ;
      RECT 74.155 3.294 74.21 3.52 ;
      RECT 74.125 3.297 74.155 3.538 ;
      RECT 74.115 3.299 74.125 3.551 ;
      RECT 74.055 3.314 74.115 3.561 ;
      RECT 74.04 3.331 74.055 3.57 ;
      RECT 74.035 3.34 74.04 3.57 ;
      RECT 74.025 3.35 74.035 3.57 ;
      RECT 74.015 3.367 74.025 3.57 ;
      RECT 73.995 3.377 74.015 3.571 ;
      RECT 73.95 3.387 73.995 3.572 ;
      RECT 73.915 3.396 73.95 3.574 ;
      RECT 73.85 3.401 73.915 3.576 ;
      RECT 73.77 3.402 73.85 3.579 ;
      RECT 73.766 3.4 73.77 3.58 ;
      RECT 73.68 3.397 73.766 3.582 ;
      RECT 73.633 3.394 73.68 3.584 ;
      RECT 73.547 3.39 73.633 3.587 ;
      RECT 73.461 3.386 73.547 3.59 ;
      RECT 73.375 3.382 73.461 3.594 ;
      RECT 76.76 5.005 76.79 5.285 ;
      RECT 76.51 4.895 76.53 5.285 ;
      RECT 76.465 4.895 76.53 5.155 ;
      RECT 76.295 3.52 76.33 3.78 ;
      RECT 76.07 3.52 76.13 3.78 ;
      RECT 76.75 4.985 76.76 5.285 ;
      RECT 76.745 4.945 76.75 5.285 ;
      RECT 76.73 4.9 76.745 5.285 ;
      RECT 76.725 4.865 76.73 5.285 ;
      RECT 76.72 4.845 76.725 5.285 ;
      RECT 76.69 4.772 76.72 5.285 ;
      RECT 76.67 4.67 76.69 5.285 ;
      RECT 76.66 4.6 76.67 5.285 ;
      RECT 76.615 4.54 76.66 5.285 ;
      RECT 76.53 4.501 76.615 5.285 ;
      RECT 76.525 4.492 76.53 4.865 ;
      RECT 76.515 4.491 76.525 4.848 ;
      RECT 76.49 4.472 76.515 4.818 ;
      RECT 76.485 4.447 76.49 4.797 ;
      RECT 76.475 4.425 76.485 4.788 ;
      RECT 76.47 4.396 76.475 4.778 ;
      RECT 76.43 4.322 76.47 4.75 ;
      RECT 76.41 4.223 76.43 4.715 ;
      RECT 76.395 4.159 76.41 4.698 ;
      RECT 76.365 4.083 76.395 4.67 ;
      RECT 76.345 3.998 76.365 4.643 ;
      RECT 76.305 3.894 76.345 4.55 ;
      RECT 76.3 3.815 76.305 4.458 ;
      RECT 76.295 3.798 76.3 4.435 ;
      RECT 76.29 3.52 76.295 4.415 ;
      RECT 76.26 3.52 76.29 4.353 ;
      RECT 76.255 3.52 76.26 4.285 ;
      RECT 76.245 3.52 76.255 4.25 ;
      RECT 76.235 3.52 76.245 4.215 ;
      RECT 76.17 3.52 76.235 4.07 ;
      RECT 76.165 3.52 76.17 3.94 ;
      RECT 76.135 3.52 76.165 3.873 ;
      RECT 76.13 3.52 76.135 3.798 ;
      RECT 75.31 4.445 75.59 4.725 ;
      RECT 75.35 4.425 75.61 4.685 ;
      RECT 75.34 4.435 75.61 4.685 ;
      RECT 75.35 4.362 75.565 4.725 ;
      RECT 75.405 4.285 75.56 4.725 ;
      RECT 75.41 4.07 75.56 4.725 ;
      RECT 75.4 3.872 75.55 4.123 ;
      RECT 75.39 3.872 75.55 3.99 ;
      RECT 75.385 3.75 75.545 3.893 ;
      RECT 75.37 3.75 75.545 3.798 ;
      RECT 75.365 3.46 75.54 3.775 ;
      RECT 75.35 3.46 75.54 3.745 ;
      RECT 75.31 3.46 75.57 3.72 ;
      RECT 75.22 4.93 75.3 5.19 ;
      RECT 74.625 3.65 74.63 3.915 ;
      RECT 74.505 3.65 74.63 3.91 ;
      RECT 75.18 4.895 75.22 5.19 ;
      RECT 75.135 4.817 75.18 5.19 ;
      RECT 75.115 4.745 75.135 5.19 ;
      RECT 75.105 4.697 75.115 5.19 ;
      RECT 75.07 4.63 75.105 5.19 ;
      RECT 75.04 4.53 75.07 5.19 ;
      RECT 75.02 4.455 75.04 4.99 ;
      RECT 75.01 4.405 75.02 4.945 ;
      RECT 75.005 4.382 75.01 4.918 ;
      RECT 75 4.367 75.005 4.905 ;
      RECT 74.995 4.352 75 4.883 ;
      RECT 74.99 4.337 74.995 4.865 ;
      RECT 74.965 4.292 74.99 4.82 ;
      RECT 74.955 4.24 74.965 4.763 ;
      RECT 74.945 4.21 74.955 4.73 ;
      RECT 74.935 4.175 74.945 4.698 ;
      RECT 74.9 4.107 74.935 4.63 ;
      RECT 74.895 4.046 74.9 4.565 ;
      RECT 74.885 4.034 74.895 4.545 ;
      RECT 74.88 4.022 74.885 4.525 ;
      RECT 74.875 4.014 74.88 4.513 ;
      RECT 74.87 4.006 74.875 4.493 ;
      RECT 74.86 3.994 74.87 4.465 ;
      RECT 74.85 3.978 74.86 4.435 ;
      RECT 74.825 3.95 74.85 4.373 ;
      RECT 74.815 3.921 74.825 4.318 ;
      RECT 74.8 3.9 74.815 4.278 ;
      RECT 74.795 3.884 74.8 4.25 ;
      RECT 74.79 3.872 74.795 4.24 ;
      RECT 74.785 3.867 74.79 4.213 ;
      RECT 74.78 3.86 74.785 4.2 ;
      RECT 74.765 3.843 74.78 4.173 ;
      RECT 74.755 3.65 74.765 4.133 ;
      RECT 74.745 3.65 74.755 4.1 ;
      RECT 74.735 3.65 74.745 4.075 ;
      RECT 74.665 3.65 74.735 4.01 ;
      RECT 74.655 3.65 74.665 3.958 ;
      RECT 74.64 3.65 74.655 3.94 ;
      RECT 74.63 3.65 74.64 3.925 ;
      RECT 74.46 4.52 74.72 4.78 ;
      RECT 72.995 4.555 73 4.762 ;
      RECT 72.63 4.445 72.705 4.76 ;
      RECT 72.445 4.5 72.6 4.76 ;
      RECT 72.63 4.445 72.735 4.725 ;
      RECT 74.445 4.617 74.46 4.778 ;
      RECT 74.42 4.625 74.445 4.783 ;
      RECT 74.395 4.632 74.42 4.788 ;
      RECT 74.332 4.643 74.395 4.797 ;
      RECT 74.246 4.662 74.332 4.814 ;
      RECT 74.16 4.684 74.246 4.833 ;
      RECT 74.145 4.697 74.16 4.844 ;
      RECT 74.105 4.705 74.145 4.851 ;
      RECT 74.085 4.71 74.105 4.858 ;
      RECT 74.047 4.711 74.085 4.861 ;
      RECT 73.961 4.714 74.047 4.862 ;
      RECT 73.875 4.718 73.961 4.863 ;
      RECT 73.826 4.72 73.875 4.865 ;
      RECT 73.74 4.72 73.826 4.867 ;
      RECT 73.7 4.715 73.74 4.869 ;
      RECT 73.69 4.709 73.7 4.87 ;
      RECT 73.65 4.704 73.69 4.867 ;
      RECT 73.64 4.697 73.65 4.863 ;
      RECT 73.625 4.693 73.64 4.861 ;
      RECT 73.608 4.689 73.625 4.859 ;
      RECT 73.522 4.679 73.608 4.851 ;
      RECT 73.436 4.661 73.522 4.837 ;
      RECT 73.35 4.644 73.436 4.823 ;
      RECT 73.325 4.632 73.35 4.814 ;
      RECT 73.255 4.622 73.325 4.807 ;
      RECT 73.21 4.61 73.255 4.798 ;
      RECT 73.15 4.597 73.21 4.79 ;
      RECT 73.145 4.589 73.15 4.785 ;
      RECT 73.11 4.584 73.145 4.783 ;
      RECT 73.055 4.575 73.11 4.776 ;
      RECT 73.015 4.564 73.055 4.768 ;
      RECT 73 4.557 73.015 4.764 ;
      RECT 72.98 4.55 72.995 4.761 ;
      RECT 72.965 4.54 72.98 4.759 ;
      RECT 72.95 4.527 72.965 4.756 ;
      RECT 72.925 4.51 72.95 4.752 ;
      RECT 72.91 4.492 72.925 4.749 ;
      RECT 72.885 4.445 72.91 4.747 ;
      RECT 72.861 4.445 72.885 4.744 ;
      RECT 72.775 4.445 72.861 4.736 ;
      RECT 72.735 4.445 72.775 4.728 ;
      RECT 72.6 4.492 72.63 4.76 ;
      RECT 74.28 4.075 74.54 4.335 ;
      RECT 74.24 4.075 74.54 4.213 ;
      RECT 74.205 4.075 74.54 4.198 ;
      RECT 74.15 4.075 74.54 4.178 ;
      RECT 74.07 3.885 74.35 4.165 ;
      RECT 74.07 4.067 74.42 4.165 ;
      RECT 74.07 4.01 74.405 4.165 ;
      RECT 74.07 3.957 74.355 4.165 ;
      RECT 71.9 3.885 72.095 4.67 ;
      RECT 71.98 2.5 72.095 4.67 ;
      RECT 71.835 4.41 71.895 4.67 ;
      RECT 73.205 3.93 73.465 4.19 ;
      RECT 71.89 3.885 72.095 4.165 ;
      RECT 73.2 3.94 73.465 4.125 ;
      RECT 72.915 3.915 72.925 4.065 ;
      RECT 72.15 2.5 72.23 2.845 ;
      RECT 71.885 2.5 72.095 2.845 ;
      RECT 73.19 3.94 73.2 4.124 ;
      RECT 73.18 3.939 73.19 4.121 ;
      RECT 73.171 3.938 73.18 4.119 ;
      RECT 73.085 3.934 73.171 4.109 ;
      RECT 73.011 3.926 73.085 4.091 ;
      RECT 72.925 3.919 73.011 4.074 ;
      RECT 72.865 3.915 72.915 4.064 ;
      RECT 72.83 3.914 72.865 4.061 ;
      RECT 72.775 3.914 72.83 4.063 ;
      RECT 72.74 3.914 72.775 4.067 ;
      RECT 72.654 3.913 72.74 4.074 ;
      RECT 72.568 3.912 72.654 4.084 ;
      RECT 72.482 3.911 72.568 4.095 ;
      RECT 72.396 3.911 72.482 4.105 ;
      RECT 72.31 3.91 72.396 4.115 ;
      RECT 72.275 3.91 72.31 4.155 ;
      RECT 72.27 3.91 72.275 4.198 ;
      RECT 72.245 3.91 72.27 4.215 ;
      RECT 72.17 3.91 72.245 4.23 ;
      RECT 72.15 3.885 72.17 4.243 ;
      RECT 72.145 2.5 72.15 4.253 ;
      RECT 72.12 2.5 72.145 4.295 ;
      RECT 72.095 2.5 72.12 4.373 ;
      RECT 71.895 4.292 71.9 4.67 ;
      RECT 71.23 4.244 71.245 4.7 ;
      RECT 71.225 4.316 71.331 4.698 ;
      RECT 71.245 3.41 71.38 4.696 ;
      RECT 71.23 4.26 71.385 4.695 ;
      RECT 71.23 4.31 71.39 4.693 ;
      RECT 71.215 4.375 71.39 4.692 ;
      RECT 71.225 4.367 71.395 4.689 ;
      RECT 71.205 4.415 71.395 4.684 ;
      RECT 71.205 4.415 71.41 4.681 ;
      RECT 71.2 4.415 71.41 4.678 ;
      RECT 71.175 4.415 71.435 4.675 ;
      RECT 71.245 3.41 71.405 4.063 ;
      RECT 71.24 3.41 71.405 4.035 ;
      RECT 71.235 3.41 71.405 3.863 ;
      RECT 71.235 3.41 71.425 3.803 ;
      RECT 71.19 3.41 71.45 3.67 ;
      RECT 70.67 3.885 70.95 4.165 ;
      RECT 70.66 3.9 70.95 4.16 ;
      RECT 70.615 3.962 70.95 4.158 ;
      RECT 70.69 3.877 70.855 4.165 ;
      RECT 70.69 3.862 70.811 4.165 ;
      RECT 70.725 3.855 70.811 4.165 ;
      RECT 70.19 5.005 70.47 5.285 ;
      RECT 70.15 4.967 70.445 5.078 ;
      RECT 70.135 4.917 70.425 4.973 ;
      RECT 70.08 4.68 70.34 4.94 ;
      RECT 70.08 4.882 70.42 4.94 ;
      RECT 70.08 4.822 70.415 4.94 ;
      RECT 70.08 4.772 70.395 4.94 ;
      RECT 70.08 4.752 70.39 4.94 ;
      RECT 70.08 4.73 70.385 4.94 ;
      RECT 70.08 4.715 70.355 4.94 ;
      RECT 65.81 8.66 66.13 8.98 ;
      RECT 65.84 8.13 66.01 8.98 ;
      RECT 65.84 8.13 66.015 8.48 ;
      RECT 65.84 8.13 66.815 8.305 ;
      RECT 66.64 3.26 66.815 8.305 ;
      RECT 66.585 3.26 66.935 3.61 ;
      RECT 66.61 9.09 66.935 9.415 ;
      RECT 65.495 9.18 66.935 9.35 ;
      RECT 65.495 3.69 65.655 9.35 ;
      RECT 65.81 3.66 66.13 3.98 ;
      RECT 65.495 3.69 66.13 3.86 ;
      RECT 64.165 2.435 64.54 2.805 ;
      RECT 56.085 2.255 56.46 2.625 ;
      RECT 54.65 2.255 55.025 2.625 ;
      RECT 54.65 2.375 64.47 2.545 ;
      RECT 60.595 5.655 64.45 5.825 ;
      RECT 64.28 4.72 64.45 5.825 ;
      RECT 60.595 4.965 60.765 5.825 ;
      RECT 60.545 5.005 60.825 5.285 ;
      RECT 60.565 4.965 60.825 5.285 ;
      RECT 60.205 4.92 60.31 5.18 ;
      RECT 64.19 4.725 64.54 5.075 ;
      RECT 60.06 3.41 60.15 3.67 ;
      RECT 60.6 4.475 60.605 4.515 ;
      RECT 60.595 4.465 60.6 4.6 ;
      RECT 60.59 4.455 60.595 4.693 ;
      RECT 60.58 4.435 60.59 4.749 ;
      RECT 60.5 4.363 60.58 4.829 ;
      RECT 60.535 5.007 60.545 5.232 ;
      RECT 60.53 5.004 60.535 5.227 ;
      RECT 60.515 5.001 60.53 5.22 ;
      RECT 60.48 4.995 60.515 5.202 ;
      RECT 60.495 4.298 60.5 4.903 ;
      RECT 60.475 4.249 60.495 4.918 ;
      RECT 60.465 4.982 60.48 5.185 ;
      RECT 60.47 4.191 60.475 4.933 ;
      RECT 60.465 4.169 60.47 4.943 ;
      RECT 60.43 4.079 60.465 5.18 ;
      RECT 60.415 3.957 60.43 5.18 ;
      RECT 60.41 3.91 60.415 5.18 ;
      RECT 60.385 3.835 60.41 5.18 ;
      RECT 60.37 3.75 60.385 5.18 ;
      RECT 60.365 3.697 60.37 5.18 ;
      RECT 60.36 3.677 60.365 5.18 ;
      RECT 60.355 3.652 60.36 4.414 ;
      RECT 60.34 4.612 60.36 5.18 ;
      RECT 60.35 3.63 60.355 4.391 ;
      RECT 60.34 3.582 60.35 4.356 ;
      RECT 60.335 3.545 60.34 4.322 ;
      RECT 60.335 4.692 60.34 5.18 ;
      RECT 60.32 3.522 60.335 4.277 ;
      RECT 60.315 4.79 60.335 5.18 ;
      RECT 60.265 3.41 60.32 4.119 ;
      RECT 60.31 4.912 60.315 5.18 ;
      RECT 60.25 3.41 60.265 3.958 ;
      RECT 60.245 3.41 60.25 3.91 ;
      RECT 60.24 3.41 60.245 3.898 ;
      RECT 60.195 3.41 60.24 3.835 ;
      RECT 60.17 3.41 60.195 3.753 ;
      RECT 60.155 3.41 60.17 3.705 ;
      RECT 60.15 3.41 60.155 3.675 ;
      RECT 62.54 3.455 62.8 3.715 ;
      RECT 62.535 3.455 62.8 3.663 ;
      RECT 62.53 3.455 62.8 3.633 ;
      RECT 62.505 3.325 62.785 3.605 ;
      RECT 51.065 9.095 51.415 9.445 ;
      RECT 62.04 9.05 62.39 9.4 ;
      RECT 51.065 9.125 62.39 9.325 ;
      RECT 61.545 5.005 61.825 5.285 ;
      RECT 61.585 4.96 61.85 5.22 ;
      RECT 61.575 4.995 61.85 5.22 ;
      RECT 61.58 4.98 61.825 5.285 ;
      RECT 61.585 4.957 61.795 5.285 ;
      RECT 61.585 4.955 61.78 5.285 ;
      RECT 61.625 4.945 61.78 5.285 ;
      RECT 61.595 4.95 61.78 5.285 ;
      RECT 61.625 4.942 61.725 5.285 ;
      RECT 61.65 4.935 61.725 5.285 ;
      RECT 61.63 4.937 61.725 5.285 ;
      RECT 60.96 4.45 61.22 4.71 ;
      RECT 61.01 4.442 61.2 4.71 ;
      RECT 61.015 4.362 61.2 4.71 ;
      RECT 61.135 3.75 61.2 4.71 ;
      RECT 61.04 4.147 61.2 4.71 ;
      RECT 61.115 3.835 61.2 4.71 ;
      RECT 61.15 3.46 61.286 4.188 ;
      RECT 61.095 3.957 61.286 4.188 ;
      RECT 61.11 3.897 61.2 4.71 ;
      RECT 61.15 3.46 61.31 3.853 ;
      RECT 61.15 3.46 61.32 3.75 ;
      RECT 61.14 3.46 61.4 3.72 ;
      RECT 59.475 4.86 59.52 5.12 ;
      RECT 59.38 3.395 59.525 3.655 ;
      RECT 59.885 4.017 59.895 4.108 ;
      RECT 59.87 3.955 59.885 4.164 ;
      RECT 59.865 3.902 59.87 4.21 ;
      RECT 59.815 3.849 59.865 4.336 ;
      RECT 59.81 3.804 59.815 4.483 ;
      RECT 59.8 3.792 59.81 4.525 ;
      RECT 59.765 3.756 59.8 4.63 ;
      RECT 59.76 3.724 59.765 4.736 ;
      RECT 59.745 3.706 59.76 4.781 ;
      RECT 59.74 3.689 59.745 4.015 ;
      RECT 59.735 4.07 59.745 4.838 ;
      RECT 59.73 3.675 59.74 3.988 ;
      RECT 59.725 4.125 59.735 5.12 ;
      RECT 59.72 3.661 59.73 3.973 ;
      RECT 59.72 4.175 59.725 5.12 ;
      RECT 59.705 3.638 59.72 3.953 ;
      RECT 59.685 4.297 59.72 5.12 ;
      RECT 59.7 3.62 59.705 3.935 ;
      RECT 59.695 3.612 59.7 3.925 ;
      RECT 59.665 3.58 59.695 3.889 ;
      RECT 59.675 4.425 59.685 5.12 ;
      RECT 59.67 4.452 59.675 5.12 ;
      RECT 59.665 4.502 59.67 5.12 ;
      RECT 59.655 3.546 59.665 3.854 ;
      RECT 59.615 4.57 59.665 5.12 ;
      RECT 59.64 3.523 59.655 3.83 ;
      RECT 59.615 3.395 59.64 3.793 ;
      RECT 59.61 3.395 59.615 3.765 ;
      RECT 59.58 4.67 59.615 5.12 ;
      RECT 59.605 3.395 59.61 3.758 ;
      RECT 59.6 3.395 59.605 3.748 ;
      RECT 59.585 3.395 59.6 3.733 ;
      RECT 59.57 3.395 59.585 3.705 ;
      RECT 59.535 4.775 59.58 5.12 ;
      RECT 59.555 3.395 59.57 3.678 ;
      RECT 59.525 3.395 59.555 3.663 ;
      RECT 59.52 4.847 59.535 5.12 ;
      RECT 59.445 3.93 59.485 4.19 ;
      RECT 59.22 3.877 59.225 4.135 ;
      RECT 55.175 3.355 55.435 3.615 ;
      RECT 55.175 3.38 55.45 3.595 ;
      RECT 57.565 3.205 57.57 3.35 ;
      RECT 59.435 3.925 59.445 4.19 ;
      RECT 59.415 3.917 59.435 4.19 ;
      RECT 59.397 3.913 59.415 4.19 ;
      RECT 59.311 3.902 59.397 4.19 ;
      RECT 59.225 3.885 59.311 4.19 ;
      RECT 59.17 3.872 59.22 4.12 ;
      RECT 59.136 3.864 59.17 4.095 ;
      RECT 59.05 3.853 59.136 4.06 ;
      RECT 59.015 3.83 59.05 4.025 ;
      RECT 59.005 3.792 59.015 4.011 ;
      RECT 59 3.765 59.005 4.007 ;
      RECT 58.995 3.752 59 4.004 ;
      RECT 58.985 3.732 58.995 4 ;
      RECT 58.98 3.707 58.985 3.996 ;
      RECT 58.955 3.662 58.98 3.99 ;
      RECT 58.945 3.603 58.955 3.982 ;
      RECT 58.935 3.571 58.945 3.973 ;
      RECT 58.915 3.523 58.935 3.953 ;
      RECT 58.91 3.483 58.915 3.923 ;
      RECT 58.895 3.457 58.91 3.897 ;
      RECT 58.89 3.435 58.895 3.873 ;
      RECT 58.875 3.407 58.89 3.849 ;
      RECT 58.86 3.38 58.875 3.813 ;
      RECT 58.845 3.357 58.86 3.775 ;
      RECT 58.84 3.347 58.845 3.75 ;
      RECT 58.83 3.34 58.84 3.733 ;
      RECT 58.815 3.327 58.83 3.703 ;
      RECT 58.81 3.317 58.815 3.678 ;
      RECT 58.805 3.312 58.81 3.665 ;
      RECT 58.795 3.305 58.805 3.645 ;
      RECT 58.79 3.298 58.795 3.63 ;
      RECT 58.765 3.291 58.79 3.588 ;
      RECT 58.75 3.281 58.765 3.538 ;
      RECT 58.74 3.276 58.75 3.508 ;
      RECT 58.73 3.272 58.74 3.483 ;
      RECT 58.715 3.269 58.73 3.473 ;
      RECT 58.665 3.266 58.715 3.458 ;
      RECT 58.645 3.264 58.665 3.443 ;
      RECT 58.596 3.262 58.645 3.438 ;
      RECT 58.51 3.258 58.596 3.433 ;
      RECT 58.471 3.255 58.51 3.429 ;
      RECT 58.385 3.251 58.471 3.424 ;
      RECT 58.335 3.248 58.385 3.418 ;
      RECT 58.286 3.245 58.335 3.413 ;
      RECT 58.2 3.242 58.286 3.408 ;
      RECT 58.196 3.24 58.2 3.405 ;
      RECT 58.11 3.237 58.196 3.4 ;
      RECT 58.061 3.233 58.11 3.393 ;
      RECT 57.975 3.23 58.061 3.388 ;
      RECT 57.951 3.227 57.975 3.384 ;
      RECT 57.865 3.225 57.951 3.379 ;
      RECT 57.8 3.221 57.865 3.372 ;
      RECT 57.797 3.22 57.8 3.369 ;
      RECT 57.711 3.217 57.797 3.366 ;
      RECT 57.625 3.211 57.711 3.359 ;
      RECT 57.595 3.207 57.625 3.355 ;
      RECT 57.57 3.205 57.595 3.353 ;
      RECT 57.515 3.202 57.565 3.35 ;
      RECT 57.435 3.201 57.515 3.35 ;
      RECT 57.38 3.203 57.435 3.353 ;
      RECT 57.365 3.204 57.38 3.357 ;
      RECT 57.31 3.212 57.365 3.367 ;
      RECT 57.28 3.22 57.31 3.38 ;
      RECT 57.261 3.221 57.28 3.386 ;
      RECT 57.175 3.224 57.261 3.391 ;
      RECT 57.105 3.229 57.175 3.4 ;
      RECT 57.086 3.232 57.105 3.406 ;
      RECT 57 3.236 57.086 3.411 ;
      RECT 56.96 3.24 57 3.418 ;
      RECT 56.951 3.242 56.96 3.421 ;
      RECT 56.865 3.246 56.951 3.426 ;
      RECT 56.862 3.249 56.865 3.43 ;
      RECT 56.776 3.252 56.862 3.434 ;
      RECT 56.69 3.258 56.776 3.442 ;
      RECT 56.666 3.262 56.69 3.446 ;
      RECT 56.58 3.266 56.666 3.451 ;
      RECT 56.535 3.271 56.58 3.458 ;
      RECT 56.455 3.276 56.535 3.465 ;
      RECT 56.375 3.282 56.455 3.48 ;
      RECT 56.35 3.286 56.375 3.493 ;
      RECT 56.285 3.289 56.35 3.505 ;
      RECT 56.23 3.294 56.285 3.52 ;
      RECT 56.2 3.297 56.23 3.538 ;
      RECT 56.19 3.299 56.2 3.551 ;
      RECT 56.13 3.314 56.19 3.561 ;
      RECT 56.115 3.331 56.13 3.57 ;
      RECT 56.11 3.34 56.115 3.57 ;
      RECT 56.1 3.35 56.11 3.57 ;
      RECT 56.09 3.367 56.1 3.57 ;
      RECT 56.07 3.377 56.09 3.571 ;
      RECT 56.025 3.387 56.07 3.572 ;
      RECT 55.99 3.396 56.025 3.574 ;
      RECT 55.925 3.401 55.99 3.576 ;
      RECT 55.845 3.402 55.925 3.579 ;
      RECT 55.841 3.4 55.845 3.58 ;
      RECT 55.755 3.397 55.841 3.582 ;
      RECT 55.708 3.394 55.755 3.584 ;
      RECT 55.622 3.39 55.708 3.587 ;
      RECT 55.536 3.386 55.622 3.59 ;
      RECT 55.45 3.382 55.536 3.594 ;
      RECT 58.835 5.005 58.865 5.285 ;
      RECT 58.585 4.895 58.605 5.285 ;
      RECT 58.54 4.895 58.605 5.155 ;
      RECT 58.37 3.52 58.405 3.78 ;
      RECT 58.145 3.52 58.205 3.78 ;
      RECT 58.825 4.985 58.835 5.285 ;
      RECT 58.82 4.945 58.825 5.285 ;
      RECT 58.805 4.9 58.82 5.285 ;
      RECT 58.8 4.865 58.805 5.285 ;
      RECT 58.795 4.845 58.8 5.285 ;
      RECT 58.765 4.772 58.795 5.285 ;
      RECT 58.745 4.67 58.765 5.285 ;
      RECT 58.735 4.6 58.745 5.285 ;
      RECT 58.69 4.54 58.735 5.285 ;
      RECT 58.605 4.501 58.69 5.285 ;
      RECT 58.6 4.492 58.605 4.865 ;
      RECT 58.59 4.491 58.6 4.848 ;
      RECT 58.565 4.472 58.59 4.818 ;
      RECT 58.56 4.447 58.565 4.797 ;
      RECT 58.55 4.425 58.56 4.788 ;
      RECT 58.545 4.396 58.55 4.778 ;
      RECT 58.505 4.322 58.545 4.75 ;
      RECT 58.485 4.223 58.505 4.715 ;
      RECT 58.47 4.159 58.485 4.698 ;
      RECT 58.44 4.083 58.47 4.67 ;
      RECT 58.42 3.998 58.44 4.643 ;
      RECT 58.38 3.894 58.42 4.55 ;
      RECT 58.375 3.815 58.38 4.458 ;
      RECT 58.37 3.798 58.375 4.435 ;
      RECT 58.365 3.52 58.37 4.415 ;
      RECT 58.335 3.52 58.365 4.353 ;
      RECT 58.33 3.52 58.335 4.285 ;
      RECT 58.32 3.52 58.33 4.25 ;
      RECT 58.31 3.52 58.32 4.215 ;
      RECT 58.245 3.52 58.31 4.07 ;
      RECT 58.24 3.52 58.245 3.94 ;
      RECT 58.21 3.52 58.24 3.873 ;
      RECT 58.205 3.52 58.21 3.798 ;
      RECT 57.385 4.445 57.665 4.725 ;
      RECT 57.425 4.425 57.685 4.685 ;
      RECT 57.415 4.435 57.685 4.685 ;
      RECT 57.425 4.362 57.64 4.725 ;
      RECT 57.48 4.285 57.635 4.725 ;
      RECT 57.485 4.07 57.635 4.725 ;
      RECT 57.475 3.872 57.625 4.123 ;
      RECT 57.465 3.872 57.625 3.99 ;
      RECT 57.46 3.75 57.62 3.893 ;
      RECT 57.445 3.75 57.62 3.798 ;
      RECT 57.44 3.46 57.615 3.775 ;
      RECT 57.425 3.46 57.615 3.745 ;
      RECT 57.385 3.46 57.645 3.72 ;
      RECT 57.295 4.93 57.375 5.19 ;
      RECT 56.7 3.65 56.705 3.915 ;
      RECT 56.58 3.65 56.705 3.91 ;
      RECT 57.255 4.895 57.295 5.19 ;
      RECT 57.21 4.817 57.255 5.19 ;
      RECT 57.19 4.745 57.21 5.19 ;
      RECT 57.18 4.697 57.19 5.19 ;
      RECT 57.145 4.63 57.18 5.19 ;
      RECT 57.115 4.53 57.145 5.19 ;
      RECT 57.095 4.455 57.115 4.99 ;
      RECT 57.085 4.405 57.095 4.945 ;
      RECT 57.08 4.382 57.085 4.918 ;
      RECT 57.075 4.367 57.08 4.905 ;
      RECT 57.07 4.352 57.075 4.883 ;
      RECT 57.065 4.337 57.07 4.865 ;
      RECT 57.04 4.292 57.065 4.82 ;
      RECT 57.03 4.24 57.04 4.763 ;
      RECT 57.02 4.21 57.03 4.73 ;
      RECT 57.01 4.175 57.02 4.698 ;
      RECT 56.975 4.107 57.01 4.63 ;
      RECT 56.97 4.046 56.975 4.565 ;
      RECT 56.96 4.034 56.97 4.545 ;
      RECT 56.955 4.022 56.96 4.525 ;
      RECT 56.95 4.014 56.955 4.513 ;
      RECT 56.945 4.006 56.95 4.493 ;
      RECT 56.935 3.994 56.945 4.465 ;
      RECT 56.925 3.978 56.935 4.435 ;
      RECT 56.9 3.95 56.925 4.373 ;
      RECT 56.89 3.921 56.9 4.318 ;
      RECT 56.875 3.9 56.89 4.278 ;
      RECT 56.87 3.884 56.875 4.25 ;
      RECT 56.865 3.872 56.87 4.24 ;
      RECT 56.86 3.867 56.865 4.213 ;
      RECT 56.855 3.86 56.86 4.2 ;
      RECT 56.84 3.843 56.855 4.173 ;
      RECT 56.83 3.65 56.84 4.133 ;
      RECT 56.82 3.65 56.83 4.1 ;
      RECT 56.81 3.65 56.82 4.075 ;
      RECT 56.74 3.65 56.81 4.01 ;
      RECT 56.73 3.65 56.74 3.958 ;
      RECT 56.715 3.65 56.73 3.94 ;
      RECT 56.705 3.65 56.715 3.925 ;
      RECT 56.535 4.52 56.795 4.78 ;
      RECT 55.07 4.555 55.075 4.762 ;
      RECT 54.705 4.445 54.78 4.76 ;
      RECT 54.52 4.5 54.675 4.76 ;
      RECT 54.705 4.445 54.81 4.725 ;
      RECT 56.52 4.617 56.535 4.778 ;
      RECT 56.495 4.625 56.52 4.783 ;
      RECT 56.47 4.632 56.495 4.788 ;
      RECT 56.407 4.643 56.47 4.797 ;
      RECT 56.321 4.662 56.407 4.814 ;
      RECT 56.235 4.684 56.321 4.833 ;
      RECT 56.22 4.697 56.235 4.844 ;
      RECT 56.18 4.705 56.22 4.851 ;
      RECT 56.16 4.71 56.18 4.858 ;
      RECT 56.122 4.711 56.16 4.861 ;
      RECT 56.036 4.714 56.122 4.862 ;
      RECT 55.95 4.718 56.036 4.863 ;
      RECT 55.901 4.72 55.95 4.865 ;
      RECT 55.815 4.72 55.901 4.867 ;
      RECT 55.775 4.715 55.815 4.869 ;
      RECT 55.765 4.709 55.775 4.87 ;
      RECT 55.725 4.704 55.765 4.867 ;
      RECT 55.715 4.697 55.725 4.863 ;
      RECT 55.7 4.693 55.715 4.861 ;
      RECT 55.683 4.689 55.7 4.859 ;
      RECT 55.597 4.679 55.683 4.851 ;
      RECT 55.511 4.661 55.597 4.837 ;
      RECT 55.425 4.644 55.511 4.823 ;
      RECT 55.4 4.632 55.425 4.814 ;
      RECT 55.33 4.622 55.4 4.807 ;
      RECT 55.285 4.61 55.33 4.798 ;
      RECT 55.225 4.597 55.285 4.79 ;
      RECT 55.22 4.589 55.225 4.785 ;
      RECT 55.185 4.584 55.22 4.783 ;
      RECT 55.13 4.575 55.185 4.776 ;
      RECT 55.09 4.564 55.13 4.768 ;
      RECT 55.075 4.557 55.09 4.764 ;
      RECT 55.055 4.55 55.07 4.761 ;
      RECT 55.04 4.54 55.055 4.759 ;
      RECT 55.025 4.527 55.04 4.756 ;
      RECT 55 4.51 55.025 4.752 ;
      RECT 54.985 4.492 55 4.749 ;
      RECT 54.96 4.445 54.985 4.747 ;
      RECT 54.936 4.445 54.96 4.744 ;
      RECT 54.85 4.445 54.936 4.736 ;
      RECT 54.81 4.445 54.85 4.728 ;
      RECT 54.675 4.492 54.705 4.76 ;
      RECT 56.355 4.075 56.615 4.335 ;
      RECT 56.315 4.075 56.615 4.213 ;
      RECT 56.28 4.075 56.615 4.198 ;
      RECT 56.225 4.075 56.615 4.178 ;
      RECT 56.145 3.885 56.425 4.165 ;
      RECT 56.145 4.067 56.495 4.165 ;
      RECT 56.145 4.01 56.48 4.165 ;
      RECT 56.145 3.957 56.43 4.165 ;
      RECT 53.975 3.885 54.17 4.67 ;
      RECT 54.055 2.5 54.17 4.67 ;
      RECT 53.91 4.41 53.97 4.67 ;
      RECT 55.28 3.93 55.54 4.19 ;
      RECT 53.965 3.885 54.17 4.165 ;
      RECT 55.275 3.94 55.54 4.125 ;
      RECT 54.99 3.915 55 4.065 ;
      RECT 54.225 2.5 54.305 2.845 ;
      RECT 53.96 2.5 54.17 2.845 ;
      RECT 55.265 3.94 55.275 4.124 ;
      RECT 55.255 3.939 55.265 4.121 ;
      RECT 55.246 3.938 55.255 4.119 ;
      RECT 55.16 3.934 55.246 4.109 ;
      RECT 55.086 3.926 55.16 4.091 ;
      RECT 55 3.919 55.086 4.074 ;
      RECT 54.94 3.915 54.99 4.064 ;
      RECT 54.905 3.914 54.94 4.061 ;
      RECT 54.85 3.914 54.905 4.063 ;
      RECT 54.815 3.914 54.85 4.067 ;
      RECT 54.729 3.913 54.815 4.074 ;
      RECT 54.643 3.912 54.729 4.084 ;
      RECT 54.557 3.911 54.643 4.095 ;
      RECT 54.471 3.911 54.557 4.105 ;
      RECT 54.385 3.91 54.471 4.115 ;
      RECT 54.35 3.91 54.385 4.155 ;
      RECT 54.345 3.91 54.35 4.198 ;
      RECT 54.32 3.91 54.345 4.215 ;
      RECT 54.245 3.91 54.32 4.23 ;
      RECT 54.225 3.885 54.245 4.243 ;
      RECT 54.22 2.5 54.225 4.253 ;
      RECT 54.195 2.5 54.22 4.295 ;
      RECT 54.17 2.5 54.195 4.373 ;
      RECT 53.97 4.292 53.975 4.67 ;
      RECT 53.305 4.244 53.32 4.7 ;
      RECT 53.3 4.316 53.406 4.698 ;
      RECT 53.32 3.41 53.455 4.696 ;
      RECT 53.305 4.26 53.46 4.695 ;
      RECT 53.305 4.31 53.465 4.693 ;
      RECT 53.29 4.375 53.465 4.692 ;
      RECT 53.3 4.367 53.47 4.689 ;
      RECT 53.28 4.415 53.47 4.684 ;
      RECT 53.28 4.415 53.485 4.681 ;
      RECT 53.275 4.415 53.485 4.678 ;
      RECT 53.25 4.415 53.51 4.675 ;
      RECT 53.32 3.41 53.48 4.063 ;
      RECT 53.315 3.41 53.48 4.035 ;
      RECT 53.31 3.41 53.48 3.863 ;
      RECT 53.31 3.41 53.5 3.803 ;
      RECT 53.265 3.41 53.525 3.67 ;
      RECT 52.745 3.885 53.025 4.165 ;
      RECT 52.735 3.9 53.025 4.16 ;
      RECT 52.69 3.962 53.025 4.158 ;
      RECT 52.765 3.877 52.93 4.165 ;
      RECT 52.765 3.862 52.886 4.165 ;
      RECT 52.8 3.855 52.886 4.165 ;
      RECT 52.265 5.005 52.545 5.285 ;
      RECT 52.225 4.967 52.52 5.078 ;
      RECT 52.21 4.917 52.5 4.973 ;
      RECT 52.155 4.68 52.415 4.94 ;
      RECT 52.155 4.882 52.495 4.94 ;
      RECT 52.155 4.822 52.49 4.94 ;
      RECT 52.155 4.772 52.47 4.94 ;
      RECT 52.155 4.752 52.465 4.94 ;
      RECT 52.155 4.73 52.46 4.94 ;
      RECT 52.155 4.715 52.43 4.94 ;
      RECT 47.885 8.66 48.205 8.98 ;
      RECT 47.915 8.13 48.085 8.98 ;
      RECT 47.915 8.13 48.09 8.48 ;
      RECT 47.915 8.13 48.89 8.305 ;
      RECT 48.715 3.26 48.89 8.305 ;
      RECT 48.66 3.26 49.01 3.61 ;
      RECT 48.685 9.09 49.01 9.415 ;
      RECT 47.57 9.18 49.01 9.35 ;
      RECT 47.57 3.69 47.73 9.35 ;
      RECT 47.885 3.66 48.205 3.98 ;
      RECT 47.57 3.69 48.205 3.86 ;
      RECT 46.24 2.435 46.615 2.805 ;
      RECT 38.16 2.255 38.535 2.625 ;
      RECT 36.725 2.255 37.1 2.625 ;
      RECT 36.725 2.375 46.545 2.545 ;
      RECT 42.67 5.655 46.525 5.825 ;
      RECT 46.355 4.72 46.525 5.825 ;
      RECT 42.67 4.965 42.84 5.825 ;
      RECT 42.62 5.005 42.9 5.285 ;
      RECT 42.64 4.965 42.9 5.285 ;
      RECT 42.28 4.92 42.385 5.18 ;
      RECT 46.265 4.725 46.615 5.075 ;
      RECT 42.135 3.41 42.225 3.67 ;
      RECT 42.675 4.475 42.68 4.515 ;
      RECT 42.67 4.465 42.675 4.6 ;
      RECT 42.665 4.455 42.67 4.693 ;
      RECT 42.655 4.435 42.665 4.749 ;
      RECT 42.575 4.363 42.655 4.829 ;
      RECT 42.61 5.007 42.62 5.232 ;
      RECT 42.605 5.004 42.61 5.227 ;
      RECT 42.59 5.001 42.605 5.22 ;
      RECT 42.555 4.995 42.59 5.202 ;
      RECT 42.57 4.298 42.575 4.903 ;
      RECT 42.55 4.249 42.57 4.918 ;
      RECT 42.54 4.982 42.555 5.185 ;
      RECT 42.545 4.191 42.55 4.933 ;
      RECT 42.54 4.169 42.545 4.943 ;
      RECT 42.505 4.079 42.54 5.18 ;
      RECT 42.49 3.957 42.505 5.18 ;
      RECT 42.485 3.91 42.49 5.18 ;
      RECT 42.46 3.835 42.485 5.18 ;
      RECT 42.445 3.75 42.46 5.18 ;
      RECT 42.44 3.697 42.445 5.18 ;
      RECT 42.435 3.677 42.44 5.18 ;
      RECT 42.43 3.652 42.435 4.414 ;
      RECT 42.415 4.612 42.435 5.18 ;
      RECT 42.425 3.63 42.43 4.391 ;
      RECT 42.415 3.582 42.425 4.356 ;
      RECT 42.41 3.545 42.415 4.322 ;
      RECT 42.41 4.692 42.415 5.18 ;
      RECT 42.395 3.522 42.41 4.277 ;
      RECT 42.39 4.79 42.41 5.18 ;
      RECT 42.34 3.41 42.395 4.119 ;
      RECT 42.385 4.912 42.39 5.18 ;
      RECT 42.325 3.41 42.34 3.958 ;
      RECT 42.32 3.41 42.325 3.91 ;
      RECT 42.315 3.41 42.32 3.898 ;
      RECT 42.27 3.41 42.315 3.835 ;
      RECT 42.245 3.41 42.27 3.753 ;
      RECT 42.23 3.41 42.245 3.705 ;
      RECT 42.225 3.41 42.23 3.675 ;
      RECT 44.615 3.455 44.875 3.715 ;
      RECT 44.61 3.455 44.875 3.663 ;
      RECT 44.605 3.455 44.875 3.633 ;
      RECT 44.58 3.325 44.86 3.605 ;
      RECT 33.14 9.09 33.49 9.44 ;
      RECT 44.11 9.045 44.46 9.395 ;
      RECT 33.14 9.12 44.46 9.32 ;
      RECT 43.62 5.005 43.9 5.285 ;
      RECT 43.66 4.96 43.925 5.22 ;
      RECT 43.65 4.995 43.925 5.22 ;
      RECT 43.655 4.98 43.9 5.285 ;
      RECT 43.66 4.957 43.87 5.285 ;
      RECT 43.66 4.955 43.855 5.285 ;
      RECT 43.7 4.945 43.855 5.285 ;
      RECT 43.67 4.95 43.855 5.285 ;
      RECT 43.7 4.942 43.8 5.285 ;
      RECT 43.725 4.935 43.8 5.285 ;
      RECT 43.705 4.937 43.8 5.285 ;
      RECT 43.035 4.45 43.295 4.71 ;
      RECT 43.085 4.442 43.275 4.71 ;
      RECT 43.09 4.362 43.275 4.71 ;
      RECT 43.21 3.75 43.275 4.71 ;
      RECT 43.115 4.147 43.275 4.71 ;
      RECT 43.19 3.835 43.275 4.71 ;
      RECT 43.225 3.46 43.361 4.188 ;
      RECT 43.17 3.957 43.361 4.188 ;
      RECT 43.185 3.897 43.275 4.71 ;
      RECT 43.225 3.46 43.385 3.853 ;
      RECT 43.225 3.46 43.395 3.75 ;
      RECT 43.215 3.46 43.475 3.72 ;
      RECT 41.55 4.86 41.595 5.12 ;
      RECT 41.455 3.395 41.6 3.655 ;
      RECT 41.96 4.017 41.97 4.108 ;
      RECT 41.945 3.955 41.96 4.164 ;
      RECT 41.94 3.902 41.945 4.21 ;
      RECT 41.89 3.849 41.94 4.336 ;
      RECT 41.885 3.804 41.89 4.483 ;
      RECT 41.875 3.792 41.885 4.525 ;
      RECT 41.84 3.756 41.875 4.63 ;
      RECT 41.835 3.724 41.84 4.736 ;
      RECT 41.82 3.706 41.835 4.781 ;
      RECT 41.815 3.689 41.82 4.015 ;
      RECT 41.81 4.07 41.82 4.838 ;
      RECT 41.805 3.675 41.815 3.988 ;
      RECT 41.8 4.125 41.81 5.12 ;
      RECT 41.795 3.661 41.805 3.973 ;
      RECT 41.795 4.175 41.8 5.12 ;
      RECT 41.78 3.638 41.795 3.953 ;
      RECT 41.76 4.297 41.795 5.12 ;
      RECT 41.775 3.62 41.78 3.935 ;
      RECT 41.77 3.612 41.775 3.925 ;
      RECT 41.74 3.58 41.77 3.889 ;
      RECT 41.75 4.425 41.76 5.12 ;
      RECT 41.745 4.452 41.75 5.12 ;
      RECT 41.74 4.502 41.745 5.12 ;
      RECT 41.73 3.546 41.74 3.854 ;
      RECT 41.69 4.57 41.74 5.12 ;
      RECT 41.715 3.523 41.73 3.83 ;
      RECT 41.69 3.395 41.715 3.793 ;
      RECT 41.685 3.395 41.69 3.765 ;
      RECT 41.655 4.67 41.69 5.12 ;
      RECT 41.68 3.395 41.685 3.758 ;
      RECT 41.675 3.395 41.68 3.748 ;
      RECT 41.66 3.395 41.675 3.733 ;
      RECT 41.645 3.395 41.66 3.705 ;
      RECT 41.61 4.775 41.655 5.12 ;
      RECT 41.63 3.395 41.645 3.678 ;
      RECT 41.6 3.395 41.63 3.663 ;
      RECT 41.595 4.847 41.61 5.12 ;
      RECT 41.52 3.93 41.56 4.19 ;
      RECT 41.295 3.877 41.3 4.135 ;
      RECT 37.25 3.355 37.51 3.615 ;
      RECT 37.25 3.38 37.525 3.595 ;
      RECT 39.64 3.205 39.645 3.35 ;
      RECT 41.51 3.925 41.52 4.19 ;
      RECT 41.49 3.917 41.51 4.19 ;
      RECT 41.472 3.913 41.49 4.19 ;
      RECT 41.386 3.902 41.472 4.19 ;
      RECT 41.3 3.885 41.386 4.19 ;
      RECT 41.245 3.872 41.295 4.12 ;
      RECT 41.211 3.864 41.245 4.095 ;
      RECT 41.125 3.853 41.211 4.06 ;
      RECT 41.09 3.83 41.125 4.025 ;
      RECT 41.08 3.792 41.09 4.011 ;
      RECT 41.075 3.765 41.08 4.007 ;
      RECT 41.07 3.752 41.075 4.004 ;
      RECT 41.06 3.732 41.07 4 ;
      RECT 41.055 3.707 41.06 3.996 ;
      RECT 41.03 3.662 41.055 3.99 ;
      RECT 41.02 3.603 41.03 3.982 ;
      RECT 41.01 3.571 41.02 3.973 ;
      RECT 40.99 3.523 41.01 3.953 ;
      RECT 40.985 3.483 40.99 3.923 ;
      RECT 40.97 3.457 40.985 3.897 ;
      RECT 40.965 3.435 40.97 3.873 ;
      RECT 40.95 3.407 40.965 3.849 ;
      RECT 40.935 3.38 40.95 3.813 ;
      RECT 40.92 3.357 40.935 3.775 ;
      RECT 40.915 3.347 40.92 3.75 ;
      RECT 40.905 3.34 40.915 3.733 ;
      RECT 40.89 3.327 40.905 3.703 ;
      RECT 40.885 3.317 40.89 3.678 ;
      RECT 40.88 3.312 40.885 3.665 ;
      RECT 40.87 3.305 40.88 3.645 ;
      RECT 40.865 3.298 40.87 3.63 ;
      RECT 40.84 3.291 40.865 3.588 ;
      RECT 40.825 3.281 40.84 3.538 ;
      RECT 40.815 3.276 40.825 3.508 ;
      RECT 40.805 3.272 40.815 3.483 ;
      RECT 40.79 3.269 40.805 3.473 ;
      RECT 40.74 3.266 40.79 3.458 ;
      RECT 40.72 3.264 40.74 3.443 ;
      RECT 40.671 3.262 40.72 3.438 ;
      RECT 40.585 3.258 40.671 3.433 ;
      RECT 40.546 3.255 40.585 3.429 ;
      RECT 40.46 3.251 40.546 3.424 ;
      RECT 40.41 3.248 40.46 3.418 ;
      RECT 40.361 3.245 40.41 3.413 ;
      RECT 40.275 3.242 40.361 3.408 ;
      RECT 40.271 3.24 40.275 3.405 ;
      RECT 40.185 3.237 40.271 3.4 ;
      RECT 40.136 3.233 40.185 3.393 ;
      RECT 40.05 3.23 40.136 3.388 ;
      RECT 40.026 3.227 40.05 3.384 ;
      RECT 39.94 3.225 40.026 3.379 ;
      RECT 39.875 3.221 39.94 3.372 ;
      RECT 39.872 3.22 39.875 3.369 ;
      RECT 39.786 3.217 39.872 3.366 ;
      RECT 39.7 3.211 39.786 3.359 ;
      RECT 39.67 3.207 39.7 3.355 ;
      RECT 39.645 3.205 39.67 3.353 ;
      RECT 39.59 3.202 39.64 3.35 ;
      RECT 39.51 3.201 39.59 3.35 ;
      RECT 39.455 3.203 39.51 3.353 ;
      RECT 39.44 3.204 39.455 3.357 ;
      RECT 39.385 3.212 39.44 3.367 ;
      RECT 39.355 3.22 39.385 3.38 ;
      RECT 39.336 3.221 39.355 3.386 ;
      RECT 39.25 3.224 39.336 3.391 ;
      RECT 39.18 3.229 39.25 3.4 ;
      RECT 39.161 3.232 39.18 3.406 ;
      RECT 39.075 3.236 39.161 3.411 ;
      RECT 39.035 3.24 39.075 3.418 ;
      RECT 39.026 3.242 39.035 3.421 ;
      RECT 38.94 3.246 39.026 3.426 ;
      RECT 38.937 3.249 38.94 3.43 ;
      RECT 38.851 3.252 38.937 3.434 ;
      RECT 38.765 3.258 38.851 3.442 ;
      RECT 38.741 3.262 38.765 3.446 ;
      RECT 38.655 3.266 38.741 3.451 ;
      RECT 38.61 3.271 38.655 3.458 ;
      RECT 38.53 3.276 38.61 3.465 ;
      RECT 38.45 3.282 38.53 3.48 ;
      RECT 38.425 3.286 38.45 3.493 ;
      RECT 38.36 3.289 38.425 3.505 ;
      RECT 38.305 3.294 38.36 3.52 ;
      RECT 38.275 3.297 38.305 3.538 ;
      RECT 38.265 3.299 38.275 3.551 ;
      RECT 38.205 3.314 38.265 3.561 ;
      RECT 38.19 3.331 38.205 3.57 ;
      RECT 38.185 3.34 38.19 3.57 ;
      RECT 38.175 3.35 38.185 3.57 ;
      RECT 38.165 3.367 38.175 3.57 ;
      RECT 38.145 3.377 38.165 3.571 ;
      RECT 38.1 3.387 38.145 3.572 ;
      RECT 38.065 3.396 38.1 3.574 ;
      RECT 38 3.401 38.065 3.576 ;
      RECT 37.92 3.402 38 3.579 ;
      RECT 37.916 3.4 37.92 3.58 ;
      RECT 37.83 3.397 37.916 3.582 ;
      RECT 37.783 3.394 37.83 3.584 ;
      RECT 37.697 3.39 37.783 3.587 ;
      RECT 37.611 3.386 37.697 3.59 ;
      RECT 37.525 3.382 37.611 3.594 ;
      RECT 40.91 5.005 40.94 5.285 ;
      RECT 40.66 4.895 40.68 5.285 ;
      RECT 40.615 4.895 40.68 5.155 ;
      RECT 40.445 3.52 40.48 3.78 ;
      RECT 40.22 3.52 40.28 3.78 ;
      RECT 40.9 4.985 40.91 5.285 ;
      RECT 40.895 4.945 40.9 5.285 ;
      RECT 40.88 4.9 40.895 5.285 ;
      RECT 40.875 4.865 40.88 5.285 ;
      RECT 40.87 4.845 40.875 5.285 ;
      RECT 40.84 4.772 40.87 5.285 ;
      RECT 40.82 4.67 40.84 5.285 ;
      RECT 40.81 4.6 40.82 5.285 ;
      RECT 40.765 4.54 40.81 5.285 ;
      RECT 40.68 4.501 40.765 5.285 ;
      RECT 40.675 4.492 40.68 4.865 ;
      RECT 40.665 4.491 40.675 4.848 ;
      RECT 40.64 4.472 40.665 4.818 ;
      RECT 40.635 4.447 40.64 4.797 ;
      RECT 40.625 4.425 40.635 4.788 ;
      RECT 40.62 4.396 40.625 4.778 ;
      RECT 40.58 4.322 40.62 4.75 ;
      RECT 40.56 4.223 40.58 4.715 ;
      RECT 40.545 4.159 40.56 4.698 ;
      RECT 40.515 4.083 40.545 4.67 ;
      RECT 40.495 3.998 40.515 4.643 ;
      RECT 40.455 3.894 40.495 4.55 ;
      RECT 40.45 3.815 40.455 4.458 ;
      RECT 40.445 3.798 40.45 4.435 ;
      RECT 40.44 3.52 40.445 4.415 ;
      RECT 40.41 3.52 40.44 4.353 ;
      RECT 40.405 3.52 40.41 4.285 ;
      RECT 40.395 3.52 40.405 4.25 ;
      RECT 40.385 3.52 40.395 4.215 ;
      RECT 40.32 3.52 40.385 4.07 ;
      RECT 40.315 3.52 40.32 3.94 ;
      RECT 40.285 3.52 40.315 3.873 ;
      RECT 40.28 3.52 40.285 3.798 ;
      RECT 39.46 4.445 39.74 4.725 ;
      RECT 39.5 4.425 39.76 4.685 ;
      RECT 39.49 4.435 39.76 4.685 ;
      RECT 39.5 4.362 39.715 4.725 ;
      RECT 39.555 4.285 39.71 4.725 ;
      RECT 39.56 4.07 39.71 4.725 ;
      RECT 39.55 3.872 39.7 4.123 ;
      RECT 39.54 3.872 39.7 3.99 ;
      RECT 39.535 3.75 39.695 3.893 ;
      RECT 39.52 3.75 39.695 3.798 ;
      RECT 39.515 3.46 39.69 3.775 ;
      RECT 39.5 3.46 39.69 3.745 ;
      RECT 39.46 3.46 39.72 3.72 ;
      RECT 39.37 4.93 39.45 5.19 ;
      RECT 38.775 3.65 38.78 3.915 ;
      RECT 38.655 3.65 38.78 3.91 ;
      RECT 39.33 4.895 39.37 5.19 ;
      RECT 39.285 4.817 39.33 5.19 ;
      RECT 39.265 4.745 39.285 5.19 ;
      RECT 39.255 4.697 39.265 5.19 ;
      RECT 39.22 4.63 39.255 5.19 ;
      RECT 39.19 4.53 39.22 5.19 ;
      RECT 39.17 4.455 39.19 4.99 ;
      RECT 39.16 4.405 39.17 4.945 ;
      RECT 39.155 4.382 39.16 4.918 ;
      RECT 39.15 4.367 39.155 4.905 ;
      RECT 39.145 4.352 39.15 4.883 ;
      RECT 39.14 4.337 39.145 4.865 ;
      RECT 39.115 4.292 39.14 4.82 ;
      RECT 39.105 4.24 39.115 4.763 ;
      RECT 39.095 4.21 39.105 4.73 ;
      RECT 39.085 4.175 39.095 4.698 ;
      RECT 39.05 4.107 39.085 4.63 ;
      RECT 39.045 4.046 39.05 4.565 ;
      RECT 39.035 4.034 39.045 4.545 ;
      RECT 39.03 4.022 39.035 4.525 ;
      RECT 39.025 4.014 39.03 4.513 ;
      RECT 39.02 4.006 39.025 4.493 ;
      RECT 39.01 3.994 39.02 4.465 ;
      RECT 39 3.978 39.01 4.435 ;
      RECT 38.975 3.95 39 4.373 ;
      RECT 38.965 3.921 38.975 4.318 ;
      RECT 38.95 3.9 38.965 4.278 ;
      RECT 38.945 3.884 38.95 4.25 ;
      RECT 38.94 3.872 38.945 4.24 ;
      RECT 38.935 3.867 38.94 4.213 ;
      RECT 38.93 3.86 38.935 4.2 ;
      RECT 38.915 3.843 38.93 4.173 ;
      RECT 38.905 3.65 38.915 4.133 ;
      RECT 38.895 3.65 38.905 4.1 ;
      RECT 38.885 3.65 38.895 4.075 ;
      RECT 38.815 3.65 38.885 4.01 ;
      RECT 38.805 3.65 38.815 3.958 ;
      RECT 38.79 3.65 38.805 3.94 ;
      RECT 38.78 3.65 38.79 3.925 ;
      RECT 38.61 4.52 38.87 4.78 ;
      RECT 37.145 4.555 37.15 4.762 ;
      RECT 36.78 4.445 36.855 4.76 ;
      RECT 36.595 4.5 36.75 4.76 ;
      RECT 36.78 4.445 36.885 4.725 ;
      RECT 38.595 4.617 38.61 4.778 ;
      RECT 38.57 4.625 38.595 4.783 ;
      RECT 38.545 4.632 38.57 4.788 ;
      RECT 38.482 4.643 38.545 4.797 ;
      RECT 38.396 4.662 38.482 4.814 ;
      RECT 38.31 4.684 38.396 4.833 ;
      RECT 38.295 4.697 38.31 4.844 ;
      RECT 38.255 4.705 38.295 4.851 ;
      RECT 38.235 4.71 38.255 4.858 ;
      RECT 38.197 4.711 38.235 4.861 ;
      RECT 38.111 4.714 38.197 4.862 ;
      RECT 38.025 4.718 38.111 4.863 ;
      RECT 37.976 4.72 38.025 4.865 ;
      RECT 37.89 4.72 37.976 4.867 ;
      RECT 37.85 4.715 37.89 4.869 ;
      RECT 37.84 4.709 37.85 4.87 ;
      RECT 37.8 4.704 37.84 4.867 ;
      RECT 37.79 4.697 37.8 4.863 ;
      RECT 37.775 4.693 37.79 4.861 ;
      RECT 37.758 4.689 37.775 4.859 ;
      RECT 37.672 4.679 37.758 4.851 ;
      RECT 37.586 4.661 37.672 4.837 ;
      RECT 37.5 4.644 37.586 4.823 ;
      RECT 37.475 4.632 37.5 4.814 ;
      RECT 37.405 4.622 37.475 4.807 ;
      RECT 37.36 4.61 37.405 4.798 ;
      RECT 37.3 4.597 37.36 4.79 ;
      RECT 37.295 4.589 37.3 4.785 ;
      RECT 37.26 4.584 37.295 4.783 ;
      RECT 37.205 4.575 37.26 4.776 ;
      RECT 37.165 4.564 37.205 4.768 ;
      RECT 37.15 4.557 37.165 4.764 ;
      RECT 37.13 4.55 37.145 4.761 ;
      RECT 37.115 4.54 37.13 4.759 ;
      RECT 37.1 4.527 37.115 4.756 ;
      RECT 37.075 4.51 37.1 4.752 ;
      RECT 37.06 4.492 37.075 4.749 ;
      RECT 37.035 4.445 37.06 4.747 ;
      RECT 37.011 4.445 37.035 4.744 ;
      RECT 36.925 4.445 37.011 4.736 ;
      RECT 36.885 4.445 36.925 4.728 ;
      RECT 36.75 4.492 36.78 4.76 ;
      RECT 38.43 4.075 38.69 4.335 ;
      RECT 38.39 4.075 38.69 4.213 ;
      RECT 38.355 4.075 38.69 4.198 ;
      RECT 38.3 4.075 38.69 4.178 ;
      RECT 38.22 3.885 38.5 4.165 ;
      RECT 38.22 4.067 38.57 4.165 ;
      RECT 38.22 4.01 38.555 4.165 ;
      RECT 38.22 3.957 38.505 4.165 ;
      RECT 36.05 3.885 36.245 4.67 ;
      RECT 36.13 2.5 36.245 4.67 ;
      RECT 35.985 4.41 36.045 4.67 ;
      RECT 37.355 3.93 37.615 4.19 ;
      RECT 36.04 3.885 36.245 4.165 ;
      RECT 37.35 3.94 37.615 4.125 ;
      RECT 37.065 3.915 37.075 4.065 ;
      RECT 36.3 2.5 36.38 2.845 ;
      RECT 36.035 2.5 36.245 2.845 ;
      RECT 37.34 3.94 37.35 4.124 ;
      RECT 37.33 3.939 37.34 4.121 ;
      RECT 37.321 3.938 37.33 4.119 ;
      RECT 37.235 3.934 37.321 4.109 ;
      RECT 37.161 3.926 37.235 4.091 ;
      RECT 37.075 3.919 37.161 4.074 ;
      RECT 37.015 3.915 37.065 4.064 ;
      RECT 36.98 3.914 37.015 4.061 ;
      RECT 36.925 3.914 36.98 4.063 ;
      RECT 36.89 3.914 36.925 4.067 ;
      RECT 36.804 3.913 36.89 4.074 ;
      RECT 36.718 3.912 36.804 4.084 ;
      RECT 36.632 3.911 36.718 4.095 ;
      RECT 36.546 3.911 36.632 4.105 ;
      RECT 36.46 3.91 36.546 4.115 ;
      RECT 36.425 3.91 36.46 4.155 ;
      RECT 36.42 3.91 36.425 4.198 ;
      RECT 36.395 3.91 36.42 4.215 ;
      RECT 36.32 3.91 36.395 4.23 ;
      RECT 36.3 3.885 36.32 4.243 ;
      RECT 36.295 2.5 36.3 4.253 ;
      RECT 36.27 2.5 36.295 4.295 ;
      RECT 36.245 2.5 36.27 4.373 ;
      RECT 36.045 4.292 36.05 4.67 ;
      RECT 35.38 4.244 35.395 4.7 ;
      RECT 35.375 4.316 35.481 4.698 ;
      RECT 35.395 3.41 35.53 4.696 ;
      RECT 35.38 4.26 35.535 4.695 ;
      RECT 35.38 4.31 35.54 4.693 ;
      RECT 35.365 4.375 35.54 4.692 ;
      RECT 35.375 4.367 35.545 4.689 ;
      RECT 35.355 4.415 35.545 4.684 ;
      RECT 35.355 4.415 35.56 4.681 ;
      RECT 35.35 4.415 35.56 4.678 ;
      RECT 35.325 4.415 35.585 4.675 ;
      RECT 35.395 3.41 35.555 4.063 ;
      RECT 35.39 3.41 35.555 4.035 ;
      RECT 35.385 3.41 35.555 3.863 ;
      RECT 35.385 3.41 35.575 3.803 ;
      RECT 35.34 3.41 35.6 3.67 ;
      RECT 34.82 3.885 35.1 4.165 ;
      RECT 34.81 3.9 35.1 4.16 ;
      RECT 34.765 3.962 35.1 4.158 ;
      RECT 34.84 3.877 35.005 4.165 ;
      RECT 34.84 3.862 34.961 4.165 ;
      RECT 34.875 3.855 34.961 4.165 ;
      RECT 34.34 5.005 34.62 5.285 ;
      RECT 34.3 4.967 34.595 5.078 ;
      RECT 34.285 4.917 34.575 4.973 ;
      RECT 34.23 4.68 34.49 4.94 ;
      RECT 34.23 4.882 34.57 4.94 ;
      RECT 34.23 4.822 34.565 4.94 ;
      RECT 34.23 4.772 34.545 4.94 ;
      RECT 34.23 4.752 34.54 4.94 ;
      RECT 34.23 4.73 34.535 4.94 ;
      RECT 34.23 4.715 34.505 4.94 ;
      RECT 29.96 8.66 30.28 8.98 ;
      RECT 29.99 8.13 30.16 8.98 ;
      RECT 29.99 8.13 30.165 8.48 ;
      RECT 29.99 8.13 30.965 8.305 ;
      RECT 30.79 3.26 30.965 8.305 ;
      RECT 30.735 3.26 31.085 3.61 ;
      RECT 30.76 9.09 31.085 9.415 ;
      RECT 29.645 9.18 31.085 9.35 ;
      RECT 29.645 3.69 29.805 9.35 ;
      RECT 29.96 3.66 30.28 3.98 ;
      RECT 29.645 3.69 30.28 3.86 ;
      RECT 28.315 2.435 28.69 2.805 ;
      RECT 20.235 2.255 20.61 2.625 ;
      RECT 18.8 2.255 19.175 2.625 ;
      RECT 18.8 2.375 28.62 2.545 ;
      RECT 24.745 5.655 28.6 5.825 ;
      RECT 28.43 4.72 28.6 5.825 ;
      RECT 24.745 4.965 24.915 5.825 ;
      RECT 24.695 5.005 24.975 5.285 ;
      RECT 24.715 4.965 24.975 5.285 ;
      RECT 24.355 4.92 24.46 5.18 ;
      RECT 28.34 4.725 28.69 5.075 ;
      RECT 24.21 3.41 24.3 3.67 ;
      RECT 24.75 4.475 24.755 4.515 ;
      RECT 24.745 4.465 24.75 4.6 ;
      RECT 24.74 4.455 24.745 4.693 ;
      RECT 24.73 4.435 24.74 4.749 ;
      RECT 24.65 4.363 24.73 4.829 ;
      RECT 24.685 5.007 24.695 5.232 ;
      RECT 24.68 5.004 24.685 5.227 ;
      RECT 24.665 5.001 24.68 5.22 ;
      RECT 24.63 4.995 24.665 5.202 ;
      RECT 24.645 4.298 24.65 4.903 ;
      RECT 24.625 4.249 24.645 4.918 ;
      RECT 24.615 4.982 24.63 5.185 ;
      RECT 24.62 4.191 24.625 4.933 ;
      RECT 24.615 4.169 24.62 4.943 ;
      RECT 24.58 4.079 24.615 5.18 ;
      RECT 24.565 3.957 24.58 5.18 ;
      RECT 24.56 3.91 24.565 5.18 ;
      RECT 24.535 3.835 24.56 5.18 ;
      RECT 24.52 3.75 24.535 5.18 ;
      RECT 24.515 3.697 24.52 5.18 ;
      RECT 24.51 3.677 24.515 5.18 ;
      RECT 24.505 3.652 24.51 4.414 ;
      RECT 24.49 4.612 24.51 5.18 ;
      RECT 24.5 3.63 24.505 4.391 ;
      RECT 24.49 3.582 24.5 4.356 ;
      RECT 24.485 3.545 24.49 4.322 ;
      RECT 24.485 4.692 24.49 5.18 ;
      RECT 24.47 3.522 24.485 4.277 ;
      RECT 24.465 4.79 24.485 5.18 ;
      RECT 24.415 3.41 24.47 4.119 ;
      RECT 24.46 4.912 24.465 5.18 ;
      RECT 24.4 3.41 24.415 3.958 ;
      RECT 24.395 3.41 24.4 3.91 ;
      RECT 24.39 3.41 24.395 3.898 ;
      RECT 24.345 3.41 24.39 3.835 ;
      RECT 24.32 3.41 24.345 3.753 ;
      RECT 24.305 3.41 24.32 3.705 ;
      RECT 24.3 3.41 24.305 3.675 ;
      RECT 26.69 3.455 26.95 3.715 ;
      RECT 26.685 3.455 26.95 3.663 ;
      RECT 26.68 3.455 26.95 3.633 ;
      RECT 26.655 3.325 26.935 3.605 ;
      RECT 14.515 9.43 14.805 9.78 ;
      RECT 14.515 9.49 15.65 9.66 ;
      RECT 15.48 9.12 15.65 9.66 ;
      RECT 26.205 9.04 26.375 9.395 ;
      RECT 26.155 9.04 26.505 9.39 ;
      RECT 15.48 9.12 26.505 9.29 ;
      RECT 25.695 5.005 25.975 5.285 ;
      RECT 25.735 4.96 26 5.22 ;
      RECT 25.725 4.995 26 5.22 ;
      RECT 25.73 4.98 25.975 5.285 ;
      RECT 25.735 4.957 25.945 5.285 ;
      RECT 25.735 4.955 25.93 5.285 ;
      RECT 25.775 4.945 25.93 5.285 ;
      RECT 25.745 4.95 25.93 5.285 ;
      RECT 25.775 4.942 25.875 5.285 ;
      RECT 25.8 4.935 25.875 5.285 ;
      RECT 25.78 4.937 25.875 5.285 ;
      RECT 25.11 4.45 25.37 4.71 ;
      RECT 25.16 4.442 25.35 4.71 ;
      RECT 25.165 4.362 25.35 4.71 ;
      RECT 25.285 3.75 25.35 4.71 ;
      RECT 25.19 4.147 25.35 4.71 ;
      RECT 25.265 3.835 25.35 4.71 ;
      RECT 25.3 3.46 25.436 4.188 ;
      RECT 25.245 3.957 25.436 4.188 ;
      RECT 25.26 3.897 25.35 4.71 ;
      RECT 25.3 3.46 25.46 3.853 ;
      RECT 25.3 3.46 25.47 3.75 ;
      RECT 25.29 3.46 25.55 3.72 ;
      RECT 23.625 4.86 23.67 5.12 ;
      RECT 23.53 3.395 23.675 3.655 ;
      RECT 24.035 4.017 24.045 4.108 ;
      RECT 24.02 3.955 24.035 4.164 ;
      RECT 24.015 3.902 24.02 4.21 ;
      RECT 23.965 3.849 24.015 4.336 ;
      RECT 23.96 3.804 23.965 4.483 ;
      RECT 23.95 3.792 23.96 4.525 ;
      RECT 23.915 3.756 23.95 4.63 ;
      RECT 23.91 3.724 23.915 4.736 ;
      RECT 23.895 3.706 23.91 4.781 ;
      RECT 23.89 3.689 23.895 4.015 ;
      RECT 23.885 4.07 23.895 4.838 ;
      RECT 23.88 3.675 23.89 3.988 ;
      RECT 23.875 4.125 23.885 5.12 ;
      RECT 23.87 3.661 23.88 3.973 ;
      RECT 23.87 4.175 23.875 5.12 ;
      RECT 23.855 3.638 23.87 3.953 ;
      RECT 23.835 4.297 23.87 5.12 ;
      RECT 23.85 3.62 23.855 3.935 ;
      RECT 23.845 3.612 23.85 3.925 ;
      RECT 23.815 3.58 23.845 3.889 ;
      RECT 23.825 4.425 23.835 5.12 ;
      RECT 23.82 4.452 23.825 5.12 ;
      RECT 23.815 4.502 23.82 5.12 ;
      RECT 23.805 3.546 23.815 3.854 ;
      RECT 23.765 4.57 23.815 5.12 ;
      RECT 23.79 3.523 23.805 3.83 ;
      RECT 23.765 3.395 23.79 3.793 ;
      RECT 23.76 3.395 23.765 3.765 ;
      RECT 23.73 4.67 23.765 5.12 ;
      RECT 23.755 3.395 23.76 3.758 ;
      RECT 23.75 3.395 23.755 3.748 ;
      RECT 23.735 3.395 23.75 3.733 ;
      RECT 23.72 3.395 23.735 3.705 ;
      RECT 23.685 4.775 23.73 5.12 ;
      RECT 23.705 3.395 23.72 3.678 ;
      RECT 23.675 3.395 23.705 3.663 ;
      RECT 23.67 4.847 23.685 5.12 ;
      RECT 23.595 3.93 23.635 4.19 ;
      RECT 23.37 3.877 23.375 4.135 ;
      RECT 19.325 3.355 19.585 3.615 ;
      RECT 19.325 3.38 19.6 3.595 ;
      RECT 21.715 3.205 21.72 3.35 ;
      RECT 23.585 3.925 23.595 4.19 ;
      RECT 23.565 3.917 23.585 4.19 ;
      RECT 23.547 3.913 23.565 4.19 ;
      RECT 23.461 3.902 23.547 4.19 ;
      RECT 23.375 3.885 23.461 4.19 ;
      RECT 23.32 3.872 23.37 4.12 ;
      RECT 23.286 3.864 23.32 4.095 ;
      RECT 23.2 3.853 23.286 4.06 ;
      RECT 23.165 3.83 23.2 4.025 ;
      RECT 23.155 3.792 23.165 4.011 ;
      RECT 23.15 3.765 23.155 4.007 ;
      RECT 23.145 3.752 23.15 4.004 ;
      RECT 23.135 3.732 23.145 4 ;
      RECT 23.13 3.707 23.135 3.996 ;
      RECT 23.105 3.662 23.13 3.99 ;
      RECT 23.095 3.603 23.105 3.982 ;
      RECT 23.085 3.571 23.095 3.973 ;
      RECT 23.065 3.523 23.085 3.953 ;
      RECT 23.06 3.483 23.065 3.923 ;
      RECT 23.045 3.457 23.06 3.897 ;
      RECT 23.04 3.435 23.045 3.873 ;
      RECT 23.025 3.407 23.04 3.849 ;
      RECT 23.01 3.38 23.025 3.813 ;
      RECT 22.995 3.357 23.01 3.775 ;
      RECT 22.99 3.347 22.995 3.75 ;
      RECT 22.98 3.34 22.99 3.733 ;
      RECT 22.965 3.327 22.98 3.703 ;
      RECT 22.96 3.317 22.965 3.678 ;
      RECT 22.955 3.312 22.96 3.665 ;
      RECT 22.945 3.305 22.955 3.645 ;
      RECT 22.94 3.298 22.945 3.63 ;
      RECT 22.915 3.291 22.94 3.588 ;
      RECT 22.9 3.281 22.915 3.538 ;
      RECT 22.89 3.276 22.9 3.508 ;
      RECT 22.88 3.272 22.89 3.483 ;
      RECT 22.865 3.269 22.88 3.473 ;
      RECT 22.815 3.266 22.865 3.458 ;
      RECT 22.795 3.264 22.815 3.443 ;
      RECT 22.746 3.262 22.795 3.438 ;
      RECT 22.66 3.258 22.746 3.433 ;
      RECT 22.621 3.255 22.66 3.429 ;
      RECT 22.535 3.251 22.621 3.424 ;
      RECT 22.485 3.248 22.535 3.418 ;
      RECT 22.436 3.245 22.485 3.413 ;
      RECT 22.35 3.242 22.436 3.408 ;
      RECT 22.346 3.24 22.35 3.405 ;
      RECT 22.26 3.237 22.346 3.4 ;
      RECT 22.211 3.233 22.26 3.393 ;
      RECT 22.125 3.23 22.211 3.388 ;
      RECT 22.101 3.227 22.125 3.384 ;
      RECT 22.015 3.225 22.101 3.379 ;
      RECT 21.95 3.221 22.015 3.372 ;
      RECT 21.947 3.22 21.95 3.369 ;
      RECT 21.861 3.217 21.947 3.366 ;
      RECT 21.775 3.211 21.861 3.359 ;
      RECT 21.745 3.207 21.775 3.355 ;
      RECT 21.72 3.205 21.745 3.353 ;
      RECT 21.665 3.202 21.715 3.35 ;
      RECT 21.585 3.201 21.665 3.35 ;
      RECT 21.53 3.203 21.585 3.353 ;
      RECT 21.515 3.204 21.53 3.357 ;
      RECT 21.46 3.212 21.515 3.367 ;
      RECT 21.43 3.22 21.46 3.38 ;
      RECT 21.411 3.221 21.43 3.386 ;
      RECT 21.325 3.224 21.411 3.391 ;
      RECT 21.255 3.229 21.325 3.4 ;
      RECT 21.236 3.232 21.255 3.406 ;
      RECT 21.15 3.236 21.236 3.411 ;
      RECT 21.11 3.24 21.15 3.418 ;
      RECT 21.101 3.242 21.11 3.421 ;
      RECT 21.015 3.246 21.101 3.426 ;
      RECT 21.012 3.249 21.015 3.43 ;
      RECT 20.926 3.252 21.012 3.434 ;
      RECT 20.84 3.258 20.926 3.442 ;
      RECT 20.816 3.262 20.84 3.446 ;
      RECT 20.73 3.266 20.816 3.451 ;
      RECT 20.685 3.271 20.73 3.458 ;
      RECT 20.605 3.276 20.685 3.465 ;
      RECT 20.525 3.282 20.605 3.48 ;
      RECT 20.5 3.286 20.525 3.493 ;
      RECT 20.435 3.289 20.5 3.505 ;
      RECT 20.38 3.294 20.435 3.52 ;
      RECT 20.35 3.297 20.38 3.538 ;
      RECT 20.34 3.299 20.35 3.551 ;
      RECT 20.28 3.314 20.34 3.561 ;
      RECT 20.265 3.331 20.28 3.57 ;
      RECT 20.26 3.34 20.265 3.57 ;
      RECT 20.25 3.35 20.26 3.57 ;
      RECT 20.24 3.367 20.25 3.57 ;
      RECT 20.22 3.377 20.24 3.571 ;
      RECT 20.175 3.387 20.22 3.572 ;
      RECT 20.14 3.396 20.175 3.574 ;
      RECT 20.075 3.401 20.14 3.576 ;
      RECT 19.995 3.402 20.075 3.579 ;
      RECT 19.991 3.4 19.995 3.58 ;
      RECT 19.905 3.397 19.991 3.582 ;
      RECT 19.858 3.394 19.905 3.584 ;
      RECT 19.772 3.39 19.858 3.587 ;
      RECT 19.686 3.386 19.772 3.59 ;
      RECT 19.6 3.382 19.686 3.594 ;
      RECT 22.985 5.005 23.015 5.285 ;
      RECT 22.735 4.895 22.755 5.285 ;
      RECT 22.69 4.895 22.755 5.155 ;
      RECT 22.52 3.52 22.555 3.78 ;
      RECT 22.295 3.52 22.355 3.78 ;
      RECT 22.975 4.985 22.985 5.285 ;
      RECT 22.97 4.945 22.975 5.285 ;
      RECT 22.955 4.9 22.97 5.285 ;
      RECT 22.95 4.865 22.955 5.285 ;
      RECT 22.945 4.845 22.95 5.285 ;
      RECT 22.915 4.772 22.945 5.285 ;
      RECT 22.895 4.67 22.915 5.285 ;
      RECT 22.885 4.6 22.895 5.285 ;
      RECT 22.84 4.54 22.885 5.285 ;
      RECT 22.755 4.501 22.84 5.285 ;
      RECT 22.75 4.492 22.755 4.865 ;
      RECT 22.74 4.491 22.75 4.848 ;
      RECT 22.715 4.472 22.74 4.818 ;
      RECT 22.71 4.447 22.715 4.797 ;
      RECT 22.7 4.425 22.71 4.788 ;
      RECT 22.695 4.396 22.7 4.778 ;
      RECT 22.655 4.322 22.695 4.75 ;
      RECT 22.635 4.223 22.655 4.715 ;
      RECT 22.62 4.159 22.635 4.698 ;
      RECT 22.59 4.083 22.62 4.67 ;
      RECT 22.57 3.998 22.59 4.643 ;
      RECT 22.53 3.894 22.57 4.55 ;
      RECT 22.525 3.815 22.53 4.458 ;
      RECT 22.52 3.798 22.525 4.435 ;
      RECT 22.515 3.52 22.52 4.415 ;
      RECT 22.485 3.52 22.515 4.353 ;
      RECT 22.48 3.52 22.485 4.285 ;
      RECT 22.47 3.52 22.48 4.25 ;
      RECT 22.46 3.52 22.47 4.215 ;
      RECT 22.395 3.52 22.46 4.07 ;
      RECT 22.39 3.52 22.395 3.94 ;
      RECT 22.36 3.52 22.39 3.873 ;
      RECT 22.355 3.52 22.36 3.798 ;
      RECT 21.535 4.445 21.815 4.725 ;
      RECT 21.575 4.425 21.835 4.685 ;
      RECT 21.565 4.435 21.835 4.685 ;
      RECT 21.575 4.362 21.79 4.725 ;
      RECT 21.63 4.285 21.785 4.725 ;
      RECT 21.635 4.07 21.785 4.725 ;
      RECT 21.625 3.872 21.775 4.123 ;
      RECT 21.615 3.872 21.775 3.99 ;
      RECT 21.61 3.75 21.77 3.893 ;
      RECT 21.595 3.75 21.77 3.798 ;
      RECT 21.59 3.46 21.765 3.775 ;
      RECT 21.575 3.46 21.765 3.745 ;
      RECT 21.535 3.46 21.795 3.72 ;
      RECT 21.445 4.93 21.525 5.19 ;
      RECT 20.85 3.65 20.855 3.915 ;
      RECT 20.73 3.65 20.855 3.91 ;
      RECT 21.405 4.895 21.445 5.19 ;
      RECT 21.36 4.817 21.405 5.19 ;
      RECT 21.34 4.745 21.36 5.19 ;
      RECT 21.33 4.697 21.34 5.19 ;
      RECT 21.295 4.63 21.33 5.19 ;
      RECT 21.265 4.53 21.295 5.19 ;
      RECT 21.245 4.455 21.265 4.99 ;
      RECT 21.235 4.405 21.245 4.945 ;
      RECT 21.23 4.382 21.235 4.918 ;
      RECT 21.225 4.367 21.23 4.905 ;
      RECT 21.22 4.352 21.225 4.883 ;
      RECT 21.215 4.337 21.22 4.865 ;
      RECT 21.19 4.292 21.215 4.82 ;
      RECT 21.18 4.24 21.19 4.763 ;
      RECT 21.17 4.21 21.18 4.73 ;
      RECT 21.16 4.175 21.17 4.698 ;
      RECT 21.125 4.107 21.16 4.63 ;
      RECT 21.12 4.046 21.125 4.565 ;
      RECT 21.11 4.034 21.12 4.545 ;
      RECT 21.105 4.022 21.11 4.525 ;
      RECT 21.1 4.014 21.105 4.513 ;
      RECT 21.095 4.006 21.1 4.493 ;
      RECT 21.085 3.994 21.095 4.465 ;
      RECT 21.075 3.978 21.085 4.435 ;
      RECT 21.05 3.95 21.075 4.373 ;
      RECT 21.04 3.921 21.05 4.318 ;
      RECT 21.025 3.9 21.04 4.278 ;
      RECT 21.02 3.884 21.025 4.25 ;
      RECT 21.015 3.872 21.02 4.24 ;
      RECT 21.01 3.867 21.015 4.213 ;
      RECT 21.005 3.86 21.01 4.2 ;
      RECT 20.99 3.843 21.005 4.173 ;
      RECT 20.98 3.65 20.99 4.133 ;
      RECT 20.97 3.65 20.98 4.1 ;
      RECT 20.96 3.65 20.97 4.075 ;
      RECT 20.89 3.65 20.96 4.01 ;
      RECT 20.88 3.65 20.89 3.958 ;
      RECT 20.865 3.65 20.88 3.94 ;
      RECT 20.855 3.65 20.865 3.925 ;
      RECT 20.685 4.52 20.945 4.78 ;
      RECT 19.22 4.555 19.225 4.762 ;
      RECT 18.855 4.445 18.93 4.76 ;
      RECT 18.67 4.5 18.825 4.76 ;
      RECT 18.855 4.445 18.96 4.725 ;
      RECT 20.67 4.617 20.685 4.778 ;
      RECT 20.645 4.625 20.67 4.783 ;
      RECT 20.62 4.632 20.645 4.788 ;
      RECT 20.557 4.643 20.62 4.797 ;
      RECT 20.471 4.662 20.557 4.814 ;
      RECT 20.385 4.684 20.471 4.833 ;
      RECT 20.37 4.697 20.385 4.844 ;
      RECT 20.33 4.705 20.37 4.851 ;
      RECT 20.31 4.71 20.33 4.858 ;
      RECT 20.272 4.711 20.31 4.861 ;
      RECT 20.186 4.714 20.272 4.862 ;
      RECT 20.1 4.718 20.186 4.863 ;
      RECT 20.051 4.72 20.1 4.865 ;
      RECT 19.965 4.72 20.051 4.867 ;
      RECT 19.925 4.715 19.965 4.869 ;
      RECT 19.915 4.709 19.925 4.87 ;
      RECT 19.875 4.704 19.915 4.867 ;
      RECT 19.865 4.697 19.875 4.863 ;
      RECT 19.85 4.693 19.865 4.861 ;
      RECT 19.833 4.689 19.85 4.859 ;
      RECT 19.747 4.679 19.833 4.851 ;
      RECT 19.661 4.661 19.747 4.837 ;
      RECT 19.575 4.644 19.661 4.823 ;
      RECT 19.55 4.632 19.575 4.814 ;
      RECT 19.48 4.622 19.55 4.807 ;
      RECT 19.435 4.61 19.48 4.798 ;
      RECT 19.375 4.597 19.435 4.79 ;
      RECT 19.37 4.589 19.375 4.785 ;
      RECT 19.335 4.584 19.37 4.783 ;
      RECT 19.28 4.575 19.335 4.776 ;
      RECT 19.24 4.564 19.28 4.768 ;
      RECT 19.225 4.557 19.24 4.764 ;
      RECT 19.205 4.55 19.22 4.761 ;
      RECT 19.19 4.54 19.205 4.759 ;
      RECT 19.175 4.527 19.19 4.756 ;
      RECT 19.15 4.51 19.175 4.752 ;
      RECT 19.135 4.492 19.15 4.749 ;
      RECT 19.11 4.445 19.135 4.747 ;
      RECT 19.086 4.445 19.11 4.744 ;
      RECT 19 4.445 19.086 4.736 ;
      RECT 18.96 4.445 19 4.728 ;
      RECT 18.825 4.492 18.855 4.76 ;
      RECT 20.505 4.075 20.765 4.335 ;
      RECT 20.465 4.075 20.765 4.213 ;
      RECT 20.43 4.075 20.765 4.198 ;
      RECT 20.375 4.075 20.765 4.178 ;
      RECT 20.295 3.885 20.575 4.165 ;
      RECT 20.295 4.067 20.645 4.165 ;
      RECT 20.295 4.01 20.63 4.165 ;
      RECT 20.295 3.957 20.58 4.165 ;
      RECT 18.125 3.885 18.32 4.67 ;
      RECT 18.205 2.5 18.32 4.67 ;
      RECT 18.06 4.41 18.12 4.67 ;
      RECT 19.43 3.93 19.69 4.19 ;
      RECT 18.115 3.885 18.32 4.165 ;
      RECT 19.425 3.94 19.69 4.125 ;
      RECT 19.14 3.915 19.15 4.065 ;
      RECT 18.375 2.5 18.455 2.845 ;
      RECT 18.11 2.5 18.32 2.845 ;
      RECT 19.415 3.94 19.425 4.124 ;
      RECT 19.405 3.939 19.415 4.121 ;
      RECT 19.396 3.938 19.405 4.119 ;
      RECT 19.31 3.934 19.396 4.109 ;
      RECT 19.236 3.926 19.31 4.091 ;
      RECT 19.15 3.919 19.236 4.074 ;
      RECT 19.09 3.915 19.14 4.064 ;
      RECT 19.055 3.914 19.09 4.061 ;
      RECT 19 3.914 19.055 4.063 ;
      RECT 18.965 3.914 19 4.067 ;
      RECT 18.879 3.913 18.965 4.074 ;
      RECT 18.793 3.912 18.879 4.084 ;
      RECT 18.707 3.911 18.793 4.095 ;
      RECT 18.621 3.911 18.707 4.105 ;
      RECT 18.535 3.91 18.621 4.115 ;
      RECT 18.5 3.91 18.535 4.155 ;
      RECT 18.495 3.91 18.5 4.198 ;
      RECT 18.47 3.91 18.495 4.215 ;
      RECT 18.395 3.91 18.47 4.23 ;
      RECT 18.375 3.885 18.395 4.243 ;
      RECT 18.37 2.5 18.375 4.253 ;
      RECT 18.345 2.5 18.37 4.295 ;
      RECT 18.32 2.5 18.345 4.373 ;
      RECT 18.12 4.292 18.125 4.67 ;
      RECT 17.455 4.244 17.47 4.7 ;
      RECT 17.45 4.316 17.556 4.698 ;
      RECT 17.47 3.41 17.605 4.696 ;
      RECT 17.455 4.26 17.61 4.695 ;
      RECT 17.455 4.31 17.615 4.693 ;
      RECT 17.44 4.375 17.615 4.692 ;
      RECT 17.45 4.367 17.62 4.689 ;
      RECT 17.43 4.415 17.62 4.684 ;
      RECT 17.43 4.415 17.635 4.681 ;
      RECT 17.425 4.415 17.635 4.678 ;
      RECT 17.4 4.415 17.66 4.675 ;
      RECT 17.47 3.41 17.63 4.063 ;
      RECT 17.465 3.41 17.63 4.035 ;
      RECT 17.46 3.41 17.63 3.863 ;
      RECT 17.46 3.41 17.65 3.803 ;
      RECT 17.415 3.41 17.675 3.67 ;
      RECT 16.895 3.885 17.175 4.165 ;
      RECT 16.885 3.9 17.175 4.16 ;
      RECT 16.84 3.962 17.175 4.158 ;
      RECT 16.915 3.877 17.08 4.165 ;
      RECT 16.915 3.862 17.036 4.165 ;
      RECT 16.95 3.855 17.036 4.165 ;
      RECT 16.415 5.005 16.695 5.285 ;
      RECT 16.375 4.967 16.67 5.078 ;
      RECT 16.36 4.917 16.65 4.973 ;
      RECT 16.305 4.68 16.565 4.94 ;
      RECT 16.305 4.882 16.645 4.94 ;
      RECT 16.305 4.822 16.64 4.94 ;
      RECT 16.305 4.772 16.62 4.94 ;
      RECT 16.305 4.752 16.615 4.94 ;
      RECT 16.305 4.73 16.61 4.94 ;
      RECT 16.305 4.715 16.58 4.94 ;
      RECT 97.195 9.49 97.57 9.86 ;
      RECT 88.53 2.225 88.905 2.595 ;
      RECT 79.27 9.49 79.645 9.86 ;
      RECT 70.605 2.225 70.98 2.595 ;
      RECT 61.345 9.49 61.72 9.86 ;
      RECT 52.68 2.225 53.055 2.595 ;
      RECT 43.42 9.49 43.795 9.86 ;
      RECT 34.755 2.225 35.13 2.595 ;
      RECT 25.495 9.49 25.87 9.86 ;
      RECT 16.83 2.225 17.205 2.595 ;
    LAYER via1 ;
      RECT 104.915 9.81 105.065 9.96 ;
      RECT 102.55 9.175 102.7 9.325 ;
      RECT 102.535 3.36 102.685 3.51 ;
      RECT 101.745 3.745 101.895 3.895 ;
      RECT 101.745 8.76 101.895 8.91 ;
      RECT 100.14 4.825 100.29 4.975 ;
      RECT 100.13 2.545 100.28 2.695 ;
      RECT 98.445 3.51 98.595 3.66 ;
      RECT 98.215 9.145 98.365 9.295 ;
      RECT 97.495 5.015 97.645 5.165 ;
      RECT 97.31 9.6 97.46 9.75 ;
      RECT 97.045 3.515 97.195 3.665 ;
      RECT 96.865 4.505 97.015 4.655 ;
      RECT 96.47 5.02 96.62 5.17 ;
      RECT 96.11 4.975 96.26 5.125 ;
      RECT 95.965 3.465 96.115 3.615 ;
      RECT 95.38 4.915 95.53 5.065 ;
      RECT 95.285 3.45 95.435 3.6 ;
      RECT 95.13 3.985 95.28 4.135 ;
      RECT 94.445 4.95 94.595 5.1 ;
      RECT 94.05 3.575 94.2 3.725 ;
      RECT 93.33 4.48 93.48 4.63 ;
      RECT 93.29 3.515 93.44 3.665 ;
      RECT 93.02 4.985 93.17 5.135 ;
      RECT 92.485 3.705 92.635 3.855 ;
      RECT 92.44 4.575 92.59 4.725 ;
      RECT 92.26 4.13 92.41 4.28 ;
      RECT 91.185 3.985 91.335 4.135 ;
      RECT 91.08 3.41 91.23 3.56 ;
      RECT 90.425 4.555 90.575 4.705 ;
      RECT 89.905 2.595 90.055 2.745 ;
      RECT 89.815 4.465 89.965 4.615 ;
      RECT 89.17 3.465 89.32 3.615 ;
      RECT 89.155 4.47 89.305 4.62 ;
      RECT 88.64 3.955 88.79 4.105 ;
      RECT 88.06 4.735 88.21 4.885 ;
      RECT 86.97 9.19 87.12 9.34 ;
      RECT 84.625 9.175 84.775 9.325 ;
      RECT 84.61 3.36 84.76 3.51 ;
      RECT 83.82 3.745 83.97 3.895 ;
      RECT 83.82 8.76 83.97 8.91 ;
      RECT 82.215 4.825 82.365 4.975 ;
      RECT 82.205 2.545 82.355 2.695 ;
      RECT 80.52 3.51 80.67 3.66 ;
      RECT 80.01 9.145 80.16 9.295 ;
      RECT 79.57 5.015 79.72 5.165 ;
      RECT 79.385 9.6 79.535 9.75 ;
      RECT 79.12 3.515 79.27 3.665 ;
      RECT 78.94 4.505 79.09 4.655 ;
      RECT 78.545 5.02 78.695 5.17 ;
      RECT 78.185 4.975 78.335 5.125 ;
      RECT 78.04 3.465 78.19 3.615 ;
      RECT 77.455 4.915 77.605 5.065 ;
      RECT 77.36 3.45 77.51 3.6 ;
      RECT 77.205 3.985 77.355 4.135 ;
      RECT 76.52 4.95 76.67 5.1 ;
      RECT 76.125 3.575 76.275 3.725 ;
      RECT 75.405 4.48 75.555 4.63 ;
      RECT 75.365 3.515 75.515 3.665 ;
      RECT 75.095 4.985 75.245 5.135 ;
      RECT 74.56 3.705 74.71 3.855 ;
      RECT 74.515 4.575 74.665 4.725 ;
      RECT 74.335 4.13 74.485 4.28 ;
      RECT 73.26 3.985 73.41 4.135 ;
      RECT 73.155 3.41 73.305 3.56 ;
      RECT 72.5 4.555 72.65 4.705 ;
      RECT 71.98 2.595 72.13 2.745 ;
      RECT 71.89 4.465 72.04 4.615 ;
      RECT 71.245 3.465 71.395 3.615 ;
      RECT 71.23 4.47 71.38 4.62 ;
      RECT 70.715 3.955 70.865 4.105 ;
      RECT 70.135 4.735 70.285 4.885 ;
      RECT 69.045 9.19 69.195 9.34 ;
      RECT 66.7 9.175 66.85 9.325 ;
      RECT 66.685 3.36 66.835 3.51 ;
      RECT 65.895 3.745 66.045 3.895 ;
      RECT 65.895 8.76 66.045 8.91 ;
      RECT 64.29 4.825 64.44 4.975 ;
      RECT 64.28 2.545 64.43 2.695 ;
      RECT 62.595 3.51 62.745 3.66 ;
      RECT 62.14 9.15 62.29 9.3 ;
      RECT 61.645 5.015 61.795 5.165 ;
      RECT 61.46 9.6 61.61 9.75 ;
      RECT 61.195 3.515 61.345 3.665 ;
      RECT 61.015 4.505 61.165 4.655 ;
      RECT 60.62 5.02 60.77 5.17 ;
      RECT 60.26 4.975 60.41 5.125 ;
      RECT 60.115 3.465 60.265 3.615 ;
      RECT 59.53 4.915 59.68 5.065 ;
      RECT 59.435 3.45 59.585 3.6 ;
      RECT 59.28 3.985 59.43 4.135 ;
      RECT 58.595 4.95 58.745 5.1 ;
      RECT 58.2 3.575 58.35 3.725 ;
      RECT 57.48 4.48 57.63 4.63 ;
      RECT 57.44 3.515 57.59 3.665 ;
      RECT 57.17 4.985 57.32 5.135 ;
      RECT 56.635 3.705 56.785 3.855 ;
      RECT 56.59 4.575 56.74 4.725 ;
      RECT 56.41 4.13 56.56 4.28 ;
      RECT 55.335 3.985 55.485 4.135 ;
      RECT 55.23 3.41 55.38 3.56 ;
      RECT 54.575 4.555 54.725 4.705 ;
      RECT 54.055 2.595 54.205 2.745 ;
      RECT 53.965 4.465 54.115 4.615 ;
      RECT 53.32 3.465 53.47 3.615 ;
      RECT 53.305 4.47 53.455 4.62 ;
      RECT 52.79 3.955 52.94 4.105 ;
      RECT 52.21 4.735 52.36 4.885 ;
      RECT 51.165 9.195 51.315 9.345 ;
      RECT 48.775 9.175 48.925 9.325 ;
      RECT 48.76 3.36 48.91 3.51 ;
      RECT 47.97 3.745 48.12 3.895 ;
      RECT 47.97 8.76 48.12 8.91 ;
      RECT 46.365 4.825 46.515 4.975 ;
      RECT 46.355 2.545 46.505 2.695 ;
      RECT 44.67 3.51 44.82 3.66 ;
      RECT 44.21 9.145 44.36 9.295 ;
      RECT 43.72 5.015 43.87 5.165 ;
      RECT 43.535 9.6 43.685 9.75 ;
      RECT 43.27 3.515 43.42 3.665 ;
      RECT 43.09 4.505 43.24 4.655 ;
      RECT 42.695 5.02 42.845 5.17 ;
      RECT 42.335 4.975 42.485 5.125 ;
      RECT 42.19 3.465 42.34 3.615 ;
      RECT 41.605 4.915 41.755 5.065 ;
      RECT 41.51 3.45 41.66 3.6 ;
      RECT 41.355 3.985 41.505 4.135 ;
      RECT 40.67 4.95 40.82 5.1 ;
      RECT 40.275 3.575 40.425 3.725 ;
      RECT 39.555 4.48 39.705 4.63 ;
      RECT 39.515 3.515 39.665 3.665 ;
      RECT 39.245 4.985 39.395 5.135 ;
      RECT 38.71 3.705 38.86 3.855 ;
      RECT 38.665 4.575 38.815 4.725 ;
      RECT 38.485 4.13 38.635 4.28 ;
      RECT 37.41 3.985 37.56 4.135 ;
      RECT 37.305 3.41 37.455 3.56 ;
      RECT 36.65 4.555 36.8 4.705 ;
      RECT 36.13 2.595 36.28 2.745 ;
      RECT 36.04 4.465 36.19 4.615 ;
      RECT 35.395 3.465 35.545 3.615 ;
      RECT 35.38 4.47 35.53 4.62 ;
      RECT 34.865 3.955 35.015 4.105 ;
      RECT 34.285 4.735 34.435 4.885 ;
      RECT 33.24 9.19 33.39 9.34 ;
      RECT 30.85 9.175 31 9.325 ;
      RECT 30.835 3.36 30.985 3.51 ;
      RECT 30.045 3.745 30.195 3.895 ;
      RECT 30.045 8.76 30.195 8.91 ;
      RECT 28.44 4.825 28.59 4.975 ;
      RECT 28.43 2.545 28.58 2.695 ;
      RECT 26.745 3.51 26.895 3.66 ;
      RECT 26.255 9.14 26.405 9.29 ;
      RECT 25.795 5.015 25.945 5.165 ;
      RECT 25.61 9.6 25.76 9.75 ;
      RECT 25.345 3.515 25.495 3.665 ;
      RECT 25.165 4.505 25.315 4.655 ;
      RECT 24.77 5.02 24.92 5.17 ;
      RECT 24.41 4.975 24.56 5.125 ;
      RECT 24.265 3.465 24.415 3.615 ;
      RECT 23.68 4.915 23.83 5.065 ;
      RECT 23.585 3.45 23.735 3.6 ;
      RECT 23.43 3.985 23.58 4.135 ;
      RECT 22.745 4.95 22.895 5.1 ;
      RECT 22.35 3.575 22.5 3.725 ;
      RECT 21.63 4.48 21.78 4.63 ;
      RECT 21.59 3.515 21.74 3.665 ;
      RECT 21.32 4.985 21.47 5.135 ;
      RECT 20.785 3.705 20.935 3.855 ;
      RECT 20.74 4.575 20.89 4.725 ;
      RECT 20.56 4.13 20.71 4.28 ;
      RECT 19.485 3.985 19.635 4.135 ;
      RECT 19.38 3.41 19.53 3.56 ;
      RECT 18.725 4.555 18.875 4.705 ;
      RECT 18.205 2.595 18.355 2.745 ;
      RECT 18.115 4.465 18.265 4.615 ;
      RECT 17.47 3.465 17.62 3.615 ;
      RECT 17.455 4.47 17.605 4.62 ;
      RECT 16.94 3.955 17.09 4.105 ;
      RECT 16.36 4.735 16.51 4.885 ;
      RECT 14.585 9.53 14.735 9.68 ;
      RECT 14.21 8.79 14.36 8.94 ;
    LAYER met1 ;
      RECT 87.84 2.58 99.8 3.185 ;
      RECT 92.265 0 99.8 3.185 ;
      RECT 69.915 2.58 81.875 3.185 ;
      RECT 74.34 0 81.875 3.185 ;
      RECT 51.99 2.58 63.95 3.185 ;
      RECT 56.415 0 63.95 3.185 ;
      RECT 34.065 2.58 46.025 3.185 ;
      RECT 38.49 0 46.025 3.185 ;
      RECT 16.14 2.58 28.1 3.185 ;
      RECT 20.565 0 28.1 3.185 ;
      RECT 87.835 0 88.58 2.975 ;
      RECT 69.91 0 70.655 2.975 ;
      RECT 51.985 0 52.73 2.975 ;
      RECT 34.06 0 34.805 2.975 ;
      RECT 16.135 0 16.88 2.975 ;
      RECT 90.83 0 91.985 3.185 ;
      RECT 87.835 2.55 90.55 2.975 ;
      RECT 88.86 0 90.55 3.185 ;
      RECT 72.905 0 74.06 3.185 ;
      RECT 69.91 2.55 72.625 2.975 ;
      RECT 70.935 0 72.625 3.185 ;
      RECT 54.98 0 56.135 3.185 ;
      RECT 51.985 2.55 54.7 2.975 ;
      RECT 53.01 0 54.7 3.185 ;
      RECT 37.055 0 38.21 3.185 ;
      RECT 34.06 2.55 36.775 2.975 ;
      RECT 35.085 0 36.775 3.185 ;
      RECT 19.13 0 20.285 3.185 ;
      RECT 16.135 2.55 18.85 2.975 ;
      RECT 17.16 0 18.85 3.185 ;
      RECT 88.86 0 99.8 2.3 ;
      RECT 70.935 0 81.875 2.3 ;
      RECT 53.01 0 63.95 2.3 ;
      RECT 35.085 0 46.025 2.3 ;
      RECT 17.16 0 28.1 2.3 ;
      RECT 87.835 0 99.8 2.27 ;
      RECT 69.91 0 81.875 2.27 ;
      RECT 51.985 0 63.95 2.27 ;
      RECT 34.06 0 46.025 2.27 ;
      RECT 16.135 0 28.1 2.27 ;
      RECT 12.97 0 105.39 1.6 ;
      RECT 104.785 10.205 105.075 10.435 ;
      RECT 104.845 8.725 105.015 10.435 ;
      RECT 104.815 9.71 105.165 10.06 ;
      RECT 104.785 8.725 105.075 8.955 ;
      RECT 104.38 3.69 104.485 4.26 ;
      RECT 104.38 4.025 104.705 4.255 ;
      RECT 104.38 4.055 104.875 4.225 ;
      RECT 104.38 3.69 104.57 4.255 ;
      RECT 103.795 3.655 104.085 3.885 ;
      RECT 103.795 3.69 104.57 3.86 ;
      RECT 103.855 2.175 104.025 3.885 ;
      RECT 103.795 2.175 104.085 2.405 ;
      RECT 103.795 10.205 104.085 10.435 ;
      RECT 103.855 8.725 104.025 10.435 ;
      RECT 103.795 8.725 104.085 8.955 ;
      RECT 103.795 8.76 104.65 8.92 ;
      RECT 104.48 8.355 104.65 8.92 ;
      RECT 103.795 8.755 104.19 8.92 ;
      RECT 104.415 8.355 104.705 8.585 ;
      RECT 104.415 8.385 104.875 8.555 ;
      RECT 103.425 4.025 103.715 4.255 ;
      RECT 103.425 4.055 103.885 4.225 ;
      RECT 103.49 2.95 103.655 4.255 ;
      RECT 102.005 2.92 102.295 3.15 ;
      RECT 102.005 2.95 103.655 3.12 ;
      RECT 102.065 2.18 102.235 3.15 ;
      RECT 102.005 2.18 102.295 2.41 ;
      RECT 102.005 10.2 102.295 10.43 ;
      RECT 102.065 9.46 102.235 10.43 ;
      RECT 102.065 9.555 103.655 9.725 ;
      RECT 103.485 8.355 103.655 9.725 ;
      RECT 102.005 9.46 102.295 9.69 ;
      RECT 103.425 8.355 103.715 8.585 ;
      RECT 103.425 8.385 103.885 8.555 ;
      RECT 100.04 4.725 100.39 5.075 ;
      RECT 100.13 3.32 100.3 5.075 ;
      RECT 102.435 3.26 102.785 3.61 ;
      RECT 100.13 3.32 101.75 3.495 ;
      RECT 100.13 3.32 102.785 3.49 ;
      RECT 102.46 9.09 102.785 9.415 ;
      RECT 98.115 9.045 98.465 9.395 ;
      RECT 102.435 9.09 102.785 9.32 ;
      RECT 97.675 9.09 97.965 9.32 ;
      RECT 97.505 9.12 102.785 9.29 ;
      RECT 101.66 3.66 101.98 3.98 ;
      RECT 101.63 3.66 101.98 3.89 ;
      RECT 101.46 3.69 101.98 3.86 ;
      RECT 101.66 8.66 101.98 8.98 ;
      RECT 101.63 8.72 101.98 8.95 ;
      RECT 101.46 8.75 101.98 8.92 ;
      RECT 97.44 4.96 97.48 5.22 ;
      RECT 97.48 4.94 97.485 4.95 ;
      RECT 98.81 4.185 98.82 4.406 ;
      RECT 98.74 4.18 98.81 4.531 ;
      RECT 98.73 4.18 98.74 4.658 ;
      RECT 98.705 4.18 98.73 4.705 ;
      RECT 98.68 4.18 98.705 4.783 ;
      RECT 98.66 4.18 98.68 4.853 ;
      RECT 98.635 4.18 98.66 4.893 ;
      RECT 98.625 4.18 98.635 4.913 ;
      RECT 98.615 4.182 98.625 4.921 ;
      RECT 98.61 4.187 98.615 4.378 ;
      RECT 98.61 4.387 98.615 4.922 ;
      RECT 98.605 4.432 98.61 4.923 ;
      RECT 98.595 4.497 98.605 4.924 ;
      RECT 98.585 4.592 98.595 4.926 ;
      RECT 98.58 4.645 98.585 4.928 ;
      RECT 98.575 4.665 98.58 4.929 ;
      RECT 98.52 4.69 98.575 4.935 ;
      RECT 98.48 4.725 98.52 4.944 ;
      RECT 98.47 4.742 98.48 4.949 ;
      RECT 98.461 4.748 98.47 4.951 ;
      RECT 98.375 4.786 98.461 4.962 ;
      RECT 98.37 4.825 98.375 4.972 ;
      RECT 98.295 4.832 98.37 4.982 ;
      RECT 98.275 4.842 98.295 4.993 ;
      RECT 98.245 4.849 98.275 5.001 ;
      RECT 98.22 4.856 98.245 5.008 ;
      RECT 98.196 4.862 98.22 5.013 ;
      RECT 98.11 4.875 98.196 5.025 ;
      RECT 98.032 4.882 98.11 5.043 ;
      RECT 97.946 4.877 98.032 5.061 ;
      RECT 97.86 4.872 97.946 5.081 ;
      RECT 97.78 4.866 97.86 5.098 ;
      RECT 97.715 4.862 97.78 5.127 ;
      RECT 97.71 4.576 97.715 4.6 ;
      RECT 97.7 4.852 97.715 5.155 ;
      RECT 97.705 4.57 97.71 4.64 ;
      RECT 97.7 4.564 97.705 4.71 ;
      RECT 97.695 4.558 97.7 4.788 ;
      RECT 97.695 4.835 97.7 5.22 ;
      RECT 97.687 4.555 97.695 5.22 ;
      RECT 97.601 4.553 97.687 5.22 ;
      RECT 97.515 4.551 97.601 5.22 ;
      RECT 97.505 4.552 97.515 5.22 ;
      RECT 97.5 4.557 97.505 5.22 ;
      RECT 97.49 4.57 97.5 5.22 ;
      RECT 97.485 4.592 97.49 5.22 ;
      RECT 97.48 4.952 97.485 5.22 ;
      RECT 98.11 4.42 98.115 4.64 ;
      RECT 98.615 3.455 98.65 3.715 ;
      RECT 98.6 3.455 98.615 3.723 ;
      RECT 98.571 3.455 98.6 3.745 ;
      RECT 98.485 3.455 98.571 3.805 ;
      RECT 98.465 3.455 98.485 3.87 ;
      RECT 98.405 3.455 98.465 4.035 ;
      RECT 98.4 3.455 98.405 4.183 ;
      RECT 98.395 3.455 98.4 4.195 ;
      RECT 98.39 3.455 98.395 4.221 ;
      RECT 98.36 3.641 98.39 4.301 ;
      RECT 98.355 3.689 98.36 4.39 ;
      RECT 98.35 3.703 98.355 4.405 ;
      RECT 98.345 3.722 98.35 4.435 ;
      RECT 98.34 3.737 98.345 4.451 ;
      RECT 98.335 3.752 98.34 4.473 ;
      RECT 98.33 3.772 98.335 4.495 ;
      RECT 98.32 3.792 98.33 4.528 ;
      RECT 98.305 3.834 98.32 4.59 ;
      RECT 98.3 3.865 98.305 4.63 ;
      RECT 98.295 3.877 98.3 4.635 ;
      RECT 98.29 3.889 98.295 4.64 ;
      RECT 98.285 3.902 98.29 4.64 ;
      RECT 98.28 3.92 98.285 4.64 ;
      RECT 98.275 3.94 98.28 4.64 ;
      RECT 98.27 3.952 98.275 4.64 ;
      RECT 98.265 3.965 98.27 4.64 ;
      RECT 98.245 4 98.265 4.64 ;
      RECT 98.195 4.102 98.245 4.64 ;
      RECT 98.19 4.187 98.195 4.64 ;
      RECT 98.185 4.195 98.19 4.64 ;
      RECT 98.18 4.212 98.185 4.64 ;
      RECT 98.175 4.227 98.18 4.64 ;
      RECT 98.14 4.292 98.175 4.64 ;
      RECT 98.125 4.357 98.14 4.64 ;
      RECT 98.12 4.387 98.125 4.64 ;
      RECT 98.115 4.412 98.12 4.64 ;
      RECT 98.1 4.422 98.11 4.64 ;
      RECT 98.085 4.435 98.1 4.633 ;
      RECT 97.83 4.025 97.9 4.235 ;
      RECT 97.62 4.002 97.625 4.195 ;
      RECT 95.075 3.93 95.335 4.19 ;
      RECT 97.91 4.212 97.915 4.215 ;
      RECT 97.9 4.03 97.91 4.23 ;
      RECT 97.801 4.023 97.83 4.235 ;
      RECT 97.715 4.015 97.801 4.235 ;
      RECT 97.7 4.009 97.715 4.233 ;
      RECT 97.68 4.008 97.7 4.22 ;
      RECT 97.675 4.007 97.68 4.203 ;
      RECT 97.625 4.004 97.675 4.198 ;
      RECT 97.595 4.001 97.62 4.193 ;
      RECT 97.575 3.999 97.595 4.188 ;
      RECT 97.56 3.997 97.575 4.185 ;
      RECT 97.53 3.995 97.56 4.183 ;
      RECT 97.465 3.991 97.53 4.175 ;
      RECT 97.435 3.986 97.465 4.17 ;
      RECT 97.415 3.984 97.435 4.168 ;
      RECT 97.385 3.981 97.415 4.163 ;
      RECT 97.325 3.977 97.385 4.155 ;
      RECT 97.32 3.974 97.325 4.15 ;
      RECT 97.25 3.972 97.32 4.145 ;
      RECT 97.221 3.968 97.25 4.138 ;
      RECT 97.135 3.963 97.221 4.13 ;
      RECT 97.101 3.958 97.135 4.122 ;
      RECT 97.015 3.95 97.101 4.114 ;
      RECT 96.976 3.943 97.015 4.106 ;
      RECT 96.89 3.938 96.976 4.098 ;
      RECT 96.825 3.932 96.89 4.088 ;
      RECT 96.805 3.927 96.825 4.083 ;
      RECT 96.796 3.924 96.805 4.082 ;
      RECT 96.71 3.92 96.796 4.076 ;
      RECT 96.67 3.916 96.71 4.068 ;
      RECT 96.65 3.912 96.67 4.066 ;
      RECT 96.59 3.912 96.65 4.063 ;
      RECT 96.57 3.915 96.59 4.061 ;
      RECT 96.549 3.915 96.57 4.061 ;
      RECT 96.463 3.917 96.549 4.065 ;
      RECT 96.377 3.919 96.463 4.071 ;
      RECT 96.291 3.921 96.377 4.078 ;
      RECT 96.205 3.924 96.291 4.084 ;
      RECT 96.171 3.925 96.205 4.089 ;
      RECT 96.085 3.928 96.171 4.094 ;
      RECT 96.056 3.935 96.085 4.099 ;
      RECT 95.97 3.935 96.056 4.104 ;
      RECT 95.937 3.935 95.97 4.109 ;
      RECT 95.851 3.937 95.937 4.114 ;
      RECT 95.765 3.939 95.851 4.121 ;
      RECT 95.701 3.941 95.765 4.127 ;
      RECT 95.615 3.943 95.701 4.133 ;
      RECT 95.612 3.945 95.615 4.136 ;
      RECT 95.526 3.946 95.612 4.14 ;
      RECT 95.44 3.949 95.526 4.147 ;
      RECT 95.421 3.951 95.44 4.151 ;
      RECT 95.335 3.953 95.421 4.156 ;
      RECT 95.065 3.965 95.075 4.16 ;
      RECT 97.245 10.2 97.535 10.43 ;
      RECT 97.305 9.46 97.475 10.43 ;
      RECT 97.195 9.49 97.57 9.86 ;
      RECT 97.245 9.46 97.535 9.86 ;
      RECT 97.3 3.545 97.485 3.755 ;
      RECT 97.295 3.546 97.49 3.753 ;
      RECT 97.29 3.551 97.5 3.748 ;
      RECT 97.285 3.527 97.29 3.745 ;
      RECT 97.255 3.524 97.285 3.738 ;
      RECT 97.25 3.52 97.255 3.729 ;
      RECT 97.215 3.551 97.5 3.724 ;
      RECT 96.99 3.46 97.25 3.72 ;
      RECT 97.29 3.529 97.295 3.748 ;
      RECT 97.295 3.53 97.3 3.753 ;
      RECT 96.99 3.542 97.37 3.72 ;
      RECT 96.99 3.54 97.355 3.72 ;
      RECT 96.99 3.535 97.345 3.72 ;
      RECT 96.945 4.45 96.995 4.735 ;
      RECT 96.89 4.42 96.895 4.735 ;
      RECT 96.86 4.4 96.865 4.735 ;
      RECT 97.01 4.45 97.07 4.71 ;
      RECT 97.005 4.45 97.01 4.718 ;
      RECT 96.995 4.45 97.005 4.73 ;
      RECT 96.91 4.44 96.945 4.735 ;
      RECT 96.905 4.427 96.91 4.735 ;
      RECT 96.895 4.422 96.905 4.735 ;
      RECT 96.875 4.412 96.89 4.735 ;
      RECT 96.865 4.405 96.875 4.735 ;
      RECT 96.855 4.397 96.86 4.735 ;
      RECT 96.825 4.387 96.855 4.735 ;
      RECT 96.81 4.375 96.825 4.735 ;
      RECT 96.795 4.365 96.81 4.73 ;
      RECT 96.775 4.355 96.795 4.705 ;
      RECT 96.765 4.347 96.775 4.682 ;
      RECT 96.735 4.33 96.765 4.672 ;
      RECT 96.73 4.307 96.735 4.663 ;
      RECT 96.725 4.294 96.73 4.661 ;
      RECT 96.71 4.27 96.725 4.655 ;
      RECT 96.705 4.246 96.71 4.649 ;
      RECT 96.695 4.235 96.705 4.644 ;
      RECT 96.69 4.225 96.695 4.64 ;
      RECT 96.685 4.217 96.69 4.637 ;
      RECT 96.675 4.212 96.685 4.633 ;
      RECT 96.67 4.207 96.675 4.629 ;
      RECT 96.585 4.205 96.67 4.604 ;
      RECT 96.555 4.205 96.585 4.57 ;
      RECT 96.54 4.205 96.555 4.553 ;
      RECT 96.485 4.205 96.54 4.498 ;
      RECT 96.48 4.21 96.485 4.447 ;
      RECT 96.47 4.215 96.48 4.437 ;
      RECT 96.465 4.225 96.47 4.423 ;
      RECT 96.415 4.965 96.675 5.225 ;
      RECT 96.335 4.98 96.675 5.201 ;
      RECT 96.315 4.98 96.675 5.196 ;
      RECT 96.291 4.98 96.675 5.194 ;
      RECT 96.205 4.98 96.675 5.189 ;
      RECT 96.055 4.92 96.315 5.185 ;
      RECT 96.01 4.98 96.675 5.18 ;
      RECT 96.005 4.987 96.675 5.175 ;
      RECT 96.02 4.975 96.335 5.185 ;
      RECT 95.91 3.41 96.17 3.67 ;
      RECT 95.91 3.467 96.175 3.663 ;
      RECT 95.91 3.497 96.18 3.595 ;
      RECT 95.97 3.928 96.085 3.93 ;
      RECT 96.056 3.925 96.085 3.93 ;
      RECT 95.08 4.929 95.105 5.169 ;
      RECT 95.065 4.932 95.155 5.163 ;
      RECT 95.06 4.937 95.241 5.158 ;
      RECT 95.055 4.945 95.305 5.156 ;
      RECT 95.055 4.945 95.315 5.155 ;
      RECT 95.05 4.952 95.325 5.148 ;
      RECT 95.05 4.952 95.411 5.137 ;
      RECT 95.045 4.987 95.411 5.133 ;
      RECT 95.045 4.987 95.42 5.122 ;
      RECT 95.325 4.86 95.585 5.12 ;
      RECT 95.035 5.037 95.585 5.118 ;
      RECT 95.305 4.905 95.325 5.153 ;
      RECT 95.241 4.908 95.305 5.157 ;
      RECT 95.155 4.913 95.241 5.162 ;
      RECT 95.085 4.924 95.585 5.12 ;
      RECT 95.105 4.918 95.155 5.167 ;
      RECT 95.23 3.395 95.24 3.657 ;
      RECT 95.22 3.452 95.23 3.66 ;
      RECT 95.195 3.457 95.22 3.666 ;
      RECT 95.17 3.461 95.195 3.678 ;
      RECT 95.16 3.464 95.17 3.688 ;
      RECT 95.155 3.465 95.16 3.693 ;
      RECT 95.15 3.466 95.155 3.698 ;
      RECT 95.145 3.467 95.15 3.7 ;
      RECT 95.12 3.47 95.145 3.703 ;
      RECT 95.09 3.476 95.12 3.706 ;
      RECT 95.025 3.487 95.09 3.709 ;
      RECT 94.98 3.495 95.025 3.713 ;
      RECT 94.965 3.495 94.98 3.721 ;
      RECT 94.96 3.496 94.965 3.728 ;
      RECT 94.955 3.498 94.96 3.731 ;
      RECT 94.95 3.502 94.955 3.734 ;
      RECT 94.94 3.51 94.95 3.738 ;
      RECT 94.935 3.523 94.94 3.743 ;
      RECT 94.93 3.531 94.935 3.745 ;
      RECT 94.925 3.537 94.93 3.745 ;
      RECT 94.92 3.541 94.925 3.748 ;
      RECT 94.915 3.543 94.92 3.751 ;
      RECT 94.91 3.546 94.915 3.754 ;
      RECT 94.9 3.551 94.91 3.758 ;
      RECT 94.895 3.557 94.9 3.763 ;
      RECT 94.885 3.563 94.895 3.767 ;
      RECT 94.87 3.57 94.885 3.773 ;
      RECT 94.841 3.584 94.87 3.783 ;
      RECT 94.755 3.619 94.841 3.815 ;
      RECT 94.735 3.652 94.755 3.844 ;
      RECT 94.715 3.665 94.735 3.855 ;
      RECT 94.695 3.677 94.715 3.866 ;
      RECT 94.645 3.699 94.695 3.886 ;
      RECT 94.63 3.717 94.645 3.903 ;
      RECT 94.625 3.723 94.63 3.906 ;
      RECT 94.62 3.727 94.625 3.909 ;
      RECT 94.615 3.731 94.62 3.913 ;
      RECT 94.61 3.733 94.615 3.916 ;
      RECT 94.6 3.74 94.61 3.919 ;
      RECT 94.595 3.745 94.6 3.923 ;
      RECT 94.59 3.747 94.595 3.926 ;
      RECT 94.585 3.751 94.59 3.929 ;
      RECT 94.58 3.753 94.585 3.933 ;
      RECT 94.565 3.758 94.58 3.938 ;
      RECT 94.56 3.763 94.565 3.941 ;
      RECT 94.555 3.771 94.56 3.944 ;
      RECT 94.55 3.773 94.555 3.947 ;
      RECT 94.545 3.775 94.55 3.95 ;
      RECT 94.535 3.777 94.545 3.956 ;
      RECT 94.5 3.791 94.535 3.968 ;
      RECT 94.49 3.806 94.5 3.978 ;
      RECT 94.415 3.835 94.49 4.002 ;
      RECT 94.41 3.86 94.415 4.025 ;
      RECT 94.395 3.864 94.41 4.031 ;
      RECT 94.385 3.872 94.395 4.036 ;
      RECT 94.355 3.885 94.385 4.04 ;
      RECT 94.345 3.9 94.355 4.045 ;
      RECT 94.335 3.905 94.345 4.048 ;
      RECT 94.33 3.907 94.335 4.05 ;
      RECT 94.315 3.91 94.33 4.053 ;
      RECT 94.31 3.912 94.315 4.056 ;
      RECT 94.29 3.917 94.31 4.06 ;
      RECT 94.26 3.922 94.29 4.068 ;
      RECT 94.235 3.929 94.26 4.076 ;
      RECT 94.23 3.934 94.235 4.081 ;
      RECT 94.2 3.937 94.23 4.085 ;
      RECT 94.16 3.94 94.2 4.095 ;
      RECT 94.125 3.937 94.16 4.107 ;
      RECT 94.115 3.933 94.125 4.114 ;
      RECT 94.09 3.929 94.115 4.12 ;
      RECT 94.085 3.925 94.09 4.125 ;
      RECT 94.045 3.922 94.085 4.125 ;
      RECT 94.03 3.907 94.045 4.126 ;
      RECT 94.007 3.895 94.03 4.126 ;
      RECT 93.921 3.895 94.007 4.127 ;
      RECT 93.835 3.895 93.921 4.129 ;
      RECT 93.815 3.895 93.835 4.126 ;
      RECT 93.81 3.9 93.815 4.121 ;
      RECT 93.805 3.905 93.81 4.119 ;
      RECT 93.795 3.915 93.805 4.117 ;
      RECT 93.79 3.921 93.795 4.11 ;
      RECT 93.785 3.923 93.79 4.095 ;
      RECT 93.78 3.927 93.785 4.085 ;
      RECT 95.24 3.395 95.49 3.655 ;
      RECT 92.965 4.93 93.225 5.19 ;
      RECT 95.26 4.42 95.265 4.63 ;
      RECT 95.265 4.425 95.275 4.625 ;
      RECT 95.215 4.42 95.26 4.645 ;
      RECT 95.205 4.42 95.215 4.665 ;
      RECT 95.186 4.42 95.205 4.67 ;
      RECT 95.1 4.42 95.186 4.667 ;
      RECT 95.07 4.422 95.1 4.665 ;
      RECT 95.015 4.432 95.07 4.663 ;
      RECT 94.95 4.446 95.015 4.661 ;
      RECT 94.945 4.454 94.95 4.66 ;
      RECT 94.93 4.457 94.945 4.658 ;
      RECT 94.865 4.467 94.93 4.654 ;
      RECT 94.817 4.481 94.865 4.655 ;
      RECT 94.731 4.498 94.817 4.669 ;
      RECT 94.645 4.519 94.731 4.686 ;
      RECT 94.625 4.532 94.645 4.696 ;
      RECT 94.58 4.54 94.625 4.703 ;
      RECT 94.545 4.548 94.58 4.711 ;
      RECT 94.511 4.556 94.545 4.719 ;
      RECT 94.425 4.57 94.511 4.731 ;
      RECT 94.39 4.587 94.425 4.743 ;
      RECT 94.381 4.596 94.39 4.747 ;
      RECT 94.295 4.614 94.381 4.764 ;
      RECT 94.236 4.641 94.295 4.791 ;
      RECT 94.15 4.668 94.236 4.819 ;
      RECT 94.13 4.69 94.15 4.839 ;
      RECT 94.07 4.705 94.13 4.855 ;
      RECT 94.06 4.717 94.07 4.868 ;
      RECT 94.055 4.722 94.06 4.871 ;
      RECT 94.045 4.725 94.055 4.874 ;
      RECT 94.04 4.727 94.045 4.877 ;
      RECT 94.01 4.735 94.04 4.884 ;
      RECT 93.995 4.742 94.01 4.892 ;
      RECT 93.985 4.747 93.995 4.896 ;
      RECT 93.98 4.75 93.985 4.899 ;
      RECT 93.97 4.752 93.98 4.902 ;
      RECT 93.935 4.762 93.97 4.911 ;
      RECT 93.86 4.785 93.935 4.933 ;
      RECT 93.84 4.803 93.86 4.951 ;
      RECT 93.81 4.81 93.84 4.961 ;
      RECT 93.79 4.818 93.81 4.971 ;
      RECT 93.78 4.824 93.79 4.978 ;
      RECT 93.761 4.829 93.78 4.984 ;
      RECT 93.675 4.849 93.761 5.004 ;
      RECT 93.66 4.869 93.675 5.023 ;
      RECT 93.615 4.881 93.66 5.034 ;
      RECT 93.55 4.902 93.615 5.057 ;
      RECT 93.51 4.922 93.55 5.078 ;
      RECT 93.5 4.932 93.51 5.088 ;
      RECT 93.45 4.944 93.5 5.099 ;
      RECT 93.43 4.96 93.45 5.111 ;
      RECT 93.4 4.97 93.43 5.117 ;
      RECT 93.39 4.975 93.4 5.119 ;
      RECT 93.321 4.976 93.39 5.125 ;
      RECT 93.235 4.978 93.321 5.135 ;
      RECT 93.225 4.979 93.235 5.14 ;
      RECT 94.495 5.005 94.685 5.215 ;
      RECT 94.485 5.01 94.695 5.208 ;
      RECT 94.47 5.01 94.695 5.173 ;
      RECT 94.39 4.895 94.65 5.155 ;
      RECT 93.305 4.425 93.49 4.72 ;
      RECT 93.295 4.425 93.49 4.718 ;
      RECT 93.28 4.425 93.495 4.713 ;
      RECT 93.28 4.425 93.5 4.71 ;
      RECT 93.275 4.425 93.5 4.708 ;
      RECT 93.27 4.68 93.5 4.698 ;
      RECT 93.275 4.425 93.535 4.685 ;
      RECT 93.235 3.46 93.495 3.72 ;
      RECT 93.045 3.385 93.131 3.718 ;
      RECT 93.02 3.389 93.175 3.714 ;
      RECT 93.131 3.381 93.175 3.714 ;
      RECT 93.131 3.382 93.18 3.713 ;
      RECT 93.045 3.387 93.195 3.712 ;
      RECT 93.02 3.395 93.235 3.711 ;
      RECT 93.015 3.39 93.195 3.706 ;
      RECT 93.005 3.405 93.235 3.613 ;
      RECT 93.005 3.457 93.435 3.613 ;
      RECT 93.005 3.45 93.415 3.613 ;
      RECT 93.005 3.437 93.385 3.613 ;
      RECT 93.005 3.425 93.325 3.613 ;
      RECT 93.005 3.41 93.3 3.613 ;
      RECT 92.205 4.04 92.34 4.335 ;
      RECT 92.465 4.063 92.47 4.25 ;
      RECT 93.185 3.96 93.33 4.195 ;
      RECT 93.345 3.96 93.35 4.185 ;
      RECT 93.38 3.971 93.385 4.165 ;
      RECT 93.375 3.963 93.38 4.17 ;
      RECT 93.355 3.96 93.375 4.175 ;
      RECT 93.35 3.96 93.355 4.183 ;
      RECT 93.34 3.96 93.345 4.188 ;
      RECT 93.33 3.96 93.34 4.193 ;
      RECT 93.16 3.962 93.185 4.195 ;
      RECT 93.11 3.969 93.16 4.195 ;
      RECT 93.105 3.974 93.11 4.195 ;
      RECT 93.066 3.979 93.105 4.196 ;
      RECT 92.98 3.991 93.066 4.197 ;
      RECT 92.971 4.001 92.98 4.197 ;
      RECT 92.885 4.01 92.971 4.199 ;
      RECT 92.861 4.02 92.885 4.201 ;
      RECT 92.775 4.031 92.861 4.202 ;
      RECT 92.745 4.042 92.775 4.204 ;
      RECT 92.715 4.047 92.745 4.206 ;
      RECT 92.69 4.053 92.715 4.209 ;
      RECT 92.675 4.058 92.69 4.21 ;
      RECT 92.63 4.064 92.675 4.21 ;
      RECT 92.625 4.069 92.63 4.211 ;
      RECT 92.605 4.069 92.625 4.213 ;
      RECT 92.585 4.067 92.605 4.218 ;
      RECT 92.55 4.066 92.585 4.225 ;
      RECT 92.52 4.065 92.55 4.235 ;
      RECT 92.47 4.064 92.52 4.245 ;
      RECT 92.38 4.061 92.465 4.335 ;
      RECT 92.355 4.055 92.38 4.335 ;
      RECT 92.34 4.045 92.355 4.335 ;
      RECT 92.155 4.04 92.205 4.255 ;
      RECT 92.145 4.045 92.155 4.245 ;
      RECT 92.385 4.52 92.645 4.78 ;
      RECT 92.385 4.52 92.675 4.673 ;
      RECT 92.385 4.52 92.71 4.658 ;
      RECT 92.64 4.44 92.83 4.65 ;
      RECT 92.63 4.445 92.84 4.643 ;
      RECT 92.595 4.515 92.84 4.643 ;
      RECT 92.625 4.457 92.645 4.78 ;
      RECT 92.61 4.505 92.84 4.643 ;
      RECT 92.615 4.477 92.645 4.78 ;
      RECT 91.695 3.545 91.765 4.65 ;
      RECT 92.43 3.65 92.69 3.91 ;
      RECT 92.01 3.696 92.025 3.905 ;
      RECT 92.346 3.709 92.43 3.86 ;
      RECT 92.26 3.706 92.346 3.86 ;
      RECT 92.221 3.704 92.26 3.86 ;
      RECT 92.135 3.702 92.221 3.86 ;
      RECT 92.075 3.7 92.135 3.871 ;
      RECT 92.04 3.698 92.075 3.889 ;
      RECT 92.025 3.696 92.04 3.9 ;
      RECT 91.995 3.696 92.01 3.913 ;
      RECT 91.985 3.696 91.995 3.918 ;
      RECT 91.96 3.695 91.985 3.923 ;
      RECT 91.945 3.69 91.96 3.929 ;
      RECT 91.94 3.683 91.945 3.934 ;
      RECT 91.915 3.674 91.94 3.94 ;
      RECT 91.87 3.653 91.915 3.953 ;
      RECT 91.86 3.637 91.87 3.963 ;
      RECT 91.845 3.63 91.86 3.973 ;
      RECT 91.835 3.623 91.845 3.99 ;
      RECT 91.83 3.62 91.835 4.02 ;
      RECT 91.825 3.618 91.83 4.05 ;
      RECT 91.82 3.616 91.825 4.087 ;
      RECT 91.805 3.612 91.82 4.154 ;
      RECT 91.805 4.445 91.815 4.645 ;
      RECT 91.8 3.608 91.805 4.28 ;
      RECT 91.8 4.432 91.805 4.65 ;
      RECT 91.795 3.606 91.8 4.365 ;
      RECT 91.795 4.422 91.8 4.65 ;
      RECT 91.78 3.577 91.795 4.65 ;
      RECT 91.765 3.55 91.78 4.65 ;
      RECT 91.69 3.545 91.695 3.9 ;
      RECT 91.69 3.955 91.695 4.65 ;
      RECT 91.675 3.545 91.69 3.878 ;
      RECT 91.685 3.977 91.69 4.65 ;
      RECT 91.675 4.017 91.685 4.65 ;
      RECT 91.64 3.545 91.675 3.82 ;
      RECT 91.67 4.052 91.675 4.65 ;
      RECT 91.655 4.107 91.67 4.65 ;
      RECT 91.65 4.172 91.655 4.65 ;
      RECT 91.635 4.22 91.65 4.65 ;
      RECT 91.61 3.545 91.64 3.775 ;
      RECT 91.63 4.275 91.635 4.65 ;
      RECT 91.615 4.335 91.63 4.65 ;
      RECT 91.61 4.383 91.615 4.648 ;
      RECT 91.605 3.545 91.61 3.768 ;
      RECT 91.605 4.415 91.61 4.643 ;
      RECT 91.58 3.545 91.605 3.76 ;
      RECT 91.57 3.55 91.58 3.75 ;
      RECT 91.785 4.825 91.805 5.065 ;
      RECT 91.015 4.755 91.02 4.965 ;
      RECT 92.295 4.828 92.305 5.023 ;
      RECT 92.29 4.818 92.295 5.026 ;
      RECT 92.21 4.815 92.29 5.049 ;
      RECT 92.206 4.815 92.21 5.071 ;
      RECT 92.12 4.815 92.206 5.081 ;
      RECT 92.105 4.815 92.12 5.089 ;
      RECT 92.076 4.816 92.105 5.087 ;
      RECT 91.99 4.821 92.076 5.083 ;
      RECT 91.977 4.825 91.99 5.079 ;
      RECT 91.891 4.825 91.977 5.075 ;
      RECT 91.805 4.825 91.891 5.069 ;
      RECT 91.721 4.825 91.785 5.063 ;
      RECT 91.635 4.825 91.721 5.058 ;
      RECT 91.615 4.825 91.635 5.054 ;
      RECT 91.555 4.82 91.615 5.051 ;
      RECT 91.527 4.814 91.555 5.048 ;
      RECT 91.441 4.809 91.527 5.044 ;
      RECT 91.355 4.803 91.441 5.038 ;
      RECT 91.28 4.785 91.355 5.033 ;
      RECT 91.245 4.762 91.28 5.029 ;
      RECT 91.235 4.752 91.245 5.028 ;
      RECT 91.18 4.75 91.235 5.027 ;
      RECT 91.105 4.75 91.18 5.023 ;
      RECT 91.095 4.75 91.105 5.018 ;
      RECT 91.08 4.75 91.095 5.01 ;
      RECT 91.03 4.752 91.08 4.988 ;
      RECT 91.02 4.755 91.03 4.968 ;
      RECT 91.01 4.76 91.015 4.963 ;
      RECT 91.005 4.765 91.01 4.958 ;
      RECT 91.13 3.93 91.39 4.19 ;
      RECT 91.13 3.945 91.41 4.155 ;
      RECT 91.13 3.95 91.42 4.15 ;
      RECT 89.115 3.41 89.375 3.67 ;
      RECT 89.105 3.44 89.375 3.65 ;
      RECT 91.025 3.355 91.285 3.615 ;
      RECT 91.02 3.43 91.025 3.616 ;
      RECT 90.995 3.435 91.02 3.618 ;
      RECT 90.98 3.442 90.995 3.621 ;
      RECT 90.92 3.46 90.98 3.626 ;
      RECT 90.89 3.48 90.92 3.633 ;
      RECT 90.865 3.488 90.89 3.638 ;
      RECT 90.84 3.496 90.865 3.64 ;
      RECT 90.822 3.5 90.84 3.639 ;
      RECT 90.736 3.498 90.822 3.639 ;
      RECT 90.65 3.496 90.736 3.639 ;
      RECT 90.564 3.494 90.65 3.638 ;
      RECT 90.478 3.492 90.564 3.638 ;
      RECT 90.392 3.49 90.478 3.638 ;
      RECT 90.306 3.488 90.392 3.638 ;
      RECT 90.22 3.486 90.306 3.637 ;
      RECT 90.202 3.485 90.22 3.637 ;
      RECT 90.116 3.484 90.202 3.637 ;
      RECT 90.03 3.482 90.116 3.637 ;
      RECT 89.944 3.481 90.03 3.636 ;
      RECT 89.858 3.48 89.944 3.636 ;
      RECT 89.772 3.478 89.858 3.636 ;
      RECT 89.686 3.477 89.772 3.636 ;
      RECT 89.6 3.475 89.686 3.635 ;
      RECT 89.576 3.473 89.6 3.635 ;
      RECT 89.49 3.466 89.576 3.635 ;
      RECT 89.461 3.458 89.49 3.635 ;
      RECT 89.375 3.45 89.461 3.635 ;
      RECT 89.095 3.447 89.105 3.645 ;
      RECT 90.6 4.41 90.605 4.76 ;
      RECT 90.37 4.5 90.51 4.76 ;
      RECT 90.845 4.185 90.89 4.395 ;
      RECT 90.9 4.196 90.91 4.39 ;
      RECT 90.89 4.188 90.9 4.395 ;
      RECT 90.825 4.185 90.845 4.4 ;
      RECT 90.795 4.185 90.825 4.423 ;
      RECT 90.785 4.185 90.795 4.448 ;
      RECT 90.78 4.185 90.785 4.458 ;
      RECT 90.725 4.185 90.78 4.498 ;
      RECT 90.72 4.185 90.725 4.538 ;
      RECT 90.715 4.187 90.72 4.543 ;
      RECT 90.7 4.197 90.715 4.554 ;
      RECT 90.655 4.255 90.7 4.59 ;
      RECT 90.645 4.31 90.655 4.624 ;
      RECT 90.63 4.337 90.645 4.64 ;
      RECT 90.62 4.364 90.63 4.76 ;
      RECT 90.605 4.387 90.62 4.76 ;
      RECT 90.595 4.427 90.6 4.76 ;
      RECT 90.59 4.437 90.595 4.76 ;
      RECT 90.585 4.452 90.59 4.76 ;
      RECT 90.575 4.457 90.585 4.76 ;
      RECT 90.51 4.48 90.575 4.76 ;
      RECT 90.01 3.975 90.2 4.185 ;
      RECT 88.585 3.9 88.845 4.16 ;
      RECT 88.935 3.895 89.03 4.105 ;
      RECT 88.91 3.91 88.92 4.105 ;
      RECT 90.2 3.982 90.21 4.18 ;
      RECT 90 3.982 90.01 4.18 ;
      RECT 89.985 3.997 90 4.17 ;
      RECT 89.98 4.005 89.985 4.163 ;
      RECT 89.97 4.008 89.98 4.16 ;
      RECT 89.935 4.007 89.97 4.158 ;
      RECT 89.906 4.003 89.935 4.155 ;
      RECT 89.82 3.998 89.906 4.152 ;
      RECT 89.76 3.992 89.82 4.148 ;
      RECT 89.731 3.988 89.76 4.145 ;
      RECT 89.645 3.98 89.731 4.142 ;
      RECT 89.636 3.974 89.645 4.14 ;
      RECT 89.55 3.969 89.636 4.138 ;
      RECT 89.527 3.964 89.55 4.135 ;
      RECT 89.441 3.958 89.527 4.132 ;
      RECT 89.355 3.949 89.441 4.127 ;
      RECT 89.345 3.944 89.355 4.125 ;
      RECT 89.326 3.943 89.345 4.124 ;
      RECT 89.24 3.938 89.326 4.12 ;
      RECT 89.22 3.933 89.24 4.116 ;
      RECT 89.16 3.928 89.22 4.113 ;
      RECT 89.135 3.918 89.16 4.111 ;
      RECT 89.13 3.911 89.135 4.11 ;
      RECT 89.12 3.902 89.13 4.109 ;
      RECT 89.116 3.895 89.12 4.109 ;
      RECT 89.03 3.895 89.116 4.107 ;
      RECT 88.92 3.902 88.935 4.105 ;
      RECT 88.905 3.912 88.91 4.105 ;
      RECT 88.885 3.915 88.905 4.102 ;
      RECT 88.855 3.915 88.885 4.098 ;
      RECT 88.845 3.915 88.855 4.098 ;
      RECT 89.76 4.41 90.02 4.67 ;
      RECT 89.69 4.42 90.02 4.63 ;
      RECT 89.68 4.427 90.02 4.625 ;
      RECT 89.1 4.415 89.36 4.675 ;
      RECT 89.1 4.455 89.465 4.665 ;
      RECT 89.1 4.457 89.47 4.664 ;
      RECT 89.1 4.465 89.475 4.661 ;
      RECT 88.025 3.54 88.125 5.065 ;
      RECT 88.215 4.68 88.265 4.94 ;
      RECT 88.21 3.553 88.215 3.74 ;
      RECT 88.205 4.661 88.215 4.94 ;
      RECT 88.205 3.55 88.21 3.748 ;
      RECT 88.19 3.544 88.205 3.755 ;
      RECT 88.2 4.649 88.205 5.023 ;
      RECT 88.19 4.637 88.2 5.06 ;
      RECT 88.18 3.54 88.19 3.762 ;
      RECT 88.18 4.622 88.19 5.065 ;
      RECT 88.175 3.54 88.18 3.77 ;
      RECT 88.155 4.592 88.18 5.065 ;
      RECT 88.135 3.54 88.175 3.818 ;
      RECT 88.145 4.552 88.155 5.065 ;
      RECT 88.135 4.507 88.145 5.065 ;
      RECT 88.13 3.54 88.135 3.888 ;
      RECT 88.13 4.465 88.135 5.065 ;
      RECT 88.125 3.54 88.13 4.365 ;
      RECT 88.125 4.447 88.13 5.065 ;
      RECT 88.015 3.543 88.025 5.065 ;
      RECT 88 3.55 88.015 5.061 ;
      RECT 87.995 3.56 88 5.056 ;
      RECT 87.99 3.76 87.995 4.948 ;
      RECT 87.985 3.845 87.99 4.5 ;
      RECT 86.86 10.205 87.15 10.435 ;
      RECT 86.92 8.725 87.09 10.435 ;
      RECT 86.87 9.09 87.22 9.44 ;
      RECT 86.86 8.725 87.15 8.955 ;
      RECT 86.455 3.69 86.56 4.26 ;
      RECT 86.455 4.025 86.78 4.255 ;
      RECT 86.455 4.055 86.95 4.225 ;
      RECT 86.455 3.69 86.645 4.255 ;
      RECT 85.87 3.655 86.16 3.885 ;
      RECT 85.87 3.69 86.645 3.86 ;
      RECT 85.93 2.175 86.1 3.885 ;
      RECT 85.87 2.175 86.16 2.405 ;
      RECT 85.87 10.205 86.16 10.435 ;
      RECT 85.93 8.725 86.1 10.435 ;
      RECT 85.87 8.725 86.16 8.955 ;
      RECT 85.87 8.76 86.725 8.92 ;
      RECT 86.555 8.355 86.725 8.92 ;
      RECT 85.87 8.755 86.265 8.92 ;
      RECT 86.49 8.355 86.78 8.585 ;
      RECT 86.49 8.385 86.95 8.555 ;
      RECT 85.5 4.025 85.79 4.255 ;
      RECT 85.5 4.055 85.96 4.225 ;
      RECT 85.565 2.95 85.73 4.255 ;
      RECT 84.08 2.92 84.37 3.15 ;
      RECT 84.08 2.95 85.73 3.12 ;
      RECT 84.14 2.18 84.31 3.15 ;
      RECT 84.08 2.18 84.37 2.41 ;
      RECT 84.08 10.2 84.37 10.43 ;
      RECT 84.14 9.46 84.31 10.43 ;
      RECT 84.14 9.555 85.73 9.725 ;
      RECT 85.56 8.355 85.73 9.725 ;
      RECT 84.08 9.46 84.37 9.69 ;
      RECT 85.5 8.355 85.79 8.585 ;
      RECT 85.5 8.385 85.96 8.555 ;
      RECT 82.115 4.725 82.465 5.075 ;
      RECT 82.205 3.32 82.375 5.075 ;
      RECT 84.51 3.26 84.86 3.61 ;
      RECT 82.205 3.32 83.825 3.495 ;
      RECT 82.205 3.32 84.86 3.49 ;
      RECT 84.535 9.09 84.86 9.415 ;
      RECT 79.91 9.045 80.26 9.395 ;
      RECT 84.51 9.09 84.86 9.32 ;
      RECT 79.75 9.09 80.26 9.32 ;
      RECT 79.58 9.12 84.86 9.29 ;
      RECT 83.735 3.66 84.055 3.98 ;
      RECT 83.705 3.66 84.055 3.89 ;
      RECT 83.535 3.69 84.055 3.86 ;
      RECT 83.735 8.66 84.055 8.98 ;
      RECT 83.705 8.72 84.055 8.95 ;
      RECT 83.535 8.75 84.055 8.92 ;
      RECT 79.515 4.96 79.555 5.22 ;
      RECT 79.555 4.94 79.56 4.95 ;
      RECT 80.885 4.185 80.895 4.406 ;
      RECT 80.815 4.18 80.885 4.531 ;
      RECT 80.805 4.18 80.815 4.658 ;
      RECT 80.78 4.18 80.805 4.705 ;
      RECT 80.755 4.18 80.78 4.783 ;
      RECT 80.735 4.18 80.755 4.853 ;
      RECT 80.71 4.18 80.735 4.893 ;
      RECT 80.7 4.18 80.71 4.913 ;
      RECT 80.69 4.182 80.7 4.921 ;
      RECT 80.685 4.187 80.69 4.378 ;
      RECT 80.685 4.387 80.69 4.922 ;
      RECT 80.68 4.432 80.685 4.923 ;
      RECT 80.67 4.497 80.68 4.924 ;
      RECT 80.66 4.592 80.67 4.926 ;
      RECT 80.655 4.645 80.66 4.928 ;
      RECT 80.65 4.665 80.655 4.929 ;
      RECT 80.595 4.69 80.65 4.935 ;
      RECT 80.555 4.725 80.595 4.944 ;
      RECT 80.545 4.742 80.555 4.949 ;
      RECT 80.536 4.748 80.545 4.951 ;
      RECT 80.45 4.786 80.536 4.962 ;
      RECT 80.445 4.825 80.45 4.972 ;
      RECT 80.37 4.832 80.445 4.982 ;
      RECT 80.35 4.842 80.37 4.993 ;
      RECT 80.32 4.849 80.35 5.001 ;
      RECT 80.295 4.856 80.32 5.008 ;
      RECT 80.271 4.862 80.295 5.013 ;
      RECT 80.185 4.875 80.271 5.025 ;
      RECT 80.107 4.882 80.185 5.043 ;
      RECT 80.021 4.877 80.107 5.061 ;
      RECT 79.935 4.872 80.021 5.081 ;
      RECT 79.855 4.866 79.935 5.098 ;
      RECT 79.79 4.862 79.855 5.127 ;
      RECT 79.785 4.576 79.79 4.6 ;
      RECT 79.775 4.852 79.79 5.155 ;
      RECT 79.78 4.57 79.785 4.64 ;
      RECT 79.775 4.564 79.78 4.71 ;
      RECT 79.77 4.558 79.775 4.788 ;
      RECT 79.77 4.835 79.775 5.22 ;
      RECT 79.762 4.555 79.77 5.22 ;
      RECT 79.676 4.553 79.762 5.22 ;
      RECT 79.59 4.551 79.676 5.22 ;
      RECT 79.58 4.552 79.59 5.22 ;
      RECT 79.575 4.557 79.58 5.22 ;
      RECT 79.565 4.57 79.575 5.22 ;
      RECT 79.56 4.592 79.565 5.22 ;
      RECT 79.555 4.952 79.56 5.22 ;
      RECT 80.185 4.42 80.19 4.64 ;
      RECT 80.69 3.455 80.725 3.715 ;
      RECT 80.675 3.455 80.69 3.723 ;
      RECT 80.646 3.455 80.675 3.745 ;
      RECT 80.56 3.455 80.646 3.805 ;
      RECT 80.54 3.455 80.56 3.87 ;
      RECT 80.48 3.455 80.54 4.035 ;
      RECT 80.475 3.455 80.48 4.183 ;
      RECT 80.47 3.455 80.475 4.195 ;
      RECT 80.465 3.455 80.47 4.221 ;
      RECT 80.435 3.641 80.465 4.301 ;
      RECT 80.43 3.689 80.435 4.39 ;
      RECT 80.425 3.703 80.43 4.405 ;
      RECT 80.42 3.722 80.425 4.435 ;
      RECT 80.415 3.737 80.42 4.451 ;
      RECT 80.41 3.752 80.415 4.473 ;
      RECT 80.405 3.772 80.41 4.495 ;
      RECT 80.395 3.792 80.405 4.528 ;
      RECT 80.38 3.834 80.395 4.59 ;
      RECT 80.375 3.865 80.38 4.63 ;
      RECT 80.37 3.877 80.375 4.635 ;
      RECT 80.365 3.889 80.37 4.64 ;
      RECT 80.36 3.902 80.365 4.64 ;
      RECT 80.355 3.92 80.36 4.64 ;
      RECT 80.35 3.94 80.355 4.64 ;
      RECT 80.345 3.952 80.35 4.64 ;
      RECT 80.34 3.965 80.345 4.64 ;
      RECT 80.32 4 80.34 4.64 ;
      RECT 80.27 4.102 80.32 4.64 ;
      RECT 80.265 4.187 80.27 4.64 ;
      RECT 80.26 4.195 80.265 4.64 ;
      RECT 80.255 4.212 80.26 4.64 ;
      RECT 80.25 4.227 80.255 4.64 ;
      RECT 80.215 4.292 80.25 4.64 ;
      RECT 80.2 4.357 80.215 4.64 ;
      RECT 80.195 4.387 80.2 4.64 ;
      RECT 80.19 4.412 80.195 4.64 ;
      RECT 80.175 4.422 80.185 4.64 ;
      RECT 80.16 4.435 80.175 4.633 ;
      RECT 79.905 4.025 79.975 4.235 ;
      RECT 79.695 4.002 79.7 4.195 ;
      RECT 77.15 3.93 77.41 4.19 ;
      RECT 79.985 4.212 79.99 4.215 ;
      RECT 79.975 4.03 79.985 4.23 ;
      RECT 79.876 4.023 79.905 4.235 ;
      RECT 79.79 4.015 79.876 4.235 ;
      RECT 79.775 4.009 79.79 4.233 ;
      RECT 79.755 4.008 79.775 4.22 ;
      RECT 79.75 4.007 79.755 4.203 ;
      RECT 79.7 4.004 79.75 4.198 ;
      RECT 79.67 4.001 79.695 4.193 ;
      RECT 79.65 3.999 79.67 4.188 ;
      RECT 79.635 3.997 79.65 4.185 ;
      RECT 79.605 3.995 79.635 4.183 ;
      RECT 79.54 3.991 79.605 4.175 ;
      RECT 79.51 3.986 79.54 4.17 ;
      RECT 79.49 3.984 79.51 4.168 ;
      RECT 79.46 3.981 79.49 4.163 ;
      RECT 79.4 3.977 79.46 4.155 ;
      RECT 79.395 3.974 79.4 4.15 ;
      RECT 79.325 3.972 79.395 4.145 ;
      RECT 79.296 3.968 79.325 4.138 ;
      RECT 79.21 3.963 79.296 4.13 ;
      RECT 79.176 3.958 79.21 4.122 ;
      RECT 79.09 3.95 79.176 4.114 ;
      RECT 79.051 3.943 79.09 4.106 ;
      RECT 78.965 3.938 79.051 4.098 ;
      RECT 78.9 3.932 78.965 4.088 ;
      RECT 78.88 3.927 78.9 4.083 ;
      RECT 78.871 3.924 78.88 4.082 ;
      RECT 78.785 3.92 78.871 4.076 ;
      RECT 78.745 3.916 78.785 4.068 ;
      RECT 78.725 3.912 78.745 4.066 ;
      RECT 78.665 3.912 78.725 4.063 ;
      RECT 78.645 3.915 78.665 4.061 ;
      RECT 78.624 3.915 78.645 4.061 ;
      RECT 78.538 3.917 78.624 4.065 ;
      RECT 78.452 3.919 78.538 4.071 ;
      RECT 78.366 3.921 78.452 4.078 ;
      RECT 78.28 3.924 78.366 4.084 ;
      RECT 78.246 3.925 78.28 4.089 ;
      RECT 78.16 3.928 78.246 4.094 ;
      RECT 78.131 3.935 78.16 4.099 ;
      RECT 78.045 3.935 78.131 4.104 ;
      RECT 78.012 3.935 78.045 4.109 ;
      RECT 77.926 3.937 78.012 4.114 ;
      RECT 77.84 3.939 77.926 4.121 ;
      RECT 77.776 3.941 77.84 4.127 ;
      RECT 77.69 3.943 77.776 4.133 ;
      RECT 77.687 3.945 77.69 4.136 ;
      RECT 77.601 3.946 77.687 4.14 ;
      RECT 77.515 3.949 77.601 4.147 ;
      RECT 77.496 3.951 77.515 4.151 ;
      RECT 77.41 3.953 77.496 4.156 ;
      RECT 77.14 3.965 77.15 4.16 ;
      RECT 79.32 10.2 79.61 10.43 ;
      RECT 79.38 9.46 79.55 10.43 ;
      RECT 79.27 9.49 79.645 9.86 ;
      RECT 79.32 9.46 79.61 9.86 ;
      RECT 79.375 3.545 79.56 3.755 ;
      RECT 79.37 3.546 79.565 3.753 ;
      RECT 79.365 3.551 79.575 3.748 ;
      RECT 79.36 3.527 79.365 3.745 ;
      RECT 79.33 3.524 79.36 3.738 ;
      RECT 79.325 3.52 79.33 3.729 ;
      RECT 79.29 3.551 79.575 3.724 ;
      RECT 79.065 3.46 79.325 3.72 ;
      RECT 79.365 3.529 79.37 3.748 ;
      RECT 79.37 3.53 79.375 3.753 ;
      RECT 79.065 3.542 79.445 3.72 ;
      RECT 79.065 3.54 79.43 3.72 ;
      RECT 79.065 3.535 79.42 3.72 ;
      RECT 79.02 4.45 79.07 4.735 ;
      RECT 78.965 4.42 78.97 4.735 ;
      RECT 78.935 4.4 78.94 4.735 ;
      RECT 79.085 4.45 79.145 4.71 ;
      RECT 79.08 4.45 79.085 4.718 ;
      RECT 79.07 4.45 79.08 4.73 ;
      RECT 78.985 4.44 79.02 4.735 ;
      RECT 78.98 4.427 78.985 4.735 ;
      RECT 78.97 4.422 78.98 4.735 ;
      RECT 78.95 4.412 78.965 4.735 ;
      RECT 78.94 4.405 78.95 4.735 ;
      RECT 78.93 4.397 78.935 4.735 ;
      RECT 78.9 4.387 78.93 4.735 ;
      RECT 78.885 4.375 78.9 4.735 ;
      RECT 78.87 4.365 78.885 4.73 ;
      RECT 78.85 4.355 78.87 4.705 ;
      RECT 78.84 4.347 78.85 4.682 ;
      RECT 78.81 4.33 78.84 4.672 ;
      RECT 78.805 4.307 78.81 4.663 ;
      RECT 78.8 4.294 78.805 4.661 ;
      RECT 78.785 4.27 78.8 4.655 ;
      RECT 78.78 4.246 78.785 4.649 ;
      RECT 78.77 4.235 78.78 4.644 ;
      RECT 78.765 4.225 78.77 4.64 ;
      RECT 78.76 4.217 78.765 4.637 ;
      RECT 78.75 4.212 78.76 4.633 ;
      RECT 78.745 4.207 78.75 4.629 ;
      RECT 78.66 4.205 78.745 4.604 ;
      RECT 78.63 4.205 78.66 4.57 ;
      RECT 78.615 4.205 78.63 4.553 ;
      RECT 78.56 4.205 78.615 4.498 ;
      RECT 78.555 4.21 78.56 4.447 ;
      RECT 78.545 4.215 78.555 4.437 ;
      RECT 78.54 4.225 78.545 4.423 ;
      RECT 78.49 4.965 78.75 5.225 ;
      RECT 78.41 4.98 78.75 5.201 ;
      RECT 78.39 4.98 78.75 5.196 ;
      RECT 78.366 4.98 78.75 5.194 ;
      RECT 78.28 4.98 78.75 5.189 ;
      RECT 78.13 4.92 78.39 5.185 ;
      RECT 78.085 4.98 78.75 5.18 ;
      RECT 78.08 4.987 78.75 5.175 ;
      RECT 78.095 4.975 78.41 5.185 ;
      RECT 77.985 3.41 78.245 3.67 ;
      RECT 77.985 3.467 78.25 3.663 ;
      RECT 77.985 3.497 78.255 3.595 ;
      RECT 78.045 3.928 78.16 3.93 ;
      RECT 78.131 3.925 78.16 3.93 ;
      RECT 77.155 4.929 77.18 5.169 ;
      RECT 77.14 4.932 77.23 5.163 ;
      RECT 77.135 4.937 77.316 5.158 ;
      RECT 77.13 4.945 77.38 5.156 ;
      RECT 77.13 4.945 77.39 5.155 ;
      RECT 77.125 4.952 77.4 5.148 ;
      RECT 77.125 4.952 77.486 5.137 ;
      RECT 77.12 4.987 77.486 5.133 ;
      RECT 77.12 4.987 77.495 5.122 ;
      RECT 77.4 4.86 77.66 5.12 ;
      RECT 77.11 5.037 77.66 5.118 ;
      RECT 77.38 4.905 77.4 5.153 ;
      RECT 77.316 4.908 77.38 5.157 ;
      RECT 77.23 4.913 77.316 5.162 ;
      RECT 77.16 4.924 77.66 5.12 ;
      RECT 77.18 4.918 77.23 5.167 ;
      RECT 77.305 3.395 77.315 3.657 ;
      RECT 77.295 3.452 77.305 3.66 ;
      RECT 77.27 3.457 77.295 3.666 ;
      RECT 77.245 3.461 77.27 3.678 ;
      RECT 77.235 3.464 77.245 3.688 ;
      RECT 77.23 3.465 77.235 3.693 ;
      RECT 77.225 3.466 77.23 3.698 ;
      RECT 77.22 3.467 77.225 3.7 ;
      RECT 77.195 3.47 77.22 3.703 ;
      RECT 77.165 3.476 77.195 3.706 ;
      RECT 77.1 3.487 77.165 3.709 ;
      RECT 77.055 3.495 77.1 3.713 ;
      RECT 77.04 3.495 77.055 3.721 ;
      RECT 77.035 3.496 77.04 3.728 ;
      RECT 77.03 3.498 77.035 3.731 ;
      RECT 77.025 3.502 77.03 3.734 ;
      RECT 77.015 3.51 77.025 3.738 ;
      RECT 77.01 3.523 77.015 3.743 ;
      RECT 77.005 3.531 77.01 3.745 ;
      RECT 77 3.537 77.005 3.745 ;
      RECT 76.995 3.541 77 3.748 ;
      RECT 76.99 3.543 76.995 3.751 ;
      RECT 76.985 3.546 76.99 3.754 ;
      RECT 76.975 3.551 76.985 3.758 ;
      RECT 76.97 3.557 76.975 3.763 ;
      RECT 76.96 3.563 76.97 3.767 ;
      RECT 76.945 3.57 76.96 3.773 ;
      RECT 76.916 3.584 76.945 3.783 ;
      RECT 76.83 3.619 76.916 3.815 ;
      RECT 76.81 3.652 76.83 3.844 ;
      RECT 76.79 3.665 76.81 3.855 ;
      RECT 76.77 3.677 76.79 3.866 ;
      RECT 76.72 3.699 76.77 3.886 ;
      RECT 76.705 3.717 76.72 3.903 ;
      RECT 76.7 3.723 76.705 3.906 ;
      RECT 76.695 3.727 76.7 3.909 ;
      RECT 76.69 3.731 76.695 3.913 ;
      RECT 76.685 3.733 76.69 3.916 ;
      RECT 76.675 3.74 76.685 3.919 ;
      RECT 76.67 3.745 76.675 3.923 ;
      RECT 76.665 3.747 76.67 3.926 ;
      RECT 76.66 3.751 76.665 3.929 ;
      RECT 76.655 3.753 76.66 3.933 ;
      RECT 76.64 3.758 76.655 3.938 ;
      RECT 76.635 3.763 76.64 3.941 ;
      RECT 76.63 3.771 76.635 3.944 ;
      RECT 76.625 3.773 76.63 3.947 ;
      RECT 76.62 3.775 76.625 3.95 ;
      RECT 76.61 3.777 76.62 3.956 ;
      RECT 76.575 3.791 76.61 3.968 ;
      RECT 76.565 3.806 76.575 3.978 ;
      RECT 76.49 3.835 76.565 4.002 ;
      RECT 76.485 3.86 76.49 4.025 ;
      RECT 76.47 3.864 76.485 4.031 ;
      RECT 76.46 3.872 76.47 4.036 ;
      RECT 76.43 3.885 76.46 4.04 ;
      RECT 76.42 3.9 76.43 4.045 ;
      RECT 76.41 3.905 76.42 4.048 ;
      RECT 76.405 3.907 76.41 4.05 ;
      RECT 76.39 3.91 76.405 4.053 ;
      RECT 76.385 3.912 76.39 4.056 ;
      RECT 76.365 3.917 76.385 4.06 ;
      RECT 76.335 3.922 76.365 4.068 ;
      RECT 76.31 3.929 76.335 4.076 ;
      RECT 76.305 3.934 76.31 4.081 ;
      RECT 76.275 3.937 76.305 4.085 ;
      RECT 76.235 3.94 76.275 4.095 ;
      RECT 76.2 3.937 76.235 4.107 ;
      RECT 76.19 3.933 76.2 4.114 ;
      RECT 76.165 3.929 76.19 4.12 ;
      RECT 76.16 3.925 76.165 4.125 ;
      RECT 76.12 3.922 76.16 4.125 ;
      RECT 76.105 3.907 76.12 4.126 ;
      RECT 76.082 3.895 76.105 4.126 ;
      RECT 75.996 3.895 76.082 4.127 ;
      RECT 75.91 3.895 75.996 4.129 ;
      RECT 75.89 3.895 75.91 4.126 ;
      RECT 75.885 3.9 75.89 4.121 ;
      RECT 75.88 3.905 75.885 4.119 ;
      RECT 75.87 3.915 75.88 4.117 ;
      RECT 75.865 3.921 75.87 4.11 ;
      RECT 75.86 3.923 75.865 4.095 ;
      RECT 75.855 3.927 75.86 4.085 ;
      RECT 77.315 3.395 77.565 3.655 ;
      RECT 75.04 4.93 75.3 5.19 ;
      RECT 77.335 4.42 77.34 4.63 ;
      RECT 77.34 4.425 77.35 4.625 ;
      RECT 77.29 4.42 77.335 4.645 ;
      RECT 77.28 4.42 77.29 4.665 ;
      RECT 77.261 4.42 77.28 4.67 ;
      RECT 77.175 4.42 77.261 4.667 ;
      RECT 77.145 4.422 77.175 4.665 ;
      RECT 77.09 4.432 77.145 4.663 ;
      RECT 77.025 4.446 77.09 4.661 ;
      RECT 77.02 4.454 77.025 4.66 ;
      RECT 77.005 4.457 77.02 4.658 ;
      RECT 76.94 4.467 77.005 4.654 ;
      RECT 76.892 4.481 76.94 4.655 ;
      RECT 76.806 4.498 76.892 4.669 ;
      RECT 76.72 4.519 76.806 4.686 ;
      RECT 76.7 4.532 76.72 4.696 ;
      RECT 76.655 4.54 76.7 4.703 ;
      RECT 76.62 4.548 76.655 4.711 ;
      RECT 76.586 4.556 76.62 4.719 ;
      RECT 76.5 4.57 76.586 4.731 ;
      RECT 76.465 4.587 76.5 4.743 ;
      RECT 76.456 4.596 76.465 4.747 ;
      RECT 76.37 4.614 76.456 4.764 ;
      RECT 76.311 4.641 76.37 4.791 ;
      RECT 76.225 4.668 76.311 4.819 ;
      RECT 76.205 4.69 76.225 4.839 ;
      RECT 76.145 4.705 76.205 4.855 ;
      RECT 76.135 4.717 76.145 4.868 ;
      RECT 76.13 4.722 76.135 4.871 ;
      RECT 76.12 4.725 76.13 4.874 ;
      RECT 76.115 4.727 76.12 4.877 ;
      RECT 76.085 4.735 76.115 4.884 ;
      RECT 76.07 4.742 76.085 4.892 ;
      RECT 76.06 4.747 76.07 4.896 ;
      RECT 76.055 4.75 76.06 4.899 ;
      RECT 76.045 4.752 76.055 4.902 ;
      RECT 76.01 4.762 76.045 4.911 ;
      RECT 75.935 4.785 76.01 4.933 ;
      RECT 75.915 4.803 75.935 4.951 ;
      RECT 75.885 4.81 75.915 4.961 ;
      RECT 75.865 4.818 75.885 4.971 ;
      RECT 75.855 4.824 75.865 4.978 ;
      RECT 75.836 4.829 75.855 4.984 ;
      RECT 75.75 4.849 75.836 5.004 ;
      RECT 75.735 4.869 75.75 5.023 ;
      RECT 75.69 4.881 75.735 5.034 ;
      RECT 75.625 4.902 75.69 5.057 ;
      RECT 75.585 4.922 75.625 5.078 ;
      RECT 75.575 4.932 75.585 5.088 ;
      RECT 75.525 4.944 75.575 5.099 ;
      RECT 75.505 4.96 75.525 5.111 ;
      RECT 75.475 4.97 75.505 5.117 ;
      RECT 75.465 4.975 75.475 5.119 ;
      RECT 75.396 4.976 75.465 5.125 ;
      RECT 75.31 4.978 75.396 5.135 ;
      RECT 75.3 4.979 75.31 5.14 ;
      RECT 76.57 5.005 76.76 5.215 ;
      RECT 76.56 5.01 76.77 5.208 ;
      RECT 76.545 5.01 76.77 5.173 ;
      RECT 76.465 4.895 76.725 5.155 ;
      RECT 75.38 4.425 75.565 4.72 ;
      RECT 75.37 4.425 75.565 4.718 ;
      RECT 75.355 4.425 75.57 4.713 ;
      RECT 75.355 4.425 75.575 4.71 ;
      RECT 75.35 4.425 75.575 4.708 ;
      RECT 75.345 4.68 75.575 4.698 ;
      RECT 75.35 4.425 75.61 4.685 ;
      RECT 75.31 3.46 75.57 3.72 ;
      RECT 75.12 3.385 75.206 3.718 ;
      RECT 75.095 3.389 75.25 3.714 ;
      RECT 75.206 3.381 75.25 3.714 ;
      RECT 75.206 3.382 75.255 3.713 ;
      RECT 75.12 3.387 75.27 3.712 ;
      RECT 75.095 3.395 75.31 3.711 ;
      RECT 75.09 3.39 75.27 3.706 ;
      RECT 75.08 3.405 75.31 3.613 ;
      RECT 75.08 3.457 75.51 3.613 ;
      RECT 75.08 3.45 75.49 3.613 ;
      RECT 75.08 3.437 75.46 3.613 ;
      RECT 75.08 3.425 75.4 3.613 ;
      RECT 75.08 3.41 75.375 3.613 ;
      RECT 74.28 4.04 74.415 4.335 ;
      RECT 74.54 4.063 74.545 4.25 ;
      RECT 75.26 3.96 75.405 4.195 ;
      RECT 75.42 3.96 75.425 4.185 ;
      RECT 75.455 3.971 75.46 4.165 ;
      RECT 75.45 3.963 75.455 4.17 ;
      RECT 75.43 3.96 75.45 4.175 ;
      RECT 75.425 3.96 75.43 4.183 ;
      RECT 75.415 3.96 75.42 4.188 ;
      RECT 75.405 3.96 75.415 4.193 ;
      RECT 75.235 3.962 75.26 4.195 ;
      RECT 75.185 3.969 75.235 4.195 ;
      RECT 75.18 3.974 75.185 4.195 ;
      RECT 75.141 3.979 75.18 4.196 ;
      RECT 75.055 3.991 75.141 4.197 ;
      RECT 75.046 4.001 75.055 4.197 ;
      RECT 74.96 4.01 75.046 4.199 ;
      RECT 74.936 4.02 74.96 4.201 ;
      RECT 74.85 4.031 74.936 4.202 ;
      RECT 74.82 4.042 74.85 4.204 ;
      RECT 74.79 4.047 74.82 4.206 ;
      RECT 74.765 4.053 74.79 4.209 ;
      RECT 74.75 4.058 74.765 4.21 ;
      RECT 74.705 4.064 74.75 4.21 ;
      RECT 74.7 4.069 74.705 4.211 ;
      RECT 74.68 4.069 74.7 4.213 ;
      RECT 74.66 4.067 74.68 4.218 ;
      RECT 74.625 4.066 74.66 4.225 ;
      RECT 74.595 4.065 74.625 4.235 ;
      RECT 74.545 4.064 74.595 4.245 ;
      RECT 74.455 4.061 74.54 4.335 ;
      RECT 74.43 4.055 74.455 4.335 ;
      RECT 74.415 4.045 74.43 4.335 ;
      RECT 74.23 4.04 74.28 4.255 ;
      RECT 74.22 4.045 74.23 4.245 ;
      RECT 74.46 4.52 74.72 4.78 ;
      RECT 74.46 4.52 74.75 4.673 ;
      RECT 74.46 4.52 74.785 4.658 ;
      RECT 74.715 4.44 74.905 4.65 ;
      RECT 74.705 4.445 74.915 4.643 ;
      RECT 74.67 4.515 74.915 4.643 ;
      RECT 74.7 4.457 74.72 4.78 ;
      RECT 74.685 4.505 74.915 4.643 ;
      RECT 74.69 4.477 74.72 4.78 ;
      RECT 73.77 3.545 73.84 4.65 ;
      RECT 74.505 3.65 74.765 3.91 ;
      RECT 74.085 3.696 74.1 3.905 ;
      RECT 74.421 3.709 74.505 3.86 ;
      RECT 74.335 3.706 74.421 3.86 ;
      RECT 74.296 3.704 74.335 3.86 ;
      RECT 74.21 3.702 74.296 3.86 ;
      RECT 74.15 3.7 74.21 3.871 ;
      RECT 74.115 3.698 74.15 3.889 ;
      RECT 74.1 3.696 74.115 3.9 ;
      RECT 74.07 3.696 74.085 3.913 ;
      RECT 74.06 3.696 74.07 3.918 ;
      RECT 74.035 3.695 74.06 3.923 ;
      RECT 74.02 3.69 74.035 3.929 ;
      RECT 74.015 3.683 74.02 3.934 ;
      RECT 73.99 3.674 74.015 3.94 ;
      RECT 73.945 3.653 73.99 3.953 ;
      RECT 73.935 3.637 73.945 3.963 ;
      RECT 73.92 3.63 73.935 3.973 ;
      RECT 73.91 3.623 73.92 3.99 ;
      RECT 73.905 3.62 73.91 4.02 ;
      RECT 73.9 3.618 73.905 4.05 ;
      RECT 73.895 3.616 73.9 4.087 ;
      RECT 73.88 3.612 73.895 4.154 ;
      RECT 73.88 4.445 73.89 4.645 ;
      RECT 73.875 3.608 73.88 4.28 ;
      RECT 73.875 4.432 73.88 4.65 ;
      RECT 73.87 3.606 73.875 4.365 ;
      RECT 73.87 4.422 73.875 4.65 ;
      RECT 73.855 3.577 73.87 4.65 ;
      RECT 73.84 3.55 73.855 4.65 ;
      RECT 73.765 3.545 73.77 3.9 ;
      RECT 73.765 3.955 73.77 4.65 ;
      RECT 73.75 3.545 73.765 3.878 ;
      RECT 73.76 3.977 73.765 4.65 ;
      RECT 73.75 4.017 73.76 4.65 ;
      RECT 73.715 3.545 73.75 3.82 ;
      RECT 73.745 4.052 73.75 4.65 ;
      RECT 73.73 4.107 73.745 4.65 ;
      RECT 73.725 4.172 73.73 4.65 ;
      RECT 73.71 4.22 73.725 4.65 ;
      RECT 73.685 3.545 73.715 3.775 ;
      RECT 73.705 4.275 73.71 4.65 ;
      RECT 73.69 4.335 73.705 4.65 ;
      RECT 73.685 4.383 73.69 4.648 ;
      RECT 73.68 3.545 73.685 3.768 ;
      RECT 73.68 4.415 73.685 4.643 ;
      RECT 73.655 3.545 73.68 3.76 ;
      RECT 73.645 3.55 73.655 3.75 ;
      RECT 73.86 4.825 73.88 5.065 ;
      RECT 73.09 4.755 73.095 4.965 ;
      RECT 74.37 4.828 74.38 5.023 ;
      RECT 74.365 4.818 74.37 5.026 ;
      RECT 74.285 4.815 74.365 5.049 ;
      RECT 74.281 4.815 74.285 5.071 ;
      RECT 74.195 4.815 74.281 5.081 ;
      RECT 74.18 4.815 74.195 5.089 ;
      RECT 74.151 4.816 74.18 5.087 ;
      RECT 74.065 4.821 74.151 5.083 ;
      RECT 74.052 4.825 74.065 5.079 ;
      RECT 73.966 4.825 74.052 5.075 ;
      RECT 73.88 4.825 73.966 5.069 ;
      RECT 73.796 4.825 73.86 5.063 ;
      RECT 73.71 4.825 73.796 5.058 ;
      RECT 73.69 4.825 73.71 5.054 ;
      RECT 73.63 4.82 73.69 5.051 ;
      RECT 73.602 4.814 73.63 5.048 ;
      RECT 73.516 4.809 73.602 5.044 ;
      RECT 73.43 4.803 73.516 5.038 ;
      RECT 73.355 4.785 73.43 5.033 ;
      RECT 73.32 4.762 73.355 5.029 ;
      RECT 73.31 4.752 73.32 5.028 ;
      RECT 73.255 4.75 73.31 5.027 ;
      RECT 73.18 4.75 73.255 5.023 ;
      RECT 73.17 4.75 73.18 5.018 ;
      RECT 73.155 4.75 73.17 5.01 ;
      RECT 73.105 4.752 73.155 4.988 ;
      RECT 73.095 4.755 73.105 4.968 ;
      RECT 73.085 4.76 73.09 4.963 ;
      RECT 73.08 4.765 73.085 4.958 ;
      RECT 73.205 3.93 73.465 4.19 ;
      RECT 73.205 3.945 73.485 4.155 ;
      RECT 73.205 3.95 73.495 4.15 ;
      RECT 71.19 3.41 71.45 3.67 ;
      RECT 71.18 3.44 71.45 3.65 ;
      RECT 73.1 3.355 73.36 3.615 ;
      RECT 73.095 3.43 73.1 3.616 ;
      RECT 73.07 3.435 73.095 3.618 ;
      RECT 73.055 3.442 73.07 3.621 ;
      RECT 72.995 3.46 73.055 3.626 ;
      RECT 72.965 3.48 72.995 3.633 ;
      RECT 72.94 3.488 72.965 3.638 ;
      RECT 72.915 3.496 72.94 3.64 ;
      RECT 72.897 3.5 72.915 3.639 ;
      RECT 72.811 3.498 72.897 3.639 ;
      RECT 72.725 3.496 72.811 3.639 ;
      RECT 72.639 3.494 72.725 3.638 ;
      RECT 72.553 3.492 72.639 3.638 ;
      RECT 72.467 3.49 72.553 3.638 ;
      RECT 72.381 3.488 72.467 3.638 ;
      RECT 72.295 3.486 72.381 3.637 ;
      RECT 72.277 3.485 72.295 3.637 ;
      RECT 72.191 3.484 72.277 3.637 ;
      RECT 72.105 3.482 72.191 3.637 ;
      RECT 72.019 3.481 72.105 3.636 ;
      RECT 71.933 3.48 72.019 3.636 ;
      RECT 71.847 3.478 71.933 3.636 ;
      RECT 71.761 3.477 71.847 3.636 ;
      RECT 71.675 3.475 71.761 3.635 ;
      RECT 71.651 3.473 71.675 3.635 ;
      RECT 71.565 3.466 71.651 3.635 ;
      RECT 71.536 3.458 71.565 3.635 ;
      RECT 71.45 3.45 71.536 3.635 ;
      RECT 71.17 3.447 71.18 3.645 ;
      RECT 72.675 4.41 72.68 4.76 ;
      RECT 72.445 4.5 72.585 4.76 ;
      RECT 72.92 4.185 72.965 4.395 ;
      RECT 72.975 4.196 72.985 4.39 ;
      RECT 72.965 4.188 72.975 4.395 ;
      RECT 72.9 4.185 72.92 4.4 ;
      RECT 72.87 4.185 72.9 4.423 ;
      RECT 72.86 4.185 72.87 4.448 ;
      RECT 72.855 4.185 72.86 4.458 ;
      RECT 72.8 4.185 72.855 4.498 ;
      RECT 72.795 4.185 72.8 4.538 ;
      RECT 72.79 4.187 72.795 4.543 ;
      RECT 72.775 4.197 72.79 4.554 ;
      RECT 72.73 4.255 72.775 4.59 ;
      RECT 72.72 4.31 72.73 4.624 ;
      RECT 72.705 4.337 72.72 4.64 ;
      RECT 72.695 4.364 72.705 4.76 ;
      RECT 72.68 4.387 72.695 4.76 ;
      RECT 72.67 4.427 72.675 4.76 ;
      RECT 72.665 4.437 72.67 4.76 ;
      RECT 72.66 4.452 72.665 4.76 ;
      RECT 72.65 4.457 72.66 4.76 ;
      RECT 72.585 4.48 72.65 4.76 ;
      RECT 72.085 3.975 72.275 4.185 ;
      RECT 70.66 3.9 70.92 4.16 ;
      RECT 71.01 3.895 71.105 4.105 ;
      RECT 70.985 3.91 70.995 4.105 ;
      RECT 72.275 3.982 72.285 4.18 ;
      RECT 72.075 3.982 72.085 4.18 ;
      RECT 72.06 3.997 72.075 4.17 ;
      RECT 72.055 4.005 72.06 4.163 ;
      RECT 72.045 4.008 72.055 4.16 ;
      RECT 72.01 4.007 72.045 4.158 ;
      RECT 71.981 4.003 72.01 4.155 ;
      RECT 71.895 3.998 71.981 4.152 ;
      RECT 71.835 3.992 71.895 4.148 ;
      RECT 71.806 3.988 71.835 4.145 ;
      RECT 71.72 3.98 71.806 4.142 ;
      RECT 71.711 3.974 71.72 4.14 ;
      RECT 71.625 3.969 71.711 4.138 ;
      RECT 71.602 3.964 71.625 4.135 ;
      RECT 71.516 3.958 71.602 4.132 ;
      RECT 71.43 3.949 71.516 4.127 ;
      RECT 71.42 3.944 71.43 4.125 ;
      RECT 71.401 3.943 71.42 4.124 ;
      RECT 71.315 3.938 71.401 4.12 ;
      RECT 71.295 3.933 71.315 4.116 ;
      RECT 71.235 3.928 71.295 4.113 ;
      RECT 71.21 3.918 71.235 4.111 ;
      RECT 71.205 3.911 71.21 4.11 ;
      RECT 71.195 3.902 71.205 4.109 ;
      RECT 71.191 3.895 71.195 4.109 ;
      RECT 71.105 3.895 71.191 4.107 ;
      RECT 70.995 3.902 71.01 4.105 ;
      RECT 70.98 3.912 70.985 4.105 ;
      RECT 70.96 3.915 70.98 4.102 ;
      RECT 70.93 3.915 70.96 4.098 ;
      RECT 70.92 3.915 70.93 4.098 ;
      RECT 71.835 4.41 72.095 4.67 ;
      RECT 71.765 4.42 72.095 4.63 ;
      RECT 71.755 4.427 72.095 4.625 ;
      RECT 71.175 4.415 71.435 4.675 ;
      RECT 71.175 4.455 71.54 4.665 ;
      RECT 71.175 4.457 71.545 4.664 ;
      RECT 71.175 4.465 71.55 4.661 ;
      RECT 70.1 3.54 70.2 5.065 ;
      RECT 70.29 4.68 70.34 4.94 ;
      RECT 70.285 3.553 70.29 3.74 ;
      RECT 70.28 4.661 70.29 4.94 ;
      RECT 70.28 3.55 70.285 3.748 ;
      RECT 70.265 3.544 70.28 3.755 ;
      RECT 70.275 4.649 70.28 5.023 ;
      RECT 70.265 4.637 70.275 5.06 ;
      RECT 70.255 3.54 70.265 3.762 ;
      RECT 70.255 4.622 70.265 5.065 ;
      RECT 70.25 3.54 70.255 3.77 ;
      RECT 70.23 4.592 70.255 5.065 ;
      RECT 70.21 3.54 70.25 3.818 ;
      RECT 70.22 4.552 70.23 5.065 ;
      RECT 70.21 4.507 70.22 5.065 ;
      RECT 70.205 3.54 70.21 3.888 ;
      RECT 70.205 4.465 70.21 5.065 ;
      RECT 70.2 3.54 70.205 4.365 ;
      RECT 70.2 4.447 70.205 5.065 ;
      RECT 70.09 3.543 70.1 5.065 ;
      RECT 70.075 3.55 70.09 5.061 ;
      RECT 70.07 3.56 70.075 5.056 ;
      RECT 70.065 3.76 70.07 4.948 ;
      RECT 70.06 3.845 70.065 4.5 ;
      RECT 68.935 10.205 69.225 10.435 ;
      RECT 68.995 8.725 69.165 10.435 ;
      RECT 68.945 9.09 69.295 9.44 ;
      RECT 68.935 8.725 69.225 8.955 ;
      RECT 68.53 3.69 68.635 4.26 ;
      RECT 68.53 4.025 68.855 4.255 ;
      RECT 68.53 4.055 69.025 4.225 ;
      RECT 68.53 3.69 68.72 4.255 ;
      RECT 67.945 3.655 68.235 3.885 ;
      RECT 67.945 3.69 68.72 3.86 ;
      RECT 68.005 2.175 68.175 3.885 ;
      RECT 67.945 2.175 68.235 2.405 ;
      RECT 67.945 10.205 68.235 10.435 ;
      RECT 68.005 8.725 68.175 10.435 ;
      RECT 67.945 8.725 68.235 8.955 ;
      RECT 67.945 8.76 68.8 8.92 ;
      RECT 68.63 8.355 68.8 8.92 ;
      RECT 67.945 8.755 68.34 8.92 ;
      RECT 68.565 8.355 68.855 8.585 ;
      RECT 68.565 8.385 69.025 8.555 ;
      RECT 67.575 4.025 67.865 4.255 ;
      RECT 67.575 4.055 68.035 4.225 ;
      RECT 67.64 2.95 67.805 4.255 ;
      RECT 66.155 2.92 66.445 3.15 ;
      RECT 66.155 2.95 67.805 3.12 ;
      RECT 66.215 2.18 66.385 3.15 ;
      RECT 66.155 2.18 66.445 2.41 ;
      RECT 66.155 10.2 66.445 10.43 ;
      RECT 66.215 9.46 66.385 10.43 ;
      RECT 66.215 9.555 67.805 9.725 ;
      RECT 67.635 8.355 67.805 9.725 ;
      RECT 66.155 9.46 66.445 9.69 ;
      RECT 67.575 8.355 67.865 8.585 ;
      RECT 67.575 8.385 68.035 8.555 ;
      RECT 64.19 4.725 64.54 5.075 ;
      RECT 64.28 3.32 64.45 5.075 ;
      RECT 66.585 3.26 66.935 3.61 ;
      RECT 64.28 3.32 65.9 3.495 ;
      RECT 64.28 3.32 66.935 3.49 ;
      RECT 66.61 9.09 66.935 9.415 ;
      RECT 62.04 9.05 62.39 9.4 ;
      RECT 66.585 9.09 66.935 9.32 ;
      RECT 61.825 9.09 62.39 9.32 ;
      RECT 61.655 9.12 66.935 9.29 ;
      RECT 65.81 3.66 66.13 3.98 ;
      RECT 65.78 3.66 66.13 3.89 ;
      RECT 65.61 3.69 66.13 3.86 ;
      RECT 65.81 8.66 66.13 8.98 ;
      RECT 65.78 8.72 66.13 8.95 ;
      RECT 65.61 8.75 66.13 8.92 ;
      RECT 61.59 4.96 61.63 5.22 ;
      RECT 61.63 4.94 61.635 4.95 ;
      RECT 62.96 4.185 62.97 4.406 ;
      RECT 62.89 4.18 62.96 4.531 ;
      RECT 62.88 4.18 62.89 4.658 ;
      RECT 62.855 4.18 62.88 4.705 ;
      RECT 62.83 4.18 62.855 4.783 ;
      RECT 62.81 4.18 62.83 4.853 ;
      RECT 62.785 4.18 62.81 4.893 ;
      RECT 62.775 4.18 62.785 4.913 ;
      RECT 62.765 4.182 62.775 4.921 ;
      RECT 62.76 4.187 62.765 4.378 ;
      RECT 62.76 4.387 62.765 4.922 ;
      RECT 62.755 4.432 62.76 4.923 ;
      RECT 62.745 4.497 62.755 4.924 ;
      RECT 62.735 4.592 62.745 4.926 ;
      RECT 62.73 4.645 62.735 4.928 ;
      RECT 62.725 4.665 62.73 4.929 ;
      RECT 62.67 4.69 62.725 4.935 ;
      RECT 62.63 4.725 62.67 4.944 ;
      RECT 62.62 4.742 62.63 4.949 ;
      RECT 62.611 4.748 62.62 4.951 ;
      RECT 62.525 4.786 62.611 4.962 ;
      RECT 62.52 4.825 62.525 4.972 ;
      RECT 62.445 4.832 62.52 4.982 ;
      RECT 62.425 4.842 62.445 4.993 ;
      RECT 62.395 4.849 62.425 5.001 ;
      RECT 62.37 4.856 62.395 5.008 ;
      RECT 62.346 4.862 62.37 5.013 ;
      RECT 62.26 4.875 62.346 5.025 ;
      RECT 62.182 4.882 62.26 5.043 ;
      RECT 62.096 4.877 62.182 5.061 ;
      RECT 62.01 4.872 62.096 5.081 ;
      RECT 61.93 4.866 62.01 5.098 ;
      RECT 61.865 4.862 61.93 5.127 ;
      RECT 61.86 4.576 61.865 4.6 ;
      RECT 61.85 4.852 61.865 5.155 ;
      RECT 61.855 4.57 61.86 4.64 ;
      RECT 61.85 4.564 61.855 4.71 ;
      RECT 61.845 4.558 61.85 4.788 ;
      RECT 61.845 4.835 61.85 5.22 ;
      RECT 61.837 4.555 61.845 5.22 ;
      RECT 61.751 4.553 61.837 5.22 ;
      RECT 61.665 4.551 61.751 5.22 ;
      RECT 61.655 4.552 61.665 5.22 ;
      RECT 61.65 4.557 61.655 5.22 ;
      RECT 61.64 4.57 61.65 5.22 ;
      RECT 61.635 4.592 61.64 5.22 ;
      RECT 61.63 4.952 61.635 5.22 ;
      RECT 62.26 4.42 62.265 4.64 ;
      RECT 62.765 3.455 62.8 3.715 ;
      RECT 62.75 3.455 62.765 3.723 ;
      RECT 62.721 3.455 62.75 3.745 ;
      RECT 62.635 3.455 62.721 3.805 ;
      RECT 62.615 3.455 62.635 3.87 ;
      RECT 62.555 3.455 62.615 4.035 ;
      RECT 62.55 3.455 62.555 4.183 ;
      RECT 62.545 3.455 62.55 4.195 ;
      RECT 62.54 3.455 62.545 4.221 ;
      RECT 62.51 3.641 62.54 4.301 ;
      RECT 62.505 3.689 62.51 4.39 ;
      RECT 62.5 3.703 62.505 4.405 ;
      RECT 62.495 3.722 62.5 4.435 ;
      RECT 62.49 3.737 62.495 4.451 ;
      RECT 62.485 3.752 62.49 4.473 ;
      RECT 62.48 3.772 62.485 4.495 ;
      RECT 62.47 3.792 62.48 4.528 ;
      RECT 62.455 3.834 62.47 4.59 ;
      RECT 62.45 3.865 62.455 4.63 ;
      RECT 62.445 3.877 62.45 4.635 ;
      RECT 62.44 3.889 62.445 4.64 ;
      RECT 62.435 3.902 62.44 4.64 ;
      RECT 62.43 3.92 62.435 4.64 ;
      RECT 62.425 3.94 62.43 4.64 ;
      RECT 62.42 3.952 62.425 4.64 ;
      RECT 62.415 3.965 62.42 4.64 ;
      RECT 62.395 4 62.415 4.64 ;
      RECT 62.345 4.102 62.395 4.64 ;
      RECT 62.34 4.187 62.345 4.64 ;
      RECT 62.335 4.195 62.34 4.64 ;
      RECT 62.33 4.212 62.335 4.64 ;
      RECT 62.325 4.227 62.33 4.64 ;
      RECT 62.29 4.292 62.325 4.64 ;
      RECT 62.275 4.357 62.29 4.64 ;
      RECT 62.27 4.387 62.275 4.64 ;
      RECT 62.265 4.412 62.27 4.64 ;
      RECT 62.25 4.422 62.26 4.64 ;
      RECT 62.235 4.435 62.25 4.633 ;
      RECT 61.98 4.025 62.05 4.235 ;
      RECT 61.77 4.002 61.775 4.195 ;
      RECT 59.225 3.93 59.485 4.19 ;
      RECT 62.06 4.212 62.065 4.215 ;
      RECT 62.05 4.03 62.06 4.23 ;
      RECT 61.951 4.023 61.98 4.235 ;
      RECT 61.865 4.015 61.951 4.235 ;
      RECT 61.85 4.009 61.865 4.233 ;
      RECT 61.83 4.008 61.85 4.22 ;
      RECT 61.825 4.007 61.83 4.203 ;
      RECT 61.775 4.004 61.825 4.198 ;
      RECT 61.745 4.001 61.77 4.193 ;
      RECT 61.725 3.999 61.745 4.188 ;
      RECT 61.71 3.997 61.725 4.185 ;
      RECT 61.68 3.995 61.71 4.183 ;
      RECT 61.615 3.991 61.68 4.175 ;
      RECT 61.585 3.986 61.615 4.17 ;
      RECT 61.565 3.984 61.585 4.168 ;
      RECT 61.535 3.981 61.565 4.163 ;
      RECT 61.475 3.977 61.535 4.155 ;
      RECT 61.47 3.974 61.475 4.15 ;
      RECT 61.4 3.972 61.47 4.145 ;
      RECT 61.371 3.968 61.4 4.138 ;
      RECT 61.285 3.963 61.371 4.13 ;
      RECT 61.251 3.958 61.285 4.122 ;
      RECT 61.165 3.95 61.251 4.114 ;
      RECT 61.126 3.943 61.165 4.106 ;
      RECT 61.04 3.938 61.126 4.098 ;
      RECT 60.975 3.932 61.04 4.088 ;
      RECT 60.955 3.927 60.975 4.083 ;
      RECT 60.946 3.924 60.955 4.082 ;
      RECT 60.86 3.92 60.946 4.076 ;
      RECT 60.82 3.916 60.86 4.068 ;
      RECT 60.8 3.912 60.82 4.066 ;
      RECT 60.74 3.912 60.8 4.063 ;
      RECT 60.72 3.915 60.74 4.061 ;
      RECT 60.699 3.915 60.72 4.061 ;
      RECT 60.613 3.917 60.699 4.065 ;
      RECT 60.527 3.919 60.613 4.071 ;
      RECT 60.441 3.921 60.527 4.078 ;
      RECT 60.355 3.924 60.441 4.084 ;
      RECT 60.321 3.925 60.355 4.089 ;
      RECT 60.235 3.928 60.321 4.094 ;
      RECT 60.206 3.935 60.235 4.099 ;
      RECT 60.12 3.935 60.206 4.104 ;
      RECT 60.087 3.935 60.12 4.109 ;
      RECT 60.001 3.937 60.087 4.114 ;
      RECT 59.915 3.939 60.001 4.121 ;
      RECT 59.851 3.941 59.915 4.127 ;
      RECT 59.765 3.943 59.851 4.133 ;
      RECT 59.762 3.945 59.765 4.136 ;
      RECT 59.676 3.946 59.762 4.14 ;
      RECT 59.59 3.949 59.676 4.147 ;
      RECT 59.571 3.951 59.59 4.151 ;
      RECT 59.485 3.953 59.571 4.156 ;
      RECT 59.215 3.965 59.225 4.16 ;
      RECT 61.395 10.2 61.685 10.43 ;
      RECT 61.455 9.46 61.625 10.43 ;
      RECT 61.345 9.49 61.72 9.86 ;
      RECT 61.395 9.46 61.685 9.86 ;
      RECT 61.45 3.545 61.635 3.755 ;
      RECT 61.445 3.546 61.64 3.753 ;
      RECT 61.44 3.551 61.65 3.748 ;
      RECT 61.435 3.527 61.44 3.745 ;
      RECT 61.405 3.524 61.435 3.738 ;
      RECT 61.4 3.52 61.405 3.729 ;
      RECT 61.365 3.551 61.65 3.724 ;
      RECT 61.14 3.46 61.4 3.72 ;
      RECT 61.44 3.529 61.445 3.748 ;
      RECT 61.445 3.53 61.45 3.753 ;
      RECT 61.14 3.542 61.52 3.72 ;
      RECT 61.14 3.54 61.505 3.72 ;
      RECT 61.14 3.535 61.495 3.72 ;
      RECT 61.095 4.45 61.145 4.735 ;
      RECT 61.04 4.42 61.045 4.735 ;
      RECT 61.01 4.4 61.015 4.735 ;
      RECT 61.16 4.45 61.22 4.71 ;
      RECT 61.155 4.45 61.16 4.718 ;
      RECT 61.145 4.45 61.155 4.73 ;
      RECT 61.06 4.44 61.095 4.735 ;
      RECT 61.055 4.427 61.06 4.735 ;
      RECT 61.045 4.422 61.055 4.735 ;
      RECT 61.025 4.412 61.04 4.735 ;
      RECT 61.015 4.405 61.025 4.735 ;
      RECT 61.005 4.397 61.01 4.735 ;
      RECT 60.975 4.387 61.005 4.735 ;
      RECT 60.96 4.375 60.975 4.735 ;
      RECT 60.945 4.365 60.96 4.73 ;
      RECT 60.925 4.355 60.945 4.705 ;
      RECT 60.915 4.347 60.925 4.682 ;
      RECT 60.885 4.33 60.915 4.672 ;
      RECT 60.88 4.307 60.885 4.663 ;
      RECT 60.875 4.294 60.88 4.661 ;
      RECT 60.86 4.27 60.875 4.655 ;
      RECT 60.855 4.246 60.86 4.649 ;
      RECT 60.845 4.235 60.855 4.644 ;
      RECT 60.84 4.225 60.845 4.64 ;
      RECT 60.835 4.217 60.84 4.637 ;
      RECT 60.825 4.212 60.835 4.633 ;
      RECT 60.82 4.207 60.825 4.629 ;
      RECT 60.735 4.205 60.82 4.604 ;
      RECT 60.705 4.205 60.735 4.57 ;
      RECT 60.69 4.205 60.705 4.553 ;
      RECT 60.635 4.205 60.69 4.498 ;
      RECT 60.63 4.21 60.635 4.447 ;
      RECT 60.62 4.215 60.63 4.437 ;
      RECT 60.615 4.225 60.62 4.423 ;
      RECT 60.565 4.965 60.825 5.225 ;
      RECT 60.485 4.98 60.825 5.201 ;
      RECT 60.465 4.98 60.825 5.196 ;
      RECT 60.441 4.98 60.825 5.194 ;
      RECT 60.355 4.98 60.825 5.189 ;
      RECT 60.205 4.92 60.465 5.185 ;
      RECT 60.16 4.98 60.825 5.18 ;
      RECT 60.155 4.987 60.825 5.175 ;
      RECT 60.17 4.975 60.485 5.185 ;
      RECT 60.06 3.41 60.32 3.67 ;
      RECT 60.06 3.467 60.325 3.663 ;
      RECT 60.06 3.497 60.33 3.595 ;
      RECT 60.12 3.928 60.235 3.93 ;
      RECT 60.206 3.925 60.235 3.93 ;
      RECT 59.23 4.929 59.255 5.169 ;
      RECT 59.215 4.932 59.305 5.163 ;
      RECT 59.21 4.937 59.391 5.158 ;
      RECT 59.205 4.945 59.455 5.156 ;
      RECT 59.205 4.945 59.465 5.155 ;
      RECT 59.2 4.952 59.475 5.148 ;
      RECT 59.2 4.952 59.561 5.137 ;
      RECT 59.195 4.987 59.561 5.133 ;
      RECT 59.195 4.987 59.57 5.122 ;
      RECT 59.475 4.86 59.735 5.12 ;
      RECT 59.185 5.037 59.735 5.118 ;
      RECT 59.455 4.905 59.475 5.153 ;
      RECT 59.391 4.908 59.455 5.157 ;
      RECT 59.305 4.913 59.391 5.162 ;
      RECT 59.235 4.924 59.735 5.12 ;
      RECT 59.255 4.918 59.305 5.167 ;
      RECT 59.38 3.395 59.39 3.657 ;
      RECT 59.37 3.452 59.38 3.66 ;
      RECT 59.345 3.457 59.37 3.666 ;
      RECT 59.32 3.461 59.345 3.678 ;
      RECT 59.31 3.464 59.32 3.688 ;
      RECT 59.305 3.465 59.31 3.693 ;
      RECT 59.3 3.466 59.305 3.698 ;
      RECT 59.295 3.467 59.3 3.7 ;
      RECT 59.27 3.47 59.295 3.703 ;
      RECT 59.24 3.476 59.27 3.706 ;
      RECT 59.175 3.487 59.24 3.709 ;
      RECT 59.13 3.495 59.175 3.713 ;
      RECT 59.115 3.495 59.13 3.721 ;
      RECT 59.11 3.496 59.115 3.728 ;
      RECT 59.105 3.498 59.11 3.731 ;
      RECT 59.1 3.502 59.105 3.734 ;
      RECT 59.09 3.51 59.1 3.738 ;
      RECT 59.085 3.523 59.09 3.743 ;
      RECT 59.08 3.531 59.085 3.745 ;
      RECT 59.075 3.537 59.08 3.745 ;
      RECT 59.07 3.541 59.075 3.748 ;
      RECT 59.065 3.543 59.07 3.751 ;
      RECT 59.06 3.546 59.065 3.754 ;
      RECT 59.05 3.551 59.06 3.758 ;
      RECT 59.045 3.557 59.05 3.763 ;
      RECT 59.035 3.563 59.045 3.767 ;
      RECT 59.02 3.57 59.035 3.773 ;
      RECT 58.991 3.584 59.02 3.783 ;
      RECT 58.905 3.619 58.991 3.815 ;
      RECT 58.885 3.652 58.905 3.844 ;
      RECT 58.865 3.665 58.885 3.855 ;
      RECT 58.845 3.677 58.865 3.866 ;
      RECT 58.795 3.699 58.845 3.886 ;
      RECT 58.78 3.717 58.795 3.903 ;
      RECT 58.775 3.723 58.78 3.906 ;
      RECT 58.77 3.727 58.775 3.909 ;
      RECT 58.765 3.731 58.77 3.913 ;
      RECT 58.76 3.733 58.765 3.916 ;
      RECT 58.75 3.74 58.76 3.919 ;
      RECT 58.745 3.745 58.75 3.923 ;
      RECT 58.74 3.747 58.745 3.926 ;
      RECT 58.735 3.751 58.74 3.929 ;
      RECT 58.73 3.753 58.735 3.933 ;
      RECT 58.715 3.758 58.73 3.938 ;
      RECT 58.71 3.763 58.715 3.941 ;
      RECT 58.705 3.771 58.71 3.944 ;
      RECT 58.7 3.773 58.705 3.947 ;
      RECT 58.695 3.775 58.7 3.95 ;
      RECT 58.685 3.777 58.695 3.956 ;
      RECT 58.65 3.791 58.685 3.968 ;
      RECT 58.64 3.806 58.65 3.978 ;
      RECT 58.565 3.835 58.64 4.002 ;
      RECT 58.56 3.86 58.565 4.025 ;
      RECT 58.545 3.864 58.56 4.031 ;
      RECT 58.535 3.872 58.545 4.036 ;
      RECT 58.505 3.885 58.535 4.04 ;
      RECT 58.495 3.9 58.505 4.045 ;
      RECT 58.485 3.905 58.495 4.048 ;
      RECT 58.48 3.907 58.485 4.05 ;
      RECT 58.465 3.91 58.48 4.053 ;
      RECT 58.46 3.912 58.465 4.056 ;
      RECT 58.44 3.917 58.46 4.06 ;
      RECT 58.41 3.922 58.44 4.068 ;
      RECT 58.385 3.929 58.41 4.076 ;
      RECT 58.38 3.934 58.385 4.081 ;
      RECT 58.35 3.937 58.38 4.085 ;
      RECT 58.31 3.94 58.35 4.095 ;
      RECT 58.275 3.937 58.31 4.107 ;
      RECT 58.265 3.933 58.275 4.114 ;
      RECT 58.24 3.929 58.265 4.12 ;
      RECT 58.235 3.925 58.24 4.125 ;
      RECT 58.195 3.922 58.235 4.125 ;
      RECT 58.18 3.907 58.195 4.126 ;
      RECT 58.157 3.895 58.18 4.126 ;
      RECT 58.071 3.895 58.157 4.127 ;
      RECT 57.985 3.895 58.071 4.129 ;
      RECT 57.965 3.895 57.985 4.126 ;
      RECT 57.96 3.9 57.965 4.121 ;
      RECT 57.955 3.905 57.96 4.119 ;
      RECT 57.945 3.915 57.955 4.117 ;
      RECT 57.94 3.921 57.945 4.11 ;
      RECT 57.935 3.923 57.94 4.095 ;
      RECT 57.93 3.927 57.935 4.085 ;
      RECT 59.39 3.395 59.64 3.655 ;
      RECT 57.115 4.93 57.375 5.19 ;
      RECT 59.41 4.42 59.415 4.63 ;
      RECT 59.415 4.425 59.425 4.625 ;
      RECT 59.365 4.42 59.41 4.645 ;
      RECT 59.355 4.42 59.365 4.665 ;
      RECT 59.336 4.42 59.355 4.67 ;
      RECT 59.25 4.42 59.336 4.667 ;
      RECT 59.22 4.422 59.25 4.665 ;
      RECT 59.165 4.432 59.22 4.663 ;
      RECT 59.1 4.446 59.165 4.661 ;
      RECT 59.095 4.454 59.1 4.66 ;
      RECT 59.08 4.457 59.095 4.658 ;
      RECT 59.015 4.467 59.08 4.654 ;
      RECT 58.967 4.481 59.015 4.655 ;
      RECT 58.881 4.498 58.967 4.669 ;
      RECT 58.795 4.519 58.881 4.686 ;
      RECT 58.775 4.532 58.795 4.696 ;
      RECT 58.73 4.54 58.775 4.703 ;
      RECT 58.695 4.548 58.73 4.711 ;
      RECT 58.661 4.556 58.695 4.719 ;
      RECT 58.575 4.57 58.661 4.731 ;
      RECT 58.54 4.587 58.575 4.743 ;
      RECT 58.531 4.596 58.54 4.747 ;
      RECT 58.445 4.614 58.531 4.764 ;
      RECT 58.386 4.641 58.445 4.791 ;
      RECT 58.3 4.668 58.386 4.819 ;
      RECT 58.28 4.69 58.3 4.839 ;
      RECT 58.22 4.705 58.28 4.855 ;
      RECT 58.21 4.717 58.22 4.868 ;
      RECT 58.205 4.722 58.21 4.871 ;
      RECT 58.195 4.725 58.205 4.874 ;
      RECT 58.19 4.727 58.195 4.877 ;
      RECT 58.16 4.735 58.19 4.884 ;
      RECT 58.145 4.742 58.16 4.892 ;
      RECT 58.135 4.747 58.145 4.896 ;
      RECT 58.13 4.75 58.135 4.899 ;
      RECT 58.12 4.752 58.13 4.902 ;
      RECT 58.085 4.762 58.12 4.911 ;
      RECT 58.01 4.785 58.085 4.933 ;
      RECT 57.99 4.803 58.01 4.951 ;
      RECT 57.96 4.81 57.99 4.961 ;
      RECT 57.94 4.818 57.96 4.971 ;
      RECT 57.93 4.824 57.94 4.978 ;
      RECT 57.911 4.829 57.93 4.984 ;
      RECT 57.825 4.849 57.911 5.004 ;
      RECT 57.81 4.869 57.825 5.023 ;
      RECT 57.765 4.881 57.81 5.034 ;
      RECT 57.7 4.902 57.765 5.057 ;
      RECT 57.66 4.922 57.7 5.078 ;
      RECT 57.65 4.932 57.66 5.088 ;
      RECT 57.6 4.944 57.65 5.099 ;
      RECT 57.58 4.96 57.6 5.111 ;
      RECT 57.55 4.97 57.58 5.117 ;
      RECT 57.54 4.975 57.55 5.119 ;
      RECT 57.471 4.976 57.54 5.125 ;
      RECT 57.385 4.978 57.471 5.135 ;
      RECT 57.375 4.979 57.385 5.14 ;
      RECT 58.645 5.005 58.835 5.215 ;
      RECT 58.635 5.01 58.845 5.208 ;
      RECT 58.62 5.01 58.845 5.173 ;
      RECT 58.54 4.895 58.8 5.155 ;
      RECT 57.455 4.425 57.64 4.72 ;
      RECT 57.445 4.425 57.64 4.718 ;
      RECT 57.43 4.425 57.645 4.713 ;
      RECT 57.43 4.425 57.65 4.71 ;
      RECT 57.425 4.425 57.65 4.708 ;
      RECT 57.42 4.68 57.65 4.698 ;
      RECT 57.425 4.425 57.685 4.685 ;
      RECT 57.385 3.46 57.645 3.72 ;
      RECT 57.195 3.385 57.281 3.718 ;
      RECT 57.17 3.389 57.325 3.714 ;
      RECT 57.281 3.381 57.325 3.714 ;
      RECT 57.281 3.382 57.33 3.713 ;
      RECT 57.195 3.387 57.345 3.712 ;
      RECT 57.17 3.395 57.385 3.711 ;
      RECT 57.165 3.39 57.345 3.706 ;
      RECT 57.155 3.405 57.385 3.613 ;
      RECT 57.155 3.457 57.585 3.613 ;
      RECT 57.155 3.45 57.565 3.613 ;
      RECT 57.155 3.437 57.535 3.613 ;
      RECT 57.155 3.425 57.475 3.613 ;
      RECT 57.155 3.41 57.45 3.613 ;
      RECT 56.355 4.04 56.49 4.335 ;
      RECT 56.615 4.063 56.62 4.25 ;
      RECT 57.335 3.96 57.48 4.195 ;
      RECT 57.495 3.96 57.5 4.185 ;
      RECT 57.53 3.971 57.535 4.165 ;
      RECT 57.525 3.963 57.53 4.17 ;
      RECT 57.505 3.96 57.525 4.175 ;
      RECT 57.5 3.96 57.505 4.183 ;
      RECT 57.49 3.96 57.495 4.188 ;
      RECT 57.48 3.96 57.49 4.193 ;
      RECT 57.31 3.962 57.335 4.195 ;
      RECT 57.26 3.969 57.31 4.195 ;
      RECT 57.255 3.974 57.26 4.195 ;
      RECT 57.216 3.979 57.255 4.196 ;
      RECT 57.13 3.991 57.216 4.197 ;
      RECT 57.121 4.001 57.13 4.197 ;
      RECT 57.035 4.01 57.121 4.199 ;
      RECT 57.011 4.02 57.035 4.201 ;
      RECT 56.925 4.031 57.011 4.202 ;
      RECT 56.895 4.042 56.925 4.204 ;
      RECT 56.865 4.047 56.895 4.206 ;
      RECT 56.84 4.053 56.865 4.209 ;
      RECT 56.825 4.058 56.84 4.21 ;
      RECT 56.78 4.064 56.825 4.21 ;
      RECT 56.775 4.069 56.78 4.211 ;
      RECT 56.755 4.069 56.775 4.213 ;
      RECT 56.735 4.067 56.755 4.218 ;
      RECT 56.7 4.066 56.735 4.225 ;
      RECT 56.67 4.065 56.7 4.235 ;
      RECT 56.62 4.064 56.67 4.245 ;
      RECT 56.53 4.061 56.615 4.335 ;
      RECT 56.505 4.055 56.53 4.335 ;
      RECT 56.49 4.045 56.505 4.335 ;
      RECT 56.305 4.04 56.355 4.255 ;
      RECT 56.295 4.045 56.305 4.245 ;
      RECT 56.535 4.52 56.795 4.78 ;
      RECT 56.535 4.52 56.825 4.673 ;
      RECT 56.535 4.52 56.86 4.658 ;
      RECT 56.79 4.44 56.98 4.65 ;
      RECT 56.78 4.445 56.99 4.643 ;
      RECT 56.745 4.515 56.99 4.643 ;
      RECT 56.775 4.457 56.795 4.78 ;
      RECT 56.76 4.505 56.99 4.643 ;
      RECT 56.765 4.477 56.795 4.78 ;
      RECT 55.845 3.545 55.915 4.65 ;
      RECT 56.58 3.65 56.84 3.91 ;
      RECT 56.16 3.696 56.175 3.905 ;
      RECT 56.496 3.709 56.58 3.86 ;
      RECT 56.41 3.706 56.496 3.86 ;
      RECT 56.371 3.704 56.41 3.86 ;
      RECT 56.285 3.702 56.371 3.86 ;
      RECT 56.225 3.7 56.285 3.871 ;
      RECT 56.19 3.698 56.225 3.889 ;
      RECT 56.175 3.696 56.19 3.9 ;
      RECT 56.145 3.696 56.16 3.913 ;
      RECT 56.135 3.696 56.145 3.918 ;
      RECT 56.11 3.695 56.135 3.923 ;
      RECT 56.095 3.69 56.11 3.929 ;
      RECT 56.09 3.683 56.095 3.934 ;
      RECT 56.065 3.674 56.09 3.94 ;
      RECT 56.02 3.653 56.065 3.953 ;
      RECT 56.01 3.637 56.02 3.963 ;
      RECT 55.995 3.63 56.01 3.973 ;
      RECT 55.985 3.623 55.995 3.99 ;
      RECT 55.98 3.62 55.985 4.02 ;
      RECT 55.975 3.618 55.98 4.05 ;
      RECT 55.97 3.616 55.975 4.087 ;
      RECT 55.955 3.612 55.97 4.154 ;
      RECT 55.955 4.445 55.965 4.645 ;
      RECT 55.95 3.608 55.955 4.28 ;
      RECT 55.95 4.432 55.955 4.65 ;
      RECT 55.945 3.606 55.95 4.365 ;
      RECT 55.945 4.422 55.95 4.65 ;
      RECT 55.93 3.577 55.945 4.65 ;
      RECT 55.915 3.55 55.93 4.65 ;
      RECT 55.84 3.545 55.845 3.9 ;
      RECT 55.84 3.955 55.845 4.65 ;
      RECT 55.825 3.545 55.84 3.878 ;
      RECT 55.835 3.977 55.84 4.65 ;
      RECT 55.825 4.017 55.835 4.65 ;
      RECT 55.79 3.545 55.825 3.82 ;
      RECT 55.82 4.052 55.825 4.65 ;
      RECT 55.805 4.107 55.82 4.65 ;
      RECT 55.8 4.172 55.805 4.65 ;
      RECT 55.785 4.22 55.8 4.65 ;
      RECT 55.76 3.545 55.79 3.775 ;
      RECT 55.78 4.275 55.785 4.65 ;
      RECT 55.765 4.335 55.78 4.65 ;
      RECT 55.76 4.383 55.765 4.648 ;
      RECT 55.755 3.545 55.76 3.768 ;
      RECT 55.755 4.415 55.76 4.643 ;
      RECT 55.73 3.545 55.755 3.76 ;
      RECT 55.72 3.55 55.73 3.75 ;
      RECT 55.935 4.825 55.955 5.065 ;
      RECT 55.165 4.755 55.17 4.965 ;
      RECT 56.445 4.828 56.455 5.023 ;
      RECT 56.44 4.818 56.445 5.026 ;
      RECT 56.36 4.815 56.44 5.049 ;
      RECT 56.356 4.815 56.36 5.071 ;
      RECT 56.27 4.815 56.356 5.081 ;
      RECT 56.255 4.815 56.27 5.089 ;
      RECT 56.226 4.816 56.255 5.087 ;
      RECT 56.14 4.821 56.226 5.083 ;
      RECT 56.127 4.825 56.14 5.079 ;
      RECT 56.041 4.825 56.127 5.075 ;
      RECT 55.955 4.825 56.041 5.069 ;
      RECT 55.871 4.825 55.935 5.063 ;
      RECT 55.785 4.825 55.871 5.058 ;
      RECT 55.765 4.825 55.785 5.054 ;
      RECT 55.705 4.82 55.765 5.051 ;
      RECT 55.677 4.814 55.705 5.048 ;
      RECT 55.591 4.809 55.677 5.044 ;
      RECT 55.505 4.803 55.591 5.038 ;
      RECT 55.43 4.785 55.505 5.033 ;
      RECT 55.395 4.762 55.43 5.029 ;
      RECT 55.385 4.752 55.395 5.028 ;
      RECT 55.33 4.75 55.385 5.027 ;
      RECT 55.255 4.75 55.33 5.023 ;
      RECT 55.245 4.75 55.255 5.018 ;
      RECT 55.23 4.75 55.245 5.01 ;
      RECT 55.18 4.752 55.23 4.988 ;
      RECT 55.17 4.755 55.18 4.968 ;
      RECT 55.16 4.76 55.165 4.963 ;
      RECT 55.155 4.765 55.16 4.958 ;
      RECT 55.28 3.93 55.54 4.19 ;
      RECT 55.28 3.945 55.56 4.155 ;
      RECT 55.28 3.95 55.57 4.15 ;
      RECT 53.265 3.41 53.525 3.67 ;
      RECT 53.255 3.44 53.525 3.65 ;
      RECT 55.175 3.355 55.435 3.615 ;
      RECT 55.17 3.43 55.175 3.616 ;
      RECT 55.145 3.435 55.17 3.618 ;
      RECT 55.13 3.442 55.145 3.621 ;
      RECT 55.07 3.46 55.13 3.626 ;
      RECT 55.04 3.48 55.07 3.633 ;
      RECT 55.015 3.488 55.04 3.638 ;
      RECT 54.99 3.496 55.015 3.64 ;
      RECT 54.972 3.5 54.99 3.639 ;
      RECT 54.886 3.498 54.972 3.639 ;
      RECT 54.8 3.496 54.886 3.639 ;
      RECT 54.714 3.494 54.8 3.638 ;
      RECT 54.628 3.492 54.714 3.638 ;
      RECT 54.542 3.49 54.628 3.638 ;
      RECT 54.456 3.488 54.542 3.638 ;
      RECT 54.37 3.486 54.456 3.637 ;
      RECT 54.352 3.485 54.37 3.637 ;
      RECT 54.266 3.484 54.352 3.637 ;
      RECT 54.18 3.482 54.266 3.637 ;
      RECT 54.094 3.481 54.18 3.636 ;
      RECT 54.008 3.48 54.094 3.636 ;
      RECT 53.922 3.478 54.008 3.636 ;
      RECT 53.836 3.477 53.922 3.636 ;
      RECT 53.75 3.475 53.836 3.635 ;
      RECT 53.726 3.473 53.75 3.635 ;
      RECT 53.64 3.466 53.726 3.635 ;
      RECT 53.611 3.458 53.64 3.635 ;
      RECT 53.525 3.45 53.611 3.635 ;
      RECT 53.245 3.447 53.255 3.645 ;
      RECT 54.75 4.41 54.755 4.76 ;
      RECT 54.52 4.5 54.66 4.76 ;
      RECT 54.995 4.185 55.04 4.395 ;
      RECT 55.05 4.196 55.06 4.39 ;
      RECT 55.04 4.188 55.05 4.395 ;
      RECT 54.975 4.185 54.995 4.4 ;
      RECT 54.945 4.185 54.975 4.423 ;
      RECT 54.935 4.185 54.945 4.448 ;
      RECT 54.93 4.185 54.935 4.458 ;
      RECT 54.875 4.185 54.93 4.498 ;
      RECT 54.87 4.185 54.875 4.538 ;
      RECT 54.865 4.187 54.87 4.543 ;
      RECT 54.85 4.197 54.865 4.554 ;
      RECT 54.805 4.255 54.85 4.59 ;
      RECT 54.795 4.31 54.805 4.624 ;
      RECT 54.78 4.337 54.795 4.64 ;
      RECT 54.77 4.364 54.78 4.76 ;
      RECT 54.755 4.387 54.77 4.76 ;
      RECT 54.745 4.427 54.75 4.76 ;
      RECT 54.74 4.437 54.745 4.76 ;
      RECT 54.735 4.452 54.74 4.76 ;
      RECT 54.725 4.457 54.735 4.76 ;
      RECT 54.66 4.48 54.725 4.76 ;
      RECT 54.16 3.975 54.35 4.185 ;
      RECT 52.735 3.9 52.995 4.16 ;
      RECT 53.085 3.895 53.18 4.105 ;
      RECT 53.06 3.91 53.07 4.105 ;
      RECT 54.35 3.982 54.36 4.18 ;
      RECT 54.15 3.982 54.16 4.18 ;
      RECT 54.135 3.997 54.15 4.17 ;
      RECT 54.13 4.005 54.135 4.163 ;
      RECT 54.12 4.008 54.13 4.16 ;
      RECT 54.085 4.007 54.12 4.158 ;
      RECT 54.056 4.003 54.085 4.155 ;
      RECT 53.97 3.998 54.056 4.152 ;
      RECT 53.91 3.992 53.97 4.148 ;
      RECT 53.881 3.988 53.91 4.145 ;
      RECT 53.795 3.98 53.881 4.142 ;
      RECT 53.786 3.974 53.795 4.14 ;
      RECT 53.7 3.969 53.786 4.138 ;
      RECT 53.677 3.964 53.7 4.135 ;
      RECT 53.591 3.958 53.677 4.132 ;
      RECT 53.505 3.949 53.591 4.127 ;
      RECT 53.495 3.944 53.505 4.125 ;
      RECT 53.476 3.943 53.495 4.124 ;
      RECT 53.39 3.938 53.476 4.12 ;
      RECT 53.37 3.933 53.39 4.116 ;
      RECT 53.31 3.928 53.37 4.113 ;
      RECT 53.285 3.918 53.31 4.111 ;
      RECT 53.28 3.911 53.285 4.11 ;
      RECT 53.27 3.902 53.28 4.109 ;
      RECT 53.266 3.895 53.27 4.109 ;
      RECT 53.18 3.895 53.266 4.107 ;
      RECT 53.07 3.902 53.085 4.105 ;
      RECT 53.055 3.912 53.06 4.105 ;
      RECT 53.035 3.915 53.055 4.102 ;
      RECT 53.005 3.915 53.035 4.098 ;
      RECT 52.995 3.915 53.005 4.098 ;
      RECT 53.91 4.41 54.17 4.67 ;
      RECT 53.84 4.42 54.17 4.63 ;
      RECT 53.83 4.427 54.17 4.625 ;
      RECT 53.25 4.415 53.51 4.675 ;
      RECT 53.25 4.455 53.615 4.665 ;
      RECT 53.25 4.457 53.62 4.664 ;
      RECT 53.25 4.465 53.625 4.661 ;
      RECT 52.175 3.54 52.275 5.065 ;
      RECT 52.365 4.68 52.415 4.94 ;
      RECT 52.36 3.553 52.365 3.74 ;
      RECT 52.355 4.661 52.365 4.94 ;
      RECT 52.355 3.55 52.36 3.748 ;
      RECT 52.34 3.544 52.355 3.755 ;
      RECT 52.35 4.649 52.355 5.023 ;
      RECT 52.34 4.637 52.35 5.06 ;
      RECT 52.33 3.54 52.34 3.762 ;
      RECT 52.33 4.622 52.34 5.065 ;
      RECT 52.325 3.54 52.33 3.77 ;
      RECT 52.305 4.592 52.33 5.065 ;
      RECT 52.285 3.54 52.325 3.818 ;
      RECT 52.295 4.552 52.305 5.065 ;
      RECT 52.285 4.507 52.295 5.065 ;
      RECT 52.28 3.54 52.285 3.888 ;
      RECT 52.28 4.465 52.285 5.065 ;
      RECT 52.275 3.54 52.28 4.365 ;
      RECT 52.275 4.447 52.28 5.065 ;
      RECT 52.165 3.543 52.175 5.065 ;
      RECT 52.15 3.55 52.165 5.061 ;
      RECT 52.145 3.56 52.15 5.056 ;
      RECT 52.14 3.76 52.145 4.948 ;
      RECT 52.135 3.845 52.14 4.5 ;
      RECT 51.01 10.205 51.3 10.435 ;
      RECT 51.07 8.725 51.24 10.435 ;
      RECT 51.06 9.095 51.415 9.45 ;
      RECT 51.01 8.725 51.3 8.955 ;
      RECT 50.605 3.69 50.71 4.26 ;
      RECT 50.605 4.025 50.93 4.255 ;
      RECT 50.605 4.055 51.1 4.225 ;
      RECT 50.605 3.69 50.795 4.255 ;
      RECT 50.02 3.655 50.31 3.885 ;
      RECT 50.02 3.69 50.795 3.86 ;
      RECT 50.08 2.175 50.25 3.885 ;
      RECT 50.02 2.175 50.31 2.405 ;
      RECT 50.02 10.205 50.31 10.435 ;
      RECT 50.08 8.725 50.25 10.435 ;
      RECT 50.02 8.725 50.31 8.955 ;
      RECT 50.02 8.76 50.875 8.92 ;
      RECT 50.705 8.355 50.875 8.92 ;
      RECT 50.02 8.755 50.415 8.92 ;
      RECT 50.64 8.355 50.93 8.585 ;
      RECT 50.64 8.385 51.1 8.555 ;
      RECT 49.65 4.025 49.94 4.255 ;
      RECT 49.65 4.055 50.11 4.225 ;
      RECT 49.715 2.95 49.88 4.255 ;
      RECT 48.23 2.92 48.52 3.15 ;
      RECT 48.23 2.95 49.88 3.12 ;
      RECT 48.29 2.18 48.46 3.15 ;
      RECT 48.23 2.18 48.52 2.41 ;
      RECT 48.23 10.2 48.52 10.43 ;
      RECT 48.29 9.46 48.46 10.43 ;
      RECT 48.29 9.555 49.88 9.725 ;
      RECT 49.71 8.355 49.88 9.725 ;
      RECT 48.23 9.46 48.52 9.69 ;
      RECT 49.65 8.355 49.94 8.585 ;
      RECT 49.65 8.385 50.11 8.555 ;
      RECT 46.265 4.725 46.615 5.075 ;
      RECT 46.355 3.32 46.525 5.075 ;
      RECT 48.66 3.26 49.01 3.61 ;
      RECT 46.355 3.32 47.975 3.495 ;
      RECT 46.355 3.32 49.01 3.49 ;
      RECT 48.685 9.09 49.01 9.415 ;
      RECT 44.11 9.045 44.46 9.395 ;
      RECT 48.66 9.09 49.01 9.32 ;
      RECT 43.9 9.09 44.46 9.32 ;
      RECT 43.73 9.12 49.01 9.29 ;
      RECT 47.885 3.66 48.205 3.98 ;
      RECT 47.855 3.66 48.205 3.89 ;
      RECT 47.685 3.69 48.205 3.86 ;
      RECT 47.885 8.66 48.205 8.98 ;
      RECT 47.855 8.72 48.205 8.95 ;
      RECT 47.685 8.75 48.205 8.92 ;
      RECT 43.665 4.96 43.705 5.22 ;
      RECT 43.705 4.94 43.71 4.95 ;
      RECT 45.035 4.185 45.045 4.406 ;
      RECT 44.965 4.18 45.035 4.531 ;
      RECT 44.955 4.18 44.965 4.658 ;
      RECT 44.93 4.18 44.955 4.705 ;
      RECT 44.905 4.18 44.93 4.783 ;
      RECT 44.885 4.18 44.905 4.853 ;
      RECT 44.86 4.18 44.885 4.893 ;
      RECT 44.85 4.18 44.86 4.913 ;
      RECT 44.84 4.182 44.85 4.921 ;
      RECT 44.835 4.187 44.84 4.378 ;
      RECT 44.835 4.387 44.84 4.922 ;
      RECT 44.83 4.432 44.835 4.923 ;
      RECT 44.82 4.497 44.83 4.924 ;
      RECT 44.81 4.592 44.82 4.926 ;
      RECT 44.805 4.645 44.81 4.928 ;
      RECT 44.8 4.665 44.805 4.929 ;
      RECT 44.745 4.69 44.8 4.935 ;
      RECT 44.705 4.725 44.745 4.944 ;
      RECT 44.695 4.742 44.705 4.949 ;
      RECT 44.686 4.748 44.695 4.951 ;
      RECT 44.6 4.786 44.686 4.962 ;
      RECT 44.595 4.825 44.6 4.972 ;
      RECT 44.52 4.832 44.595 4.982 ;
      RECT 44.5 4.842 44.52 4.993 ;
      RECT 44.47 4.849 44.5 5.001 ;
      RECT 44.445 4.856 44.47 5.008 ;
      RECT 44.421 4.862 44.445 5.013 ;
      RECT 44.335 4.875 44.421 5.025 ;
      RECT 44.257 4.882 44.335 5.043 ;
      RECT 44.171 4.877 44.257 5.061 ;
      RECT 44.085 4.872 44.171 5.081 ;
      RECT 44.005 4.866 44.085 5.098 ;
      RECT 43.94 4.862 44.005 5.127 ;
      RECT 43.935 4.576 43.94 4.6 ;
      RECT 43.925 4.852 43.94 5.155 ;
      RECT 43.93 4.57 43.935 4.64 ;
      RECT 43.925 4.564 43.93 4.71 ;
      RECT 43.92 4.558 43.925 4.788 ;
      RECT 43.92 4.835 43.925 5.22 ;
      RECT 43.912 4.555 43.92 5.22 ;
      RECT 43.826 4.553 43.912 5.22 ;
      RECT 43.74 4.551 43.826 5.22 ;
      RECT 43.73 4.552 43.74 5.22 ;
      RECT 43.725 4.557 43.73 5.22 ;
      RECT 43.715 4.57 43.725 5.22 ;
      RECT 43.71 4.592 43.715 5.22 ;
      RECT 43.705 4.952 43.71 5.22 ;
      RECT 44.335 4.42 44.34 4.64 ;
      RECT 44.84 3.455 44.875 3.715 ;
      RECT 44.825 3.455 44.84 3.723 ;
      RECT 44.796 3.455 44.825 3.745 ;
      RECT 44.71 3.455 44.796 3.805 ;
      RECT 44.69 3.455 44.71 3.87 ;
      RECT 44.63 3.455 44.69 4.035 ;
      RECT 44.625 3.455 44.63 4.183 ;
      RECT 44.62 3.455 44.625 4.195 ;
      RECT 44.615 3.455 44.62 4.221 ;
      RECT 44.585 3.641 44.615 4.301 ;
      RECT 44.58 3.689 44.585 4.39 ;
      RECT 44.575 3.703 44.58 4.405 ;
      RECT 44.57 3.722 44.575 4.435 ;
      RECT 44.565 3.737 44.57 4.451 ;
      RECT 44.56 3.752 44.565 4.473 ;
      RECT 44.555 3.772 44.56 4.495 ;
      RECT 44.545 3.792 44.555 4.528 ;
      RECT 44.53 3.834 44.545 4.59 ;
      RECT 44.525 3.865 44.53 4.63 ;
      RECT 44.52 3.877 44.525 4.635 ;
      RECT 44.515 3.889 44.52 4.64 ;
      RECT 44.51 3.902 44.515 4.64 ;
      RECT 44.505 3.92 44.51 4.64 ;
      RECT 44.5 3.94 44.505 4.64 ;
      RECT 44.495 3.952 44.5 4.64 ;
      RECT 44.49 3.965 44.495 4.64 ;
      RECT 44.47 4 44.49 4.64 ;
      RECT 44.42 4.102 44.47 4.64 ;
      RECT 44.415 4.187 44.42 4.64 ;
      RECT 44.41 4.195 44.415 4.64 ;
      RECT 44.405 4.212 44.41 4.64 ;
      RECT 44.4 4.227 44.405 4.64 ;
      RECT 44.365 4.292 44.4 4.64 ;
      RECT 44.35 4.357 44.365 4.64 ;
      RECT 44.345 4.387 44.35 4.64 ;
      RECT 44.34 4.412 44.345 4.64 ;
      RECT 44.325 4.422 44.335 4.64 ;
      RECT 44.31 4.435 44.325 4.633 ;
      RECT 44.055 4.025 44.125 4.235 ;
      RECT 43.845 4.002 43.85 4.195 ;
      RECT 41.3 3.93 41.56 4.19 ;
      RECT 44.135 4.212 44.14 4.215 ;
      RECT 44.125 4.03 44.135 4.23 ;
      RECT 44.026 4.023 44.055 4.235 ;
      RECT 43.94 4.015 44.026 4.235 ;
      RECT 43.925 4.009 43.94 4.233 ;
      RECT 43.905 4.008 43.925 4.22 ;
      RECT 43.9 4.007 43.905 4.203 ;
      RECT 43.85 4.004 43.9 4.198 ;
      RECT 43.82 4.001 43.845 4.193 ;
      RECT 43.8 3.999 43.82 4.188 ;
      RECT 43.785 3.997 43.8 4.185 ;
      RECT 43.755 3.995 43.785 4.183 ;
      RECT 43.69 3.991 43.755 4.175 ;
      RECT 43.66 3.986 43.69 4.17 ;
      RECT 43.64 3.984 43.66 4.168 ;
      RECT 43.61 3.981 43.64 4.163 ;
      RECT 43.55 3.977 43.61 4.155 ;
      RECT 43.545 3.974 43.55 4.15 ;
      RECT 43.475 3.972 43.545 4.145 ;
      RECT 43.446 3.968 43.475 4.138 ;
      RECT 43.36 3.963 43.446 4.13 ;
      RECT 43.326 3.958 43.36 4.122 ;
      RECT 43.24 3.95 43.326 4.114 ;
      RECT 43.201 3.943 43.24 4.106 ;
      RECT 43.115 3.938 43.201 4.098 ;
      RECT 43.05 3.932 43.115 4.088 ;
      RECT 43.03 3.927 43.05 4.083 ;
      RECT 43.021 3.924 43.03 4.082 ;
      RECT 42.935 3.92 43.021 4.076 ;
      RECT 42.895 3.916 42.935 4.068 ;
      RECT 42.875 3.912 42.895 4.066 ;
      RECT 42.815 3.912 42.875 4.063 ;
      RECT 42.795 3.915 42.815 4.061 ;
      RECT 42.774 3.915 42.795 4.061 ;
      RECT 42.688 3.917 42.774 4.065 ;
      RECT 42.602 3.919 42.688 4.071 ;
      RECT 42.516 3.921 42.602 4.078 ;
      RECT 42.43 3.924 42.516 4.084 ;
      RECT 42.396 3.925 42.43 4.089 ;
      RECT 42.31 3.928 42.396 4.094 ;
      RECT 42.281 3.935 42.31 4.099 ;
      RECT 42.195 3.935 42.281 4.104 ;
      RECT 42.162 3.935 42.195 4.109 ;
      RECT 42.076 3.937 42.162 4.114 ;
      RECT 41.99 3.939 42.076 4.121 ;
      RECT 41.926 3.941 41.99 4.127 ;
      RECT 41.84 3.943 41.926 4.133 ;
      RECT 41.837 3.945 41.84 4.136 ;
      RECT 41.751 3.946 41.837 4.14 ;
      RECT 41.665 3.949 41.751 4.147 ;
      RECT 41.646 3.951 41.665 4.151 ;
      RECT 41.56 3.953 41.646 4.156 ;
      RECT 41.29 3.965 41.3 4.16 ;
      RECT 43.47 10.2 43.76 10.43 ;
      RECT 43.53 9.46 43.7 10.43 ;
      RECT 43.42 9.49 43.795 9.86 ;
      RECT 43.47 9.46 43.76 9.86 ;
      RECT 43.525 3.545 43.71 3.755 ;
      RECT 43.52 3.546 43.715 3.753 ;
      RECT 43.515 3.551 43.725 3.748 ;
      RECT 43.51 3.527 43.515 3.745 ;
      RECT 43.48 3.524 43.51 3.738 ;
      RECT 43.475 3.52 43.48 3.729 ;
      RECT 43.44 3.551 43.725 3.724 ;
      RECT 43.215 3.46 43.475 3.72 ;
      RECT 43.515 3.529 43.52 3.748 ;
      RECT 43.52 3.53 43.525 3.753 ;
      RECT 43.215 3.542 43.595 3.72 ;
      RECT 43.215 3.54 43.58 3.72 ;
      RECT 43.215 3.535 43.57 3.72 ;
      RECT 43.17 4.45 43.22 4.735 ;
      RECT 43.115 4.42 43.12 4.735 ;
      RECT 43.085 4.4 43.09 4.735 ;
      RECT 43.235 4.45 43.295 4.71 ;
      RECT 43.23 4.45 43.235 4.718 ;
      RECT 43.22 4.45 43.23 4.73 ;
      RECT 43.135 4.44 43.17 4.735 ;
      RECT 43.13 4.427 43.135 4.735 ;
      RECT 43.12 4.422 43.13 4.735 ;
      RECT 43.1 4.412 43.115 4.735 ;
      RECT 43.09 4.405 43.1 4.735 ;
      RECT 43.08 4.397 43.085 4.735 ;
      RECT 43.05 4.387 43.08 4.735 ;
      RECT 43.035 4.375 43.05 4.735 ;
      RECT 43.02 4.365 43.035 4.73 ;
      RECT 43 4.355 43.02 4.705 ;
      RECT 42.99 4.347 43 4.682 ;
      RECT 42.96 4.33 42.99 4.672 ;
      RECT 42.955 4.307 42.96 4.663 ;
      RECT 42.95 4.294 42.955 4.661 ;
      RECT 42.935 4.27 42.95 4.655 ;
      RECT 42.93 4.246 42.935 4.649 ;
      RECT 42.92 4.235 42.93 4.644 ;
      RECT 42.915 4.225 42.92 4.64 ;
      RECT 42.91 4.217 42.915 4.637 ;
      RECT 42.9 4.212 42.91 4.633 ;
      RECT 42.895 4.207 42.9 4.629 ;
      RECT 42.81 4.205 42.895 4.604 ;
      RECT 42.78 4.205 42.81 4.57 ;
      RECT 42.765 4.205 42.78 4.553 ;
      RECT 42.71 4.205 42.765 4.498 ;
      RECT 42.705 4.21 42.71 4.447 ;
      RECT 42.695 4.215 42.705 4.437 ;
      RECT 42.69 4.225 42.695 4.423 ;
      RECT 42.64 4.965 42.9 5.225 ;
      RECT 42.56 4.98 42.9 5.201 ;
      RECT 42.54 4.98 42.9 5.196 ;
      RECT 42.516 4.98 42.9 5.194 ;
      RECT 42.43 4.98 42.9 5.189 ;
      RECT 42.28 4.92 42.54 5.185 ;
      RECT 42.235 4.98 42.9 5.18 ;
      RECT 42.23 4.987 42.9 5.175 ;
      RECT 42.245 4.975 42.56 5.185 ;
      RECT 42.135 3.41 42.395 3.67 ;
      RECT 42.135 3.467 42.4 3.663 ;
      RECT 42.135 3.497 42.405 3.595 ;
      RECT 42.195 3.928 42.31 3.93 ;
      RECT 42.281 3.925 42.31 3.93 ;
      RECT 41.305 4.929 41.33 5.169 ;
      RECT 41.29 4.932 41.38 5.163 ;
      RECT 41.285 4.937 41.466 5.158 ;
      RECT 41.28 4.945 41.53 5.156 ;
      RECT 41.28 4.945 41.54 5.155 ;
      RECT 41.275 4.952 41.55 5.148 ;
      RECT 41.275 4.952 41.636 5.137 ;
      RECT 41.27 4.987 41.636 5.133 ;
      RECT 41.27 4.987 41.645 5.122 ;
      RECT 41.55 4.86 41.81 5.12 ;
      RECT 41.26 5.037 41.81 5.118 ;
      RECT 41.53 4.905 41.55 5.153 ;
      RECT 41.466 4.908 41.53 5.157 ;
      RECT 41.38 4.913 41.466 5.162 ;
      RECT 41.31 4.924 41.81 5.12 ;
      RECT 41.33 4.918 41.38 5.167 ;
      RECT 41.455 3.395 41.465 3.657 ;
      RECT 41.445 3.452 41.455 3.66 ;
      RECT 41.42 3.457 41.445 3.666 ;
      RECT 41.395 3.461 41.42 3.678 ;
      RECT 41.385 3.464 41.395 3.688 ;
      RECT 41.38 3.465 41.385 3.693 ;
      RECT 41.375 3.466 41.38 3.698 ;
      RECT 41.37 3.467 41.375 3.7 ;
      RECT 41.345 3.47 41.37 3.703 ;
      RECT 41.315 3.476 41.345 3.706 ;
      RECT 41.25 3.487 41.315 3.709 ;
      RECT 41.205 3.495 41.25 3.713 ;
      RECT 41.19 3.495 41.205 3.721 ;
      RECT 41.185 3.496 41.19 3.728 ;
      RECT 41.18 3.498 41.185 3.731 ;
      RECT 41.175 3.502 41.18 3.734 ;
      RECT 41.165 3.51 41.175 3.738 ;
      RECT 41.16 3.523 41.165 3.743 ;
      RECT 41.155 3.531 41.16 3.745 ;
      RECT 41.15 3.537 41.155 3.745 ;
      RECT 41.145 3.541 41.15 3.748 ;
      RECT 41.14 3.543 41.145 3.751 ;
      RECT 41.135 3.546 41.14 3.754 ;
      RECT 41.125 3.551 41.135 3.758 ;
      RECT 41.12 3.557 41.125 3.763 ;
      RECT 41.11 3.563 41.12 3.767 ;
      RECT 41.095 3.57 41.11 3.773 ;
      RECT 41.066 3.584 41.095 3.783 ;
      RECT 40.98 3.619 41.066 3.815 ;
      RECT 40.96 3.652 40.98 3.844 ;
      RECT 40.94 3.665 40.96 3.855 ;
      RECT 40.92 3.677 40.94 3.866 ;
      RECT 40.87 3.699 40.92 3.886 ;
      RECT 40.855 3.717 40.87 3.903 ;
      RECT 40.85 3.723 40.855 3.906 ;
      RECT 40.845 3.727 40.85 3.909 ;
      RECT 40.84 3.731 40.845 3.913 ;
      RECT 40.835 3.733 40.84 3.916 ;
      RECT 40.825 3.74 40.835 3.919 ;
      RECT 40.82 3.745 40.825 3.923 ;
      RECT 40.815 3.747 40.82 3.926 ;
      RECT 40.81 3.751 40.815 3.929 ;
      RECT 40.805 3.753 40.81 3.933 ;
      RECT 40.79 3.758 40.805 3.938 ;
      RECT 40.785 3.763 40.79 3.941 ;
      RECT 40.78 3.771 40.785 3.944 ;
      RECT 40.775 3.773 40.78 3.947 ;
      RECT 40.77 3.775 40.775 3.95 ;
      RECT 40.76 3.777 40.77 3.956 ;
      RECT 40.725 3.791 40.76 3.968 ;
      RECT 40.715 3.806 40.725 3.978 ;
      RECT 40.64 3.835 40.715 4.002 ;
      RECT 40.635 3.86 40.64 4.025 ;
      RECT 40.62 3.864 40.635 4.031 ;
      RECT 40.61 3.872 40.62 4.036 ;
      RECT 40.58 3.885 40.61 4.04 ;
      RECT 40.57 3.9 40.58 4.045 ;
      RECT 40.56 3.905 40.57 4.048 ;
      RECT 40.555 3.907 40.56 4.05 ;
      RECT 40.54 3.91 40.555 4.053 ;
      RECT 40.535 3.912 40.54 4.056 ;
      RECT 40.515 3.917 40.535 4.06 ;
      RECT 40.485 3.922 40.515 4.068 ;
      RECT 40.46 3.929 40.485 4.076 ;
      RECT 40.455 3.934 40.46 4.081 ;
      RECT 40.425 3.937 40.455 4.085 ;
      RECT 40.385 3.94 40.425 4.095 ;
      RECT 40.35 3.937 40.385 4.107 ;
      RECT 40.34 3.933 40.35 4.114 ;
      RECT 40.315 3.929 40.34 4.12 ;
      RECT 40.31 3.925 40.315 4.125 ;
      RECT 40.27 3.922 40.31 4.125 ;
      RECT 40.255 3.907 40.27 4.126 ;
      RECT 40.232 3.895 40.255 4.126 ;
      RECT 40.146 3.895 40.232 4.127 ;
      RECT 40.06 3.895 40.146 4.129 ;
      RECT 40.04 3.895 40.06 4.126 ;
      RECT 40.035 3.9 40.04 4.121 ;
      RECT 40.03 3.905 40.035 4.119 ;
      RECT 40.02 3.915 40.03 4.117 ;
      RECT 40.015 3.921 40.02 4.11 ;
      RECT 40.01 3.923 40.015 4.095 ;
      RECT 40.005 3.927 40.01 4.085 ;
      RECT 41.465 3.395 41.715 3.655 ;
      RECT 39.19 4.93 39.45 5.19 ;
      RECT 41.485 4.42 41.49 4.63 ;
      RECT 41.49 4.425 41.5 4.625 ;
      RECT 41.44 4.42 41.485 4.645 ;
      RECT 41.43 4.42 41.44 4.665 ;
      RECT 41.411 4.42 41.43 4.67 ;
      RECT 41.325 4.42 41.411 4.667 ;
      RECT 41.295 4.422 41.325 4.665 ;
      RECT 41.24 4.432 41.295 4.663 ;
      RECT 41.175 4.446 41.24 4.661 ;
      RECT 41.17 4.454 41.175 4.66 ;
      RECT 41.155 4.457 41.17 4.658 ;
      RECT 41.09 4.467 41.155 4.654 ;
      RECT 41.042 4.481 41.09 4.655 ;
      RECT 40.956 4.498 41.042 4.669 ;
      RECT 40.87 4.519 40.956 4.686 ;
      RECT 40.85 4.532 40.87 4.696 ;
      RECT 40.805 4.54 40.85 4.703 ;
      RECT 40.77 4.548 40.805 4.711 ;
      RECT 40.736 4.556 40.77 4.719 ;
      RECT 40.65 4.57 40.736 4.731 ;
      RECT 40.615 4.587 40.65 4.743 ;
      RECT 40.606 4.596 40.615 4.747 ;
      RECT 40.52 4.614 40.606 4.764 ;
      RECT 40.461 4.641 40.52 4.791 ;
      RECT 40.375 4.668 40.461 4.819 ;
      RECT 40.355 4.69 40.375 4.839 ;
      RECT 40.295 4.705 40.355 4.855 ;
      RECT 40.285 4.717 40.295 4.868 ;
      RECT 40.28 4.722 40.285 4.871 ;
      RECT 40.27 4.725 40.28 4.874 ;
      RECT 40.265 4.727 40.27 4.877 ;
      RECT 40.235 4.735 40.265 4.884 ;
      RECT 40.22 4.742 40.235 4.892 ;
      RECT 40.21 4.747 40.22 4.896 ;
      RECT 40.205 4.75 40.21 4.899 ;
      RECT 40.195 4.752 40.205 4.902 ;
      RECT 40.16 4.762 40.195 4.911 ;
      RECT 40.085 4.785 40.16 4.933 ;
      RECT 40.065 4.803 40.085 4.951 ;
      RECT 40.035 4.81 40.065 4.961 ;
      RECT 40.015 4.818 40.035 4.971 ;
      RECT 40.005 4.824 40.015 4.978 ;
      RECT 39.986 4.829 40.005 4.984 ;
      RECT 39.9 4.849 39.986 5.004 ;
      RECT 39.885 4.869 39.9 5.023 ;
      RECT 39.84 4.881 39.885 5.034 ;
      RECT 39.775 4.902 39.84 5.057 ;
      RECT 39.735 4.922 39.775 5.078 ;
      RECT 39.725 4.932 39.735 5.088 ;
      RECT 39.675 4.944 39.725 5.099 ;
      RECT 39.655 4.96 39.675 5.111 ;
      RECT 39.625 4.97 39.655 5.117 ;
      RECT 39.615 4.975 39.625 5.119 ;
      RECT 39.546 4.976 39.615 5.125 ;
      RECT 39.46 4.978 39.546 5.135 ;
      RECT 39.45 4.979 39.46 5.14 ;
      RECT 40.72 5.005 40.91 5.215 ;
      RECT 40.71 5.01 40.92 5.208 ;
      RECT 40.695 5.01 40.92 5.173 ;
      RECT 40.615 4.895 40.875 5.155 ;
      RECT 39.53 4.425 39.715 4.72 ;
      RECT 39.52 4.425 39.715 4.718 ;
      RECT 39.505 4.425 39.72 4.713 ;
      RECT 39.505 4.425 39.725 4.71 ;
      RECT 39.5 4.425 39.725 4.708 ;
      RECT 39.495 4.68 39.725 4.698 ;
      RECT 39.5 4.425 39.76 4.685 ;
      RECT 39.46 3.46 39.72 3.72 ;
      RECT 39.27 3.385 39.356 3.718 ;
      RECT 39.245 3.389 39.4 3.714 ;
      RECT 39.356 3.381 39.4 3.714 ;
      RECT 39.356 3.382 39.405 3.713 ;
      RECT 39.27 3.387 39.42 3.712 ;
      RECT 39.245 3.395 39.46 3.711 ;
      RECT 39.24 3.39 39.42 3.706 ;
      RECT 39.23 3.405 39.46 3.613 ;
      RECT 39.23 3.457 39.66 3.613 ;
      RECT 39.23 3.45 39.64 3.613 ;
      RECT 39.23 3.437 39.61 3.613 ;
      RECT 39.23 3.425 39.55 3.613 ;
      RECT 39.23 3.41 39.525 3.613 ;
      RECT 38.43 4.04 38.565 4.335 ;
      RECT 38.69 4.063 38.695 4.25 ;
      RECT 39.41 3.96 39.555 4.195 ;
      RECT 39.57 3.96 39.575 4.185 ;
      RECT 39.605 3.971 39.61 4.165 ;
      RECT 39.6 3.963 39.605 4.17 ;
      RECT 39.58 3.96 39.6 4.175 ;
      RECT 39.575 3.96 39.58 4.183 ;
      RECT 39.565 3.96 39.57 4.188 ;
      RECT 39.555 3.96 39.565 4.193 ;
      RECT 39.385 3.962 39.41 4.195 ;
      RECT 39.335 3.969 39.385 4.195 ;
      RECT 39.33 3.974 39.335 4.195 ;
      RECT 39.291 3.979 39.33 4.196 ;
      RECT 39.205 3.991 39.291 4.197 ;
      RECT 39.196 4.001 39.205 4.197 ;
      RECT 39.11 4.01 39.196 4.199 ;
      RECT 39.086 4.02 39.11 4.201 ;
      RECT 39 4.031 39.086 4.202 ;
      RECT 38.97 4.042 39 4.204 ;
      RECT 38.94 4.047 38.97 4.206 ;
      RECT 38.915 4.053 38.94 4.209 ;
      RECT 38.9 4.058 38.915 4.21 ;
      RECT 38.855 4.064 38.9 4.21 ;
      RECT 38.85 4.069 38.855 4.211 ;
      RECT 38.83 4.069 38.85 4.213 ;
      RECT 38.81 4.067 38.83 4.218 ;
      RECT 38.775 4.066 38.81 4.225 ;
      RECT 38.745 4.065 38.775 4.235 ;
      RECT 38.695 4.064 38.745 4.245 ;
      RECT 38.605 4.061 38.69 4.335 ;
      RECT 38.58 4.055 38.605 4.335 ;
      RECT 38.565 4.045 38.58 4.335 ;
      RECT 38.38 4.04 38.43 4.255 ;
      RECT 38.37 4.045 38.38 4.245 ;
      RECT 38.61 4.52 38.87 4.78 ;
      RECT 38.61 4.52 38.9 4.673 ;
      RECT 38.61 4.52 38.935 4.658 ;
      RECT 38.865 4.44 39.055 4.65 ;
      RECT 38.855 4.445 39.065 4.643 ;
      RECT 38.82 4.515 39.065 4.643 ;
      RECT 38.85 4.457 38.87 4.78 ;
      RECT 38.835 4.505 39.065 4.643 ;
      RECT 38.84 4.477 38.87 4.78 ;
      RECT 37.92 3.545 37.99 4.65 ;
      RECT 38.655 3.65 38.915 3.91 ;
      RECT 38.235 3.696 38.25 3.905 ;
      RECT 38.571 3.709 38.655 3.86 ;
      RECT 38.485 3.706 38.571 3.86 ;
      RECT 38.446 3.704 38.485 3.86 ;
      RECT 38.36 3.702 38.446 3.86 ;
      RECT 38.3 3.7 38.36 3.871 ;
      RECT 38.265 3.698 38.3 3.889 ;
      RECT 38.25 3.696 38.265 3.9 ;
      RECT 38.22 3.696 38.235 3.913 ;
      RECT 38.21 3.696 38.22 3.918 ;
      RECT 38.185 3.695 38.21 3.923 ;
      RECT 38.17 3.69 38.185 3.929 ;
      RECT 38.165 3.683 38.17 3.934 ;
      RECT 38.14 3.674 38.165 3.94 ;
      RECT 38.095 3.653 38.14 3.953 ;
      RECT 38.085 3.637 38.095 3.963 ;
      RECT 38.07 3.63 38.085 3.973 ;
      RECT 38.06 3.623 38.07 3.99 ;
      RECT 38.055 3.62 38.06 4.02 ;
      RECT 38.05 3.618 38.055 4.05 ;
      RECT 38.045 3.616 38.05 4.087 ;
      RECT 38.03 3.612 38.045 4.154 ;
      RECT 38.03 4.445 38.04 4.645 ;
      RECT 38.025 3.608 38.03 4.28 ;
      RECT 38.025 4.432 38.03 4.65 ;
      RECT 38.02 3.606 38.025 4.365 ;
      RECT 38.02 4.422 38.025 4.65 ;
      RECT 38.005 3.577 38.02 4.65 ;
      RECT 37.99 3.55 38.005 4.65 ;
      RECT 37.915 3.545 37.92 3.9 ;
      RECT 37.915 3.955 37.92 4.65 ;
      RECT 37.9 3.545 37.915 3.878 ;
      RECT 37.91 3.977 37.915 4.65 ;
      RECT 37.9 4.017 37.91 4.65 ;
      RECT 37.865 3.545 37.9 3.82 ;
      RECT 37.895 4.052 37.9 4.65 ;
      RECT 37.88 4.107 37.895 4.65 ;
      RECT 37.875 4.172 37.88 4.65 ;
      RECT 37.86 4.22 37.875 4.65 ;
      RECT 37.835 3.545 37.865 3.775 ;
      RECT 37.855 4.275 37.86 4.65 ;
      RECT 37.84 4.335 37.855 4.65 ;
      RECT 37.835 4.383 37.84 4.648 ;
      RECT 37.83 3.545 37.835 3.768 ;
      RECT 37.83 4.415 37.835 4.643 ;
      RECT 37.805 3.545 37.83 3.76 ;
      RECT 37.795 3.55 37.805 3.75 ;
      RECT 38.01 4.825 38.03 5.065 ;
      RECT 37.24 4.755 37.245 4.965 ;
      RECT 38.52 4.828 38.53 5.023 ;
      RECT 38.515 4.818 38.52 5.026 ;
      RECT 38.435 4.815 38.515 5.049 ;
      RECT 38.431 4.815 38.435 5.071 ;
      RECT 38.345 4.815 38.431 5.081 ;
      RECT 38.33 4.815 38.345 5.089 ;
      RECT 38.301 4.816 38.33 5.087 ;
      RECT 38.215 4.821 38.301 5.083 ;
      RECT 38.202 4.825 38.215 5.079 ;
      RECT 38.116 4.825 38.202 5.075 ;
      RECT 38.03 4.825 38.116 5.069 ;
      RECT 37.946 4.825 38.01 5.063 ;
      RECT 37.86 4.825 37.946 5.058 ;
      RECT 37.84 4.825 37.86 5.054 ;
      RECT 37.78 4.82 37.84 5.051 ;
      RECT 37.752 4.814 37.78 5.048 ;
      RECT 37.666 4.809 37.752 5.044 ;
      RECT 37.58 4.803 37.666 5.038 ;
      RECT 37.505 4.785 37.58 5.033 ;
      RECT 37.47 4.762 37.505 5.029 ;
      RECT 37.46 4.752 37.47 5.028 ;
      RECT 37.405 4.75 37.46 5.027 ;
      RECT 37.33 4.75 37.405 5.023 ;
      RECT 37.32 4.75 37.33 5.018 ;
      RECT 37.305 4.75 37.32 5.01 ;
      RECT 37.255 4.752 37.305 4.988 ;
      RECT 37.245 4.755 37.255 4.968 ;
      RECT 37.235 4.76 37.24 4.963 ;
      RECT 37.23 4.765 37.235 4.958 ;
      RECT 37.355 3.93 37.615 4.19 ;
      RECT 37.355 3.945 37.635 4.155 ;
      RECT 37.355 3.95 37.645 4.15 ;
      RECT 35.34 3.41 35.6 3.67 ;
      RECT 35.33 3.44 35.6 3.65 ;
      RECT 37.25 3.355 37.51 3.615 ;
      RECT 37.245 3.43 37.25 3.616 ;
      RECT 37.22 3.435 37.245 3.618 ;
      RECT 37.205 3.442 37.22 3.621 ;
      RECT 37.145 3.46 37.205 3.626 ;
      RECT 37.115 3.48 37.145 3.633 ;
      RECT 37.09 3.488 37.115 3.638 ;
      RECT 37.065 3.496 37.09 3.64 ;
      RECT 37.047 3.5 37.065 3.639 ;
      RECT 36.961 3.498 37.047 3.639 ;
      RECT 36.875 3.496 36.961 3.639 ;
      RECT 36.789 3.494 36.875 3.638 ;
      RECT 36.703 3.492 36.789 3.638 ;
      RECT 36.617 3.49 36.703 3.638 ;
      RECT 36.531 3.488 36.617 3.638 ;
      RECT 36.445 3.486 36.531 3.637 ;
      RECT 36.427 3.485 36.445 3.637 ;
      RECT 36.341 3.484 36.427 3.637 ;
      RECT 36.255 3.482 36.341 3.637 ;
      RECT 36.169 3.481 36.255 3.636 ;
      RECT 36.083 3.48 36.169 3.636 ;
      RECT 35.997 3.478 36.083 3.636 ;
      RECT 35.911 3.477 35.997 3.636 ;
      RECT 35.825 3.475 35.911 3.635 ;
      RECT 35.801 3.473 35.825 3.635 ;
      RECT 35.715 3.466 35.801 3.635 ;
      RECT 35.686 3.458 35.715 3.635 ;
      RECT 35.6 3.45 35.686 3.635 ;
      RECT 35.32 3.447 35.33 3.645 ;
      RECT 36.825 4.41 36.83 4.76 ;
      RECT 36.595 4.5 36.735 4.76 ;
      RECT 37.07 4.185 37.115 4.395 ;
      RECT 37.125 4.196 37.135 4.39 ;
      RECT 37.115 4.188 37.125 4.395 ;
      RECT 37.05 4.185 37.07 4.4 ;
      RECT 37.02 4.185 37.05 4.423 ;
      RECT 37.01 4.185 37.02 4.448 ;
      RECT 37.005 4.185 37.01 4.458 ;
      RECT 36.95 4.185 37.005 4.498 ;
      RECT 36.945 4.185 36.95 4.538 ;
      RECT 36.94 4.187 36.945 4.543 ;
      RECT 36.925 4.197 36.94 4.554 ;
      RECT 36.88 4.255 36.925 4.59 ;
      RECT 36.87 4.31 36.88 4.624 ;
      RECT 36.855 4.337 36.87 4.64 ;
      RECT 36.845 4.364 36.855 4.76 ;
      RECT 36.83 4.387 36.845 4.76 ;
      RECT 36.82 4.427 36.825 4.76 ;
      RECT 36.815 4.437 36.82 4.76 ;
      RECT 36.81 4.452 36.815 4.76 ;
      RECT 36.8 4.457 36.81 4.76 ;
      RECT 36.735 4.48 36.8 4.76 ;
      RECT 36.235 3.975 36.425 4.185 ;
      RECT 34.81 3.9 35.07 4.16 ;
      RECT 35.16 3.895 35.255 4.105 ;
      RECT 35.135 3.91 35.145 4.105 ;
      RECT 36.425 3.982 36.435 4.18 ;
      RECT 36.225 3.982 36.235 4.18 ;
      RECT 36.21 3.997 36.225 4.17 ;
      RECT 36.205 4.005 36.21 4.163 ;
      RECT 36.195 4.008 36.205 4.16 ;
      RECT 36.16 4.007 36.195 4.158 ;
      RECT 36.131 4.003 36.16 4.155 ;
      RECT 36.045 3.998 36.131 4.152 ;
      RECT 35.985 3.992 36.045 4.148 ;
      RECT 35.956 3.988 35.985 4.145 ;
      RECT 35.87 3.98 35.956 4.142 ;
      RECT 35.861 3.974 35.87 4.14 ;
      RECT 35.775 3.969 35.861 4.138 ;
      RECT 35.752 3.964 35.775 4.135 ;
      RECT 35.666 3.958 35.752 4.132 ;
      RECT 35.58 3.949 35.666 4.127 ;
      RECT 35.57 3.944 35.58 4.125 ;
      RECT 35.551 3.943 35.57 4.124 ;
      RECT 35.465 3.938 35.551 4.12 ;
      RECT 35.445 3.933 35.465 4.116 ;
      RECT 35.385 3.928 35.445 4.113 ;
      RECT 35.36 3.918 35.385 4.111 ;
      RECT 35.355 3.911 35.36 4.11 ;
      RECT 35.345 3.902 35.355 4.109 ;
      RECT 35.341 3.895 35.345 4.109 ;
      RECT 35.255 3.895 35.341 4.107 ;
      RECT 35.145 3.902 35.16 4.105 ;
      RECT 35.13 3.912 35.135 4.105 ;
      RECT 35.11 3.915 35.13 4.102 ;
      RECT 35.08 3.915 35.11 4.098 ;
      RECT 35.07 3.915 35.08 4.098 ;
      RECT 35.985 4.41 36.245 4.67 ;
      RECT 35.915 4.42 36.245 4.63 ;
      RECT 35.905 4.427 36.245 4.625 ;
      RECT 35.325 4.415 35.585 4.675 ;
      RECT 35.325 4.455 35.69 4.665 ;
      RECT 35.325 4.457 35.695 4.664 ;
      RECT 35.325 4.465 35.7 4.661 ;
      RECT 34.25 3.54 34.35 5.065 ;
      RECT 34.44 4.68 34.49 4.94 ;
      RECT 34.435 3.553 34.44 3.74 ;
      RECT 34.43 4.661 34.44 4.94 ;
      RECT 34.43 3.55 34.435 3.748 ;
      RECT 34.415 3.544 34.43 3.755 ;
      RECT 34.425 4.649 34.43 5.023 ;
      RECT 34.415 4.637 34.425 5.06 ;
      RECT 34.405 3.54 34.415 3.762 ;
      RECT 34.405 4.622 34.415 5.065 ;
      RECT 34.4 3.54 34.405 3.77 ;
      RECT 34.38 4.592 34.405 5.065 ;
      RECT 34.36 3.54 34.4 3.818 ;
      RECT 34.37 4.552 34.38 5.065 ;
      RECT 34.36 4.507 34.37 5.065 ;
      RECT 34.355 3.54 34.36 3.888 ;
      RECT 34.355 4.465 34.36 5.065 ;
      RECT 34.35 3.54 34.355 4.365 ;
      RECT 34.35 4.447 34.355 5.065 ;
      RECT 34.24 3.543 34.25 5.065 ;
      RECT 34.225 3.55 34.24 5.061 ;
      RECT 34.22 3.56 34.225 5.056 ;
      RECT 34.215 3.76 34.22 4.948 ;
      RECT 34.21 3.845 34.215 4.5 ;
      RECT 33.085 10.205 33.375 10.435 ;
      RECT 33.145 8.725 33.315 10.435 ;
      RECT 33.14 9.09 33.49 9.44 ;
      RECT 33.085 8.725 33.375 8.955 ;
      RECT 32.68 3.69 32.785 4.26 ;
      RECT 32.68 4.025 33.005 4.255 ;
      RECT 32.68 4.055 33.175 4.225 ;
      RECT 32.68 3.69 32.87 4.255 ;
      RECT 32.095 3.655 32.385 3.885 ;
      RECT 32.095 3.69 32.87 3.86 ;
      RECT 32.155 2.175 32.325 3.885 ;
      RECT 32.095 2.175 32.385 2.405 ;
      RECT 32.095 10.205 32.385 10.435 ;
      RECT 32.155 8.725 32.325 10.435 ;
      RECT 32.095 8.725 32.385 8.955 ;
      RECT 32.095 8.76 32.95 8.92 ;
      RECT 32.78 8.355 32.95 8.92 ;
      RECT 32.095 8.755 32.49 8.92 ;
      RECT 32.715 8.355 33.005 8.585 ;
      RECT 32.715 8.385 33.175 8.555 ;
      RECT 31.725 4.025 32.015 4.255 ;
      RECT 31.725 4.055 32.185 4.225 ;
      RECT 31.79 2.95 31.955 4.255 ;
      RECT 30.305 2.92 30.595 3.15 ;
      RECT 30.305 2.95 31.955 3.12 ;
      RECT 30.365 2.18 30.535 3.15 ;
      RECT 30.305 2.18 30.595 2.41 ;
      RECT 30.305 10.2 30.595 10.43 ;
      RECT 30.365 9.46 30.535 10.43 ;
      RECT 30.365 9.555 31.955 9.725 ;
      RECT 31.785 8.355 31.955 9.725 ;
      RECT 30.305 9.46 30.595 9.69 ;
      RECT 31.725 8.355 32.015 8.585 ;
      RECT 31.725 8.385 32.185 8.555 ;
      RECT 28.34 4.725 28.69 5.075 ;
      RECT 28.43 3.32 28.6 5.075 ;
      RECT 30.735 3.26 31.085 3.61 ;
      RECT 28.43 3.32 30.05 3.495 ;
      RECT 28.43 3.32 31.085 3.49 ;
      RECT 30.76 9.09 31.085 9.415 ;
      RECT 26.155 9.04 26.505 9.39 ;
      RECT 30.735 9.09 31.085 9.32 ;
      RECT 25.975 9.09 26.505 9.32 ;
      RECT 25.805 9.12 31.085 9.29 ;
      RECT 29.96 3.66 30.28 3.98 ;
      RECT 29.93 3.66 30.28 3.89 ;
      RECT 29.76 3.69 30.28 3.86 ;
      RECT 29.96 8.66 30.28 8.98 ;
      RECT 29.93 8.72 30.28 8.95 ;
      RECT 29.76 8.75 30.28 8.92 ;
      RECT 25.74 4.96 25.78 5.22 ;
      RECT 25.78 4.94 25.785 4.95 ;
      RECT 27.11 4.185 27.12 4.406 ;
      RECT 27.04 4.18 27.11 4.531 ;
      RECT 27.03 4.18 27.04 4.658 ;
      RECT 27.005 4.18 27.03 4.705 ;
      RECT 26.98 4.18 27.005 4.783 ;
      RECT 26.96 4.18 26.98 4.853 ;
      RECT 26.935 4.18 26.96 4.893 ;
      RECT 26.925 4.18 26.935 4.913 ;
      RECT 26.915 4.182 26.925 4.921 ;
      RECT 26.91 4.187 26.915 4.378 ;
      RECT 26.91 4.387 26.915 4.922 ;
      RECT 26.905 4.432 26.91 4.923 ;
      RECT 26.895 4.497 26.905 4.924 ;
      RECT 26.885 4.592 26.895 4.926 ;
      RECT 26.88 4.645 26.885 4.928 ;
      RECT 26.875 4.665 26.88 4.929 ;
      RECT 26.82 4.69 26.875 4.935 ;
      RECT 26.78 4.725 26.82 4.944 ;
      RECT 26.77 4.742 26.78 4.949 ;
      RECT 26.761 4.748 26.77 4.951 ;
      RECT 26.675 4.786 26.761 4.962 ;
      RECT 26.67 4.825 26.675 4.972 ;
      RECT 26.595 4.832 26.67 4.982 ;
      RECT 26.575 4.842 26.595 4.993 ;
      RECT 26.545 4.849 26.575 5.001 ;
      RECT 26.52 4.856 26.545 5.008 ;
      RECT 26.496 4.862 26.52 5.013 ;
      RECT 26.41 4.875 26.496 5.025 ;
      RECT 26.332 4.882 26.41 5.043 ;
      RECT 26.246 4.877 26.332 5.061 ;
      RECT 26.16 4.872 26.246 5.081 ;
      RECT 26.08 4.866 26.16 5.098 ;
      RECT 26.015 4.862 26.08 5.127 ;
      RECT 26.01 4.576 26.015 4.6 ;
      RECT 26 4.852 26.015 5.155 ;
      RECT 26.005 4.57 26.01 4.64 ;
      RECT 26 4.564 26.005 4.71 ;
      RECT 25.995 4.558 26 4.788 ;
      RECT 25.995 4.835 26 5.22 ;
      RECT 25.987 4.555 25.995 5.22 ;
      RECT 25.901 4.553 25.987 5.22 ;
      RECT 25.815 4.551 25.901 5.22 ;
      RECT 25.805 4.552 25.815 5.22 ;
      RECT 25.8 4.557 25.805 5.22 ;
      RECT 25.79 4.57 25.8 5.22 ;
      RECT 25.785 4.592 25.79 5.22 ;
      RECT 25.78 4.952 25.785 5.22 ;
      RECT 26.41 4.42 26.415 4.64 ;
      RECT 26.915 3.455 26.95 3.715 ;
      RECT 26.9 3.455 26.915 3.723 ;
      RECT 26.871 3.455 26.9 3.745 ;
      RECT 26.785 3.455 26.871 3.805 ;
      RECT 26.765 3.455 26.785 3.87 ;
      RECT 26.705 3.455 26.765 4.035 ;
      RECT 26.7 3.455 26.705 4.183 ;
      RECT 26.695 3.455 26.7 4.195 ;
      RECT 26.69 3.455 26.695 4.221 ;
      RECT 26.66 3.641 26.69 4.301 ;
      RECT 26.655 3.689 26.66 4.39 ;
      RECT 26.65 3.703 26.655 4.405 ;
      RECT 26.645 3.722 26.65 4.435 ;
      RECT 26.64 3.737 26.645 4.451 ;
      RECT 26.635 3.752 26.64 4.473 ;
      RECT 26.63 3.772 26.635 4.495 ;
      RECT 26.62 3.792 26.63 4.528 ;
      RECT 26.605 3.834 26.62 4.59 ;
      RECT 26.6 3.865 26.605 4.63 ;
      RECT 26.595 3.877 26.6 4.635 ;
      RECT 26.59 3.889 26.595 4.64 ;
      RECT 26.585 3.902 26.59 4.64 ;
      RECT 26.58 3.92 26.585 4.64 ;
      RECT 26.575 3.94 26.58 4.64 ;
      RECT 26.57 3.952 26.575 4.64 ;
      RECT 26.565 3.965 26.57 4.64 ;
      RECT 26.545 4 26.565 4.64 ;
      RECT 26.495 4.102 26.545 4.64 ;
      RECT 26.49 4.187 26.495 4.64 ;
      RECT 26.485 4.195 26.49 4.64 ;
      RECT 26.48 4.212 26.485 4.64 ;
      RECT 26.475 4.227 26.48 4.64 ;
      RECT 26.44 4.292 26.475 4.64 ;
      RECT 26.425 4.357 26.44 4.64 ;
      RECT 26.42 4.387 26.425 4.64 ;
      RECT 26.415 4.412 26.42 4.64 ;
      RECT 26.4 4.422 26.41 4.64 ;
      RECT 26.385 4.435 26.4 4.633 ;
      RECT 26.13 4.025 26.2 4.235 ;
      RECT 25.92 4.002 25.925 4.195 ;
      RECT 23.375 3.93 23.635 4.19 ;
      RECT 26.21 4.212 26.215 4.215 ;
      RECT 26.2 4.03 26.21 4.23 ;
      RECT 26.101 4.023 26.13 4.235 ;
      RECT 26.015 4.015 26.101 4.235 ;
      RECT 26 4.009 26.015 4.233 ;
      RECT 25.98 4.008 26 4.22 ;
      RECT 25.975 4.007 25.98 4.203 ;
      RECT 25.925 4.004 25.975 4.198 ;
      RECT 25.895 4.001 25.92 4.193 ;
      RECT 25.875 3.999 25.895 4.188 ;
      RECT 25.86 3.997 25.875 4.185 ;
      RECT 25.83 3.995 25.86 4.183 ;
      RECT 25.765 3.991 25.83 4.175 ;
      RECT 25.735 3.986 25.765 4.17 ;
      RECT 25.715 3.984 25.735 4.168 ;
      RECT 25.685 3.981 25.715 4.163 ;
      RECT 25.625 3.977 25.685 4.155 ;
      RECT 25.62 3.974 25.625 4.15 ;
      RECT 25.55 3.972 25.62 4.145 ;
      RECT 25.521 3.968 25.55 4.138 ;
      RECT 25.435 3.963 25.521 4.13 ;
      RECT 25.401 3.958 25.435 4.122 ;
      RECT 25.315 3.95 25.401 4.114 ;
      RECT 25.276 3.943 25.315 4.106 ;
      RECT 25.19 3.938 25.276 4.098 ;
      RECT 25.125 3.932 25.19 4.088 ;
      RECT 25.105 3.927 25.125 4.083 ;
      RECT 25.096 3.924 25.105 4.082 ;
      RECT 25.01 3.92 25.096 4.076 ;
      RECT 24.97 3.916 25.01 4.068 ;
      RECT 24.95 3.912 24.97 4.066 ;
      RECT 24.89 3.912 24.95 4.063 ;
      RECT 24.87 3.915 24.89 4.061 ;
      RECT 24.849 3.915 24.87 4.061 ;
      RECT 24.763 3.917 24.849 4.065 ;
      RECT 24.677 3.919 24.763 4.071 ;
      RECT 24.591 3.921 24.677 4.078 ;
      RECT 24.505 3.924 24.591 4.084 ;
      RECT 24.471 3.925 24.505 4.089 ;
      RECT 24.385 3.928 24.471 4.094 ;
      RECT 24.356 3.935 24.385 4.099 ;
      RECT 24.27 3.935 24.356 4.104 ;
      RECT 24.237 3.935 24.27 4.109 ;
      RECT 24.151 3.937 24.237 4.114 ;
      RECT 24.065 3.939 24.151 4.121 ;
      RECT 24.001 3.941 24.065 4.127 ;
      RECT 23.915 3.943 24.001 4.133 ;
      RECT 23.912 3.945 23.915 4.136 ;
      RECT 23.826 3.946 23.912 4.14 ;
      RECT 23.74 3.949 23.826 4.147 ;
      RECT 23.721 3.951 23.74 4.151 ;
      RECT 23.635 3.953 23.721 4.156 ;
      RECT 23.365 3.965 23.375 4.16 ;
      RECT 25.545 10.2 25.835 10.43 ;
      RECT 25.605 9.46 25.775 10.43 ;
      RECT 25.495 9.49 25.87 9.86 ;
      RECT 25.545 9.46 25.835 9.86 ;
      RECT 25.6 3.545 25.785 3.755 ;
      RECT 25.595 3.546 25.79 3.753 ;
      RECT 25.59 3.551 25.8 3.748 ;
      RECT 25.585 3.527 25.59 3.745 ;
      RECT 25.555 3.524 25.585 3.738 ;
      RECT 25.55 3.52 25.555 3.729 ;
      RECT 25.515 3.551 25.8 3.724 ;
      RECT 25.29 3.46 25.55 3.72 ;
      RECT 25.59 3.529 25.595 3.748 ;
      RECT 25.595 3.53 25.6 3.753 ;
      RECT 25.29 3.542 25.67 3.72 ;
      RECT 25.29 3.54 25.655 3.72 ;
      RECT 25.29 3.535 25.645 3.72 ;
      RECT 25.245 4.45 25.295 4.735 ;
      RECT 25.19 4.42 25.195 4.735 ;
      RECT 25.16 4.4 25.165 4.735 ;
      RECT 25.31 4.45 25.37 4.71 ;
      RECT 25.305 4.45 25.31 4.718 ;
      RECT 25.295 4.45 25.305 4.73 ;
      RECT 25.21 4.44 25.245 4.735 ;
      RECT 25.205 4.427 25.21 4.735 ;
      RECT 25.195 4.422 25.205 4.735 ;
      RECT 25.175 4.412 25.19 4.735 ;
      RECT 25.165 4.405 25.175 4.735 ;
      RECT 25.155 4.397 25.16 4.735 ;
      RECT 25.125 4.387 25.155 4.735 ;
      RECT 25.11 4.375 25.125 4.735 ;
      RECT 25.095 4.365 25.11 4.73 ;
      RECT 25.075 4.355 25.095 4.705 ;
      RECT 25.065 4.347 25.075 4.682 ;
      RECT 25.035 4.33 25.065 4.672 ;
      RECT 25.03 4.307 25.035 4.663 ;
      RECT 25.025 4.294 25.03 4.661 ;
      RECT 25.01 4.27 25.025 4.655 ;
      RECT 25.005 4.246 25.01 4.649 ;
      RECT 24.995 4.235 25.005 4.644 ;
      RECT 24.99 4.225 24.995 4.64 ;
      RECT 24.985 4.217 24.99 4.637 ;
      RECT 24.975 4.212 24.985 4.633 ;
      RECT 24.97 4.207 24.975 4.629 ;
      RECT 24.885 4.205 24.97 4.604 ;
      RECT 24.855 4.205 24.885 4.57 ;
      RECT 24.84 4.205 24.855 4.553 ;
      RECT 24.785 4.205 24.84 4.498 ;
      RECT 24.78 4.21 24.785 4.447 ;
      RECT 24.77 4.215 24.78 4.437 ;
      RECT 24.765 4.225 24.77 4.423 ;
      RECT 24.715 4.965 24.975 5.225 ;
      RECT 24.635 4.98 24.975 5.201 ;
      RECT 24.615 4.98 24.975 5.196 ;
      RECT 24.591 4.98 24.975 5.194 ;
      RECT 24.505 4.98 24.975 5.189 ;
      RECT 24.355 4.92 24.615 5.185 ;
      RECT 24.31 4.98 24.975 5.18 ;
      RECT 24.305 4.987 24.975 5.175 ;
      RECT 24.32 4.975 24.635 5.185 ;
      RECT 24.21 3.41 24.47 3.67 ;
      RECT 24.21 3.467 24.475 3.663 ;
      RECT 24.21 3.497 24.48 3.595 ;
      RECT 24.27 3.928 24.385 3.93 ;
      RECT 24.356 3.925 24.385 3.93 ;
      RECT 23.38 4.929 23.405 5.169 ;
      RECT 23.365 4.932 23.455 5.163 ;
      RECT 23.36 4.937 23.541 5.158 ;
      RECT 23.355 4.945 23.605 5.156 ;
      RECT 23.355 4.945 23.615 5.155 ;
      RECT 23.35 4.952 23.625 5.148 ;
      RECT 23.35 4.952 23.711 5.137 ;
      RECT 23.345 4.987 23.711 5.133 ;
      RECT 23.345 4.987 23.72 5.122 ;
      RECT 23.625 4.86 23.885 5.12 ;
      RECT 23.335 5.037 23.885 5.118 ;
      RECT 23.605 4.905 23.625 5.153 ;
      RECT 23.541 4.908 23.605 5.157 ;
      RECT 23.455 4.913 23.541 5.162 ;
      RECT 23.385 4.924 23.885 5.12 ;
      RECT 23.405 4.918 23.455 5.167 ;
      RECT 23.53 3.395 23.54 3.657 ;
      RECT 23.52 3.452 23.53 3.66 ;
      RECT 23.495 3.457 23.52 3.666 ;
      RECT 23.47 3.461 23.495 3.678 ;
      RECT 23.46 3.464 23.47 3.688 ;
      RECT 23.455 3.465 23.46 3.693 ;
      RECT 23.45 3.466 23.455 3.698 ;
      RECT 23.445 3.467 23.45 3.7 ;
      RECT 23.42 3.47 23.445 3.703 ;
      RECT 23.39 3.476 23.42 3.706 ;
      RECT 23.325 3.487 23.39 3.709 ;
      RECT 23.28 3.495 23.325 3.713 ;
      RECT 23.265 3.495 23.28 3.721 ;
      RECT 23.26 3.496 23.265 3.728 ;
      RECT 23.255 3.498 23.26 3.731 ;
      RECT 23.25 3.502 23.255 3.734 ;
      RECT 23.24 3.51 23.25 3.738 ;
      RECT 23.235 3.523 23.24 3.743 ;
      RECT 23.23 3.531 23.235 3.745 ;
      RECT 23.225 3.537 23.23 3.745 ;
      RECT 23.22 3.541 23.225 3.748 ;
      RECT 23.215 3.543 23.22 3.751 ;
      RECT 23.21 3.546 23.215 3.754 ;
      RECT 23.2 3.551 23.21 3.758 ;
      RECT 23.195 3.557 23.2 3.763 ;
      RECT 23.185 3.563 23.195 3.767 ;
      RECT 23.17 3.57 23.185 3.773 ;
      RECT 23.141 3.584 23.17 3.783 ;
      RECT 23.055 3.619 23.141 3.815 ;
      RECT 23.035 3.652 23.055 3.844 ;
      RECT 23.015 3.665 23.035 3.855 ;
      RECT 22.995 3.677 23.015 3.866 ;
      RECT 22.945 3.699 22.995 3.886 ;
      RECT 22.93 3.717 22.945 3.903 ;
      RECT 22.925 3.723 22.93 3.906 ;
      RECT 22.92 3.727 22.925 3.909 ;
      RECT 22.915 3.731 22.92 3.913 ;
      RECT 22.91 3.733 22.915 3.916 ;
      RECT 22.9 3.74 22.91 3.919 ;
      RECT 22.895 3.745 22.9 3.923 ;
      RECT 22.89 3.747 22.895 3.926 ;
      RECT 22.885 3.751 22.89 3.929 ;
      RECT 22.88 3.753 22.885 3.933 ;
      RECT 22.865 3.758 22.88 3.938 ;
      RECT 22.86 3.763 22.865 3.941 ;
      RECT 22.855 3.771 22.86 3.944 ;
      RECT 22.85 3.773 22.855 3.947 ;
      RECT 22.845 3.775 22.85 3.95 ;
      RECT 22.835 3.777 22.845 3.956 ;
      RECT 22.8 3.791 22.835 3.968 ;
      RECT 22.79 3.806 22.8 3.978 ;
      RECT 22.715 3.835 22.79 4.002 ;
      RECT 22.71 3.86 22.715 4.025 ;
      RECT 22.695 3.864 22.71 4.031 ;
      RECT 22.685 3.872 22.695 4.036 ;
      RECT 22.655 3.885 22.685 4.04 ;
      RECT 22.645 3.9 22.655 4.045 ;
      RECT 22.635 3.905 22.645 4.048 ;
      RECT 22.63 3.907 22.635 4.05 ;
      RECT 22.615 3.91 22.63 4.053 ;
      RECT 22.61 3.912 22.615 4.056 ;
      RECT 22.59 3.917 22.61 4.06 ;
      RECT 22.56 3.922 22.59 4.068 ;
      RECT 22.535 3.929 22.56 4.076 ;
      RECT 22.53 3.934 22.535 4.081 ;
      RECT 22.5 3.937 22.53 4.085 ;
      RECT 22.46 3.94 22.5 4.095 ;
      RECT 22.425 3.937 22.46 4.107 ;
      RECT 22.415 3.933 22.425 4.114 ;
      RECT 22.39 3.929 22.415 4.12 ;
      RECT 22.385 3.925 22.39 4.125 ;
      RECT 22.345 3.922 22.385 4.125 ;
      RECT 22.33 3.907 22.345 4.126 ;
      RECT 22.307 3.895 22.33 4.126 ;
      RECT 22.221 3.895 22.307 4.127 ;
      RECT 22.135 3.895 22.221 4.129 ;
      RECT 22.115 3.895 22.135 4.126 ;
      RECT 22.11 3.9 22.115 4.121 ;
      RECT 22.105 3.905 22.11 4.119 ;
      RECT 22.095 3.915 22.105 4.117 ;
      RECT 22.09 3.921 22.095 4.11 ;
      RECT 22.085 3.923 22.09 4.095 ;
      RECT 22.08 3.927 22.085 4.085 ;
      RECT 23.54 3.395 23.79 3.655 ;
      RECT 21.265 4.93 21.525 5.19 ;
      RECT 23.56 4.42 23.565 4.63 ;
      RECT 23.565 4.425 23.575 4.625 ;
      RECT 23.515 4.42 23.56 4.645 ;
      RECT 23.505 4.42 23.515 4.665 ;
      RECT 23.486 4.42 23.505 4.67 ;
      RECT 23.4 4.42 23.486 4.667 ;
      RECT 23.37 4.422 23.4 4.665 ;
      RECT 23.315 4.432 23.37 4.663 ;
      RECT 23.25 4.446 23.315 4.661 ;
      RECT 23.245 4.454 23.25 4.66 ;
      RECT 23.23 4.457 23.245 4.658 ;
      RECT 23.165 4.467 23.23 4.654 ;
      RECT 23.117 4.481 23.165 4.655 ;
      RECT 23.031 4.498 23.117 4.669 ;
      RECT 22.945 4.519 23.031 4.686 ;
      RECT 22.925 4.532 22.945 4.696 ;
      RECT 22.88 4.54 22.925 4.703 ;
      RECT 22.845 4.548 22.88 4.711 ;
      RECT 22.811 4.556 22.845 4.719 ;
      RECT 22.725 4.57 22.811 4.731 ;
      RECT 22.69 4.587 22.725 4.743 ;
      RECT 22.681 4.596 22.69 4.747 ;
      RECT 22.595 4.614 22.681 4.764 ;
      RECT 22.536 4.641 22.595 4.791 ;
      RECT 22.45 4.668 22.536 4.819 ;
      RECT 22.43 4.69 22.45 4.839 ;
      RECT 22.37 4.705 22.43 4.855 ;
      RECT 22.36 4.717 22.37 4.868 ;
      RECT 22.355 4.722 22.36 4.871 ;
      RECT 22.345 4.725 22.355 4.874 ;
      RECT 22.34 4.727 22.345 4.877 ;
      RECT 22.31 4.735 22.34 4.884 ;
      RECT 22.295 4.742 22.31 4.892 ;
      RECT 22.285 4.747 22.295 4.896 ;
      RECT 22.28 4.75 22.285 4.899 ;
      RECT 22.27 4.752 22.28 4.902 ;
      RECT 22.235 4.762 22.27 4.911 ;
      RECT 22.16 4.785 22.235 4.933 ;
      RECT 22.14 4.803 22.16 4.951 ;
      RECT 22.11 4.81 22.14 4.961 ;
      RECT 22.09 4.818 22.11 4.971 ;
      RECT 22.08 4.824 22.09 4.978 ;
      RECT 22.061 4.829 22.08 4.984 ;
      RECT 21.975 4.849 22.061 5.004 ;
      RECT 21.96 4.869 21.975 5.023 ;
      RECT 21.915 4.881 21.96 5.034 ;
      RECT 21.85 4.902 21.915 5.057 ;
      RECT 21.81 4.922 21.85 5.078 ;
      RECT 21.8 4.932 21.81 5.088 ;
      RECT 21.75 4.944 21.8 5.099 ;
      RECT 21.73 4.96 21.75 5.111 ;
      RECT 21.7 4.97 21.73 5.117 ;
      RECT 21.69 4.975 21.7 5.119 ;
      RECT 21.621 4.976 21.69 5.125 ;
      RECT 21.535 4.978 21.621 5.135 ;
      RECT 21.525 4.979 21.535 5.14 ;
      RECT 22.795 5.005 22.985 5.215 ;
      RECT 22.785 5.01 22.995 5.208 ;
      RECT 22.77 5.01 22.995 5.173 ;
      RECT 22.69 4.895 22.95 5.155 ;
      RECT 21.605 4.425 21.79 4.72 ;
      RECT 21.595 4.425 21.79 4.718 ;
      RECT 21.58 4.425 21.795 4.713 ;
      RECT 21.58 4.425 21.8 4.71 ;
      RECT 21.575 4.425 21.8 4.708 ;
      RECT 21.57 4.68 21.8 4.698 ;
      RECT 21.575 4.425 21.835 4.685 ;
      RECT 21.535 3.46 21.795 3.72 ;
      RECT 21.345 3.385 21.431 3.718 ;
      RECT 21.32 3.389 21.475 3.714 ;
      RECT 21.431 3.381 21.475 3.714 ;
      RECT 21.431 3.382 21.48 3.713 ;
      RECT 21.345 3.387 21.495 3.712 ;
      RECT 21.32 3.395 21.535 3.711 ;
      RECT 21.315 3.39 21.495 3.706 ;
      RECT 21.305 3.405 21.535 3.613 ;
      RECT 21.305 3.457 21.735 3.613 ;
      RECT 21.305 3.45 21.715 3.613 ;
      RECT 21.305 3.437 21.685 3.613 ;
      RECT 21.305 3.425 21.625 3.613 ;
      RECT 21.305 3.41 21.6 3.613 ;
      RECT 20.505 4.04 20.64 4.335 ;
      RECT 20.765 4.063 20.77 4.25 ;
      RECT 21.485 3.96 21.63 4.195 ;
      RECT 21.645 3.96 21.65 4.185 ;
      RECT 21.68 3.971 21.685 4.165 ;
      RECT 21.675 3.963 21.68 4.17 ;
      RECT 21.655 3.96 21.675 4.175 ;
      RECT 21.65 3.96 21.655 4.183 ;
      RECT 21.64 3.96 21.645 4.188 ;
      RECT 21.63 3.96 21.64 4.193 ;
      RECT 21.46 3.962 21.485 4.195 ;
      RECT 21.41 3.969 21.46 4.195 ;
      RECT 21.405 3.974 21.41 4.195 ;
      RECT 21.366 3.979 21.405 4.196 ;
      RECT 21.28 3.991 21.366 4.197 ;
      RECT 21.271 4.001 21.28 4.197 ;
      RECT 21.185 4.01 21.271 4.199 ;
      RECT 21.161 4.02 21.185 4.201 ;
      RECT 21.075 4.031 21.161 4.202 ;
      RECT 21.045 4.042 21.075 4.204 ;
      RECT 21.015 4.047 21.045 4.206 ;
      RECT 20.99 4.053 21.015 4.209 ;
      RECT 20.975 4.058 20.99 4.21 ;
      RECT 20.93 4.064 20.975 4.21 ;
      RECT 20.925 4.069 20.93 4.211 ;
      RECT 20.905 4.069 20.925 4.213 ;
      RECT 20.885 4.067 20.905 4.218 ;
      RECT 20.85 4.066 20.885 4.225 ;
      RECT 20.82 4.065 20.85 4.235 ;
      RECT 20.77 4.064 20.82 4.245 ;
      RECT 20.68 4.061 20.765 4.335 ;
      RECT 20.655 4.055 20.68 4.335 ;
      RECT 20.64 4.045 20.655 4.335 ;
      RECT 20.455 4.04 20.505 4.255 ;
      RECT 20.445 4.045 20.455 4.245 ;
      RECT 20.685 4.52 20.945 4.78 ;
      RECT 20.685 4.52 20.975 4.673 ;
      RECT 20.685 4.52 21.01 4.658 ;
      RECT 20.94 4.44 21.13 4.65 ;
      RECT 20.93 4.445 21.14 4.643 ;
      RECT 20.895 4.515 21.14 4.643 ;
      RECT 20.925 4.457 20.945 4.78 ;
      RECT 20.91 4.505 21.14 4.643 ;
      RECT 20.915 4.477 20.945 4.78 ;
      RECT 19.995 3.545 20.065 4.65 ;
      RECT 20.73 3.65 20.99 3.91 ;
      RECT 20.31 3.696 20.325 3.905 ;
      RECT 20.646 3.709 20.73 3.86 ;
      RECT 20.56 3.706 20.646 3.86 ;
      RECT 20.521 3.704 20.56 3.86 ;
      RECT 20.435 3.702 20.521 3.86 ;
      RECT 20.375 3.7 20.435 3.871 ;
      RECT 20.34 3.698 20.375 3.889 ;
      RECT 20.325 3.696 20.34 3.9 ;
      RECT 20.295 3.696 20.31 3.913 ;
      RECT 20.285 3.696 20.295 3.918 ;
      RECT 20.26 3.695 20.285 3.923 ;
      RECT 20.245 3.69 20.26 3.929 ;
      RECT 20.24 3.683 20.245 3.934 ;
      RECT 20.215 3.674 20.24 3.94 ;
      RECT 20.17 3.653 20.215 3.953 ;
      RECT 20.16 3.637 20.17 3.963 ;
      RECT 20.145 3.63 20.16 3.973 ;
      RECT 20.135 3.623 20.145 3.99 ;
      RECT 20.13 3.62 20.135 4.02 ;
      RECT 20.125 3.618 20.13 4.05 ;
      RECT 20.12 3.616 20.125 4.087 ;
      RECT 20.105 3.612 20.12 4.154 ;
      RECT 20.105 4.445 20.115 4.645 ;
      RECT 20.1 3.608 20.105 4.28 ;
      RECT 20.1 4.432 20.105 4.65 ;
      RECT 20.095 3.606 20.1 4.365 ;
      RECT 20.095 4.422 20.1 4.65 ;
      RECT 20.08 3.577 20.095 4.65 ;
      RECT 20.065 3.55 20.08 4.65 ;
      RECT 19.99 3.545 19.995 3.9 ;
      RECT 19.99 3.955 19.995 4.65 ;
      RECT 19.975 3.545 19.99 3.878 ;
      RECT 19.985 3.977 19.99 4.65 ;
      RECT 19.975 4.017 19.985 4.65 ;
      RECT 19.94 3.545 19.975 3.82 ;
      RECT 19.97 4.052 19.975 4.65 ;
      RECT 19.955 4.107 19.97 4.65 ;
      RECT 19.95 4.172 19.955 4.65 ;
      RECT 19.935 4.22 19.95 4.65 ;
      RECT 19.91 3.545 19.94 3.775 ;
      RECT 19.93 4.275 19.935 4.65 ;
      RECT 19.915 4.335 19.93 4.65 ;
      RECT 19.91 4.383 19.915 4.648 ;
      RECT 19.905 3.545 19.91 3.768 ;
      RECT 19.905 4.415 19.91 4.643 ;
      RECT 19.88 3.545 19.905 3.76 ;
      RECT 19.87 3.55 19.88 3.75 ;
      RECT 20.085 4.825 20.105 5.065 ;
      RECT 19.315 4.755 19.32 4.965 ;
      RECT 20.595 4.828 20.605 5.023 ;
      RECT 20.59 4.818 20.595 5.026 ;
      RECT 20.51 4.815 20.59 5.049 ;
      RECT 20.506 4.815 20.51 5.071 ;
      RECT 20.42 4.815 20.506 5.081 ;
      RECT 20.405 4.815 20.42 5.089 ;
      RECT 20.376 4.816 20.405 5.087 ;
      RECT 20.29 4.821 20.376 5.083 ;
      RECT 20.277 4.825 20.29 5.079 ;
      RECT 20.191 4.825 20.277 5.075 ;
      RECT 20.105 4.825 20.191 5.069 ;
      RECT 20.021 4.825 20.085 5.063 ;
      RECT 19.935 4.825 20.021 5.058 ;
      RECT 19.915 4.825 19.935 5.054 ;
      RECT 19.855 4.82 19.915 5.051 ;
      RECT 19.827 4.814 19.855 5.048 ;
      RECT 19.741 4.809 19.827 5.044 ;
      RECT 19.655 4.803 19.741 5.038 ;
      RECT 19.58 4.785 19.655 5.033 ;
      RECT 19.545 4.762 19.58 5.029 ;
      RECT 19.535 4.752 19.545 5.028 ;
      RECT 19.48 4.75 19.535 5.027 ;
      RECT 19.405 4.75 19.48 5.023 ;
      RECT 19.395 4.75 19.405 5.018 ;
      RECT 19.38 4.75 19.395 5.01 ;
      RECT 19.33 4.752 19.38 4.988 ;
      RECT 19.32 4.755 19.33 4.968 ;
      RECT 19.31 4.76 19.315 4.963 ;
      RECT 19.305 4.765 19.31 4.958 ;
      RECT 19.43 3.93 19.69 4.19 ;
      RECT 19.43 3.945 19.71 4.155 ;
      RECT 19.43 3.95 19.72 4.15 ;
      RECT 17.415 3.41 17.675 3.67 ;
      RECT 17.405 3.44 17.675 3.65 ;
      RECT 19.325 3.355 19.585 3.615 ;
      RECT 19.32 3.43 19.325 3.616 ;
      RECT 19.295 3.435 19.32 3.618 ;
      RECT 19.28 3.442 19.295 3.621 ;
      RECT 19.22 3.46 19.28 3.626 ;
      RECT 19.19 3.48 19.22 3.633 ;
      RECT 19.165 3.488 19.19 3.638 ;
      RECT 19.14 3.496 19.165 3.64 ;
      RECT 19.122 3.5 19.14 3.639 ;
      RECT 19.036 3.498 19.122 3.639 ;
      RECT 18.95 3.496 19.036 3.639 ;
      RECT 18.864 3.494 18.95 3.638 ;
      RECT 18.778 3.492 18.864 3.638 ;
      RECT 18.692 3.49 18.778 3.638 ;
      RECT 18.606 3.488 18.692 3.638 ;
      RECT 18.52 3.486 18.606 3.637 ;
      RECT 18.502 3.485 18.52 3.637 ;
      RECT 18.416 3.484 18.502 3.637 ;
      RECT 18.33 3.482 18.416 3.637 ;
      RECT 18.244 3.481 18.33 3.636 ;
      RECT 18.158 3.48 18.244 3.636 ;
      RECT 18.072 3.478 18.158 3.636 ;
      RECT 17.986 3.477 18.072 3.636 ;
      RECT 17.9 3.475 17.986 3.635 ;
      RECT 17.876 3.473 17.9 3.635 ;
      RECT 17.79 3.466 17.876 3.635 ;
      RECT 17.761 3.458 17.79 3.635 ;
      RECT 17.675 3.45 17.761 3.635 ;
      RECT 17.395 3.447 17.405 3.645 ;
      RECT 18.9 4.41 18.905 4.76 ;
      RECT 18.67 4.5 18.81 4.76 ;
      RECT 19.145 4.185 19.19 4.395 ;
      RECT 19.2 4.196 19.21 4.39 ;
      RECT 19.19 4.188 19.2 4.395 ;
      RECT 19.125 4.185 19.145 4.4 ;
      RECT 19.095 4.185 19.125 4.423 ;
      RECT 19.085 4.185 19.095 4.448 ;
      RECT 19.08 4.185 19.085 4.458 ;
      RECT 19.025 4.185 19.08 4.498 ;
      RECT 19.02 4.185 19.025 4.538 ;
      RECT 19.015 4.187 19.02 4.543 ;
      RECT 19 4.197 19.015 4.554 ;
      RECT 18.955 4.255 19 4.59 ;
      RECT 18.945 4.31 18.955 4.624 ;
      RECT 18.93 4.337 18.945 4.64 ;
      RECT 18.92 4.364 18.93 4.76 ;
      RECT 18.905 4.387 18.92 4.76 ;
      RECT 18.895 4.427 18.9 4.76 ;
      RECT 18.89 4.437 18.895 4.76 ;
      RECT 18.885 4.452 18.89 4.76 ;
      RECT 18.875 4.457 18.885 4.76 ;
      RECT 18.81 4.48 18.875 4.76 ;
      RECT 18.31 3.975 18.5 4.185 ;
      RECT 16.885 3.9 17.145 4.16 ;
      RECT 17.235 3.895 17.33 4.105 ;
      RECT 17.21 3.91 17.22 4.105 ;
      RECT 18.5 3.982 18.51 4.18 ;
      RECT 18.3 3.982 18.31 4.18 ;
      RECT 18.285 3.997 18.3 4.17 ;
      RECT 18.28 4.005 18.285 4.163 ;
      RECT 18.27 4.008 18.28 4.16 ;
      RECT 18.235 4.007 18.27 4.158 ;
      RECT 18.206 4.003 18.235 4.155 ;
      RECT 18.12 3.998 18.206 4.152 ;
      RECT 18.06 3.992 18.12 4.148 ;
      RECT 18.031 3.988 18.06 4.145 ;
      RECT 17.945 3.98 18.031 4.142 ;
      RECT 17.936 3.974 17.945 4.14 ;
      RECT 17.85 3.969 17.936 4.138 ;
      RECT 17.827 3.964 17.85 4.135 ;
      RECT 17.741 3.958 17.827 4.132 ;
      RECT 17.655 3.949 17.741 4.127 ;
      RECT 17.645 3.944 17.655 4.125 ;
      RECT 17.626 3.943 17.645 4.124 ;
      RECT 17.54 3.938 17.626 4.12 ;
      RECT 17.52 3.933 17.54 4.116 ;
      RECT 17.46 3.928 17.52 4.113 ;
      RECT 17.435 3.918 17.46 4.111 ;
      RECT 17.43 3.911 17.435 4.11 ;
      RECT 17.42 3.902 17.43 4.109 ;
      RECT 17.416 3.895 17.42 4.109 ;
      RECT 17.33 3.895 17.416 4.107 ;
      RECT 17.22 3.902 17.235 4.105 ;
      RECT 17.205 3.912 17.21 4.105 ;
      RECT 17.185 3.915 17.205 4.102 ;
      RECT 17.155 3.915 17.185 4.098 ;
      RECT 17.145 3.915 17.155 4.098 ;
      RECT 18.06 4.41 18.32 4.67 ;
      RECT 17.99 4.42 18.32 4.63 ;
      RECT 17.98 4.427 18.32 4.625 ;
      RECT 17.4 4.415 17.66 4.675 ;
      RECT 17.4 4.455 17.765 4.665 ;
      RECT 17.4 4.457 17.77 4.664 ;
      RECT 17.4 4.465 17.775 4.661 ;
      RECT 16.325 3.54 16.425 5.065 ;
      RECT 16.515 4.68 16.565 4.94 ;
      RECT 16.51 3.553 16.515 3.74 ;
      RECT 16.505 4.661 16.515 4.94 ;
      RECT 16.505 3.55 16.51 3.748 ;
      RECT 16.49 3.544 16.505 3.755 ;
      RECT 16.5 4.649 16.505 5.023 ;
      RECT 16.49 4.637 16.5 5.06 ;
      RECT 16.48 3.54 16.49 3.762 ;
      RECT 16.48 4.622 16.49 5.065 ;
      RECT 16.475 3.54 16.48 3.77 ;
      RECT 16.455 4.592 16.48 5.065 ;
      RECT 16.435 3.54 16.475 3.818 ;
      RECT 16.445 4.552 16.455 5.065 ;
      RECT 16.435 4.507 16.445 5.065 ;
      RECT 16.43 3.54 16.435 3.888 ;
      RECT 16.43 4.465 16.435 5.065 ;
      RECT 16.425 3.54 16.43 4.365 ;
      RECT 16.425 4.447 16.43 5.065 ;
      RECT 16.315 3.543 16.325 5.065 ;
      RECT 16.3 3.55 16.315 5.061 ;
      RECT 16.295 3.56 16.3 5.056 ;
      RECT 16.29 3.76 16.295 4.948 ;
      RECT 16.285 3.845 16.29 4.5 ;
      RECT 14.515 10.2 14.805 10.43 ;
      RECT 14.575 9.46 14.745 10.43 ;
      RECT 14.485 9.46 14.835 9.75 ;
      RECT 14.11 8.72 14.46 9.01 ;
      RECT 13.97 8.75 14.46 8.92 ;
      RECT 100.015 2.435 100.39 2.805 ;
      RECT 93.995 3.52 94.255 3.78 ;
      RECT 82.09 2.435 82.465 2.805 ;
      RECT 76.07 3.52 76.33 3.78 ;
      RECT 64.165 2.435 64.54 2.805 ;
      RECT 58.145 3.52 58.405 3.78 ;
      RECT 46.24 2.435 46.615 2.805 ;
      RECT 40.22 3.52 40.48 3.78 ;
      RECT 28.315 2.435 28.69 2.805 ;
      RECT 22.295 3.52 22.555 3.78 ;
    LAYER mcon ;
      RECT 104.845 8.755 105.015 8.925 ;
      RECT 104.845 10.235 105.015 10.405 ;
      RECT 104.495 1.395 104.665 1.565 ;
      RECT 104.475 4.055 104.645 4.225 ;
      RECT 104.475 8.385 104.645 8.555 ;
      RECT 103.855 2.205 104.025 2.375 ;
      RECT 103.855 3.685 104.025 3.855 ;
      RECT 103.855 8.755 104.025 8.925 ;
      RECT 103.855 10.235 104.025 10.405 ;
      RECT 103.505 1.395 103.675 1.565 ;
      RECT 103.485 4.055 103.655 4.225 ;
      RECT 103.485 8.385 103.655 8.555 ;
      RECT 102.805 1.4 102.975 1.57 ;
      RECT 102.495 3.32 102.665 3.49 ;
      RECT 102.495 9.12 102.665 9.29 ;
      RECT 102.125 1.4 102.295 1.57 ;
      RECT 102.065 2.21 102.235 2.38 ;
      RECT 102.065 2.95 102.235 3.12 ;
      RECT 102.065 9.49 102.235 9.66 ;
      RECT 102.065 10.23 102.235 10.4 ;
      RECT 101.69 3.69 101.86 3.86 ;
      RECT 101.69 8.75 101.86 8.92 ;
      RECT 101.445 1.4 101.615 1.57 ;
      RECT 100.765 1.4 100.935 1.57 ;
      RECT 99.485 2.86 99.655 3.03 ;
      RECT 99.025 2.86 99.195 3.03 ;
      RECT 98.63 4.2 98.8 4.37 ;
      RECT 98.565 2.86 98.735 3.03 ;
      RECT 98.42 3.54 98.59 3.71 ;
      RECT 98.105 2.86 98.275 3.03 ;
      RECT 98.105 4.45 98.275 4.62 ;
      RECT 97.735 9.12 97.905 9.29 ;
      RECT 97.72 4.045 97.89 4.215 ;
      RECT 97.645 2.86 97.815 3.03 ;
      RECT 97.505 4.61 97.675 4.78 ;
      RECT 97.485 5.01 97.655 5.18 ;
      RECT 97.31 3.565 97.48 3.735 ;
      RECT 97.305 9.49 97.475 9.66 ;
      RECT 97.305 10.23 97.475 10.4 ;
      RECT 97.185 2.86 97.355 3.03 ;
      RECT 96.815 4.545 96.985 4.715 ;
      RECT 96.725 2.86 96.895 3.03 ;
      RECT 96.49 4.23 96.66 4.4 ;
      RECT 96.425 5.01 96.595 5.18 ;
      RECT 96.265 2.86 96.435 3.03 ;
      RECT 96.025 4.995 96.195 5.165 ;
      RECT 95.985 3.48 96.155 3.65 ;
      RECT 95.805 2.86 95.975 3.03 ;
      RECT 95.345 2.86 95.515 3.03 ;
      RECT 95.085 3.98 95.255 4.15 ;
      RECT 95.085 4.44 95.255 4.61 ;
      RECT 95.085 4.955 95.255 5.125 ;
      RECT 94.97 3.515 95.14 3.685 ;
      RECT 94.885 2.86 95.055 3.03 ;
      RECT 94.505 5.025 94.675 5.195 ;
      RECT 94.425 2.86 94.595 3.03 ;
      RECT 94.025 3.555 94.195 3.725 ;
      RECT 93.965 2.86 94.135 3.03 ;
      RECT 93.81 3.93 93.98 4.1 ;
      RECT 93.505 2.86 93.675 3.03 ;
      RECT 93.31 4.53 93.48 4.7 ;
      RECT 93.195 3.98 93.365 4.15 ;
      RECT 93.045 2.86 93.215 3.03 ;
      RECT 93.025 3.43 93.195 3.6 ;
      RECT 92.65 4.46 92.82 4.63 ;
      RECT 92.585 2.86 92.755 3.03 ;
      RECT 92.165 4.06 92.335 4.23 ;
      RECT 92.125 2.86 92.295 3.03 ;
      RECT 92.115 4.835 92.285 5.005 ;
      RECT 91.665 2.86 91.835 3.03 ;
      RECT 91.625 4.46 91.795 4.63 ;
      RECT 91.59 3.565 91.76 3.735 ;
      RECT 91.23 3.965 91.4 4.135 ;
      RECT 91.205 2.86 91.375 3.03 ;
      RECT 91.025 4.775 91.195 4.945 ;
      RECT 90.745 2.86 90.915 3.03 ;
      RECT 90.72 4.205 90.89 4.375 ;
      RECT 90.285 2.86 90.455 3.03 ;
      RECT 90.02 3.995 90.19 4.165 ;
      RECT 89.825 2.86 89.995 3.03 ;
      RECT 89.7 4.44 89.87 4.61 ;
      RECT 89.365 2.86 89.535 3.03 ;
      RECT 89.285 4.475 89.455 4.645 ;
      RECT 89.115 3.46 89.285 3.63 ;
      RECT 88.94 3.915 89.11 4.085 ;
      RECT 88.905 2.86 89.075 3.03 ;
      RECT 88.445 2.86 88.615 3.03 ;
      RECT 88.02 3.565 88.19 3.735 ;
      RECT 88.015 4.88 88.185 5.05 ;
      RECT 87.985 2.86 88.155 3.03 ;
      RECT 86.92 8.755 87.09 8.925 ;
      RECT 86.92 10.235 87.09 10.405 ;
      RECT 86.57 1.395 86.74 1.565 ;
      RECT 86.55 4.055 86.72 4.225 ;
      RECT 86.55 8.385 86.72 8.555 ;
      RECT 85.93 2.205 86.1 2.375 ;
      RECT 85.93 3.685 86.1 3.855 ;
      RECT 85.93 8.755 86.1 8.925 ;
      RECT 85.93 10.235 86.1 10.405 ;
      RECT 85.58 1.395 85.75 1.565 ;
      RECT 85.56 4.055 85.73 4.225 ;
      RECT 85.56 8.385 85.73 8.555 ;
      RECT 84.88 1.4 85.05 1.57 ;
      RECT 84.57 3.32 84.74 3.49 ;
      RECT 84.57 9.12 84.74 9.29 ;
      RECT 84.2 1.4 84.37 1.57 ;
      RECT 84.14 2.21 84.31 2.38 ;
      RECT 84.14 2.95 84.31 3.12 ;
      RECT 84.14 9.49 84.31 9.66 ;
      RECT 84.14 10.23 84.31 10.4 ;
      RECT 83.765 3.69 83.935 3.86 ;
      RECT 83.765 8.75 83.935 8.92 ;
      RECT 83.52 1.4 83.69 1.57 ;
      RECT 82.84 1.4 83.01 1.57 ;
      RECT 81.56 2.86 81.73 3.03 ;
      RECT 81.1 2.86 81.27 3.03 ;
      RECT 80.705 4.2 80.875 4.37 ;
      RECT 80.64 2.86 80.81 3.03 ;
      RECT 80.495 3.54 80.665 3.71 ;
      RECT 80.18 2.86 80.35 3.03 ;
      RECT 80.18 4.45 80.35 4.62 ;
      RECT 79.81 9.12 79.98 9.29 ;
      RECT 79.795 4.045 79.965 4.215 ;
      RECT 79.72 2.86 79.89 3.03 ;
      RECT 79.58 4.61 79.75 4.78 ;
      RECT 79.56 5.01 79.73 5.18 ;
      RECT 79.385 3.565 79.555 3.735 ;
      RECT 79.38 9.49 79.55 9.66 ;
      RECT 79.38 10.23 79.55 10.4 ;
      RECT 79.26 2.86 79.43 3.03 ;
      RECT 78.89 4.545 79.06 4.715 ;
      RECT 78.8 2.86 78.97 3.03 ;
      RECT 78.565 4.23 78.735 4.4 ;
      RECT 78.5 5.01 78.67 5.18 ;
      RECT 78.34 2.86 78.51 3.03 ;
      RECT 78.1 4.995 78.27 5.165 ;
      RECT 78.06 3.48 78.23 3.65 ;
      RECT 77.88 2.86 78.05 3.03 ;
      RECT 77.42 2.86 77.59 3.03 ;
      RECT 77.16 3.98 77.33 4.15 ;
      RECT 77.16 4.44 77.33 4.61 ;
      RECT 77.16 4.955 77.33 5.125 ;
      RECT 77.045 3.515 77.215 3.685 ;
      RECT 76.96 2.86 77.13 3.03 ;
      RECT 76.58 5.025 76.75 5.195 ;
      RECT 76.5 2.86 76.67 3.03 ;
      RECT 76.1 3.555 76.27 3.725 ;
      RECT 76.04 2.86 76.21 3.03 ;
      RECT 75.885 3.93 76.055 4.1 ;
      RECT 75.58 2.86 75.75 3.03 ;
      RECT 75.385 4.53 75.555 4.7 ;
      RECT 75.27 3.98 75.44 4.15 ;
      RECT 75.12 2.86 75.29 3.03 ;
      RECT 75.1 3.43 75.27 3.6 ;
      RECT 74.725 4.46 74.895 4.63 ;
      RECT 74.66 2.86 74.83 3.03 ;
      RECT 74.24 4.06 74.41 4.23 ;
      RECT 74.2 2.86 74.37 3.03 ;
      RECT 74.19 4.835 74.36 5.005 ;
      RECT 73.74 2.86 73.91 3.03 ;
      RECT 73.7 4.46 73.87 4.63 ;
      RECT 73.665 3.565 73.835 3.735 ;
      RECT 73.305 3.965 73.475 4.135 ;
      RECT 73.28 2.86 73.45 3.03 ;
      RECT 73.1 4.775 73.27 4.945 ;
      RECT 72.82 2.86 72.99 3.03 ;
      RECT 72.795 4.205 72.965 4.375 ;
      RECT 72.36 2.86 72.53 3.03 ;
      RECT 72.095 3.995 72.265 4.165 ;
      RECT 71.9 2.86 72.07 3.03 ;
      RECT 71.775 4.44 71.945 4.61 ;
      RECT 71.44 2.86 71.61 3.03 ;
      RECT 71.36 4.475 71.53 4.645 ;
      RECT 71.19 3.46 71.36 3.63 ;
      RECT 71.015 3.915 71.185 4.085 ;
      RECT 70.98 2.86 71.15 3.03 ;
      RECT 70.52 2.86 70.69 3.03 ;
      RECT 70.095 3.565 70.265 3.735 ;
      RECT 70.09 4.88 70.26 5.05 ;
      RECT 70.06 2.86 70.23 3.03 ;
      RECT 68.995 8.755 69.165 8.925 ;
      RECT 68.995 10.235 69.165 10.405 ;
      RECT 68.645 1.395 68.815 1.565 ;
      RECT 68.625 4.055 68.795 4.225 ;
      RECT 68.625 8.385 68.795 8.555 ;
      RECT 68.005 2.205 68.175 2.375 ;
      RECT 68.005 3.685 68.175 3.855 ;
      RECT 68.005 8.755 68.175 8.925 ;
      RECT 68.005 10.235 68.175 10.405 ;
      RECT 67.655 1.395 67.825 1.565 ;
      RECT 67.635 4.055 67.805 4.225 ;
      RECT 67.635 8.385 67.805 8.555 ;
      RECT 66.955 1.4 67.125 1.57 ;
      RECT 66.645 3.32 66.815 3.49 ;
      RECT 66.645 9.12 66.815 9.29 ;
      RECT 66.275 1.4 66.445 1.57 ;
      RECT 66.215 2.21 66.385 2.38 ;
      RECT 66.215 2.95 66.385 3.12 ;
      RECT 66.215 9.49 66.385 9.66 ;
      RECT 66.215 10.23 66.385 10.4 ;
      RECT 65.84 3.69 66.01 3.86 ;
      RECT 65.84 8.75 66.01 8.92 ;
      RECT 65.595 1.4 65.765 1.57 ;
      RECT 64.915 1.4 65.085 1.57 ;
      RECT 63.635 2.86 63.805 3.03 ;
      RECT 63.175 2.86 63.345 3.03 ;
      RECT 62.78 4.2 62.95 4.37 ;
      RECT 62.715 2.86 62.885 3.03 ;
      RECT 62.57 3.54 62.74 3.71 ;
      RECT 62.255 2.86 62.425 3.03 ;
      RECT 62.255 4.45 62.425 4.62 ;
      RECT 61.885 9.12 62.055 9.29 ;
      RECT 61.87 4.045 62.04 4.215 ;
      RECT 61.795 2.86 61.965 3.03 ;
      RECT 61.655 4.61 61.825 4.78 ;
      RECT 61.635 5.01 61.805 5.18 ;
      RECT 61.46 3.565 61.63 3.735 ;
      RECT 61.455 9.49 61.625 9.66 ;
      RECT 61.455 10.23 61.625 10.4 ;
      RECT 61.335 2.86 61.505 3.03 ;
      RECT 60.965 4.545 61.135 4.715 ;
      RECT 60.875 2.86 61.045 3.03 ;
      RECT 60.64 4.23 60.81 4.4 ;
      RECT 60.575 5.01 60.745 5.18 ;
      RECT 60.415 2.86 60.585 3.03 ;
      RECT 60.175 4.995 60.345 5.165 ;
      RECT 60.135 3.48 60.305 3.65 ;
      RECT 59.955 2.86 60.125 3.03 ;
      RECT 59.495 2.86 59.665 3.03 ;
      RECT 59.235 3.98 59.405 4.15 ;
      RECT 59.235 4.44 59.405 4.61 ;
      RECT 59.235 4.955 59.405 5.125 ;
      RECT 59.12 3.515 59.29 3.685 ;
      RECT 59.035 2.86 59.205 3.03 ;
      RECT 58.655 5.025 58.825 5.195 ;
      RECT 58.575 2.86 58.745 3.03 ;
      RECT 58.175 3.555 58.345 3.725 ;
      RECT 58.115 2.86 58.285 3.03 ;
      RECT 57.96 3.93 58.13 4.1 ;
      RECT 57.655 2.86 57.825 3.03 ;
      RECT 57.46 4.53 57.63 4.7 ;
      RECT 57.345 3.98 57.515 4.15 ;
      RECT 57.195 2.86 57.365 3.03 ;
      RECT 57.175 3.43 57.345 3.6 ;
      RECT 56.8 4.46 56.97 4.63 ;
      RECT 56.735 2.86 56.905 3.03 ;
      RECT 56.315 4.06 56.485 4.23 ;
      RECT 56.275 2.86 56.445 3.03 ;
      RECT 56.265 4.835 56.435 5.005 ;
      RECT 55.815 2.86 55.985 3.03 ;
      RECT 55.775 4.46 55.945 4.63 ;
      RECT 55.74 3.565 55.91 3.735 ;
      RECT 55.38 3.965 55.55 4.135 ;
      RECT 55.355 2.86 55.525 3.03 ;
      RECT 55.175 4.775 55.345 4.945 ;
      RECT 54.895 2.86 55.065 3.03 ;
      RECT 54.87 4.205 55.04 4.375 ;
      RECT 54.435 2.86 54.605 3.03 ;
      RECT 54.17 3.995 54.34 4.165 ;
      RECT 53.975 2.86 54.145 3.03 ;
      RECT 53.85 4.44 54.02 4.61 ;
      RECT 53.515 2.86 53.685 3.03 ;
      RECT 53.435 4.475 53.605 4.645 ;
      RECT 53.265 3.46 53.435 3.63 ;
      RECT 53.09 3.915 53.26 4.085 ;
      RECT 53.055 2.86 53.225 3.03 ;
      RECT 52.595 2.86 52.765 3.03 ;
      RECT 52.17 3.565 52.34 3.735 ;
      RECT 52.165 4.88 52.335 5.05 ;
      RECT 52.135 2.86 52.305 3.03 ;
      RECT 51.07 8.755 51.24 8.925 ;
      RECT 51.07 10.235 51.24 10.405 ;
      RECT 50.72 1.395 50.89 1.565 ;
      RECT 50.7 4.055 50.87 4.225 ;
      RECT 50.7 8.385 50.87 8.555 ;
      RECT 50.08 2.205 50.25 2.375 ;
      RECT 50.08 3.685 50.25 3.855 ;
      RECT 50.08 8.755 50.25 8.925 ;
      RECT 50.08 10.235 50.25 10.405 ;
      RECT 49.73 1.395 49.9 1.565 ;
      RECT 49.71 4.055 49.88 4.225 ;
      RECT 49.71 8.385 49.88 8.555 ;
      RECT 49.03 1.4 49.2 1.57 ;
      RECT 48.72 3.32 48.89 3.49 ;
      RECT 48.72 9.12 48.89 9.29 ;
      RECT 48.35 1.4 48.52 1.57 ;
      RECT 48.29 2.21 48.46 2.38 ;
      RECT 48.29 2.95 48.46 3.12 ;
      RECT 48.29 9.49 48.46 9.66 ;
      RECT 48.29 10.23 48.46 10.4 ;
      RECT 47.915 3.69 48.085 3.86 ;
      RECT 47.915 8.75 48.085 8.92 ;
      RECT 47.67 1.4 47.84 1.57 ;
      RECT 46.99 1.4 47.16 1.57 ;
      RECT 45.71 2.86 45.88 3.03 ;
      RECT 45.25 2.86 45.42 3.03 ;
      RECT 44.855 4.2 45.025 4.37 ;
      RECT 44.79 2.86 44.96 3.03 ;
      RECT 44.645 3.54 44.815 3.71 ;
      RECT 44.33 2.86 44.5 3.03 ;
      RECT 44.33 4.45 44.5 4.62 ;
      RECT 43.96 9.12 44.13 9.29 ;
      RECT 43.945 4.045 44.115 4.215 ;
      RECT 43.87 2.86 44.04 3.03 ;
      RECT 43.73 4.61 43.9 4.78 ;
      RECT 43.71 5.01 43.88 5.18 ;
      RECT 43.535 3.565 43.705 3.735 ;
      RECT 43.53 9.49 43.7 9.66 ;
      RECT 43.53 10.23 43.7 10.4 ;
      RECT 43.41 2.86 43.58 3.03 ;
      RECT 43.04 4.545 43.21 4.715 ;
      RECT 42.95 2.86 43.12 3.03 ;
      RECT 42.715 4.23 42.885 4.4 ;
      RECT 42.65 5.01 42.82 5.18 ;
      RECT 42.49 2.86 42.66 3.03 ;
      RECT 42.25 4.995 42.42 5.165 ;
      RECT 42.21 3.48 42.38 3.65 ;
      RECT 42.03 2.86 42.2 3.03 ;
      RECT 41.57 2.86 41.74 3.03 ;
      RECT 41.31 3.98 41.48 4.15 ;
      RECT 41.31 4.44 41.48 4.61 ;
      RECT 41.31 4.955 41.48 5.125 ;
      RECT 41.195 3.515 41.365 3.685 ;
      RECT 41.11 2.86 41.28 3.03 ;
      RECT 40.73 5.025 40.9 5.195 ;
      RECT 40.65 2.86 40.82 3.03 ;
      RECT 40.25 3.555 40.42 3.725 ;
      RECT 40.19 2.86 40.36 3.03 ;
      RECT 40.035 3.93 40.205 4.1 ;
      RECT 39.73 2.86 39.9 3.03 ;
      RECT 39.535 4.53 39.705 4.7 ;
      RECT 39.42 3.98 39.59 4.15 ;
      RECT 39.27 2.86 39.44 3.03 ;
      RECT 39.25 3.43 39.42 3.6 ;
      RECT 38.875 4.46 39.045 4.63 ;
      RECT 38.81 2.86 38.98 3.03 ;
      RECT 38.39 4.06 38.56 4.23 ;
      RECT 38.35 2.86 38.52 3.03 ;
      RECT 38.34 4.835 38.51 5.005 ;
      RECT 37.89 2.86 38.06 3.03 ;
      RECT 37.85 4.46 38.02 4.63 ;
      RECT 37.815 3.565 37.985 3.735 ;
      RECT 37.455 3.965 37.625 4.135 ;
      RECT 37.43 2.86 37.6 3.03 ;
      RECT 37.25 4.775 37.42 4.945 ;
      RECT 36.97 2.86 37.14 3.03 ;
      RECT 36.945 4.205 37.115 4.375 ;
      RECT 36.51 2.86 36.68 3.03 ;
      RECT 36.245 3.995 36.415 4.165 ;
      RECT 36.05 2.86 36.22 3.03 ;
      RECT 35.925 4.44 36.095 4.61 ;
      RECT 35.59 2.86 35.76 3.03 ;
      RECT 35.51 4.475 35.68 4.645 ;
      RECT 35.34 3.46 35.51 3.63 ;
      RECT 35.165 3.915 35.335 4.085 ;
      RECT 35.13 2.86 35.3 3.03 ;
      RECT 34.67 2.86 34.84 3.03 ;
      RECT 34.245 3.565 34.415 3.735 ;
      RECT 34.24 4.88 34.41 5.05 ;
      RECT 34.21 2.86 34.38 3.03 ;
      RECT 33.145 8.755 33.315 8.925 ;
      RECT 33.145 10.235 33.315 10.405 ;
      RECT 32.795 1.395 32.965 1.565 ;
      RECT 32.775 4.055 32.945 4.225 ;
      RECT 32.775 8.385 32.945 8.555 ;
      RECT 32.155 2.205 32.325 2.375 ;
      RECT 32.155 3.685 32.325 3.855 ;
      RECT 32.155 8.755 32.325 8.925 ;
      RECT 32.155 10.235 32.325 10.405 ;
      RECT 31.805 1.395 31.975 1.565 ;
      RECT 31.785 4.055 31.955 4.225 ;
      RECT 31.785 8.385 31.955 8.555 ;
      RECT 31.105 1.4 31.275 1.57 ;
      RECT 30.795 3.32 30.965 3.49 ;
      RECT 30.795 9.12 30.965 9.29 ;
      RECT 30.425 1.4 30.595 1.57 ;
      RECT 30.365 2.21 30.535 2.38 ;
      RECT 30.365 2.95 30.535 3.12 ;
      RECT 30.365 9.49 30.535 9.66 ;
      RECT 30.365 10.23 30.535 10.4 ;
      RECT 29.99 3.69 30.16 3.86 ;
      RECT 29.99 8.75 30.16 8.92 ;
      RECT 29.745 1.4 29.915 1.57 ;
      RECT 29.065 1.4 29.235 1.57 ;
      RECT 27.785 2.86 27.955 3.03 ;
      RECT 27.325 2.86 27.495 3.03 ;
      RECT 26.93 4.2 27.1 4.37 ;
      RECT 26.865 2.86 27.035 3.03 ;
      RECT 26.72 3.54 26.89 3.71 ;
      RECT 26.405 2.86 26.575 3.03 ;
      RECT 26.405 4.45 26.575 4.62 ;
      RECT 26.035 9.12 26.205 9.29 ;
      RECT 26.02 4.045 26.19 4.215 ;
      RECT 25.945 2.86 26.115 3.03 ;
      RECT 25.805 4.61 25.975 4.78 ;
      RECT 25.785 5.01 25.955 5.18 ;
      RECT 25.61 3.565 25.78 3.735 ;
      RECT 25.605 9.49 25.775 9.66 ;
      RECT 25.605 10.23 25.775 10.4 ;
      RECT 25.485 2.86 25.655 3.03 ;
      RECT 25.115 4.545 25.285 4.715 ;
      RECT 25.025 2.86 25.195 3.03 ;
      RECT 24.79 4.23 24.96 4.4 ;
      RECT 24.725 5.01 24.895 5.18 ;
      RECT 24.565 2.86 24.735 3.03 ;
      RECT 24.325 4.995 24.495 5.165 ;
      RECT 24.285 3.48 24.455 3.65 ;
      RECT 24.105 2.86 24.275 3.03 ;
      RECT 23.645 2.86 23.815 3.03 ;
      RECT 23.385 3.98 23.555 4.15 ;
      RECT 23.385 4.44 23.555 4.61 ;
      RECT 23.385 4.955 23.555 5.125 ;
      RECT 23.27 3.515 23.44 3.685 ;
      RECT 23.185 2.86 23.355 3.03 ;
      RECT 22.805 5.025 22.975 5.195 ;
      RECT 22.725 2.86 22.895 3.03 ;
      RECT 22.325 3.555 22.495 3.725 ;
      RECT 22.265 2.86 22.435 3.03 ;
      RECT 22.11 3.93 22.28 4.1 ;
      RECT 21.805 2.86 21.975 3.03 ;
      RECT 21.61 4.53 21.78 4.7 ;
      RECT 21.495 3.98 21.665 4.15 ;
      RECT 21.345 2.86 21.515 3.03 ;
      RECT 21.325 3.43 21.495 3.6 ;
      RECT 20.95 4.46 21.12 4.63 ;
      RECT 20.885 2.86 21.055 3.03 ;
      RECT 20.465 4.06 20.635 4.23 ;
      RECT 20.425 2.86 20.595 3.03 ;
      RECT 20.415 4.835 20.585 5.005 ;
      RECT 19.965 2.86 20.135 3.03 ;
      RECT 19.925 4.46 20.095 4.63 ;
      RECT 19.89 3.565 20.06 3.735 ;
      RECT 19.53 3.965 19.7 4.135 ;
      RECT 19.505 2.86 19.675 3.03 ;
      RECT 19.325 4.775 19.495 4.945 ;
      RECT 19.045 2.86 19.215 3.03 ;
      RECT 19.02 4.205 19.19 4.375 ;
      RECT 18.585 2.86 18.755 3.03 ;
      RECT 18.32 3.995 18.49 4.165 ;
      RECT 18.125 2.86 18.295 3.03 ;
      RECT 18 4.44 18.17 4.61 ;
      RECT 17.665 2.86 17.835 3.03 ;
      RECT 17.585 4.475 17.755 4.645 ;
      RECT 17.415 3.46 17.585 3.63 ;
      RECT 17.24 3.915 17.41 4.085 ;
      RECT 17.205 2.86 17.375 3.03 ;
      RECT 16.745 2.86 16.915 3.03 ;
      RECT 16.32 3.565 16.49 3.735 ;
      RECT 16.315 4.88 16.485 5.05 ;
      RECT 16.285 2.86 16.455 3.03 ;
      RECT 14.575 9.49 14.745 9.66 ;
      RECT 14.575 10.23 14.745 10.4 ;
      RECT 14.2 8.75 14.37 8.92 ;
    LAYER li1 ;
      RECT 98.89 0 99.06 3.53 ;
      RECT 97.93 0 98.1 3.53 ;
      RECT 96.97 0 97.14 3.53 ;
      RECT 96.45 0 96.62 3.53 ;
      RECT 95.49 0 95.66 3.53 ;
      RECT 94.49 0 94.66 3.53 ;
      RECT 93.53 0 93.7 3.53 ;
      RECT 92.05 0 92.22 3.53 ;
      RECT 90.13 0 90.3 3.53 ;
      RECT 88.65 0 88.82 3.53 ;
      RECT 80.965 0 81.135 3.53 ;
      RECT 80.005 0 80.175 3.53 ;
      RECT 79.045 0 79.215 3.53 ;
      RECT 78.525 0 78.695 3.53 ;
      RECT 77.565 0 77.735 3.53 ;
      RECT 76.565 0 76.735 3.53 ;
      RECT 75.605 0 75.775 3.53 ;
      RECT 74.125 0 74.295 3.53 ;
      RECT 72.205 0 72.375 3.53 ;
      RECT 70.725 0 70.895 3.53 ;
      RECT 63.04 0 63.21 3.53 ;
      RECT 62.08 0 62.25 3.53 ;
      RECT 61.12 0 61.29 3.53 ;
      RECT 60.6 0 60.77 3.53 ;
      RECT 59.64 0 59.81 3.53 ;
      RECT 58.64 0 58.81 3.53 ;
      RECT 57.68 0 57.85 3.53 ;
      RECT 56.2 0 56.37 3.53 ;
      RECT 54.28 0 54.45 3.53 ;
      RECT 52.8 0 52.97 3.53 ;
      RECT 45.115 0 45.285 3.53 ;
      RECT 44.155 0 44.325 3.53 ;
      RECT 43.195 0 43.365 3.53 ;
      RECT 42.675 0 42.845 3.53 ;
      RECT 41.715 0 41.885 3.53 ;
      RECT 40.715 0 40.885 3.53 ;
      RECT 39.755 0 39.925 3.53 ;
      RECT 38.275 0 38.445 3.53 ;
      RECT 36.355 0 36.525 3.53 ;
      RECT 34.875 0 35.045 3.53 ;
      RECT 27.19 0 27.36 3.53 ;
      RECT 26.23 0 26.4 3.53 ;
      RECT 25.27 0 25.44 3.53 ;
      RECT 24.75 0 24.92 3.53 ;
      RECT 23.79 0 23.96 3.53 ;
      RECT 22.79 0 22.96 3.53 ;
      RECT 21.83 0 22 3.53 ;
      RECT 20.35 0 20.52 3.53 ;
      RECT 18.43 0 18.6 3.53 ;
      RECT 16.95 0 17.12 3.53 ;
      RECT 87.84 0 99.8 3.03 ;
      RECT 69.915 0 81.875 3.03 ;
      RECT 51.99 0 63.95 3.03 ;
      RECT 34.065 0 46.025 3.03 ;
      RECT 16.14 0 28.1 3.03 ;
      RECT 87.835 0 99.8 2.975 ;
      RECT 69.91 0 81.875 2.975 ;
      RECT 51.985 0 63.95 2.975 ;
      RECT 34.06 0 46.025 2.975 ;
      RECT 16.135 0 28.1 2.975 ;
      RECT 100.685 0 100.855 2.23 ;
      RECT 82.76 0 82.93 2.23 ;
      RECT 64.835 0 65.005 2.23 ;
      RECT 46.91 0 47.08 2.23 ;
      RECT 28.985 0 29.155 2.23 ;
      RECT 104.415 0 104.585 2.225 ;
      RECT 103.425 0 103.595 2.225 ;
      RECT 86.49 0 86.66 2.225 ;
      RECT 85.5 0 85.67 2.225 ;
      RECT 68.565 0 68.735 2.225 ;
      RECT 67.575 0 67.745 2.225 ;
      RECT 50.64 0 50.81 2.225 ;
      RECT 49.65 0 49.82 2.225 ;
      RECT 32.715 0 32.885 2.225 ;
      RECT 31.725 0 31.895 2.225 ;
      RECT 12.97 0 105.39 1.6 ;
      RECT 104.475 3.035 104.645 4.225 ;
      RECT 104.475 3.035 104.945 3.205 ;
      RECT 104.475 9.405 104.945 9.575 ;
      RECT 104.475 8.385 104.645 9.575 ;
      RECT 103.485 3.035 103.655 4.225 ;
      RECT 103.485 3.035 103.955 3.205 ;
      RECT 103.485 9.405 103.955 9.575 ;
      RECT 103.485 8.385 103.655 9.575 ;
      RECT 101.635 3.93 101.805 5.16 ;
      RECT 101.69 2.15 101.86 4.1 ;
      RECT 101.635 1.87 101.805 2.32 ;
      RECT 101.635 10.29 101.805 10.74 ;
      RECT 101.69 8.51 101.86 10.46 ;
      RECT 101.635 7.45 101.805 8.68 ;
      RECT 101.115 1.87 101.285 5.16 ;
      RECT 101.115 3.37 101.52 3.7 ;
      RECT 101.115 2.53 101.52 2.86 ;
      RECT 101.115 7.45 101.285 10.74 ;
      RECT 101.115 9.75 101.52 10.08 ;
      RECT 101.115 8.91 101.52 9.24 ;
      RECT 99.215 4.687 99.23 4.738 ;
      RECT 99.21 4.667 99.215 4.785 ;
      RECT 99.195 4.657 99.21 4.853 ;
      RECT 99.17 4.637 99.195 4.908 ;
      RECT 99.13 4.622 99.17 4.928 ;
      RECT 99.085 4.616 99.13 4.956 ;
      RECT 99.015 4.606 99.085 4.973 ;
      RECT 98.995 4.598 99.015 4.973 ;
      RECT 98.935 4.592 98.995 4.965 ;
      RECT 98.876 4.583 98.935 4.953 ;
      RECT 98.79 4.572 98.876 4.936 ;
      RECT 98.768 4.563 98.79 4.924 ;
      RECT 98.682 4.556 98.768 4.911 ;
      RECT 98.596 4.543 98.682 4.892 ;
      RECT 98.51 4.531 98.596 4.872 ;
      RECT 98.48 4.52 98.51 4.859 ;
      RECT 98.43 4.506 98.48 4.851 ;
      RECT 98.41 4.495 98.43 4.843 ;
      RECT 98.361 4.484 98.41 4.835 ;
      RECT 98.275 4.463 98.361 4.82 ;
      RECT 98.23 4.45 98.275 4.805 ;
      RECT 98.185 4.45 98.23 4.785 ;
      RECT 98.13 4.45 98.185 4.72 ;
      RECT 98.105 4.45 98.13 4.643 ;
      RECT 98.63 4.187 98.8 4.37 ;
      RECT 98.63 4.187 98.815 4.328 ;
      RECT 98.63 4.187 98.82 4.27 ;
      RECT 98.69 3.955 98.825 4.246 ;
      RECT 98.69 3.959 98.83 4.229 ;
      RECT 98.635 4.122 98.83 4.229 ;
      RECT 98.66 3.967 98.8 4.37 ;
      RECT 98.66 3.971 98.84 4.17 ;
      RECT 98.645 4.057 98.84 4.17 ;
      RECT 98.655 3.987 98.8 4.37 ;
      RECT 98.655 3.99 98.85 4.083 ;
      RECT 98.65 4.007 98.85 4.083 ;
      RECT 98.42 3.227 98.59 3.71 ;
      RECT 98.415 3.222 98.565 3.7 ;
      RECT 98.415 3.229 98.595 3.694 ;
      RECT 98.405 3.223 98.565 3.673 ;
      RECT 98.405 3.239 98.61 3.632 ;
      RECT 98.375 3.224 98.565 3.595 ;
      RECT 98.375 3.254 98.62 3.535 ;
      RECT 98.37 3.226 98.565 3.533 ;
      RECT 98.35 3.235 98.595 3.49 ;
      RECT 98.325 3.251 98.61 3.402 ;
      RECT 98.325 3.27 98.635 3.393 ;
      RECT 98.32 3.307 98.635 3.345 ;
      RECT 98.325 3.287 98.64 3.313 ;
      RECT 98.42 3.221 98.53 3.71 ;
      RECT 98.506 3.22 98.53 3.71 ;
      RECT 97.74 4.005 97.745 4.216 ;
      RECT 98.34 4.005 98.345 4.19 ;
      RECT 98.405 4.045 98.41 4.158 ;
      RECT 98.4 4.037 98.405 4.164 ;
      RECT 98.395 4.027 98.4 4.172 ;
      RECT 98.39 4.017 98.395 4.181 ;
      RECT 98.385 4.007 98.39 4.185 ;
      RECT 98.345 4.005 98.385 4.188 ;
      RECT 98.317 4.004 98.34 4.192 ;
      RECT 98.231 4.001 98.317 4.199 ;
      RECT 98.145 3.997 98.231 4.21 ;
      RECT 98.125 3.995 98.145 4.216 ;
      RECT 98.107 3.994 98.125 4.219 ;
      RECT 98.021 3.992 98.107 4.226 ;
      RECT 97.935 3.987 98.021 4.239 ;
      RECT 97.916 3.984 97.935 4.244 ;
      RECT 97.83 3.982 97.916 4.235 ;
      RECT 97.82 3.982 97.83 4.228 ;
      RECT 97.745 3.995 97.82 4.222 ;
      RECT 97.73 4.006 97.74 4.216 ;
      RECT 97.72 4.008 97.73 4.215 ;
      RECT 97.71 4.012 97.72 4.211 ;
      RECT 97.705 4.015 97.71 4.205 ;
      RECT 97.695 4.017 97.705 4.199 ;
      RECT 97.69 4.02 97.695 4.193 ;
      RECT 97.67 4.606 97.675 4.81 ;
      RECT 97.655 4.593 97.67 4.903 ;
      RECT 97.64 4.574 97.655 5.18 ;
      RECT 97.605 4.54 97.64 5.18 ;
      RECT 97.601 4.51 97.605 5.18 ;
      RECT 97.515 4.392 97.601 5.18 ;
      RECT 97.505 4.267 97.515 5.18 ;
      RECT 97.49 4.235 97.505 5.18 ;
      RECT 97.485 4.21 97.49 5.18 ;
      RECT 97.48 4.2 97.485 5.136 ;
      RECT 97.465 4.172 97.48 5.041 ;
      RECT 97.45 4.138 97.465 4.94 ;
      RECT 97.445 4.116 97.45 4.893 ;
      RECT 97.44 4.105 97.445 4.863 ;
      RECT 97.435 4.095 97.44 4.829 ;
      RECT 97.425 4.082 97.435 4.797 ;
      RECT 97.4 4.058 97.425 4.723 ;
      RECT 97.395 4.038 97.4 4.648 ;
      RECT 97.39 4.032 97.395 4.623 ;
      RECT 97.385 4.027 97.39 4.588 ;
      RECT 97.38 4.022 97.385 4.563 ;
      RECT 97.375 4.02 97.38 4.543 ;
      RECT 97.37 4.02 97.375 4.528 ;
      RECT 97.365 4.02 97.37 4.488 ;
      RECT 97.355 4.02 97.365 4.46 ;
      RECT 97.345 4.02 97.355 4.405 ;
      RECT 97.33 4.02 97.345 4.343 ;
      RECT 97.325 4.019 97.33 4.288 ;
      RECT 97.31 4.018 97.325 4.268 ;
      RECT 97.25 4.016 97.31 4.242 ;
      RECT 97.215 4.017 97.25 4.222 ;
      RECT 97.21 4.019 97.215 4.212 ;
      RECT 97.2 4.038 97.21 4.202 ;
      RECT 97.195 4.065 97.2 4.133 ;
      RECT 97.31 3.49 97.48 3.735 ;
      RECT 97.345 3.261 97.48 3.735 ;
      RECT 97.345 3.263 97.49 3.73 ;
      RECT 97.345 3.265 97.515 3.718 ;
      RECT 97.345 3.268 97.54 3.7 ;
      RECT 97.345 3.273 97.59 3.673 ;
      RECT 97.345 3.278 97.61 3.638 ;
      RECT 97.325 3.28 97.62 3.613 ;
      RECT 97.315 3.375 97.62 3.613 ;
      RECT 97.345 3.26 97.455 3.735 ;
      RECT 97.355 3.257 97.45 3.735 ;
      RECT 96.875 4.522 97.065 4.88 ;
      RECT 96.875 4.534 97.1 4.879 ;
      RECT 96.875 4.562 97.12 4.877 ;
      RECT 96.875 4.587 97.125 4.876 ;
      RECT 96.875 4.645 97.14 4.875 ;
      RECT 96.86 4.518 97.02 4.86 ;
      RECT 96.84 4.527 97.065 4.813 ;
      RECT 96.815 4.538 97.1 4.75 ;
      RECT 96.815 4.622 97.135 4.75 ;
      RECT 96.815 4.597 97.13 4.75 ;
      RECT 96.875 4.513 97.02 4.88 ;
      RECT 96.961 4.512 97.02 4.88 ;
      RECT 96.961 4.511 97.005 4.88 ;
      RECT 96.355 7.45 96.525 10.74 ;
      RECT 96.355 9.75 96.76 10.08 ;
      RECT 96.355 8.91 96.76 9.24 ;
      RECT 96.66 4.027 96.665 4.405 ;
      RECT 96.655 3.995 96.66 4.405 ;
      RECT 96.65 3.967 96.655 4.405 ;
      RECT 96.645 3.947 96.65 4.405 ;
      RECT 96.59 3.93 96.645 4.405 ;
      RECT 96.55 3.915 96.59 4.405 ;
      RECT 96.495 3.902 96.55 4.405 ;
      RECT 96.46 3.893 96.495 4.405 ;
      RECT 96.456 3.891 96.46 4.404 ;
      RECT 96.37 3.887 96.456 4.387 ;
      RECT 96.285 3.879 96.37 4.35 ;
      RECT 96.275 3.875 96.285 4.323 ;
      RECT 96.265 3.875 96.275 4.305 ;
      RECT 96.255 3.877 96.265 4.288 ;
      RECT 96.25 3.882 96.255 4.274 ;
      RECT 96.245 3.886 96.25 4.261 ;
      RECT 96.235 3.891 96.245 4.245 ;
      RECT 96.22 3.905 96.235 4.22 ;
      RECT 96.215 3.911 96.22 4.2 ;
      RECT 96.21 3.913 96.215 4.193 ;
      RECT 96.205 3.917 96.21 4.068 ;
      RECT 96.385 4.717 96.63 5.18 ;
      RECT 96.305 4.69 96.625 5.176 ;
      RECT 96.235 4.725 96.63 5.169 ;
      RECT 96.025 4.98 96.63 5.165 ;
      RECT 96.205 4.748 96.63 5.165 ;
      RECT 96.045 4.94 96.63 5.165 ;
      RECT 96.195 4.76 96.63 5.165 ;
      RECT 96.08 4.877 96.63 5.165 ;
      RECT 96.135 4.802 96.63 5.165 ;
      RECT 96.385 4.667 96.625 5.18 ;
      RECT 96.415 4.66 96.625 5.18 ;
      RECT 96.405 4.662 96.625 5.18 ;
      RECT 96.415 4.657 96.545 5.18 ;
      RECT 95.97 3.22 96.056 3.659 ;
      RECT 95.965 3.22 96.056 3.657 ;
      RECT 95.965 3.22 96.125 3.656 ;
      RECT 95.965 3.22 96.155 3.653 ;
      RECT 95.95 3.227 96.155 3.644 ;
      RECT 95.95 3.227 96.16 3.64 ;
      RECT 95.945 3.237 96.16 3.633 ;
      RECT 95.94 3.242 96.16 3.608 ;
      RECT 95.94 3.242 96.175 3.59 ;
      RECT 95.965 3.22 96.195 3.505 ;
      RECT 95.935 3.247 96.195 3.503 ;
      RECT 95.945 3.24 96.2 3.441 ;
      RECT 95.935 3.362 96.205 3.424 ;
      RECT 95.92 3.257 96.2 3.375 ;
      RECT 95.915 3.267 96.2 3.275 ;
      RECT 95.995 4.038 96 4.115 ;
      RECT 95.985 4.032 95.995 4.305 ;
      RECT 95.975 4.024 95.985 4.326 ;
      RECT 95.965 4.015 95.975 4.348 ;
      RECT 95.96 4.01 95.965 4.365 ;
      RECT 95.92 4.01 95.96 4.405 ;
      RECT 95.9 4.01 95.92 4.46 ;
      RECT 95.895 4.01 95.9 4.488 ;
      RECT 95.885 4.01 95.895 4.503 ;
      RECT 95.85 4.01 95.885 4.545 ;
      RECT 95.845 4.01 95.85 4.588 ;
      RECT 95.835 4.01 95.845 4.603 ;
      RECT 95.82 4.01 95.835 4.623 ;
      RECT 95.805 4.01 95.82 4.65 ;
      RECT 95.8 4.011 95.805 4.668 ;
      RECT 95.78 4.012 95.8 4.675 ;
      RECT 95.725 4.013 95.78 4.695 ;
      RECT 95.715 4.014 95.725 4.709 ;
      RECT 95.71 4.017 95.715 4.708 ;
      RECT 95.67 4.09 95.71 4.706 ;
      RECT 95.655 4.17 95.67 4.704 ;
      RECT 95.63 4.225 95.655 4.702 ;
      RECT 95.615 4.29 95.63 4.701 ;
      RECT 95.57 4.322 95.615 4.698 ;
      RECT 95.485 4.345 95.57 4.693 ;
      RECT 95.46 4.365 95.485 4.688 ;
      RECT 95.39 4.37 95.46 4.684 ;
      RECT 95.37 4.372 95.39 4.681 ;
      RECT 95.285 4.383 95.37 4.675 ;
      RECT 95.28 4.394 95.285 4.67 ;
      RECT 95.27 4.396 95.28 4.67 ;
      RECT 95.235 4.4 95.27 4.668 ;
      RECT 95.185 4.41 95.235 4.655 ;
      RECT 95.165 4.418 95.185 4.64 ;
      RECT 95.085 4.43 95.165 4.623 ;
      RECT 95.25 3.98 95.42 4.19 ;
      RECT 95.366 3.976 95.42 4.19 ;
      RECT 95.171 3.98 95.42 4.181 ;
      RECT 95.171 3.98 95.425 4.17 ;
      RECT 95.085 3.98 95.425 4.161 ;
      RECT 95.085 3.988 95.435 4.105 ;
      RECT 95.085 4 95.44 4.018 ;
      RECT 95.085 4.007 95.445 4.01 ;
      RECT 95.28 3.978 95.42 4.19 ;
      RECT 95.035 4.923 95.28 5.255 ;
      RECT 95.03 4.915 95.035 5.252 ;
      RECT 95 4.935 95.28 5.233 ;
      RECT 94.98 4.967 95.28 5.206 ;
      RECT 95.03 4.92 95.207 5.252 ;
      RECT 95.03 4.917 95.121 5.252 ;
      RECT 94.97 3.265 95.14 3.685 ;
      RECT 94.965 3.265 95.14 3.683 ;
      RECT 94.965 3.265 95.165 3.673 ;
      RECT 94.965 3.265 95.185 3.648 ;
      RECT 94.96 3.265 95.185 3.643 ;
      RECT 94.96 3.265 95.195 3.633 ;
      RECT 94.96 3.265 95.2 3.628 ;
      RECT 94.96 3.27 95.205 3.623 ;
      RECT 94.96 3.302 95.22 3.613 ;
      RECT 94.96 3.372 95.245 3.596 ;
      RECT 94.94 3.372 95.245 3.588 ;
      RECT 94.94 3.432 95.255 3.565 ;
      RECT 94.94 3.472 95.265 3.51 ;
      RECT 94.925 3.265 95.2 3.49 ;
      RECT 94.915 3.28 95.205 3.388 ;
      RECT 94.505 4.67 94.675 5.195 ;
      RECT 94.5 4.67 94.675 5.188 ;
      RECT 94.49 4.67 94.68 5.153 ;
      RECT 94.485 4.68 94.68 5.125 ;
      RECT 94.48 4.7 94.68 5.108 ;
      RECT 94.49 4.675 94.685 5.098 ;
      RECT 94.475 4.72 94.685 5.09 ;
      RECT 94.47 4.74 94.685 5.075 ;
      RECT 94.465 4.77 94.685 5.065 ;
      RECT 94.455 4.815 94.685 5.04 ;
      RECT 94.485 4.685 94.69 5.023 ;
      RECT 94.45 4.867 94.69 5.018 ;
      RECT 94.485 4.695 94.695 4.988 ;
      RECT 94.445 4.9 94.695 4.985 ;
      RECT 94.44 4.925 94.695 4.965 ;
      RECT 94.48 4.712 94.705 4.905 ;
      RECT 94.475 4.734 94.715 4.798 ;
      RECT 94.425 3.981 94.44 4.25 ;
      RECT 94.38 3.965 94.425 4.295 ;
      RECT 94.375 3.953 94.38 4.345 ;
      RECT 94.365 3.949 94.375 4.378 ;
      RECT 94.36 3.946 94.365 4.406 ;
      RECT 94.345 3.948 94.36 4.448 ;
      RECT 94.34 3.952 94.345 4.488 ;
      RECT 94.32 3.957 94.34 4.54 ;
      RECT 94.316 3.962 94.32 4.597 ;
      RECT 94.23 3.981 94.316 4.634 ;
      RECT 94.22 4.002 94.23 4.67 ;
      RECT 94.215 4.01 94.22 4.671 ;
      RECT 94.21 4.052 94.215 4.672 ;
      RECT 94.195 4.14 94.21 4.673 ;
      RECT 94.185 4.29 94.195 4.675 ;
      RECT 94.18 4.335 94.185 4.677 ;
      RECT 94.145 4.377 94.18 4.68 ;
      RECT 94.14 4.395 94.145 4.683 ;
      RECT 94.063 4.401 94.14 4.689 ;
      RECT 93.977 4.415 94.063 4.702 ;
      RECT 93.891 4.429 93.977 4.716 ;
      RECT 93.805 4.443 93.891 4.729 ;
      RECT 93.745 4.455 93.805 4.741 ;
      RECT 93.72 4.462 93.745 4.748 ;
      RECT 93.706 4.465 93.72 4.753 ;
      RECT 93.62 4.473 93.706 4.769 ;
      RECT 93.615 4.48 93.62 4.784 ;
      RECT 93.591 4.48 93.615 4.791 ;
      RECT 93.505 4.483 93.591 4.819 ;
      RECT 93.42 4.487 93.505 4.863 ;
      RECT 93.355 4.491 93.42 4.9 ;
      RECT 93.33 4.494 93.355 4.916 ;
      RECT 93.255 4.507 93.33 4.92 ;
      RECT 93.23 4.525 93.255 4.924 ;
      RECT 93.22 4.532 93.23 4.926 ;
      RECT 93.205 4.535 93.22 4.927 ;
      RECT 93.145 4.547 93.205 4.931 ;
      RECT 93.135 4.561 93.145 4.935 ;
      RECT 93.08 4.571 93.135 4.923 ;
      RECT 93.055 4.592 93.08 4.906 ;
      RECT 93.035 4.612 93.055 4.897 ;
      RECT 93.03 4.625 93.035 4.892 ;
      RECT 93.015 4.637 93.03 4.888 ;
      RECT 94.25 3.292 94.255 3.315 ;
      RECT 94.245 3.283 94.25 3.355 ;
      RECT 94.24 3.281 94.245 3.398 ;
      RECT 94.235 3.272 94.24 3.433 ;
      RECT 94.23 3.262 94.235 3.505 ;
      RECT 94.225 3.252 94.23 3.57 ;
      RECT 94.22 3.249 94.225 3.61 ;
      RECT 94.195 3.243 94.22 3.7 ;
      RECT 94.16 3.231 94.195 3.725 ;
      RECT 94.15 3.222 94.16 3.725 ;
      RECT 94.015 3.22 94.025 3.708 ;
      RECT 94.005 3.22 94.015 3.675 ;
      RECT 94 3.22 94.005 3.65 ;
      RECT 93.995 3.22 94 3.638 ;
      RECT 93.99 3.22 93.995 3.62 ;
      RECT 93.98 3.22 93.99 3.585 ;
      RECT 93.975 3.222 93.98 3.563 ;
      RECT 93.97 3.228 93.975 3.548 ;
      RECT 93.965 3.234 93.97 3.533 ;
      RECT 93.95 3.246 93.965 3.506 ;
      RECT 93.945 3.257 93.95 3.474 ;
      RECT 93.94 3.267 93.945 3.458 ;
      RECT 93.93 3.275 93.94 3.427 ;
      RECT 93.925 3.285 93.93 3.401 ;
      RECT 93.92 3.342 93.925 3.384 ;
      RECT 94.025 3.22 94.15 3.725 ;
      RECT 93.74 3.907 94 4.205 ;
      RECT 93.735 3.914 94 4.203 ;
      RECT 93.74 3.909 94.015 4.198 ;
      RECT 93.73 3.922 94.015 4.195 ;
      RECT 93.73 3.927 94.02 4.188 ;
      RECT 93.725 3.935 94.02 4.185 ;
      RECT 93.725 3.952 94.025 3.983 ;
      RECT 93.74 3.904 93.971 4.205 ;
      RECT 93.795 3.903 93.971 4.205 ;
      RECT 93.795 3.9 93.885 4.205 ;
      RECT 93.795 3.897 93.881 4.205 ;
      RECT 93.485 4.17 93.49 4.183 ;
      RECT 93.48 4.137 93.485 4.188 ;
      RECT 93.475 4.092 93.48 4.195 ;
      RECT 93.47 4.047 93.475 4.203 ;
      RECT 93.465 4.015 93.47 4.211 ;
      RECT 93.46 3.975 93.465 4.212 ;
      RECT 93.445 3.955 93.46 4.214 ;
      RECT 93.37 3.937 93.445 4.226 ;
      RECT 93.36 3.93 93.37 4.237 ;
      RECT 93.355 3.93 93.36 4.239 ;
      RECT 93.325 3.936 93.355 4.243 ;
      RECT 93.285 3.949 93.325 4.243 ;
      RECT 93.26 3.96 93.285 4.229 ;
      RECT 93.245 3.966 93.26 4.212 ;
      RECT 93.235 3.968 93.245 4.203 ;
      RECT 93.23 3.969 93.235 4.198 ;
      RECT 93.225 3.97 93.23 4.193 ;
      RECT 93.22 3.971 93.225 4.19 ;
      RECT 93.195 3.976 93.22 4.18 ;
      RECT 93.185 3.992 93.195 4.167 ;
      RECT 93.18 4.012 93.185 4.162 ;
      RECT 93.19 3.405 93.195 3.601 ;
      RECT 93.175 3.369 93.19 3.603 ;
      RECT 93.165 3.351 93.175 3.608 ;
      RECT 93.155 3.337 93.165 3.612 ;
      RECT 93.11 3.321 93.155 3.622 ;
      RECT 93.105 3.311 93.11 3.631 ;
      RECT 93.06 3.3 93.105 3.637 ;
      RECT 93.055 3.288 93.06 3.644 ;
      RECT 93.04 3.283 93.055 3.648 ;
      RECT 93.025 3.275 93.04 3.653 ;
      RECT 93.015 3.268 93.025 3.658 ;
      RECT 93.005 3.265 93.015 3.663 ;
      RECT 92.995 3.265 93.005 3.664 ;
      RECT 92.99 3.262 92.995 3.663 ;
      RECT 92.955 3.257 92.98 3.662 ;
      RECT 92.931 3.253 92.955 3.661 ;
      RECT 92.845 3.244 92.931 3.658 ;
      RECT 92.83 3.236 92.845 3.655 ;
      RECT 92.808 3.235 92.83 3.654 ;
      RECT 92.722 3.235 92.808 3.652 ;
      RECT 92.636 3.235 92.722 3.65 ;
      RECT 92.55 3.235 92.636 3.647 ;
      RECT 92.54 3.235 92.55 3.638 ;
      RECT 92.51 3.235 92.54 3.598 ;
      RECT 92.5 3.245 92.51 3.553 ;
      RECT 92.495 3.285 92.5 3.538 ;
      RECT 92.49 3.3 92.495 3.525 ;
      RECT 92.46 3.38 92.49 3.487 ;
      RECT 92.98 3.26 92.99 3.663 ;
      RECT 92.805 4.025 92.82 4.63 ;
      RECT 92.81 4.02 92.82 4.63 ;
      RECT 92.975 4.02 92.98 4.203 ;
      RECT 92.965 4.02 92.975 4.233 ;
      RECT 92.95 4.02 92.965 4.293 ;
      RECT 92.945 4.02 92.95 4.338 ;
      RECT 92.94 4.02 92.945 4.368 ;
      RECT 92.935 4.02 92.94 4.388 ;
      RECT 92.925 4.02 92.935 4.423 ;
      RECT 92.91 4.02 92.925 4.455 ;
      RECT 92.865 4.02 92.91 4.483 ;
      RECT 92.86 4.02 92.865 4.513 ;
      RECT 92.855 4.02 92.86 4.525 ;
      RECT 92.85 4.02 92.855 4.533 ;
      RECT 92.84 4.02 92.85 4.548 ;
      RECT 92.835 4.02 92.84 4.57 ;
      RECT 92.825 4.02 92.835 4.593 ;
      RECT 92.82 4.02 92.825 4.613 ;
      RECT 92.785 4.035 92.805 4.63 ;
      RECT 92.76 4.052 92.785 4.63 ;
      RECT 92.755 4.062 92.76 4.63 ;
      RECT 92.725 4.077 92.755 4.63 ;
      RECT 92.65 4.119 92.725 4.63 ;
      RECT 92.645 4.15 92.65 4.613 ;
      RECT 92.64 4.154 92.645 4.595 ;
      RECT 92.635 4.158 92.64 4.558 ;
      RECT 92.63 4.342 92.635 4.525 ;
      RECT 92.115 4.531 92.201 5.096 ;
      RECT 92.07 4.533 92.235 5.09 ;
      RECT 92.201 4.53 92.235 5.09 ;
      RECT 92.115 4.532 92.32 5.084 ;
      RECT 92.07 4.542 92.33 5.08 ;
      RECT 92.045 4.534 92.32 5.076 ;
      RECT 92.04 4.537 92.32 5.071 ;
      RECT 92.015 4.552 92.33 5.065 ;
      RECT 92.015 4.577 92.37 5.06 ;
      RECT 91.975 4.585 92.37 5.035 ;
      RECT 91.975 4.612 92.385 5.033 ;
      RECT 91.975 4.642 92.395 5.02 ;
      RECT 91.97 4.787 92.395 5.008 ;
      RECT 91.975 4.716 92.415 5.005 ;
      RECT 91.975 4.773 92.42 4.813 ;
      RECT 92.165 4.052 92.335 4.23 ;
      RECT 92.115 3.991 92.165 4.215 ;
      RECT 91.85 3.971 92.115 4.2 ;
      RECT 91.81 4.035 92.285 4.2 ;
      RECT 91.81 4.025 92.24 4.2 ;
      RECT 91.81 4.022 92.23 4.2 ;
      RECT 91.81 4.01 92.22 4.2 ;
      RECT 91.81 3.995 92.165 4.2 ;
      RECT 91.85 3.967 92.051 4.2 ;
      RECT 91.86 3.945 92.051 4.2 ;
      RECT 91.885 3.93 91.965 4.2 ;
      RECT 91.64 4.46 91.76 4.905 ;
      RECT 91.625 4.46 91.76 4.904 ;
      RECT 91.58 4.482 91.76 4.899 ;
      RECT 91.54 4.531 91.76 4.893 ;
      RECT 91.54 4.531 91.765 4.868 ;
      RECT 91.54 4.531 91.785 4.758 ;
      RECT 91.535 4.561 91.785 4.755 ;
      RECT 91.625 4.46 91.795 4.65 ;
      RECT 91.285 3.245 91.29 3.69 ;
      RECT 91.095 3.245 91.115 3.655 ;
      RECT 91.065 3.245 91.07 3.63 ;
      RECT 91.745 3.552 91.76 3.74 ;
      RECT 91.74 3.537 91.745 3.746 ;
      RECT 91.72 3.51 91.74 3.749 ;
      RECT 91.67 3.477 91.72 3.758 ;
      RECT 91.64 3.457 91.67 3.762 ;
      RECT 91.621 3.445 91.64 3.758 ;
      RECT 91.535 3.417 91.621 3.748 ;
      RECT 91.525 3.392 91.535 3.738 ;
      RECT 91.455 3.36 91.525 3.73 ;
      RECT 91.43 3.32 91.455 3.722 ;
      RECT 91.41 3.302 91.43 3.716 ;
      RECT 91.4 3.292 91.41 3.713 ;
      RECT 91.39 3.285 91.4 3.711 ;
      RECT 91.37 3.272 91.39 3.708 ;
      RECT 91.36 3.262 91.37 3.705 ;
      RECT 91.35 3.255 91.36 3.703 ;
      RECT 91.3 3.247 91.35 3.697 ;
      RECT 91.29 3.245 91.3 3.691 ;
      RECT 91.26 3.245 91.285 3.688 ;
      RECT 91.231 3.245 91.26 3.683 ;
      RECT 91.145 3.245 91.231 3.673 ;
      RECT 91.115 3.245 91.145 3.66 ;
      RECT 91.07 3.245 91.095 3.643 ;
      RECT 91.055 3.245 91.065 3.625 ;
      RECT 91.035 3.252 91.055 3.61 ;
      RECT 91.03 3.267 91.035 3.598 ;
      RECT 91.025 3.272 91.03 3.538 ;
      RECT 91.02 3.277 91.025 3.38 ;
      RECT 91.015 3.28 91.02 3.298 ;
      RECT 91.28 3.965 91.366 4.286 ;
      RECT 91.28 3.965 91.4 4.279 ;
      RECT 91.23 3.965 91.4 4.275 ;
      RECT 91.23 3.967 91.486 4.273 ;
      RECT 91.23 3.969 91.51 4.267 ;
      RECT 91.23 3.976 91.52 4.266 ;
      RECT 91.23 3.985 91.525 4.263 ;
      RECT 91.23 3.991 91.53 4.258 ;
      RECT 91.23 4.035 91.535 4.255 ;
      RECT 91.23 4.127 91.54 4.252 ;
      RECT 90.755 4.57 90.79 4.89 ;
      RECT 91.34 4.755 91.345 4.937 ;
      RECT 91.295 4.637 91.34 4.956 ;
      RECT 91.28 4.614 91.295 4.979 ;
      RECT 91.27 4.604 91.28 4.989 ;
      RECT 91.25 4.599 91.27 5.002 ;
      RECT 91.225 4.597 91.25 5.023 ;
      RECT 91.206 4.596 91.225 5.035 ;
      RECT 91.12 4.593 91.206 5.035 ;
      RECT 91.05 4.588 91.12 5.023 ;
      RECT 90.975 4.584 91.05 4.998 ;
      RECT 90.91 4.58 90.975 4.965 ;
      RECT 90.84 4.577 90.91 4.925 ;
      RECT 90.81 4.573 90.84 4.9 ;
      RECT 90.79 4.571 90.81 4.893 ;
      RECT 90.706 4.569 90.755 4.891 ;
      RECT 90.62 4.566 90.706 4.892 ;
      RECT 90.545 4.565 90.62 4.894 ;
      RECT 90.46 4.565 90.545 4.92 ;
      RECT 90.383 4.566 90.46 4.945 ;
      RECT 90.297 4.567 90.383 4.945 ;
      RECT 90.211 4.567 90.297 4.945 ;
      RECT 90.125 4.568 90.211 4.945 ;
      RECT 90.105 4.569 90.125 4.937 ;
      RECT 90.09 4.575 90.105 4.922 ;
      RECT 90.055 4.595 90.09 4.902 ;
      RECT 90.045 4.615 90.055 4.884 ;
      RECT 91.015 3.92 91.02 4.19 ;
      RECT 91.01 3.911 91.015 4.195 ;
      RECT 91 3.901 91.01 4.207 ;
      RECT 90.995 3.89 91 4.218 ;
      RECT 90.975 3.884 90.995 4.236 ;
      RECT 90.93 3.881 90.975 4.285 ;
      RECT 90.915 3.88 90.93 4.33 ;
      RECT 90.91 3.88 90.915 4.343 ;
      RECT 90.9 3.88 90.91 4.355 ;
      RECT 90.895 3.881 90.9 4.37 ;
      RECT 90.875 3.889 90.895 4.375 ;
      RECT 90.845 3.905 90.875 4.375 ;
      RECT 90.835 3.917 90.84 4.375 ;
      RECT 90.8 3.932 90.835 4.375 ;
      RECT 90.77 3.952 90.8 4.375 ;
      RECT 90.76 3.977 90.77 4.375 ;
      RECT 90.755 4.005 90.76 4.375 ;
      RECT 90.75 4.035 90.755 4.375 ;
      RECT 90.745 4.052 90.75 4.375 ;
      RECT 90.735 4.08 90.745 4.375 ;
      RECT 90.725 4.115 90.735 4.375 ;
      RECT 90.72 4.15 90.725 4.375 ;
      RECT 90.84 3.915 90.845 4.375 ;
      RECT 90.355 4.017 90.54 4.19 ;
      RECT 90.315 3.935 90.5 4.188 ;
      RECT 90.276 3.94 90.5 4.184 ;
      RECT 90.19 3.949 90.5 4.179 ;
      RECT 90.106 3.965 90.505 4.174 ;
      RECT 90.02 3.985 90.53 4.168 ;
      RECT 90.02 4.005 90.535 4.168 ;
      RECT 90.106 3.975 90.53 4.174 ;
      RECT 90.19 3.95 90.505 4.179 ;
      RECT 90.355 3.932 90.5 4.19 ;
      RECT 90.355 3.927 90.455 4.19 ;
      RECT 90.441 3.921 90.455 4.19 ;
      RECT 89.83 3.245 89.835 3.644 ;
      RECT 89.575 3.245 89.61 3.642 ;
      RECT 89.17 3.28 89.175 3.636 ;
      RECT 89.915 3.283 89.92 3.538 ;
      RECT 89.91 3.281 89.915 3.544 ;
      RECT 89.905 3.28 89.91 3.551 ;
      RECT 89.88 3.273 89.905 3.575 ;
      RECT 89.875 3.266 89.88 3.599 ;
      RECT 89.87 3.262 89.875 3.608 ;
      RECT 89.86 3.257 89.87 3.621 ;
      RECT 89.855 3.254 89.86 3.63 ;
      RECT 89.85 3.252 89.855 3.635 ;
      RECT 89.835 3.248 89.85 3.645 ;
      RECT 89.82 3.242 89.83 3.644 ;
      RECT 89.782 3.24 89.82 3.644 ;
      RECT 89.696 3.242 89.782 3.644 ;
      RECT 89.61 3.244 89.696 3.643 ;
      RECT 89.539 3.245 89.575 3.642 ;
      RECT 89.453 3.247 89.539 3.642 ;
      RECT 89.367 3.249 89.453 3.641 ;
      RECT 89.281 3.251 89.367 3.641 ;
      RECT 89.195 3.254 89.281 3.64 ;
      RECT 89.185 3.26 89.195 3.639 ;
      RECT 89.175 3.272 89.185 3.637 ;
      RECT 89.115 3.307 89.17 3.633 ;
      RECT 89.11 3.337 89.115 3.395 ;
      RECT 89.855 4.417 89.87 4.61 ;
      RECT 89.85 4.385 89.855 4.61 ;
      RECT 89.84 4.36 89.85 4.61 ;
      RECT 89.835 4.332 89.84 4.61 ;
      RECT 89.805 4.255 89.835 4.61 ;
      RECT 89.78 4.137 89.805 4.61 ;
      RECT 89.775 4.075 89.78 4.61 ;
      RECT 89.765 4.062 89.775 4.61 ;
      RECT 89.745 4.052 89.765 4.61 ;
      RECT 89.73 4.035 89.745 4.61 ;
      RECT 89.7 4.023 89.73 4.61 ;
      RECT 89.695 4.022 89.7 4.555 ;
      RECT 89.69 4.022 89.695 4.513 ;
      RECT 89.675 4.021 89.69 4.465 ;
      RECT 89.66 4.021 89.675 4.403 ;
      RECT 89.64 4.021 89.66 4.363 ;
      RECT 89.635 4.021 89.64 4.348 ;
      RECT 89.61 4.02 89.635 4.343 ;
      RECT 89.54 4.019 89.61 4.33 ;
      RECT 89.525 4.018 89.54 4.315 ;
      RECT 89.495 4.017 89.525 4.298 ;
      RECT 89.49 4.017 89.495 4.283 ;
      RECT 89.44 4.016 89.49 4.263 ;
      RECT 89.375 4.015 89.44 4.218 ;
      RECT 89.37 4.015 89.375 4.19 ;
      RECT 89.455 4.552 89.46 4.809 ;
      RECT 89.435 4.471 89.455 4.826 ;
      RECT 89.415 4.465 89.435 4.855 ;
      RECT 89.355 4.452 89.415 4.875 ;
      RECT 89.31 4.436 89.355 4.876 ;
      RECT 89.226 4.424 89.31 4.864 ;
      RECT 89.14 4.411 89.226 4.848 ;
      RECT 89.13 4.404 89.14 4.84 ;
      RECT 89.085 4.401 89.13 4.78 ;
      RECT 89.065 4.397 89.085 4.695 ;
      RECT 89.05 4.395 89.065 4.648 ;
      RECT 89.02 4.392 89.05 4.618 ;
      RECT 88.985 4.388 89.02 4.595 ;
      RECT 88.942 4.383 88.985 4.583 ;
      RECT 88.856 4.374 88.942 4.592 ;
      RECT 88.77 4.363 88.856 4.604 ;
      RECT 88.705 4.354 88.77 4.613 ;
      RECT 88.685 4.345 88.705 4.618 ;
      RECT 88.68 4.338 88.685 4.62 ;
      RECT 88.64 4.323 88.68 4.617 ;
      RECT 88.62 4.302 88.64 4.612 ;
      RECT 88.605 4.29 88.62 4.605 ;
      RECT 88.6 4.282 88.605 4.598 ;
      RECT 88.585 4.262 88.6 4.591 ;
      RECT 88.58 4.125 88.585 4.585 ;
      RECT 88.5 4.014 88.58 4.557 ;
      RECT 88.491 4.007 88.5 4.523 ;
      RECT 88.405 4.001 88.491 4.448 ;
      RECT 88.38 3.992 88.405 4.36 ;
      RECT 88.35 3.987 88.38 4.335 ;
      RECT 88.285 3.996 88.35 4.32 ;
      RECT 88.265 4.012 88.285 4.295 ;
      RECT 88.255 4.018 88.265 4.243 ;
      RECT 88.235 4.04 88.255 4.125 ;
      RECT 88.89 4.005 89.06 4.19 ;
      RECT 88.89 4.005 89.095 4.188 ;
      RECT 88.94 3.915 89.11 4.179 ;
      RECT 88.89 4.072 89.115 4.172 ;
      RECT 88.905 3.95 89.11 4.179 ;
      RECT 88.105 4.683 88.17 5.126 ;
      RECT 88.045 4.708 88.17 5.124 ;
      RECT 88.045 4.708 88.225 5.118 ;
      RECT 88.03 4.733 88.225 5.117 ;
      RECT 88.17 4.67 88.245 5.114 ;
      RECT 88.105 4.695 88.325 5.108 ;
      RECT 88.03 4.734 88.37 5.102 ;
      RECT 88.015 4.761 88.37 5.093 ;
      RECT 88.03 4.754 88.39 5.085 ;
      RECT 88.015 4.763 88.395 5.068 ;
      RECT 88.01 4.78 88.395 4.895 ;
      RECT 88.015 3.502 88.05 3.74 ;
      RECT 88.015 3.502 88.08 3.739 ;
      RECT 88.015 3.502 88.195 3.735 ;
      RECT 88.015 3.502 88.25 3.713 ;
      RECT 88.025 3.445 88.305 3.613 ;
      RECT 88.13 3.285 88.16 3.736 ;
      RECT 88.16 3.28 88.34 3.493 ;
      RECT 88.03 3.421 88.34 3.493 ;
      RECT 88.08 3.317 88.13 3.737 ;
      RECT 88.05 3.373 88.34 3.493 ;
      RECT 86.55 3.035 86.72 4.225 ;
      RECT 86.55 3.035 87.02 3.205 ;
      RECT 86.55 9.405 87.02 9.575 ;
      RECT 86.55 8.385 86.72 9.575 ;
      RECT 85.56 3.035 85.73 4.225 ;
      RECT 85.56 3.035 86.03 3.205 ;
      RECT 85.56 9.405 86.03 9.575 ;
      RECT 85.56 8.385 85.73 9.575 ;
      RECT 83.71 3.93 83.88 5.16 ;
      RECT 83.765 2.15 83.935 4.1 ;
      RECT 83.71 1.87 83.88 2.32 ;
      RECT 83.71 10.29 83.88 10.74 ;
      RECT 83.765 8.51 83.935 10.46 ;
      RECT 83.71 7.45 83.88 8.68 ;
      RECT 83.19 1.87 83.36 5.16 ;
      RECT 83.19 3.37 83.595 3.7 ;
      RECT 83.19 2.53 83.595 2.86 ;
      RECT 83.19 7.45 83.36 10.74 ;
      RECT 83.19 9.75 83.595 10.08 ;
      RECT 83.19 8.91 83.595 9.24 ;
      RECT 81.29 4.687 81.305 4.738 ;
      RECT 81.285 4.667 81.29 4.785 ;
      RECT 81.27 4.657 81.285 4.853 ;
      RECT 81.245 4.637 81.27 4.908 ;
      RECT 81.205 4.622 81.245 4.928 ;
      RECT 81.16 4.616 81.205 4.956 ;
      RECT 81.09 4.606 81.16 4.973 ;
      RECT 81.07 4.598 81.09 4.973 ;
      RECT 81.01 4.592 81.07 4.965 ;
      RECT 80.951 4.583 81.01 4.953 ;
      RECT 80.865 4.572 80.951 4.936 ;
      RECT 80.843 4.563 80.865 4.924 ;
      RECT 80.757 4.556 80.843 4.911 ;
      RECT 80.671 4.543 80.757 4.892 ;
      RECT 80.585 4.531 80.671 4.872 ;
      RECT 80.555 4.52 80.585 4.859 ;
      RECT 80.505 4.506 80.555 4.851 ;
      RECT 80.485 4.495 80.505 4.843 ;
      RECT 80.436 4.484 80.485 4.835 ;
      RECT 80.35 4.463 80.436 4.82 ;
      RECT 80.305 4.45 80.35 4.805 ;
      RECT 80.26 4.45 80.305 4.785 ;
      RECT 80.205 4.45 80.26 4.72 ;
      RECT 80.18 4.45 80.205 4.643 ;
      RECT 80.705 4.187 80.875 4.37 ;
      RECT 80.705 4.187 80.89 4.328 ;
      RECT 80.705 4.187 80.895 4.27 ;
      RECT 80.765 3.955 80.9 4.246 ;
      RECT 80.765 3.959 80.905 4.229 ;
      RECT 80.71 4.122 80.905 4.229 ;
      RECT 80.735 3.967 80.875 4.37 ;
      RECT 80.735 3.971 80.915 4.17 ;
      RECT 80.72 4.057 80.915 4.17 ;
      RECT 80.73 3.987 80.875 4.37 ;
      RECT 80.73 3.99 80.925 4.083 ;
      RECT 80.725 4.007 80.925 4.083 ;
      RECT 80.495 3.227 80.665 3.71 ;
      RECT 80.49 3.222 80.64 3.7 ;
      RECT 80.49 3.229 80.67 3.694 ;
      RECT 80.48 3.223 80.64 3.673 ;
      RECT 80.48 3.239 80.685 3.632 ;
      RECT 80.45 3.224 80.64 3.595 ;
      RECT 80.45 3.254 80.695 3.535 ;
      RECT 80.445 3.226 80.64 3.533 ;
      RECT 80.425 3.235 80.67 3.49 ;
      RECT 80.4 3.251 80.685 3.402 ;
      RECT 80.4 3.27 80.71 3.393 ;
      RECT 80.395 3.307 80.71 3.345 ;
      RECT 80.4 3.287 80.715 3.313 ;
      RECT 80.495 3.221 80.605 3.71 ;
      RECT 80.581 3.22 80.605 3.71 ;
      RECT 79.815 4.005 79.82 4.216 ;
      RECT 80.415 4.005 80.42 4.19 ;
      RECT 80.48 4.045 80.485 4.158 ;
      RECT 80.475 4.037 80.48 4.164 ;
      RECT 80.47 4.027 80.475 4.172 ;
      RECT 80.465 4.017 80.47 4.181 ;
      RECT 80.46 4.007 80.465 4.185 ;
      RECT 80.42 4.005 80.46 4.188 ;
      RECT 80.392 4.004 80.415 4.192 ;
      RECT 80.306 4.001 80.392 4.199 ;
      RECT 80.22 3.997 80.306 4.21 ;
      RECT 80.2 3.995 80.22 4.216 ;
      RECT 80.182 3.994 80.2 4.219 ;
      RECT 80.096 3.992 80.182 4.226 ;
      RECT 80.01 3.987 80.096 4.239 ;
      RECT 79.991 3.984 80.01 4.244 ;
      RECT 79.905 3.982 79.991 4.235 ;
      RECT 79.895 3.982 79.905 4.228 ;
      RECT 79.82 3.995 79.895 4.222 ;
      RECT 79.805 4.006 79.815 4.216 ;
      RECT 79.795 4.008 79.805 4.215 ;
      RECT 79.785 4.012 79.795 4.211 ;
      RECT 79.78 4.015 79.785 4.205 ;
      RECT 79.77 4.017 79.78 4.199 ;
      RECT 79.765 4.02 79.77 4.193 ;
      RECT 79.745 4.606 79.75 4.81 ;
      RECT 79.73 4.593 79.745 4.903 ;
      RECT 79.715 4.574 79.73 5.18 ;
      RECT 79.68 4.54 79.715 5.18 ;
      RECT 79.676 4.51 79.68 5.18 ;
      RECT 79.59 4.392 79.676 5.18 ;
      RECT 79.58 4.267 79.59 5.18 ;
      RECT 79.565 4.235 79.58 5.18 ;
      RECT 79.56 4.21 79.565 5.18 ;
      RECT 79.555 4.2 79.56 5.136 ;
      RECT 79.54 4.172 79.555 5.041 ;
      RECT 79.525 4.138 79.54 4.94 ;
      RECT 79.52 4.116 79.525 4.893 ;
      RECT 79.515 4.105 79.52 4.863 ;
      RECT 79.51 4.095 79.515 4.829 ;
      RECT 79.5 4.082 79.51 4.797 ;
      RECT 79.475 4.058 79.5 4.723 ;
      RECT 79.47 4.038 79.475 4.648 ;
      RECT 79.465 4.032 79.47 4.623 ;
      RECT 79.46 4.027 79.465 4.588 ;
      RECT 79.455 4.022 79.46 4.563 ;
      RECT 79.45 4.02 79.455 4.543 ;
      RECT 79.445 4.02 79.45 4.528 ;
      RECT 79.44 4.02 79.445 4.488 ;
      RECT 79.43 4.02 79.44 4.46 ;
      RECT 79.42 4.02 79.43 4.405 ;
      RECT 79.405 4.02 79.42 4.343 ;
      RECT 79.4 4.019 79.405 4.288 ;
      RECT 79.385 4.018 79.4 4.268 ;
      RECT 79.325 4.016 79.385 4.242 ;
      RECT 79.29 4.017 79.325 4.222 ;
      RECT 79.285 4.019 79.29 4.212 ;
      RECT 79.275 4.038 79.285 4.202 ;
      RECT 79.27 4.065 79.275 4.133 ;
      RECT 79.385 3.49 79.555 3.735 ;
      RECT 79.42 3.261 79.555 3.735 ;
      RECT 79.42 3.263 79.565 3.73 ;
      RECT 79.42 3.265 79.59 3.718 ;
      RECT 79.42 3.268 79.615 3.7 ;
      RECT 79.42 3.273 79.665 3.673 ;
      RECT 79.42 3.278 79.685 3.638 ;
      RECT 79.4 3.28 79.695 3.613 ;
      RECT 79.39 3.375 79.695 3.613 ;
      RECT 79.42 3.26 79.53 3.735 ;
      RECT 79.43 3.257 79.525 3.735 ;
      RECT 78.95 4.522 79.14 4.88 ;
      RECT 78.95 4.534 79.175 4.879 ;
      RECT 78.95 4.562 79.195 4.877 ;
      RECT 78.95 4.587 79.2 4.876 ;
      RECT 78.95 4.645 79.215 4.875 ;
      RECT 78.935 4.518 79.095 4.86 ;
      RECT 78.915 4.527 79.14 4.813 ;
      RECT 78.89 4.538 79.175 4.75 ;
      RECT 78.89 4.622 79.21 4.75 ;
      RECT 78.89 4.597 79.205 4.75 ;
      RECT 78.95 4.513 79.095 4.88 ;
      RECT 79.036 4.512 79.095 4.88 ;
      RECT 79.036 4.511 79.08 4.88 ;
      RECT 78.43 7.45 78.6 10.74 ;
      RECT 78.43 9.75 78.835 10.08 ;
      RECT 78.43 8.91 78.835 9.24 ;
      RECT 78.735 4.027 78.74 4.405 ;
      RECT 78.73 3.995 78.735 4.405 ;
      RECT 78.725 3.967 78.73 4.405 ;
      RECT 78.72 3.947 78.725 4.405 ;
      RECT 78.665 3.93 78.72 4.405 ;
      RECT 78.625 3.915 78.665 4.405 ;
      RECT 78.57 3.902 78.625 4.405 ;
      RECT 78.535 3.893 78.57 4.405 ;
      RECT 78.531 3.891 78.535 4.404 ;
      RECT 78.445 3.887 78.531 4.387 ;
      RECT 78.36 3.879 78.445 4.35 ;
      RECT 78.35 3.875 78.36 4.323 ;
      RECT 78.34 3.875 78.35 4.305 ;
      RECT 78.33 3.877 78.34 4.288 ;
      RECT 78.325 3.882 78.33 4.274 ;
      RECT 78.32 3.886 78.325 4.261 ;
      RECT 78.31 3.891 78.32 4.245 ;
      RECT 78.295 3.905 78.31 4.22 ;
      RECT 78.29 3.911 78.295 4.2 ;
      RECT 78.285 3.913 78.29 4.193 ;
      RECT 78.28 3.917 78.285 4.068 ;
      RECT 78.46 4.717 78.705 5.18 ;
      RECT 78.38 4.69 78.7 5.176 ;
      RECT 78.31 4.725 78.705 5.169 ;
      RECT 78.1 4.98 78.705 5.165 ;
      RECT 78.28 4.748 78.705 5.165 ;
      RECT 78.12 4.94 78.705 5.165 ;
      RECT 78.27 4.76 78.705 5.165 ;
      RECT 78.155 4.877 78.705 5.165 ;
      RECT 78.21 4.802 78.705 5.165 ;
      RECT 78.46 4.667 78.7 5.18 ;
      RECT 78.49 4.66 78.7 5.18 ;
      RECT 78.48 4.662 78.7 5.18 ;
      RECT 78.49 4.657 78.62 5.18 ;
      RECT 78.045 3.22 78.131 3.659 ;
      RECT 78.04 3.22 78.131 3.657 ;
      RECT 78.04 3.22 78.2 3.656 ;
      RECT 78.04 3.22 78.23 3.653 ;
      RECT 78.025 3.227 78.23 3.644 ;
      RECT 78.025 3.227 78.235 3.64 ;
      RECT 78.02 3.237 78.235 3.633 ;
      RECT 78.015 3.242 78.235 3.608 ;
      RECT 78.015 3.242 78.25 3.59 ;
      RECT 78.04 3.22 78.27 3.505 ;
      RECT 78.01 3.247 78.27 3.503 ;
      RECT 78.02 3.24 78.275 3.441 ;
      RECT 78.01 3.362 78.28 3.424 ;
      RECT 77.995 3.257 78.275 3.375 ;
      RECT 77.99 3.267 78.275 3.275 ;
      RECT 78.07 4.038 78.075 4.115 ;
      RECT 78.06 4.032 78.07 4.305 ;
      RECT 78.05 4.024 78.06 4.326 ;
      RECT 78.04 4.015 78.05 4.348 ;
      RECT 78.035 4.01 78.04 4.365 ;
      RECT 77.995 4.01 78.035 4.405 ;
      RECT 77.975 4.01 77.995 4.46 ;
      RECT 77.97 4.01 77.975 4.488 ;
      RECT 77.96 4.01 77.97 4.503 ;
      RECT 77.925 4.01 77.96 4.545 ;
      RECT 77.92 4.01 77.925 4.588 ;
      RECT 77.91 4.01 77.92 4.603 ;
      RECT 77.895 4.01 77.91 4.623 ;
      RECT 77.88 4.01 77.895 4.65 ;
      RECT 77.875 4.011 77.88 4.668 ;
      RECT 77.855 4.012 77.875 4.675 ;
      RECT 77.8 4.013 77.855 4.695 ;
      RECT 77.79 4.014 77.8 4.709 ;
      RECT 77.785 4.017 77.79 4.708 ;
      RECT 77.745 4.09 77.785 4.706 ;
      RECT 77.73 4.17 77.745 4.704 ;
      RECT 77.705 4.225 77.73 4.702 ;
      RECT 77.69 4.29 77.705 4.701 ;
      RECT 77.645 4.322 77.69 4.698 ;
      RECT 77.56 4.345 77.645 4.693 ;
      RECT 77.535 4.365 77.56 4.688 ;
      RECT 77.465 4.37 77.535 4.684 ;
      RECT 77.445 4.372 77.465 4.681 ;
      RECT 77.36 4.383 77.445 4.675 ;
      RECT 77.355 4.394 77.36 4.67 ;
      RECT 77.345 4.396 77.355 4.67 ;
      RECT 77.31 4.4 77.345 4.668 ;
      RECT 77.26 4.41 77.31 4.655 ;
      RECT 77.24 4.418 77.26 4.64 ;
      RECT 77.16 4.43 77.24 4.623 ;
      RECT 77.325 3.98 77.495 4.19 ;
      RECT 77.441 3.976 77.495 4.19 ;
      RECT 77.246 3.98 77.495 4.181 ;
      RECT 77.246 3.98 77.5 4.17 ;
      RECT 77.16 3.98 77.5 4.161 ;
      RECT 77.16 3.988 77.51 4.105 ;
      RECT 77.16 4 77.515 4.018 ;
      RECT 77.16 4.007 77.52 4.01 ;
      RECT 77.355 3.978 77.495 4.19 ;
      RECT 77.11 4.923 77.355 5.255 ;
      RECT 77.105 4.915 77.11 5.252 ;
      RECT 77.075 4.935 77.355 5.233 ;
      RECT 77.055 4.967 77.355 5.206 ;
      RECT 77.105 4.92 77.282 5.252 ;
      RECT 77.105 4.917 77.196 5.252 ;
      RECT 77.045 3.265 77.215 3.685 ;
      RECT 77.04 3.265 77.215 3.683 ;
      RECT 77.04 3.265 77.24 3.673 ;
      RECT 77.04 3.265 77.26 3.648 ;
      RECT 77.035 3.265 77.26 3.643 ;
      RECT 77.035 3.265 77.27 3.633 ;
      RECT 77.035 3.265 77.275 3.628 ;
      RECT 77.035 3.27 77.28 3.623 ;
      RECT 77.035 3.302 77.295 3.613 ;
      RECT 77.035 3.372 77.32 3.596 ;
      RECT 77.015 3.372 77.32 3.588 ;
      RECT 77.015 3.432 77.33 3.565 ;
      RECT 77.015 3.472 77.34 3.51 ;
      RECT 77 3.265 77.275 3.49 ;
      RECT 76.99 3.28 77.28 3.388 ;
      RECT 76.58 4.67 76.75 5.195 ;
      RECT 76.575 4.67 76.75 5.188 ;
      RECT 76.565 4.67 76.755 5.153 ;
      RECT 76.56 4.68 76.755 5.125 ;
      RECT 76.555 4.7 76.755 5.108 ;
      RECT 76.565 4.675 76.76 5.098 ;
      RECT 76.55 4.72 76.76 5.09 ;
      RECT 76.545 4.74 76.76 5.075 ;
      RECT 76.54 4.77 76.76 5.065 ;
      RECT 76.53 4.815 76.76 5.04 ;
      RECT 76.56 4.685 76.765 5.023 ;
      RECT 76.525 4.867 76.765 5.018 ;
      RECT 76.56 4.695 76.77 4.988 ;
      RECT 76.52 4.9 76.77 4.985 ;
      RECT 76.515 4.925 76.77 4.965 ;
      RECT 76.555 4.712 76.78 4.905 ;
      RECT 76.55 4.734 76.79 4.798 ;
      RECT 76.5 3.981 76.515 4.25 ;
      RECT 76.455 3.965 76.5 4.295 ;
      RECT 76.45 3.953 76.455 4.345 ;
      RECT 76.44 3.949 76.45 4.378 ;
      RECT 76.435 3.946 76.44 4.406 ;
      RECT 76.42 3.948 76.435 4.448 ;
      RECT 76.415 3.952 76.42 4.488 ;
      RECT 76.395 3.957 76.415 4.54 ;
      RECT 76.391 3.962 76.395 4.597 ;
      RECT 76.305 3.981 76.391 4.634 ;
      RECT 76.295 4.002 76.305 4.67 ;
      RECT 76.29 4.01 76.295 4.671 ;
      RECT 76.285 4.052 76.29 4.672 ;
      RECT 76.27 4.14 76.285 4.673 ;
      RECT 76.26 4.29 76.27 4.675 ;
      RECT 76.255 4.335 76.26 4.677 ;
      RECT 76.22 4.377 76.255 4.68 ;
      RECT 76.215 4.395 76.22 4.683 ;
      RECT 76.138 4.401 76.215 4.689 ;
      RECT 76.052 4.415 76.138 4.702 ;
      RECT 75.966 4.429 76.052 4.716 ;
      RECT 75.88 4.443 75.966 4.729 ;
      RECT 75.82 4.455 75.88 4.741 ;
      RECT 75.795 4.462 75.82 4.748 ;
      RECT 75.781 4.465 75.795 4.753 ;
      RECT 75.695 4.473 75.781 4.769 ;
      RECT 75.69 4.48 75.695 4.784 ;
      RECT 75.666 4.48 75.69 4.791 ;
      RECT 75.58 4.483 75.666 4.819 ;
      RECT 75.495 4.487 75.58 4.863 ;
      RECT 75.43 4.491 75.495 4.9 ;
      RECT 75.405 4.494 75.43 4.916 ;
      RECT 75.33 4.507 75.405 4.92 ;
      RECT 75.305 4.525 75.33 4.924 ;
      RECT 75.295 4.532 75.305 4.926 ;
      RECT 75.28 4.535 75.295 4.927 ;
      RECT 75.22 4.547 75.28 4.931 ;
      RECT 75.21 4.561 75.22 4.935 ;
      RECT 75.155 4.571 75.21 4.923 ;
      RECT 75.13 4.592 75.155 4.906 ;
      RECT 75.11 4.612 75.13 4.897 ;
      RECT 75.105 4.625 75.11 4.892 ;
      RECT 75.09 4.637 75.105 4.888 ;
      RECT 76.325 3.292 76.33 3.315 ;
      RECT 76.32 3.283 76.325 3.355 ;
      RECT 76.315 3.281 76.32 3.398 ;
      RECT 76.31 3.272 76.315 3.433 ;
      RECT 76.305 3.262 76.31 3.505 ;
      RECT 76.3 3.252 76.305 3.57 ;
      RECT 76.295 3.249 76.3 3.61 ;
      RECT 76.27 3.243 76.295 3.7 ;
      RECT 76.235 3.231 76.27 3.725 ;
      RECT 76.225 3.222 76.235 3.725 ;
      RECT 76.09 3.22 76.1 3.708 ;
      RECT 76.08 3.22 76.09 3.675 ;
      RECT 76.075 3.22 76.08 3.65 ;
      RECT 76.07 3.22 76.075 3.638 ;
      RECT 76.065 3.22 76.07 3.62 ;
      RECT 76.055 3.22 76.065 3.585 ;
      RECT 76.05 3.222 76.055 3.563 ;
      RECT 76.045 3.228 76.05 3.548 ;
      RECT 76.04 3.234 76.045 3.533 ;
      RECT 76.025 3.246 76.04 3.506 ;
      RECT 76.02 3.257 76.025 3.474 ;
      RECT 76.015 3.267 76.02 3.458 ;
      RECT 76.005 3.275 76.015 3.427 ;
      RECT 76 3.285 76.005 3.401 ;
      RECT 75.995 3.342 76 3.384 ;
      RECT 76.1 3.22 76.225 3.725 ;
      RECT 75.815 3.907 76.075 4.205 ;
      RECT 75.81 3.914 76.075 4.203 ;
      RECT 75.815 3.909 76.09 4.198 ;
      RECT 75.805 3.922 76.09 4.195 ;
      RECT 75.805 3.927 76.095 4.188 ;
      RECT 75.8 3.935 76.095 4.185 ;
      RECT 75.8 3.952 76.1 3.983 ;
      RECT 75.815 3.904 76.046 4.205 ;
      RECT 75.87 3.903 76.046 4.205 ;
      RECT 75.87 3.9 75.96 4.205 ;
      RECT 75.87 3.897 75.956 4.205 ;
      RECT 75.56 4.17 75.565 4.183 ;
      RECT 75.555 4.137 75.56 4.188 ;
      RECT 75.55 4.092 75.555 4.195 ;
      RECT 75.545 4.047 75.55 4.203 ;
      RECT 75.54 4.015 75.545 4.211 ;
      RECT 75.535 3.975 75.54 4.212 ;
      RECT 75.52 3.955 75.535 4.214 ;
      RECT 75.445 3.937 75.52 4.226 ;
      RECT 75.435 3.93 75.445 4.237 ;
      RECT 75.43 3.93 75.435 4.239 ;
      RECT 75.4 3.936 75.43 4.243 ;
      RECT 75.36 3.949 75.4 4.243 ;
      RECT 75.335 3.96 75.36 4.229 ;
      RECT 75.32 3.966 75.335 4.212 ;
      RECT 75.31 3.968 75.32 4.203 ;
      RECT 75.305 3.969 75.31 4.198 ;
      RECT 75.3 3.97 75.305 4.193 ;
      RECT 75.295 3.971 75.3 4.19 ;
      RECT 75.27 3.976 75.295 4.18 ;
      RECT 75.26 3.992 75.27 4.167 ;
      RECT 75.255 4.012 75.26 4.162 ;
      RECT 75.265 3.405 75.27 3.601 ;
      RECT 75.25 3.369 75.265 3.603 ;
      RECT 75.24 3.351 75.25 3.608 ;
      RECT 75.23 3.337 75.24 3.612 ;
      RECT 75.185 3.321 75.23 3.622 ;
      RECT 75.18 3.311 75.185 3.631 ;
      RECT 75.135 3.3 75.18 3.637 ;
      RECT 75.13 3.288 75.135 3.644 ;
      RECT 75.115 3.283 75.13 3.648 ;
      RECT 75.1 3.275 75.115 3.653 ;
      RECT 75.09 3.268 75.1 3.658 ;
      RECT 75.08 3.265 75.09 3.663 ;
      RECT 75.07 3.265 75.08 3.664 ;
      RECT 75.065 3.262 75.07 3.663 ;
      RECT 75.03 3.257 75.055 3.662 ;
      RECT 75.006 3.253 75.03 3.661 ;
      RECT 74.92 3.244 75.006 3.658 ;
      RECT 74.905 3.236 74.92 3.655 ;
      RECT 74.883 3.235 74.905 3.654 ;
      RECT 74.797 3.235 74.883 3.652 ;
      RECT 74.711 3.235 74.797 3.65 ;
      RECT 74.625 3.235 74.711 3.647 ;
      RECT 74.615 3.235 74.625 3.638 ;
      RECT 74.585 3.235 74.615 3.598 ;
      RECT 74.575 3.245 74.585 3.553 ;
      RECT 74.57 3.285 74.575 3.538 ;
      RECT 74.565 3.3 74.57 3.525 ;
      RECT 74.535 3.38 74.565 3.487 ;
      RECT 75.055 3.26 75.065 3.663 ;
      RECT 74.88 4.025 74.895 4.63 ;
      RECT 74.885 4.02 74.895 4.63 ;
      RECT 75.05 4.02 75.055 4.203 ;
      RECT 75.04 4.02 75.05 4.233 ;
      RECT 75.025 4.02 75.04 4.293 ;
      RECT 75.02 4.02 75.025 4.338 ;
      RECT 75.015 4.02 75.02 4.368 ;
      RECT 75.01 4.02 75.015 4.388 ;
      RECT 75 4.02 75.01 4.423 ;
      RECT 74.985 4.02 75 4.455 ;
      RECT 74.94 4.02 74.985 4.483 ;
      RECT 74.935 4.02 74.94 4.513 ;
      RECT 74.93 4.02 74.935 4.525 ;
      RECT 74.925 4.02 74.93 4.533 ;
      RECT 74.915 4.02 74.925 4.548 ;
      RECT 74.91 4.02 74.915 4.57 ;
      RECT 74.9 4.02 74.91 4.593 ;
      RECT 74.895 4.02 74.9 4.613 ;
      RECT 74.86 4.035 74.88 4.63 ;
      RECT 74.835 4.052 74.86 4.63 ;
      RECT 74.83 4.062 74.835 4.63 ;
      RECT 74.8 4.077 74.83 4.63 ;
      RECT 74.725 4.119 74.8 4.63 ;
      RECT 74.72 4.15 74.725 4.613 ;
      RECT 74.715 4.154 74.72 4.595 ;
      RECT 74.71 4.158 74.715 4.558 ;
      RECT 74.705 4.342 74.71 4.525 ;
      RECT 74.19 4.531 74.276 5.096 ;
      RECT 74.145 4.533 74.31 5.09 ;
      RECT 74.276 4.53 74.31 5.09 ;
      RECT 74.19 4.532 74.395 5.084 ;
      RECT 74.145 4.542 74.405 5.08 ;
      RECT 74.12 4.534 74.395 5.076 ;
      RECT 74.115 4.537 74.395 5.071 ;
      RECT 74.09 4.552 74.405 5.065 ;
      RECT 74.09 4.577 74.445 5.06 ;
      RECT 74.05 4.585 74.445 5.035 ;
      RECT 74.05 4.612 74.46 5.033 ;
      RECT 74.05 4.642 74.47 5.02 ;
      RECT 74.045 4.787 74.47 5.008 ;
      RECT 74.05 4.716 74.49 5.005 ;
      RECT 74.05 4.773 74.495 4.813 ;
      RECT 74.24 4.052 74.41 4.23 ;
      RECT 74.19 3.991 74.24 4.215 ;
      RECT 73.925 3.971 74.19 4.2 ;
      RECT 73.885 4.035 74.36 4.2 ;
      RECT 73.885 4.025 74.315 4.2 ;
      RECT 73.885 4.022 74.305 4.2 ;
      RECT 73.885 4.01 74.295 4.2 ;
      RECT 73.885 3.995 74.24 4.2 ;
      RECT 73.925 3.967 74.126 4.2 ;
      RECT 73.935 3.945 74.126 4.2 ;
      RECT 73.96 3.93 74.04 4.2 ;
      RECT 73.715 4.46 73.835 4.905 ;
      RECT 73.7 4.46 73.835 4.904 ;
      RECT 73.655 4.482 73.835 4.899 ;
      RECT 73.615 4.531 73.835 4.893 ;
      RECT 73.615 4.531 73.84 4.868 ;
      RECT 73.615 4.531 73.86 4.758 ;
      RECT 73.61 4.561 73.86 4.755 ;
      RECT 73.7 4.46 73.87 4.65 ;
      RECT 73.36 3.245 73.365 3.69 ;
      RECT 73.17 3.245 73.19 3.655 ;
      RECT 73.14 3.245 73.145 3.63 ;
      RECT 73.82 3.552 73.835 3.74 ;
      RECT 73.815 3.537 73.82 3.746 ;
      RECT 73.795 3.51 73.815 3.749 ;
      RECT 73.745 3.477 73.795 3.758 ;
      RECT 73.715 3.457 73.745 3.762 ;
      RECT 73.696 3.445 73.715 3.758 ;
      RECT 73.61 3.417 73.696 3.748 ;
      RECT 73.6 3.392 73.61 3.738 ;
      RECT 73.53 3.36 73.6 3.73 ;
      RECT 73.505 3.32 73.53 3.722 ;
      RECT 73.485 3.302 73.505 3.716 ;
      RECT 73.475 3.292 73.485 3.713 ;
      RECT 73.465 3.285 73.475 3.711 ;
      RECT 73.445 3.272 73.465 3.708 ;
      RECT 73.435 3.262 73.445 3.705 ;
      RECT 73.425 3.255 73.435 3.703 ;
      RECT 73.375 3.247 73.425 3.697 ;
      RECT 73.365 3.245 73.375 3.691 ;
      RECT 73.335 3.245 73.36 3.688 ;
      RECT 73.306 3.245 73.335 3.683 ;
      RECT 73.22 3.245 73.306 3.673 ;
      RECT 73.19 3.245 73.22 3.66 ;
      RECT 73.145 3.245 73.17 3.643 ;
      RECT 73.13 3.245 73.14 3.625 ;
      RECT 73.11 3.252 73.13 3.61 ;
      RECT 73.105 3.267 73.11 3.598 ;
      RECT 73.1 3.272 73.105 3.538 ;
      RECT 73.095 3.277 73.1 3.38 ;
      RECT 73.09 3.28 73.095 3.298 ;
      RECT 73.355 3.965 73.441 4.286 ;
      RECT 73.355 3.965 73.475 4.279 ;
      RECT 73.305 3.965 73.475 4.275 ;
      RECT 73.305 3.967 73.561 4.273 ;
      RECT 73.305 3.969 73.585 4.267 ;
      RECT 73.305 3.976 73.595 4.266 ;
      RECT 73.305 3.985 73.6 4.263 ;
      RECT 73.305 3.991 73.605 4.258 ;
      RECT 73.305 4.035 73.61 4.255 ;
      RECT 73.305 4.127 73.615 4.252 ;
      RECT 72.83 4.57 72.865 4.89 ;
      RECT 73.415 4.755 73.42 4.937 ;
      RECT 73.37 4.637 73.415 4.956 ;
      RECT 73.355 4.614 73.37 4.979 ;
      RECT 73.345 4.604 73.355 4.989 ;
      RECT 73.325 4.599 73.345 5.002 ;
      RECT 73.3 4.597 73.325 5.023 ;
      RECT 73.281 4.596 73.3 5.035 ;
      RECT 73.195 4.593 73.281 5.035 ;
      RECT 73.125 4.588 73.195 5.023 ;
      RECT 73.05 4.584 73.125 4.998 ;
      RECT 72.985 4.58 73.05 4.965 ;
      RECT 72.915 4.577 72.985 4.925 ;
      RECT 72.885 4.573 72.915 4.9 ;
      RECT 72.865 4.571 72.885 4.893 ;
      RECT 72.781 4.569 72.83 4.891 ;
      RECT 72.695 4.566 72.781 4.892 ;
      RECT 72.62 4.565 72.695 4.894 ;
      RECT 72.535 4.565 72.62 4.92 ;
      RECT 72.458 4.566 72.535 4.945 ;
      RECT 72.372 4.567 72.458 4.945 ;
      RECT 72.286 4.567 72.372 4.945 ;
      RECT 72.2 4.568 72.286 4.945 ;
      RECT 72.18 4.569 72.2 4.937 ;
      RECT 72.165 4.575 72.18 4.922 ;
      RECT 72.13 4.595 72.165 4.902 ;
      RECT 72.12 4.615 72.13 4.884 ;
      RECT 73.09 3.92 73.095 4.19 ;
      RECT 73.085 3.911 73.09 4.195 ;
      RECT 73.075 3.901 73.085 4.207 ;
      RECT 73.07 3.89 73.075 4.218 ;
      RECT 73.05 3.884 73.07 4.236 ;
      RECT 73.005 3.881 73.05 4.285 ;
      RECT 72.99 3.88 73.005 4.33 ;
      RECT 72.985 3.88 72.99 4.343 ;
      RECT 72.975 3.88 72.985 4.355 ;
      RECT 72.97 3.881 72.975 4.37 ;
      RECT 72.95 3.889 72.97 4.375 ;
      RECT 72.92 3.905 72.95 4.375 ;
      RECT 72.91 3.917 72.915 4.375 ;
      RECT 72.875 3.932 72.91 4.375 ;
      RECT 72.845 3.952 72.875 4.375 ;
      RECT 72.835 3.977 72.845 4.375 ;
      RECT 72.83 4.005 72.835 4.375 ;
      RECT 72.825 4.035 72.83 4.375 ;
      RECT 72.82 4.052 72.825 4.375 ;
      RECT 72.81 4.08 72.82 4.375 ;
      RECT 72.8 4.115 72.81 4.375 ;
      RECT 72.795 4.15 72.8 4.375 ;
      RECT 72.915 3.915 72.92 4.375 ;
      RECT 72.43 4.017 72.615 4.19 ;
      RECT 72.39 3.935 72.575 4.188 ;
      RECT 72.351 3.94 72.575 4.184 ;
      RECT 72.265 3.949 72.575 4.179 ;
      RECT 72.181 3.965 72.58 4.174 ;
      RECT 72.095 3.985 72.605 4.168 ;
      RECT 72.095 4.005 72.61 4.168 ;
      RECT 72.181 3.975 72.605 4.174 ;
      RECT 72.265 3.95 72.58 4.179 ;
      RECT 72.43 3.932 72.575 4.19 ;
      RECT 72.43 3.927 72.53 4.19 ;
      RECT 72.516 3.921 72.53 4.19 ;
      RECT 71.905 3.245 71.91 3.644 ;
      RECT 71.65 3.245 71.685 3.642 ;
      RECT 71.245 3.28 71.25 3.636 ;
      RECT 71.99 3.283 71.995 3.538 ;
      RECT 71.985 3.281 71.99 3.544 ;
      RECT 71.98 3.28 71.985 3.551 ;
      RECT 71.955 3.273 71.98 3.575 ;
      RECT 71.95 3.266 71.955 3.599 ;
      RECT 71.945 3.262 71.95 3.608 ;
      RECT 71.935 3.257 71.945 3.621 ;
      RECT 71.93 3.254 71.935 3.63 ;
      RECT 71.925 3.252 71.93 3.635 ;
      RECT 71.91 3.248 71.925 3.645 ;
      RECT 71.895 3.242 71.905 3.644 ;
      RECT 71.857 3.24 71.895 3.644 ;
      RECT 71.771 3.242 71.857 3.644 ;
      RECT 71.685 3.244 71.771 3.643 ;
      RECT 71.614 3.245 71.65 3.642 ;
      RECT 71.528 3.247 71.614 3.642 ;
      RECT 71.442 3.249 71.528 3.641 ;
      RECT 71.356 3.251 71.442 3.641 ;
      RECT 71.27 3.254 71.356 3.64 ;
      RECT 71.26 3.26 71.27 3.639 ;
      RECT 71.25 3.272 71.26 3.637 ;
      RECT 71.19 3.307 71.245 3.633 ;
      RECT 71.185 3.337 71.19 3.395 ;
      RECT 71.93 4.417 71.945 4.61 ;
      RECT 71.925 4.385 71.93 4.61 ;
      RECT 71.915 4.36 71.925 4.61 ;
      RECT 71.91 4.332 71.915 4.61 ;
      RECT 71.88 4.255 71.91 4.61 ;
      RECT 71.855 4.137 71.88 4.61 ;
      RECT 71.85 4.075 71.855 4.61 ;
      RECT 71.84 4.062 71.85 4.61 ;
      RECT 71.82 4.052 71.84 4.61 ;
      RECT 71.805 4.035 71.82 4.61 ;
      RECT 71.775 4.023 71.805 4.61 ;
      RECT 71.77 4.022 71.775 4.555 ;
      RECT 71.765 4.022 71.77 4.513 ;
      RECT 71.75 4.021 71.765 4.465 ;
      RECT 71.735 4.021 71.75 4.403 ;
      RECT 71.715 4.021 71.735 4.363 ;
      RECT 71.71 4.021 71.715 4.348 ;
      RECT 71.685 4.02 71.71 4.343 ;
      RECT 71.615 4.019 71.685 4.33 ;
      RECT 71.6 4.018 71.615 4.315 ;
      RECT 71.57 4.017 71.6 4.298 ;
      RECT 71.565 4.017 71.57 4.283 ;
      RECT 71.515 4.016 71.565 4.263 ;
      RECT 71.45 4.015 71.515 4.218 ;
      RECT 71.445 4.015 71.45 4.19 ;
      RECT 71.53 4.552 71.535 4.809 ;
      RECT 71.51 4.471 71.53 4.826 ;
      RECT 71.49 4.465 71.51 4.855 ;
      RECT 71.43 4.452 71.49 4.875 ;
      RECT 71.385 4.436 71.43 4.876 ;
      RECT 71.301 4.424 71.385 4.864 ;
      RECT 71.215 4.411 71.301 4.848 ;
      RECT 71.205 4.404 71.215 4.84 ;
      RECT 71.16 4.401 71.205 4.78 ;
      RECT 71.14 4.397 71.16 4.695 ;
      RECT 71.125 4.395 71.14 4.648 ;
      RECT 71.095 4.392 71.125 4.618 ;
      RECT 71.06 4.388 71.095 4.595 ;
      RECT 71.017 4.383 71.06 4.583 ;
      RECT 70.931 4.374 71.017 4.592 ;
      RECT 70.845 4.363 70.931 4.604 ;
      RECT 70.78 4.354 70.845 4.613 ;
      RECT 70.76 4.345 70.78 4.618 ;
      RECT 70.755 4.338 70.76 4.62 ;
      RECT 70.715 4.323 70.755 4.617 ;
      RECT 70.695 4.302 70.715 4.612 ;
      RECT 70.68 4.29 70.695 4.605 ;
      RECT 70.675 4.282 70.68 4.598 ;
      RECT 70.66 4.262 70.675 4.591 ;
      RECT 70.655 4.125 70.66 4.585 ;
      RECT 70.575 4.014 70.655 4.557 ;
      RECT 70.566 4.007 70.575 4.523 ;
      RECT 70.48 4.001 70.566 4.448 ;
      RECT 70.455 3.992 70.48 4.36 ;
      RECT 70.425 3.987 70.455 4.335 ;
      RECT 70.36 3.996 70.425 4.32 ;
      RECT 70.34 4.012 70.36 4.295 ;
      RECT 70.33 4.018 70.34 4.243 ;
      RECT 70.31 4.04 70.33 4.125 ;
      RECT 70.965 4.005 71.135 4.19 ;
      RECT 70.965 4.005 71.17 4.188 ;
      RECT 71.015 3.915 71.185 4.179 ;
      RECT 70.965 4.072 71.19 4.172 ;
      RECT 70.98 3.95 71.185 4.179 ;
      RECT 70.18 4.683 70.245 5.126 ;
      RECT 70.12 4.708 70.245 5.124 ;
      RECT 70.12 4.708 70.3 5.118 ;
      RECT 70.105 4.733 70.3 5.117 ;
      RECT 70.245 4.67 70.32 5.114 ;
      RECT 70.18 4.695 70.4 5.108 ;
      RECT 70.105 4.734 70.445 5.102 ;
      RECT 70.09 4.761 70.445 5.093 ;
      RECT 70.105 4.754 70.465 5.085 ;
      RECT 70.09 4.763 70.47 5.068 ;
      RECT 70.085 4.78 70.47 4.895 ;
      RECT 70.09 3.502 70.125 3.74 ;
      RECT 70.09 3.502 70.155 3.739 ;
      RECT 70.09 3.502 70.27 3.735 ;
      RECT 70.09 3.502 70.325 3.713 ;
      RECT 70.1 3.445 70.38 3.613 ;
      RECT 70.205 3.285 70.235 3.736 ;
      RECT 70.235 3.28 70.415 3.493 ;
      RECT 70.105 3.421 70.415 3.493 ;
      RECT 70.155 3.317 70.205 3.737 ;
      RECT 70.125 3.373 70.415 3.493 ;
      RECT 68.625 3.035 68.795 4.225 ;
      RECT 68.625 3.035 69.095 3.205 ;
      RECT 68.625 9.405 69.095 9.575 ;
      RECT 68.625 8.385 68.795 9.575 ;
      RECT 67.635 3.035 67.805 4.225 ;
      RECT 67.635 3.035 68.105 3.205 ;
      RECT 67.635 9.405 68.105 9.575 ;
      RECT 67.635 8.385 67.805 9.575 ;
      RECT 65.785 3.93 65.955 5.16 ;
      RECT 65.84 2.15 66.01 4.1 ;
      RECT 65.785 1.87 65.955 2.32 ;
      RECT 65.785 10.29 65.955 10.74 ;
      RECT 65.84 8.51 66.01 10.46 ;
      RECT 65.785 7.45 65.955 8.68 ;
      RECT 65.265 1.87 65.435 5.16 ;
      RECT 65.265 3.37 65.67 3.7 ;
      RECT 65.265 2.53 65.67 2.86 ;
      RECT 65.265 7.45 65.435 10.74 ;
      RECT 65.265 9.75 65.67 10.08 ;
      RECT 65.265 8.91 65.67 9.24 ;
      RECT 63.365 4.687 63.38 4.738 ;
      RECT 63.36 4.667 63.365 4.785 ;
      RECT 63.345 4.657 63.36 4.853 ;
      RECT 63.32 4.637 63.345 4.908 ;
      RECT 63.28 4.622 63.32 4.928 ;
      RECT 63.235 4.616 63.28 4.956 ;
      RECT 63.165 4.606 63.235 4.973 ;
      RECT 63.145 4.598 63.165 4.973 ;
      RECT 63.085 4.592 63.145 4.965 ;
      RECT 63.026 4.583 63.085 4.953 ;
      RECT 62.94 4.572 63.026 4.936 ;
      RECT 62.918 4.563 62.94 4.924 ;
      RECT 62.832 4.556 62.918 4.911 ;
      RECT 62.746 4.543 62.832 4.892 ;
      RECT 62.66 4.531 62.746 4.872 ;
      RECT 62.63 4.52 62.66 4.859 ;
      RECT 62.58 4.506 62.63 4.851 ;
      RECT 62.56 4.495 62.58 4.843 ;
      RECT 62.511 4.484 62.56 4.835 ;
      RECT 62.425 4.463 62.511 4.82 ;
      RECT 62.38 4.45 62.425 4.805 ;
      RECT 62.335 4.45 62.38 4.785 ;
      RECT 62.28 4.45 62.335 4.72 ;
      RECT 62.255 4.45 62.28 4.643 ;
      RECT 62.78 4.187 62.95 4.37 ;
      RECT 62.78 4.187 62.965 4.328 ;
      RECT 62.78 4.187 62.97 4.27 ;
      RECT 62.84 3.955 62.975 4.246 ;
      RECT 62.84 3.959 62.98 4.229 ;
      RECT 62.785 4.122 62.98 4.229 ;
      RECT 62.81 3.967 62.95 4.37 ;
      RECT 62.81 3.971 62.99 4.17 ;
      RECT 62.795 4.057 62.99 4.17 ;
      RECT 62.805 3.987 62.95 4.37 ;
      RECT 62.805 3.99 63 4.083 ;
      RECT 62.8 4.007 63 4.083 ;
      RECT 62.57 3.227 62.74 3.71 ;
      RECT 62.565 3.222 62.715 3.7 ;
      RECT 62.565 3.229 62.745 3.694 ;
      RECT 62.555 3.223 62.715 3.673 ;
      RECT 62.555 3.239 62.76 3.632 ;
      RECT 62.525 3.224 62.715 3.595 ;
      RECT 62.525 3.254 62.77 3.535 ;
      RECT 62.52 3.226 62.715 3.533 ;
      RECT 62.5 3.235 62.745 3.49 ;
      RECT 62.475 3.251 62.76 3.402 ;
      RECT 62.475 3.27 62.785 3.393 ;
      RECT 62.47 3.307 62.785 3.345 ;
      RECT 62.475 3.287 62.79 3.313 ;
      RECT 62.57 3.221 62.68 3.71 ;
      RECT 62.656 3.22 62.68 3.71 ;
      RECT 61.89 4.005 61.895 4.216 ;
      RECT 62.49 4.005 62.495 4.19 ;
      RECT 62.555 4.045 62.56 4.158 ;
      RECT 62.55 4.037 62.555 4.164 ;
      RECT 62.545 4.027 62.55 4.172 ;
      RECT 62.54 4.017 62.545 4.181 ;
      RECT 62.535 4.007 62.54 4.185 ;
      RECT 62.495 4.005 62.535 4.188 ;
      RECT 62.467 4.004 62.49 4.192 ;
      RECT 62.381 4.001 62.467 4.199 ;
      RECT 62.295 3.997 62.381 4.21 ;
      RECT 62.275 3.995 62.295 4.216 ;
      RECT 62.257 3.994 62.275 4.219 ;
      RECT 62.171 3.992 62.257 4.226 ;
      RECT 62.085 3.987 62.171 4.239 ;
      RECT 62.066 3.984 62.085 4.244 ;
      RECT 61.98 3.982 62.066 4.235 ;
      RECT 61.97 3.982 61.98 4.228 ;
      RECT 61.895 3.995 61.97 4.222 ;
      RECT 61.88 4.006 61.89 4.216 ;
      RECT 61.87 4.008 61.88 4.215 ;
      RECT 61.86 4.012 61.87 4.211 ;
      RECT 61.855 4.015 61.86 4.205 ;
      RECT 61.845 4.017 61.855 4.199 ;
      RECT 61.84 4.02 61.845 4.193 ;
      RECT 61.82 4.606 61.825 4.81 ;
      RECT 61.805 4.593 61.82 4.903 ;
      RECT 61.79 4.574 61.805 5.18 ;
      RECT 61.755 4.54 61.79 5.18 ;
      RECT 61.751 4.51 61.755 5.18 ;
      RECT 61.665 4.392 61.751 5.18 ;
      RECT 61.655 4.267 61.665 5.18 ;
      RECT 61.64 4.235 61.655 5.18 ;
      RECT 61.635 4.21 61.64 5.18 ;
      RECT 61.63 4.2 61.635 5.136 ;
      RECT 61.615 4.172 61.63 5.041 ;
      RECT 61.6 4.138 61.615 4.94 ;
      RECT 61.595 4.116 61.6 4.893 ;
      RECT 61.59 4.105 61.595 4.863 ;
      RECT 61.585 4.095 61.59 4.829 ;
      RECT 61.575 4.082 61.585 4.797 ;
      RECT 61.55 4.058 61.575 4.723 ;
      RECT 61.545 4.038 61.55 4.648 ;
      RECT 61.54 4.032 61.545 4.623 ;
      RECT 61.535 4.027 61.54 4.588 ;
      RECT 61.53 4.022 61.535 4.563 ;
      RECT 61.525 4.02 61.53 4.543 ;
      RECT 61.52 4.02 61.525 4.528 ;
      RECT 61.515 4.02 61.52 4.488 ;
      RECT 61.505 4.02 61.515 4.46 ;
      RECT 61.495 4.02 61.505 4.405 ;
      RECT 61.48 4.02 61.495 4.343 ;
      RECT 61.475 4.019 61.48 4.288 ;
      RECT 61.46 4.018 61.475 4.268 ;
      RECT 61.4 4.016 61.46 4.242 ;
      RECT 61.365 4.017 61.4 4.222 ;
      RECT 61.36 4.019 61.365 4.212 ;
      RECT 61.35 4.038 61.36 4.202 ;
      RECT 61.345 4.065 61.35 4.133 ;
      RECT 61.46 3.49 61.63 3.735 ;
      RECT 61.495 3.261 61.63 3.735 ;
      RECT 61.495 3.263 61.64 3.73 ;
      RECT 61.495 3.265 61.665 3.718 ;
      RECT 61.495 3.268 61.69 3.7 ;
      RECT 61.495 3.273 61.74 3.673 ;
      RECT 61.495 3.278 61.76 3.638 ;
      RECT 61.475 3.28 61.77 3.613 ;
      RECT 61.465 3.375 61.77 3.613 ;
      RECT 61.495 3.26 61.605 3.735 ;
      RECT 61.505 3.257 61.6 3.735 ;
      RECT 61.025 4.522 61.215 4.88 ;
      RECT 61.025 4.534 61.25 4.879 ;
      RECT 61.025 4.562 61.27 4.877 ;
      RECT 61.025 4.587 61.275 4.876 ;
      RECT 61.025 4.645 61.29 4.875 ;
      RECT 61.01 4.518 61.17 4.86 ;
      RECT 60.99 4.527 61.215 4.813 ;
      RECT 60.965 4.538 61.25 4.75 ;
      RECT 60.965 4.622 61.285 4.75 ;
      RECT 60.965 4.597 61.28 4.75 ;
      RECT 61.025 4.513 61.17 4.88 ;
      RECT 61.111 4.512 61.17 4.88 ;
      RECT 61.111 4.511 61.155 4.88 ;
      RECT 60.505 7.45 60.675 10.74 ;
      RECT 60.505 9.75 60.91 10.08 ;
      RECT 60.505 8.91 60.91 9.24 ;
      RECT 60.81 4.027 60.815 4.405 ;
      RECT 60.805 3.995 60.81 4.405 ;
      RECT 60.8 3.967 60.805 4.405 ;
      RECT 60.795 3.947 60.8 4.405 ;
      RECT 60.74 3.93 60.795 4.405 ;
      RECT 60.7 3.915 60.74 4.405 ;
      RECT 60.645 3.902 60.7 4.405 ;
      RECT 60.61 3.893 60.645 4.405 ;
      RECT 60.606 3.891 60.61 4.404 ;
      RECT 60.52 3.887 60.606 4.387 ;
      RECT 60.435 3.879 60.52 4.35 ;
      RECT 60.425 3.875 60.435 4.323 ;
      RECT 60.415 3.875 60.425 4.305 ;
      RECT 60.405 3.877 60.415 4.288 ;
      RECT 60.4 3.882 60.405 4.274 ;
      RECT 60.395 3.886 60.4 4.261 ;
      RECT 60.385 3.891 60.395 4.245 ;
      RECT 60.37 3.905 60.385 4.22 ;
      RECT 60.365 3.911 60.37 4.2 ;
      RECT 60.36 3.913 60.365 4.193 ;
      RECT 60.355 3.917 60.36 4.068 ;
      RECT 60.535 4.717 60.78 5.18 ;
      RECT 60.455 4.69 60.775 5.176 ;
      RECT 60.385 4.725 60.78 5.169 ;
      RECT 60.175 4.98 60.78 5.165 ;
      RECT 60.355 4.748 60.78 5.165 ;
      RECT 60.195 4.94 60.78 5.165 ;
      RECT 60.345 4.76 60.78 5.165 ;
      RECT 60.23 4.877 60.78 5.165 ;
      RECT 60.285 4.802 60.78 5.165 ;
      RECT 60.535 4.667 60.775 5.18 ;
      RECT 60.565 4.66 60.775 5.18 ;
      RECT 60.555 4.662 60.775 5.18 ;
      RECT 60.565 4.657 60.695 5.18 ;
      RECT 60.12 3.22 60.206 3.659 ;
      RECT 60.115 3.22 60.206 3.657 ;
      RECT 60.115 3.22 60.275 3.656 ;
      RECT 60.115 3.22 60.305 3.653 ;
      RECT 60.1 3.227 60.305 3.644 ;
      RECT 60.1 3.227 60.31 3.64 ;
      RECT 60.095 3.237 60.31 3.633 ;
      RECT 60.09 3.242 60.31 3.608 ;
      RECT 60.09 3.242 60.325 3.59 ;
      RECT 60.115 3.22 60.345 3.505 ;
      RECT 60.085 3.247 60.345 3.503 ;
      RECT 60.095 3.24 60.35 3.441 ;
      RECT 60.085 3.362 60.355 3.424 ;
      RECT 60.07 3.257 60.35 3.375 ;
      RECT 60.065 3.267 60.35 3.275 ;
      RECT 60.145 4.038 60.15 4.115 ;
      RECT 60.135 4.032 60.145 4.305 ;
      RECT 60.125 4.024 60.135 4.326 ;
      RECT 60.115 4.015 60.125 4.348 ;
      RECT 60.11 4.01 60.115 4.365 ;
      RECT 60.07 4.01 60.11 4.405 ;
      RECT 60.05 4.01 60.07 4.46 ;
      RECT 60.045 4.01 60.05 4.488 ;
      RECT 60.035 4.01 60.045 4.503 ;
      RECT 60 4.01 60.035 4.545 ;
      RECT 59.995 4.01 60 4.588 ;
      RECT 59.985 4.01 59.995 4.603 ;
      RECT 59.97 4.01 59.985 4.623 ;
      RECT 59.955 4.01 59.97 4.65 ;
      RECT 59.95 4.011 59.955 4.668 ;
      RECT 59.93 4.012 59.95 4.675 ;
      RECT 59.875 4.013 59.93 4.695 ;
      RECT 59.865 4.014 59.875 4.709 ;
      RECT 59.86 4.017 59.865 4.708 ;
      RECT 59.82 4.09 59.86 4.706 ;
      RECT 59.805 4.17 59.82 4.704 ;
      RECT 59.78 4.225 59.805 4.702 ;
      RECT 59.765 4.29 59.78 4.701 ;
      RECT 59.72 4.322 59.765 4.698 ;
      RECT 59.635 4.345 59.72 4.693 ;
      RECT 59.61 4.365 59.635 4.688 ;
      RECT 59.54 4.37 59.61 4.684 ;
      RECT 59.52 4.372 59.54 4.681 ;
      RECT 59.435 4.383 59.52 4.675 ;
      RECT 59.43 4.394 59.435 4.67 ;
      RECT 59.42 4.396 59.43 4.67 ;
      RECT 59.385 4.4 59.42 4.668 ;
      RECT 59.335 4.41 59.385 4.655 ;
      RECT 59.315 4.418 59.335 4.64 ;
      RECT 59.235 4.43 59.315 4.623 ;
      RECT 59.4 3.98 59.57 4.19 ;
      RECT 59.516 3.976 59.57 4.19 ;
      RECT 59.321 3.98 59.57 4.181 ;
      RECT 59.321 3.98 59.575 4.17 ;
      RECT 59.235 3.98 59.575 4.161 ;
      RECT 59.235 3.988 59.585 4.105 ;
      RECT 59.235 4 59.59 4.018 ;
      RECT 59.235 4.007 59.595 4.01 ;
      RECT 59.43 3.978 59.57 4.19 ;
      RECT 59.185 4.923 59.43 5.255 ;
      RECT 59.18 4.915 59.185 5.252 ;
      RECT 59.15 4.935 59.43 5.233 ;
      RECT 59.13 4.967 59.43 5.206 ;
      RECT 59.18 4.92 59.357 5.252 ;
      RECT 59.18 4.917 59.271 5.252 ;
      RECT 59.12 3.265 59.29 3.685 ;
      RECT 59.115 3.265 59.29 3.683 ;
      RECT 59.115 3.265 59.315 3.673 ;
      RECT 59.115 3.265 59.335 3.648 ;
      RECT 59.11 3.265 59.335 3.643 ;
      RECT 59.11 3.265 59.345 3.633 ;
      RECT 59.11 3.265 59.35 3.628 ;
      RECT 59.11 3.27 59.355 3.623 ;
      RECT 59.11 3.302 59.37 3.613 ;
      RECT 59.11 3.372 59.395 3.596 ;
      RECT 59.09 3.372 59.395 3.588 ;
      RECT 59.09 3.432 59.405 3.565 ;
      RECT 59.09 3.472 59.415 3.51 ;
      RECT 59.075 3.265 59.35 3.49 ;
      RECT 59.065 3.28 59.355 3.388 ;
      RECT 58.655 4.67 58.825 5.195 ;
      RECT 58.65 4.67 58.825 5.188 ;
      RECT 58.64 4.67 58.83 5.153 ;
      RECT 58.635 4.68 58.83 5.125 ;
      RECT 58.63 4.7 58.83 5.108 ;
      RECT 58.64 4.675 58.835 5.098 ;
      RECT 58.625 4.72 58.835 5.09 ;
      RECT 58.62 4.74 58.835 5.075 ;
      RECT 58.615 4.77 58.835 5.065 ;
      RECT 58.605 4.815 58.835 5.04 ;
      RECT 58.635 4.685 58.84 5.023 ;
      RECT 58.6 4.867 58.84 5.018 ;
      RECT 58.635 4.695 58.845 4.988 ;
      RECT 58.595 4.9 58.845 4.985 ;
      RECT 58.59 4.925 58.845 4.965 ;
      RECT 58.63 4.712 58.855 4.905 ;
      RECT 58.625 4.734 58.865 4.798 ;
      RECT 58.575 3.981 58.59 4.25 ;
      RECT 58.53 3.965 58.575 4.295 ;
      RECT 58.525 3.953 58.53 4.345 ;
      RECT 58.515 3.949 58.525 4.378 ;
      RECT 58.51 3.946 58.515 4.406 ;
      RECT 58.495 3.948 58.51 4.448 ;
      RECT 58.49 3.952 58.495 4.488 ;
      RECT 58.47 3.957 58.49 4.54 ;
      RECT 58.466 3.962 58.47 4.597 ;
      RECT 58.38 3.981 58.466 4.634 ;
      RECT 58.37 4.002 58.38 4.67 ;
      RECT 58.365 4.01 58.37 4.671 ;
      RECT 58.36 4.052 58.365 4.672 ;
      RECT 58.345 4.14 58.36 4.673 ;
      RECT 58.335 4.29 58.345 4.675 ;
      RECT 58.33 4.335 58.335 4.677 ;
      RECT 58.295 4.377 58.33 4.68 ;
      RECT 58.29 4.395 58.295 4.683 ;
      RECT 58.213 4.401 58.29 4.689 ;
      RECT 58.127 4.415 58.213 4.702 ;
      RECT 58.041 4.429 58.127 4.716 ;
      RECT 57.955 4.443 58.041 4.729 ;
      RECT 57.895 4.455 57.955 4.741 ;
      RECT 57.87 4.462 57.895 4.748 ;
      RECT 57.856 4.465 57.87 4.753 ;
      RECT 57.77 4.473 57.856 4.769 ;
      RECT 57.765 4.48 57.77 4.784 ;
      RECT 57.741 4.48 57.765 4.791 ;
      RECT 57.655 4.483 57.741 4.819 ;
      RECT 57.57 4.487 57.655 4.863 ;
      RECT 57.505 4.491 57.57 4.9 ;
      RECT 57.48 4.494 57.505 4.916 ;
      RECT 57.405 4.507 57.48 4.92 ;
      RECT 57.38 4.525 57.405 4.924 ;
      RECT 57.37 4.532 57.38 4.926 ;
      RECT 57.355 4.535 57.37 4.927 ;
      RECT 57.295 4.547 57.355 4.931 ;
      RECT 57.285 4.561 57.295 4.935 ;
      RECT 57.23 4.571 57.285 4.923 ;
      RECT 57.205 4.592 57.23 4.906 ;
      RECT 57.185 4.612 57.205 4.897 ;
      RECT 57.18 4.625 57.185 4.892 ;
      RECT 57.165 4.637 57.18 4.888 ;
      RECT 58.4 3.292 58.405 3.315 ;
      RECT 58.395 3.283 58.4 3.355 ;
      RECT 58.39 3.281 58.395 3.398 ;
      RECT 58.385 3.272 58.39 3.433 ;
      RECT 58.38 3.262 58.385 3.505 ;
      RECT 58.375 3.252 58.38 3.57 ;
      RECT 58.37 3.249 58.375 3.61 ;
      RECT 58.345 3.243 58.37 3.7 ;
      RECT 58.31 3.231 58.345 3.725 ;
      RECT 58.3 3.222 58.31 3.725 ;
      RECT 58.165 3.22 58.175 3.708 ;
      RECT 58.155 3.22 58.165 3.675 ;
      RECT 58.15 3.22 58.155 3.65 ;
      RECT 58.145 3.22 58.15 3.638 ;
      RECT 58.14 3.22 58.145 3.62 ;
      RECT 58.13 3.22 58.14 3.585 ;
      RECT 58.125 3.222 58.13 3.563 ;
      RECT 58.12 3.228 58.125 3.548 ;
      RECT 58.115 3.234 58.12 3.533 ;
      RECT 58.1 3.246 58.115 3.506 ;
      RECT 58.095 3.257 58.1 3.474 ;
      RECT 58.09 3.267 58.095 3.458 ;
      RECT 58.08 3.275 58.09 3.427 ;
      RECT 58.075 3.285 58.08 3.401 ;
      RECT 58.07 3.342 58.075 3.384 ;
      RECT 58.175 3.22 58.3 3.725 ;
      RECT 57.89 3.907 58.15 4.205 ;
      RECT 57.885 3.914 58.15 4.203 ;
      RECT 57.89 3.909 58.165 4.198 ;
      RECT 57.88 3.922 58.165 4.195 ;
      RECT 57.88 3.927 58.17 4.188 ;
      RECT 57.875 3.935 58.17 4.185 ;
      RECT 57.875 3.952 58.175 3.983 ;
      RECT 57.89 3.904 58.121 4.205 ;
      RECT 57.945 3.903 58.121 4.205 ;
      RECT 57.945 3.9 58.035 4.205 ;
      RECT 57.945 3.897 58.031 4.205 ;
      RECT 57.635 4.17 57.64 4.183 ;
      RECT 57.63 4.137 57.635 4.188 ;
      RECT 57.625 4.092 57.63 4.195 ;
      RECT 57.62 4.047 57.625 4.203 ;
      RECT 57.615 4.015 57.62 4.211 ;
      RECT 57.61 3.975 57.615 4.212 ;
      RECT 57.595 3.955 57.61 4.214 ;
      RECT 57.52 3.937 57.595 4.226 ;
      RECT 57.51 3.93 57.52 4.237 ;
      RECT 57.505 3.93 57.51 4.239 ;
      RECT 57.475 3.936 57.505 4.243 ;
      RECT 57.435 3.949 57.475 4.243 ;
      RECT 57.41 3.96 57.435 4.229 ;
      RECT 57.395 3.966 57.41 4.212 ;
      RECT 57.385 3.968 57.395 4.203 ;
      RECT 57.38 3.969 57.385 4.198 ;
      RECT 57.375 3.97 57.38 4.193 ;
      RECT 57.37 3.971 57.375 4.19 ;
      RECT 57.345 3.976 57.37 4.18 ;
      RECT 57.335 3.992 57.345 4.167 ;
      RECT 57.33 4.012 57.335 4.162 ;
      RECT 57.34 3.405 57.345 3.601 ;
      RECT 57.325 3.369 57.34 3.603 ;
      RECT 57.315 3.351 57.325 3.608 ;
      RECT 57.305 3.337 57.315 3.612 ;
      RECT 57.26 3.321 57.305 3.622 ;
      RECT 57.255 3.311 57.26 3.631 ;
      RECT 57.21 3.3 57.255 3.637 ;
      RECT 57.205 3.288 57.21 3.644 ;
      RECT 57.19 3.283 57.205 3.648 ;
      RECT 57.175 3.275 57.19 3.653 ;
      RECT 57.165 3.268 57.175 3.658 ;
      RECT 57.155 3.265 57.165 3.663 ;
      RECT 57.145 3.265 57.155 3.664 ;
      RECT 57.14 3.262 57.145 3.663 ;
      RECT 57.105 3.257 57.13 3.662 ;
      RECT 57.081 3.253 57.105 3.661 ;
      RECT 56.995 3.244 57.081 3.658 ;
      RECT 56.98 3.236 56.995 3.655 ;
      RECT 56.958 3.235 56.98 3.654 ;
      RECT 56.872 3.235 56.958 3.652 ;
      RECT 56.786 3.235 56.872 3.65 ;
      RECT 56.7 3.235 56.786 3.647 ;
      RECT 56.69 3.235 56.7 3.638 ;
      RECT 56.66 3.235 56.69 3.598 ;
      RECT 56.65 3.245 56.66 3.553 ;
      RECT 56.645 3.285 56.65 3.538 ;
      RECT 56.64 3.3 56.645 3.525 ;
      RECT 56.61 3.38 56.64 3.487 ;
      RECT 57.13 3.26 57.14 3.663 ;
      RECT 56.955 4.025 56.97 4.63 ;
      RECT 56.96 4.02 56.97 4.63 ;
      RECT 57.125 4.02 57.13 4.203 ;
      RECT 57.115 4.02 57.125 4.233 ;
      RECT 57.1 4.02 57.115 4.293 ;
      RECT 57.095 4.02 57.1 4.338 ;
      RECT 57.09 4.02 57.095 4.368 ;
      RECT 57.085 4.02 57.09 4.388 ;
      RECT 57.075 4.02 57.085 4.423 ;
      RECT 57.06 4.02 57.075 4.455 ;
      RECT 57.015 4.02 57.06 4.483 ;
      RECT 57.01 4.02 57.015 4.513 ;
      RECT 57.005 4.02 57.01 4.525 ;
      RECT 57 4.02 57.005 4.533 ;
      RECT 56.99 4.02 57 4.548 ;
      RECT 56.985 4.02 56.99 4.57 ;
      RECT 56.975 4.02 56.985 4.593 ;
      RECT 56.97 4.02 56.975 4.613 ;
      RECT 56.935 4.035 56.955 4.63 ;
      RECT 56.91 4.052 56.935 4.63 ;
      RECT 56.905 4.062 56.91 4.63 ;
      RECT 56.875 4.077 56.905 4.63 ;
      RECT 56.8 4.119 56.875 4.63 ;
      RECT 56.795 4.15 56.8 4.613 ;
      RECT 56.79 4.154 56.795 4.595 ;
      RECT 56.785 4.158 56.79 4.558 ;
      RECT 56.78 4.342 56.785 4.525 ;
      RECT 56.265 4.531 56.351 5.096 ;
      RECT 56.22 4.533 56.385 5.09 ;
      RECT 56.351 4.53 56.385 5.09 ;
      RECT 56.265 4.532 56.47 5.084 ;
      RECT 56.22 4.542 56.48 5.08 ;
      RECT 56.195 4.534 56.47 5.076 ;
      RECT 56.19 4.537 56.47 5.071 ;
      RECT 56.165 4.552 56.48 5.065 ;
      RECT 56.165 4.577 56.52 5.06 ;
      RECT 56.125 4.585 56.52 5.035 ;
      RECT 56.125 4.612 56.535 5.033 ;
      RECT 56.125 4.642 56.545 5.02 ;
      RECT 56.12 4.787 56.545 5.008 ;
      RECT 56.125 4.716 56.565 5.005 ;
      RECT 56.125 4.773 56.57 4.813 ;
      RECT 56.315 4.052 56.485 4.23 ;
      RECT 56.265 3.991 56.315 4.215 ;
      RECT 56 3.971 56.265 4.2 ;
      RECT 55.96 4.035 56.435 4.2 ;
      RECT 55.96 4.025 56.39 4.2 ;
      RECT 55.96 4.022 56.38 4.2 ;
      RECT 55.96 4.01 56.37 4.2 ;
      RECT 55.96 3.995 56.315 4.2 ;
      RECT 56 3.967 56.201 4.2 ;
      RECT 56.01 3.945 56.201 4.2 ;
      RECT 56.035 3.93 56.115 4.2 ;
      RECT 55.79 4.46 55.91 4.905 ;
      RECT 55.775 4.46 55.91 4.904 ;
      RECT 55.73 4.482 55.91 4.899 ;
      RECT 55.69 4.531 55.91 4.893 ;
      RECT 55.69 4.531 55.915 4.868 ;
      RECT 55.69 4.531 55.935 4.758 ;
      RECT 55.685 4.561 55.935 4.755 ;
      RECT 55.775 4.46 55.945 4.65 ;
      RECT 55.435 3.245 55.44 3.69 ;
      RECT 55.245 3.245 55.265 3.655 ;
      RECT 55.215 3.245 55.22 3.63 ;
      RECT 55.895 3.552 55.91 3.74 ;
      RECT 55.89 3.537 55.895 3.746 ;
      RECT 55.87 3.51 55.89 3.749 ;
      RECT 55.82 3.477 55.87 3.758 ;
      RECT 55.79 3.457 55.82 3.762 ;
      RECT 55.771 3.445 55.79 3.758 ;
      RECT 55.685 3.417 55.771 3.748 ;
      RECT 55.675 3.392 55.685 3.738 ;
      RECT 55.605 3.36 55.675 3.73 ;
      RECT 55.58 3.32 55.605 3.722 ;
      RECT 55.56 3.302 55.58 3.716 ;
      RECT 55.55 3.292 55.56 3.713 ;
      RECT 55.54 3.285 55.55 3.711 ;
      RECT 55.52 3.272 55.54 3.708 ;
      RECT 55.51 3.262 55.52 3.705 ;
      RECT 55.5 3.255 55.51 3.703 ;
      RECT 55.45 3.247 55.5 3.697 ;
      RECT 55.44 3.245 55.45 3.691 ;
      RECT 55.41 3.245 55.435 3.688 ;
      RECT 55.381 3.245 55.41 3.683 ;
      RECT 55.295 3.245 55.381 3.673 ;
      RECT 55.265 3.245 55.295 3.66 ;
      RECT 55.22 3.245 55.245 3.643 ;
      RECT 55.205 3.245 55.215 3.625 ;
      RECT 55.185 3.252 55.205 3.61 ;
      RECT 55.18 3.267 55.185 3.598 ;
      RECT 55.175 3.272 55.18 3.538 ;
      RECT 55.17 3.277 55.175 3.38 ;
      RECT 55.165 3.28 55.17 3.298 ;
      RECT 55.43 3.965 55.516 4.286 ;
      RECT 55.43 3.965 55.55 4.279 ;
      RECT 55.38 3.965 55.55 4.275 ;
      RECT 55.38 3.967 55.636 4.273 ;
      RECT 55.38 3.969 55.66 4.267 ;
      RECT 55.38 3.976 55.67 4.266 ;
      RECT 55.38 3.985 55.675 4.263 ;
      RECT 55.38 3.991 55.68 4.258 ;
      RECT 55.38 4.035 55.685 4.255 ;
      RECT 55.38 4.127 55.69 4.252 ;
      RECT 54.905 4.57 54.94 4.89 ;
      RECT 55.49 4.755 55.495 4.937 ;
      RECT 55.445 4.637 55.49 4.956 ;
      RECT 55.43 4.614 55.445 4.979 ;
      RECT 55.42 4.604 55.43 4.989 ;
      RECT 55.4 4.599 55.42 5.002 ;
      RECT 55.375 4.597 55.4 5.023 ;
      RECT 55.356 4.596 55.375 5.035 ;
      RECT 55.27 4.593 55.356 5.035 ;
      RECT 55.2 4.588 55.27 5.023 ;
      RECT 55.125 4.584 55.2 4.998 ;
      RECT 55.06 4.58 55.125 4.965 ;
      RECT 54.99 4.577 55.06 4.925 ;
      RECT 54.96 4.573 54.99 4.9 ;
      RECT 54.94 4.571 54.96 4.893 ;
      RECT 54.856 4.569 54.905 4.891 ;
      RECT 54.77 4.566 54.856 4.892 ;
      RECT 54.695 4.565 54.77 4.894 ;
      RECT 54.61 4.565 54.695 4.92 ;
      RECT 54.533 4.566 54.61 4.945 ;
      RECT 54.447 4.567 54.533 4.945 ;
      RECT 54.361 4.567 54.447 4.945 ;
      RECT 54.275 4.568 54.361 4.945 ;
      RECT 54.255 4.569 54.275 4.937 ;
      RECT 54.24 4.575 54.255 4.922 ;
      RECT 54.205 4.595 54.24 4.902 ;
      RECT 54.195 4.615 54.205 4.884 ;
      RECT 55.165 3.92 55.17 4.19 ;
      RECT 55.16 3.911 55.165 4.195 ;
      RECT 55.15 3.901 55.16 4.207 ;
      RECT 55.145 3.89 55.15 4.218 ;
      RECT 55.125 3.884 55.145 4.236 ;
      RECT 55.08 3.881 55.125 4.285 ;
      RECT 55.065 3.88 55.08 4.33 ;
      RECT 55.06 3.88 55.065 4.343 ;
      RECT 55.05 3.88 55.06 4.355 ;
      RECT 55.045 3.881 55.05 4.37 ;
      RECT 55.025 3.889 55.045 4.375 ;
      RECT 54.995 3.905 55.025 4.375 ;
      RECT 54.985 3.917 54.99 4.375 ;
      RECT 54.95 3.932 54.985 4.375 ;
      RECT 54.92 3.952 54.95 4.375 ;
      RECT 54.91 3.977 54.92 4.375 ;
      RECT 54.905 4.005 54.91 4.375 ;
      RECT 54.9 4.035 54.905 4.375 ;
      RECT 54.895 4.052 54.9 4.375 ;
      RECT 54.885 4.08 54.895 4.375 ;
      RECT 54.875 4.115 54.885 4.375 ;
      RECT 54.87 4.15 54.875 4.375 ;
      RECT 54.99 3.915 54.995 4.375 ;
      RECT 54.505 4.017 54.69 4.19 ;
      RECT 54.465 3.935 54.65 4.188 ;
      RECT 54.426 3.94 54.65 4.184 ;
      RECT 54.34 3.949 54.65 4.179 ;
      RECT 54.256 3.965 54.655 4.174 ;
      RECT 54.17 3.985 54.68 4.168 ;
      RECT 54.17 4.005 54.685 4.168 ;
      RECT 54.256 3.975 54.68 4.174 ;
      RECT 54.34 3.95 54.655 4.179 ;
      RECT 54.505 3.932 54.65 4.19 ;
      RECT 54.505 3.927 54.605 4.19 ;
      RECT 54.591 3.921 54.605 4.19 ;
      RECT 53.98 3.245 53.985 3.644 ;
      RECT 53.725 3.245 53.76 3.642 ;
      RECT 53.32 3.28 53.325 3.636 ;
      RECT 54.065 3.283 54.07 3.538 ;
      RECT 54.06 3.281 54.065 3.544 ;
      RECT 54.055 3.28 54.06 3.551 ;
      RECT 54.03 3.273 54.055 3.575 ;
      RECT 54.025 3.266 54.03 3.599 ;
      RECT 54.02 3.262 54.025 3.608 ;
      RECT 54.01 3.257 54.02 3.621 ;
      RECT 54.005 3.254 54.01 3.63 ;
      RECT 54 3.252 54.005 3.635 ;
      RECT 53.985 3.248 54 3.645 ;
      RECT 53.97 3.242 53.98 3.644 ;
      RECT 53.932 3.24 53.97 3.644 ;
      RECT 53.846 3.242 53.932 3.644 ;
      RECT 53.76 3.244 53.846 3.643 ;
      RECT 53.689 3.245 53.725 3.642 ;
      RECT 53.603 3.247 53.689 3.642 ;
      RECT 53.517 3.249 53.603 3.641 ;
      RECT 53.431 3.251 53.517 3.641 ;
      RECT 53.345 3.254 53.431 3.64 ;
      RECT 53.335 3.26 53.345 3.639 ;
      RECT 53.325 3.272 53.335 3.637 ;
      RECT 53.265 3.307 53.32 3.633 ;
      RECT 53.26 3.337 53.265 3.395 ;
      RECT 54.005 4.417 54.02 4.61 ;
      RECT 54 4.385 54.005 4.61 ;
      RECT 53.99 4.36 54 4.61 ;
      RECT 53.985 4.332 53.99 4.61 ;
      RECT 53.955 4.255 53.985 4.61 ;
      RECT 53.93 4.137 53.955 4.61 ;
      RECT 53.925 4.075 53.93 4.61 ;
      RECT 53.915 4.062 53.925 4.61 ;
      RECT 53.895 4.052 53.915 4.61 ;
      RECT 53.88 4.035 53.895 4.61 ;
      RECT 53.85 4.023 53.88 4.61 ;
      RECT 53.845 4.022 53.85 4.555 ;
      RECT 53.84 4.022 53.845 4.513 ;
      RECT 53.825 4.021 53.84 4.465 ;
      RECT 53.81 4.021 53.825 4.403 ;
      RECT 53.79 4.021 53.81 4.363 ;
      RECT 53.785 4.021 53.79 4.348 ;
      RECT 53.76 4.02 53.785 4.343 ;
      RECT 53.69 4.019 53.76 4.33 ;
      RECT 53.675 4.018 53.69 4.315 ;
      RECT 53.645 4.017 53.675 4.298 ;
      RECT 53.64 4.017 53.645 4.283 ;
      RECT 53.59 4.016 53.64 4.263 ;
      RECT 53.525 4.015 53.59 4.218 ;
      RECT 53.52 4.015 53.525 4.19 ;
      RECT 53.605 4.552 53.61 4.809 ;
      RECT 53.585 4.471 53.605 4.826 ;
      RECT 53.565 4.465 53.585 4.855 ;
      RECT 53.505 4.452 53.565 4.875 ;
      RECT 53.46 4.436 53.505 4.876 ;
      RECT 53.376 4.424 53.46 4.864 ;
      RECT 53.29 4.411 53.376 4.848 ;
      RECT 53.28 4.404 53.29 4.84 ;
      RECT 53.235 4.401 53.28 4.78 ;
      RECT 53.215 4.397 53.235 4.695 ;
      RECT 53.2 4.395 53.215 4.648 ;
      RECT 53.17 4.392 53.2 4.618 ;
      RECT 53.135 4.388 53.17 4.595 ;
      RECT 53.092 4.383 53.135 4.583 ;
      RECT 53.006 4.374 53.092 4.592 ;
      RECT 52.92 4.363 53.006 4.604 ;
      RECT 52.855 4.354 52.92 4.613 ;
      RECT 52.835 4.345 52.855 4.618 ;
      RECT 52.83 4.338 52.835 4.62 ;
      RECT 52.79 4.323 52.83 4.617 ;
      RECT 52.77 4.302 52.79 4.612 ;
      RECT 52.755 4.29 52.77 4.605 ;
      RECT 52.75 4.282 52.755 4.598 ;
      RECT 52.735 4.262 52.75 4.591 ;
      RECT 52.73 4.125 52.735 4.585 ;
      RECT 52.65 4.014 52.73 4.557 ;
      RECT 52.641 4.007 52.65 4.523 ;
      RECT 52.555 4.001 52.641 4.448 ;
      RECT 52.53 3.992 52.555 4.36 ;
      RECT 52.5 3.987 52.53 4.335 ;
      RECT 52.435 3.996 52.5 4.32 ;
      RECT 52.415 4.012 52.435 4.295 ;
      RECT 52.405 4.018 52.415 4.243 ;
      RECT 52.385 4.04 52.405 4.125 ;
      RECT 53.04 4.005 53.21 4.19 ;
      RECT 53.04 4.005 53.245 4.188 ;
      RECT 53.09 3.915 53.26 4.179 ;
      RECT 53.04 4.072 53.265 4.172 ;
      RECT 53.055 3.95 53.26 4.179 ;
      RECT 52.255 4.683 52.32 5.126 ;
      RECT 52.195 4.708 52.32 5.124 ;
      RECT 52.195 4.708 52.375 5.118 ;
      RECT 52.18 4.733 52.375 5.117 ;
      RECT 52.32 4.67 52.395 5.114 ;
      RECT 52.255 4.695 52.475 5.108 ;
      RECT 52.18 4.734 52.52 5.102 ;
      RECT 52.165 4.761 52.52 5.093 ;
      RECT 52.18 4.754 52.54 5.085 ;
      RECT 52.165 4.763 52.545 5.068 ;
      RECT 52.16 4.78 52.545 4.895 ;
      RECT 52.165 3.502 52.2 3.74 ;
      RECT 52.165 3.502 52.23 3.739 ;
      RECT 52.165 3.502 52.345 3.735 ;
      RECT 52.165 3.502 52.4 3.713 ;
      RECT 52.175 3.445 52.455 3.613 ;
      RECT 52.28 3.285 52.31 3.736 ;
      RECT 52.31 3.28 52.49 3.493 ;
      RECT 52.18 3.421 52.49 3.493 ;
      RECT 52.23 3.317 52.28 3.737 ;
      RECT 52.2 3.373 52.49 3.493 ;
      RECT 50.7 3.035 50.87 4.225 ;
      RECT 50.7 3.035 51.17 3.205 ;
      RECT 50.7 9.405 51.17 9.575 ;
      RECT 50.7 8.385 50.87 9.575 ;
      RECT 49.71 3.035 49.88 4.225 ;
      RECT 49.71 3.035 50.18 3.205 ;
      RECT 49.71 9.405 50.18 9.575 ;
      RECT 49.71 8.385 49.88 9.575 ;
      RECT 47.86 3.93 48.03 5.16 ;
      RECT 47.915 2.15 48.085 4.1 ;
      RECT 47.86 1.87 48.03 2.32 ;
      RECT 47.86 10.29 48.03 10.74 ;
      RECT 47.915 8.51 48.085 10.46 ;
      RECT 47.86 7.45 48.03 8.68 ;
      RECT 47.34 1.87 47.51 5.16 ;
      RECT 47.34 3.37 47.745 3.7 ;
      RECT 47.34 2.53 47.745 2.86 ;
      RECT 47.34 7.45 47.51 10.74 ;
      RECT 47.34 9.75 47.745 10.08 ;
      RECT 47.34 8.91 47.745 9.24 ;
      RECT 45.44 4.687 45.455 4.738 ;
      RECT 45.435 4.667 45.44 4.785 ;
      RECT 45.42 4.657 45.435 4.853 ;
      RECT 45.395 4.637 45.42 4.908 ;
      RECT 45.355 4.622 45.395 4.928 ;
      RECT 45.31 4.616 45.355 4.956 ;
      RECT 45.24 4.606 45.31 4.973 ;
      RECT 45.22 4.598 45.24 4.973 ;
      RECT 45.16 4.592 45.22 4.965 ;
      RECT 45.101 4.583 45.16 4.953 ;
      RECT 45.015 4.572 45.101 4.936 ;
      RECT 44.993 4.563 45.015 4.924 ;
      RECT 44.907 4.556 44.993 4.911 ;
      RECT 44.821 4.543 44.907 4.892 ;
      RECT 44.735 4.531 44.821 4.872 ;
      RECT 44.705 4.52 44.735 4.859 ;
      RECT 44.655 4.506 44.705 4.851 ;
      RECT 44.635 4.495 44.655 4.843 ;
      RECT 44.586 4.484 44.635 4.835 ;
      RECT 44.5 4.463 44.586 4.82 ;
      RECT 44.455 4.45 44.5 4.805 ;
      RECT 44.41 4.45 44.455 4.785 ;
      RECT 44.355 4.45 44.41 4.72 ;
      RECT 44.33 4.45 44.355 4.643 ;
      RECT 44.855 4.187 45.025 4.37 ;
      RECT 44.855 4.187 45.04 4.328 ;
      RECT 44.855 4.187 45.045 4.27 ;
      RECT 44.915 3.955 45.05 4.246 ;
      RECT 44.915 3.959 45.055 4.229 ;
      RECT 44.86 4.122 45.055 4.229 ;
      RECT 44.885 3.967 45.025 4.37 ;
      RECT 44.885 3.971 45.065 4.17 ;
      RECT 44.87 4.057 45.065 4.17 ;
      RECT 44.88 3.987 45.025 4.37 ;
      RECT 44.88 3.99 45.075 4.083 ;
      RECT 44.875 4.007 45.075 4.083 ;
      RECT 44.645 3.227 44.815 3.71 ;
      RECT 44.64 3.222 44.79 3.7 ;
      RECT 44.64 3.229 44.82 3.694 ;
      RECT 44.63 3.223 44.79 3.673 ;
      RECT 44.63 3.239 44.835 3.632 ;
      RECT 44.6 3.224 44.79 3.595 ;
      RECT 44.6 3.254 44.845 3.535 ;
      RECT 44.595 3.226 44.79 3.533 ;
      RECT 44.575 3.235 44.82 3.49 ;
      RECT 44.55 3.251 44.835 3.402 ;
      RECT 44.55 3.27 44.86 3.393 ;
      RECT 44.545 3.307 44.86 3.345 ;
      RECT 44.55 3.287 44.865 3.313 ;
      RECT 44.645 3.221 44.755 3.71 ;
      RECT 44.731 3.22 44.755 3.71 ;
      RECT 43.965 4.005 43.97 4.216 ;
      RECT 44.565 4.005 44.57 4.19 ;
      RECT 44.63 4.045 44.635 4.158 ;
      RECT 44.625 4.037 44.63 4.164 ;
      RECT 44.62 4.027 44.625 4.172 ;
      RECT 44.615 4.017 44.62 4.181 ;
      RECT 44.61 4.007 44.615 4.185 ;
      RECT 44.57 4.005 44.61 4.188 ;
      RECT 44.542 4.004 44.565 4.192 ;
      RECT 44.456 4.001 44.542 4.199 ;
      RECT 44.37 3.997 44.456 4.21 ;
      RECT 44.35 3.995 44.37 4.216 ;
      RECT 44.332 3.994 44.35 4.219 ;
      RECT 44.246 3.992 44.332 4.226 ;
      RECT 44.16 3.987 44.246 4.239 ;
      RECT 44.141 3.984 44.16 4.244 ;
      RECT 44.055 3.982 44.141 4.235 ;
      RECT 44.045 3.982 44.055 4.228 ;
      RECT 43.97 3.995 44.045 4.222 ;
      RECT 43.955 4.006 43.965 4.216 ;
      RECT 43.945 4.008 43.955 4.215 ;
      RECT 43.935 4.012 43.945 4.211 ;
      RECT 43.93 4.015 43.935 4.205 ;
      RECT 43.92 4.017 43.93 4.199 ;
      RECT 43.915 4.02 43.92 4.193 ;
      RECT 43.895 4.606 43.9 4.81 ;
      RECT 43.88 4.593 43.895 4.903 ;
      RECT 43.865 4.574 43.88 5.18 ;
      RECT 43.83 4.54 43.865 5.18 ;
      RECT 43.826 4.51 43.83 5.18 ;
      RECT 43.74 4.392 43.826 5.18 ;
      RECT 43.73 4.267 43.74 5.18 ;
      RECT 43.715 4.235 43.73 5.18 ;
      RECT 43.71 4.21 43.715 5.18 ;
      RECT 43.705 4.2 43.71 5.136 ;
      RECT 43.69 4.172 43.705 5.041 ;
      RECT 43.675 4.138 43.69 4.94 ;
      RECT 43.67 4.116 43.675 4.893 ;
      RECT 43.665 4.105 43.67 4.863 ;
      RECT 43.66 4.095 43.665 4.829 ;
      RECT 43.65 4.082 43.66 4.797 ;
      RECT 43.625 4.058 43.65 4.723 ;
      RECT 43.62 4.038 43.625 4.648 ;
      RECT 43.615 4.032 43.62 4.623 ;
      RECT 43.61 4.027 43.615 4.588 ;
      RECT 43.605 4.022 43.61 4.563 ;
      RECT 43.6 4.02 43.605 4.543 ;
      RECT 43.595 4.02 43.6 4.528 ;
      RECT 43.59 4.02 43.595 4.488 ;
      RECT 43.58 4.02 43.59 4.46 ;
      RECT 43.57 4.02 43.58 4.405 ;
      RECT 43.555 4.02 43.57 4.343 ;
      RECT 43.55 4.019 43.555 4.288 ;
      RECT 43.535 4.018 43.55 4.268 ;
      RECT 43.475 4.016 43.535 4.242 ;
      RECT 43.44 4.017 43.475 4.222 ;
      RECT 43.435 4.019 43.44 4.212 ;
      RECT 43.425 4.038 43.435 4.202 ;
      RECT 43.42 4.065 43.425 4.133 ;
      RECT 43.535 3.49 43.705 3.735 ;
      RECT 43.57 3.261 43.705 3.735 ;
      RECT 43.57 3.263 43.715 3.73 ;
      RECT 43.57 3.265 43.74 3.718 ;
      RECT 43.57 3.268 43.765 3.7 ;
      RECT 43.57 3.273 43.815 3.673 ;
      RECT 43.57 3.278 43.835 3.638 ;
      RECT 43.55 3.28 43.845 3.613 ;
      RECT 43.54 3.375 43.845 3.613 ;
      RECT 43.57 3.26 43.68 3.735 ;
      RECT 43.58 3.257 43.675 3.735 ;
      RECT 43.1 4.522 43.29 4.88 ;
      RECT 43.1 4.534 43.325 4.879 ;
      RECT 43.1 4.562 43.345 4.877 ;
      RECT 43.1 4.587 43.35 4.876 ;
      RECT 43.1 4.645 43.365 4.875 ;
      RECT 43.085 4.518 43.245 4.86 ;
      RECT 43.065 4.527 43.29 4.813 ;
      RECT 43.04 4.538 43.325 4.75 ;
      RECT 43.04 4.622 43.36 4.75 ;
      RECT 43.04 4.597 43.355 4.75 ;
      RECT 43.1 4.513 43.245 4.88 ;
      RECT 43.186 4.512 43.245 4.88 ;
      RECT 43.186 4.511 43.23 4.88 ;
      RECT 42.58 7.45 42.75 10.74 ;
      RECT 42.58 9.75 42.985 10.08 ;
      RECT 42.58 8.91 42.985 9.24 ;
      RECT 42.885 4.027 42.89 4.405 ;
      RECT 42.88 3.995 42.885 4.405 ;
      RECT 42.875 3.967 42.88 4.405 ;
      RECT 42.87 3.947 42.875 4.405 ;
      RECT 42.815 3.93 42.87 4.405 ;
      RECT 42.775 3.915 42.815 4.405 ;
      RECT 42.72 3.902 42.775 4.405 ;
      RECT 42.685 3.893 42.72 4.405 ;
      RECT 42.681 3.891 42.685 4.404 ;
      RECT 42.595 3.887 42.681 4.387 ;
      RECT 42.51 3.879 42.595 4.35 ;
      RECT 42.5 3.875 42.51 4.323 ;
      RECT 42.49 3.875 42.5 4.305 ;
      RECT 42.48 3.877 42.49 4.288 ;
      RECT 42.475 3.882 42.48 4.274 ;
      RECT 42.47 3.886 42.475 4.261 ;
      RECT 42.46 3.891 42.47 4.245 ;
      RECT 42.445 3.905 42.46 4.22 ;
      RECT 42.44 3.911 42.445 4.2 ;
      RECT 42.435 3.913 42.44 4.193 ;
      RECT 42.43 3.917 42.435 4.068 ;
      RECT 42.61 4.717 42.855 5.18 ;
      RECT 42.53 4.69 42.85 5.176 ;
      RECT 42.46 4.725 42.855 5.169 ;
      RECT 42.25 4.98 42.855 5.165 ;
      RECT 42.43 4.748 42.855 5.165 ;
      RECT 42.27 4.94 42.855 5.165 ;
      RECT 42.42 4.76 42.855 5.165 ;
      RECT 42.305 4.877 42.855 5.165 ;
      RECT 42.36 4.802 42.855 5.165 ;
      RECT 42.61 4.667 42.85 5.18 ;
      RECT 42.64 4.66 42.85 5.18 ;
      RECT 42.63 4.662 42.85 5.18 ;
      RECT 42.64 4.657 42.77 5.18 ;
      RECT 42.195 3.22 42.281 3.659 ;
      RECT 42.19 3.22 42.281 3.657 ;
      RECT 42.19 3.22 42.35 3.656 ;
      RECT 42.19 3.22 42.38 3.653 ;
      RECT 42.175 3.227 42.38 3.644 ;
      RECT 42.175 3.227 42.385 3.64 ;
      RECT 42.17 3.237 42.385 3.633 ;
      RECT 42.165 3.242 42.385 3.608 ;
      RECT 42.165 3.242 42.4 3.59 ;
      RECT 42.19 3.22 42.42 3.505 ;
      RECT 42.16 3.247 42.42 3.503 ;
      RECT 42.17 3.24 42.425 3.441 ;
      RECT 42.16 3.362 42.43 3.424 ;
      RECT 42.145 3.257 42.425 3.375 ;
      RECT 42.14 3.267 42.425 3.275 ;
      RECT 42.22 4.038 42.225 4.115 ;
      RECT 42.21 4.032 42.22 4.305 ;
      RECT 42.2 4.024 42.21 4.326 ;
      RECT 42.19 4.015 42.2 4.348 ;
      RECT 42.185 4.01 42.19 4.365 ;
      RECT 42.145 4.01 42.185 4.405 ;
      RECT 42.125 4.01 42.145 4.46 ;
      RECT 42.12 4.01 42.125 4.488 ;
      RECT 42.11 4.01 42.12 4.503 ;
      RECT 42.075 4.01 42.11 4.545 ;
      RECT 42.07 4.01 42.075 4.588 ;
      RECT 42.06 4.01 42.07 4.603 ;
      RECT 42.045 4.01 42.06 4.623 ;
      RECT 42.03 4.01 42.045 4.65 ;
      RECT 42.025 4.011 42.03 4.668 ;
      RECT 42.005 4.012 42.025 4.675 ;
      RECT 41.95 4.013 42.005 4.695 ;
      RECT 41.94 4.014 41.95 4.709 ;
      RECT 41.935 4.017 41.94 4.708 ;
      RECT 41.895 4.09 41.935 4.706 ;
      RECT 41.88 4.17 41.895 4.704 ;
      RECT 41.855 4.225 41.88 4.702 ;
      RECT 41.84 4.29 41.855 4.701 ;
      RECT 41.795 4.322 41.84 4.698 ;
      RECT 41.71 4.345 41.795 4.693 ;
      RECT 41.685 4.365 41.71 4.688 ;
      RECT 41.615 4.37 41.685 4.684 ;
      RECT 41.595 4.372 41.615 4.681 ;
      RECT 41.51 4.383 41.595 4.675 ;
      RECT 41.505 4.394 41.51 4.67 ;
      RECT 41.495 4.396 41.505 4.67 ;
      RECT 41.46 4.4 41.495 4.668 ;
      RECT 41.41 4.41 41.46 4.655 ;
      RECT 41.39 4.418 41.41 4.64 ;
      RECT 41.31 4.43 41.39 4.623 ;
      RECT 41.475 3.98 41.645 4.19 ;
      RECT 41.591 3.976 41.645 4.19 ;
      RECT 41.396 3.98 41.645 4.181 ;
      RECT 41.396 3.98 41.65 4.17 ;
      RECT 41.31 3.98 41.65 4.161 ;
      RECT 41.31 3.988 41.66 4.105 ;
      RECT 41.31 4 41.665 4.018 ;
      RECT 41.31 4.007 41.67 4.01 ;
      RECT 41.505 3.978 41.645 4.19 ;
      RECT 41.26 4.923 41.505 5.255 ;
      RECT 41.255 4.915 41.26 5.252 ;
      RECT 41.225 4.935 41.505 5.233 ;
      RECT 41.205 4.967 41.505 5.206 ;
      RECT 41.255 4.92 41.432 5.252 ;
      RECT 41.255 4.917 41.346 5.252 ;
      RECT 41.195 3.265 41.365 3.685 ;
      RECT 41.19 3.265 41.365 3.683 ;
      RECT 41.19 3.265 41.39 3.673 ;
      RECT 41.19 3.265 41.41 3.648 ;
      RECT 41.185 3.265 41.41 3.643 ;
      RECT 41.185 3.265 41.42 3.633 ;
      RECT 41.185 3.265 41.425 3.628 ;
      RECT 41.185 3.27 41.43 3.623 ;
      RECT 41.185 3.302 41.445 3.613 ;
      RECT 41.185 3.372 41.47 3.596 ;
      RECT 41.165 3.372 41.47 3.588 ;
      RECT 41.165 3.432 41.48 3.565 ;
      RECT 41.165 3.472 41.49 3.51 ;
      RECT 41.15 3.265 41.425 3.49 ;
      RECT 41.14 3.28 41.43 3.388 ;
      RECT 40.73 4.67 40.9 5.195 ;
      RECT 40.725 4.67 40.9 5.188 ;
      RECT 40.715 4.67 40.905 5.153 ;
      RECT 40.71 4.68 40.905 5.125 ;
      RECT 40.705 4.7 40.905 5.108 ;
      RECT 40.715 4.675 40.91 5.098 ;
      RECT 40.7 4.72 40.91 5.09 ;
      RECT 40.695 4.74 40.91 5.075 ;
      RECT 40.69 4.77 40.91 5.065 ;
      RECT 40.68 4.815 40.91 5.04 ;
      RECT 40.71 4.685 40.915 5.023 ;
      RECT 40.675 4.867 40.915 5.018 ;
      RECT 40.71 4.695 40.92 4.988 ;
      RECT 40.67 4.9 40.92 4.985 ;
      RECT 40.665 4.925 40.92 4.965 ;
      RECT 40.705 4.712 40.93 4.905 ;
      RECT 40.7 4.734 40.94 4.798 ;
      RECT 40.65 3.981 40.665 4.25 ;
      RECT 40.605 3.965 40.65 4.295 ;
      RECT 40.6 3.953 40.605 4.345 ;
      RECT 40.59 3.949 40.6 4.378 ;
      RECT 40.585 3.946 40.59 4.406 ;
      RECT 40.57 3.948 40.585 4.448 ;
      RECT 40.565 3.952 40.57 4.488 ;
      RECT 40.545 3.957 40.565 4.54 ;
      RECT 40.541 3.962 40.545 4.597 ;
      RECT 40.455 3.981 40.541 4.634 ;
      RECT 40.445 4.002 40.455 4.67 ;
      RECT 40.44 4.01 40.445 4.671 ;
      RECT 40.435 4.052 40.44 4.672 ;
      RECT 40.42 4.14 40.435 4.673 ;
      RECT 40.41 4.29 40.42 4.675 ;
      RECT 40.405 4.335 40.41 4.677 ;
      RECT 40.37 4.377 40.405 4.68 ;
      RECT 40.365 4.395 40.37 4.683 ;
      RECT 40.288 4.401 40.365 4.689 ;
      RECT 40.202 4.415 40.288 4.702 ;
      RECT 40.116 4.429 40.202 4.716 ;
      RECT 40.03 4.443 40.116 4.729 ;
      RECT 39.97 4.455 40.03 4.741 ;
      RECT 39.945 4.462 39.97 4.748 ;
      RECT 39.931 4.465 39.945 4.753 ;
      RECT 39.845 4.473 39.931 4.769 ;
      RECT 39.84 4.48 39.845 4.784 ;
      RECT 39.816 4.48 39.84 4.791 ;
      RECT 39.73 4.483 39.816 4.819 ;
      RECT 39.645 4.487 39.73 4.863 ;
      RECT 39.58 4.491 39.645 4.9 ;
      RECT 39.555 4.494 39.58 4.916 ;
      RECT 39.48 4.507 39.555 4.92 ;
      RECT 39.455 4.525 39.48 4.924 ;
      RECT 39.445 4.532 39.455 4.926 ;
      RECT 39.43 4.535 39.445 4.927 ;
      RECT 39.37 4.547 39.43 4.931 ;
      RECT 39.36 4.561 39.37 4.935 ;
      RECT 39.305 4.571 39.36 4.923 ;
      RECT 39.28 4.592 39.305 4.906 ;
      RECT 39.26 4.612 39.28 4.897 ;
      RECT 39.255 4.625 39.26 4.892 ;
      RECT 39.24 4.637 39.255 4.888 ;
      RECT 40.475 3.292 40.48 3.315 ;
      RECT 40.47 3.283 40.475 3.355 ;
      RECT 40.465 3.281 40.47 3.398 ;
      RECT 40.46 3.272 40.465 3.433 ;
      RECT 40.455 3.262 40.46 3.505 ;
      RECT 40.45 3.252 40.455 3.57 ;
      RECT 40.445 3.249 40.45 3.61 ;
      RECT 40.42 3.243 40.445 3.7 ;
      RECT 40.385 3.231 40.42 3.725 ;
      RECT 40.375 3.222 40.385 3.725 ;
      RECT 40.24 3.22 40.25 3.708 ;
      RECT 40.23 3.22 40.24 3.675 ;
      RECT 40.225 3.22 40.23 3.65 ;
      RECT 40.22 3.22 40.225 3.638 ;
      RECT 40.215 3.22 40.22 3.62 ;
      RECT 40.205 3.22 40.215 3.585 ;
      RECT 40.2 3.222 40.205 3.563 ;
      RECT 40.195 3.228 40.2 3.548 ;
      RECT 40.19 3.234 40.195 3.533 ;
      RECT 40.175 3.246 40.19 3.506 ;
      RECT 40.17 3.257 40.175 3.474 ;
      RECT 40.165 3.267 40.17 3.458 ;
      RECT 40.155 3.275 40.165 3.427 ;
      RECT 40.15 3.285 40.155 3.401 ;
      RECT 40.145 3.342 40.15 3.384 ;
      RECT 40.25 3.22 40.375 3.725 ;
      RECT 39.965 3.907 40.225 4.205 ;
      RECT 39.96 3.914 40.225 4.203 ;
      RECT 39.965 3.909 40.24 4.198 ;
      RECT 39.955 3.922 40.24 4.195 ;
      RECT 39.955 3.927 40.245 4.188 ;
      RECT 39.95 3.935 40.245 4.185 ;
      RECT 39.95 3.952 40.25 3.983 ;
      RECT 39.965 3.904 40.196 4.205 ;
      RECT 40.02 3.903 40.196 4.205 ;
      RECT 40.02 3.9 40.11 4.205 ;
      RECT 40.02 3.897 40.106 4.205 ;
      RECT 39.71 4.17 39.715 4.183 ;
      RECT 39.705 4.137 39.71 4.188 ;
      RECT 39.7 4.092 39.705 4.195 ;
      RECT 39.695 4.047 39.7 4.203 ;
      RECT 39.69 4.015 39.695 4.211 ;
      RECT 39.685 3.975 39.69 4.212 ;
      RECT 39.67 3.955 39.685 4.214 ;
      RECT 39.595 3.937 39.67 4.226 ;
      RECT 39.585 3.93 39.595 4.237 ;
      RECT 39.58 3.93 39.585 4.239 ;
      RECT 39.55 3.936 39.58 4.243 ;
      RECT 39.51 3.949 39.55 4.243 ;
      RECT 39.485 3.96 39.51 4.229 ;
      RECT 39.47 3.966 39.485 4.212 ;
      RECT 39.46 3.968 39.47 4.203 ;
      RECT 39.455 3.969 39.46 4.198 ;
      RECT 39.45 3.97 39.455 4.193 ;
      RECT 39.445 3.971 39.45 4.19 ;
      RECT 39.42 3.976 39.445 4.18 ;
      RECT 39.41 3.992 39.42 4.167 ;
      RECT 39.405 4.012 39.41 4.162 ;
      RECT 39.415 3.405 39.42 3.601 ;
      RECT 39.4 3.369 39.415 3.603 ;
      RECT 39.39 3.351 39.4 3.608 ;
      RECT 39.38 3.337 39.39 3.612 ;
      RECT 39.335 3.321 39.38 3.622 ;
      RECT 39.33 3.311 39.335 3.631 ;
      RECT 39.285 3.3 39.33 3.637 ;
      RECT 39.28 3.288 39.285 3.644 ;
      RECT 39.265 3.283 39.28 3.648 ;
      RECT 39.25 3.275 39.265 3.653 ;
      RECT 39.24 3.268 39.25 3.658 ;
      RECT 39.23 3.265 39.24 3.663 ;
      RECT 39.22 3.265 39.23 3.664 ;
      RECT 39.215 3.262 39.22 3.663 ;
      RECT 39.18 3.257 39.205 3.662 ;
      RECT 39.156 3.253 39.18 3.661 ;
      RECT 39.07 3.244 39.156 3.658 ;
      RECT 39.055 3.236 39.07 3.655 ;
      RECT 39.033 3.235 39.055 3.654 ;
      RECT 38.947 3.235 39.033 3.652 ;
      RECT 38.861 3.235 38.947 3.65 ;
      RECT 38.775 3.235 38.861 3.647 ;
      RECT 38.765 3.235 38.775 3.638 ;
      RECT 38.735 3.235 38.765 3.598 ;
      RECT 38.725 3.245 38.735 3.553 ;
      RECT 38.72 3.285 38.725 3.538 ;
      RECT 38.715 3.3 38.72 3.525 ;
      RECT 38.685 3.38 38.715 3.487 ;
      RECT 39.205 3.26 39.215 3.663 ;
      RECT 39.03 4.025 39.045 4.63 ;
      RECT 39.035 4.02 39.045 4.63 ;
      RECT 39.2 4.02 39.205 4.203 ;
      RECT 39.19 4.02 39.2 4.233 ;
      RECT 39.175 4.02 39.19 4.293 ;
      RECT 39.17 4.02 39.175 4.338 ;
      RECT 39.165 4.02 39.17 4.368 ;
      RECT 39.16 4.02 39.165 4.388 ;
      RECT 39.15 4.02 39.16 4.423 ;
      RECT 39.135 4.02 39.15 4.455 ;
      RECT 39.09 4.02 39.135 4.483 ;
      RECT 39.085 4.02 39.09 4.513 ;
      RECT 39.08 4.02 39.085 4.525 ;
      RECT 39.075 4.02 39.08 4.533 ;
      RECT 39.065 4.02 39.075 4.548 ;
      RECT 39.06 4.02 39.065 4.57 ;
      RECT 39.05 4.02 39.06 4.593 ;
      RECT 39.045 4.02 39.05 4.613 ;
      RECT 39.01 4.035 39.03 4.63 ;
      RECT 38.985 4.052 39.01 4.63 ;
      RECT 38.98 4.062 38.985 4.63 ;
      RECT 38.95 4.077 38.98 4.63 ;
      RECT 38.875 4.119 38.95 4.63 ;
      RECT 38.87 4.15 38.875 4.613 ;
      RECT 38.865 4.154 38.87 4.595 ;
      RECT 38.86 4.158 38.865 4.558 ;
      RECT 38.855 4.342 38.86 4.525 ;
      RECT 38.34 4.531 38.426 5.096 ;
      RECT 38.295 4.533 38.46 5.09 ;
      RECT 38.426 4.53 38.46 5.09 ;
      RECT 38.34 4.532 38.545 5.084 ;
      RECT 38.295 4.542 38.555 5.08 ;
      RECT 38.27 4.534 38.545 5.076 ;
      RECT 38.265 4.537 38.545 5.071 ;
      RECT 38.24 4.552 38.555 5.065 ;
      RECT 38.24 4.577 38.595 5.06 ;
      RECT 38.2 4.585 38.595 5.035 ;
      RECT 38.2 4.612 38.61 5.033 ;
      RECT 38.2 4.642 38.62 5.02 ;
      RECT 38.195 4.787 38.62 5.008 ;
      RECT 38.2 4.716 38.64 5.005 ;
      RECT 38.2 4.773 38.645 4.813 ;
      RECT 38.39 4.052 38.56 4.23 ;
      RECT 38.34 3.991 38.39 4.215 ;
      RECT 38.075 3.971 38.34 4.2 ;
      RECT 38.035 4.035 38.51 4.2 ;
      RECT 38.035 4.025 38.465 4.2 ;
      RECT 38.035 4.022 38.455 4.2 ;
      RECT 38.035 4.01 38.445 4.2 ;
      RECT 38.035 3.995 38.39 4.2 ;
      RECT 38.075 3.967 38.276 4.2 ;
      RECT 38.085 3.945 38.276 4.2 ;
      RECT 38.11 3.93 38.19 4.2 ;
      RECT 37.865 4.46 37.985 4.905 ;
      RECT 37.85 4.46 37.985 4.904 ;
      RECT 37.805 4.482 37.985 4.899 ;
      RECT 37.765 4.531 37.985 4.893 ;
      RECT 37.765 4.531 37.99 4.868 ;
      RECT 37.765 4.531 38.01 4.758 ;
      RECT 37.76 4.561 38.01 4.755 ;
      RECT 37.85 4.46 38.02 4.65 ;
      RECT 37.51 3.245 37.515 3.69 ;
      RECT 37.32 3.245 37.34 3.655 ;
      RECT 37.29 3.245 37.295 3.63 ;
      RECT 37.97 3.552 37.985 3.74 ;
      RECT 37.965 3.537 37.97 3.746 ;
      RECT 37.945 3.51 37.965 3.749 ;
      RECT 37.895 3.477 37.945 3.758 ;
      RECT 37.865 3.457 37.895 3.762 ;
      RECT 37.846 3.445 37.865 3.758 ;
      RECT 37.76 3.417 37.846 3.748 ;
      RECT 37.75 3.392 37.76 3.738 ;
      RECT 37.68 3.36 37.75 3.73 ;
      RECT 37.655 3.32 37.68 3.722 ;
      RECT 37.635 3.302 37.655 3.716 ;
      RECT 37.625 3.292 37.635 3.713 ;
      RECT 37.615 3.285 37.625 3.711 ;
      RECT 37.595 3.272 37.615 3.708 ;
      RECT 37.585 3.262 37.595 3.705 ;
      RECT 37.575 3.255 37.585 3.703 ;
      RECT 37.525 3.247 37.575 3.697 ;
      RECT 37.515 3.245 37.525 3.691 ;
      RECT 37.485 3.245 37.51 3.688 ;
      RECT 37.456 3.245 37.485 3.683 ;
      RECT 37.37 3.245 37.456 3.673 ;
      RECT 37.34 3.245 37.37 3.66 ;
      RECT 37.295 3.245 37.32 3.643 ;
      RECT 37.28 3.245 37.29 3.625 ;
      RECT 37.26 3.252 37.28 3.61 ;
      RECT 37.255 3.267 37.26 3.598 ;
      RECT 37.25 3.272 37.255 3.538 ;
      RECT 37.245 3.277 37.25 3.38 ;
      RECT 37.24 3.28 37.245 3.298 ;
      RECT 37.505 3.965 37.591 4.286 ;
      RECT 37.505 3.965 37.625 4.279 ;
      RECT 37.455 3.965 37.625 4.275 ;
      RECT 37.455 3.967 37.711 4.273 ;
      RECT 37.455 3.969 37.735 4.267 ;
      RECT 37.455 3.976 37.745 4.266 ;
      RECT 37.455 3.985 37.75 4.263 ;
      RECT 37.455 3.991 37.755 4.258 ;
      RECT 37.455 4.035 37.76 4.255 ;
      RECT 37.455 4.127 37.765 4.252 ;
      RECT 36.98 4.57 37.015 4.89 ;
      RECT 37.565 4.755 37.57 4.937 ;
      RECT 37.52 4.637 37.565 4.956 ;
      RECT 37.505 4.614 37.52 4.979 ;
      RECT 37.495 4.604 37.505 4.989 ;
      RECT 37.475 4.599 37.495 5.002 ;
      RECT 37.45 4.597 37.475 5.023 ;
      RECT 37.431 4.596 37.45 5.035 ;
      RECT 37.345 4.593 37.431 5.035 ;
      RECT 37.275 4.588 37.345 5.023 ;
      RECT 37.2 4.584 37.275 4.998 ;
      RECT 37.135 4.58 37.2 4.965 ;
      RECT 37.065 4.577 37.135 4.925 ;
      RECT 37.035 4.573 37.065 4.9 ;
      RECT 37.015 4.571 37.035 4.893 ;
      RECT 36.931 4.569 36.98 4.891 ;
      RECT 36.845 4.566 36.931 4.892 ;
      RECT 36.77 4.565 36.845 4.894 ;
      RECT 36.685 4.565 36.77 4.92 ;
      RECT 36.608 4.566 36.685 4.945 ;
      RECT 36.522 4.567 36.608 4.945 ;
      RECT 36.436 4.567 36.522 4.945 ;
      RECT 36.35 4.568 36.436 4.945 ;
      RECT 36.33 4.569 36.35 4.937 ;
      RECT 36.315 4.575 36.33 4.922 ;
      RECT 36.28 4.595 36.315 4.902 ;
      RECT 36.27 4.615 36.28 4.884 ;
      RECT 37.24 3.92 37.245 4.19 ;
      RECT 37.235 3.911 37.24 4.195 ;
      RECT 37.225 3.901 37.235 4.207 ;
      RECT 37.22 3.89 37.225 4.218 ;
      RECT 37.2 3.884 37.22 4.236 ;
      RECT 37.155 3.881 37.2 4.285 ;
      RECT 37.14 3.88 37.155 4.33 ;
      RECT 37.135 3.88 37.14 4.343 ;
      RECT 37.125 3.88 37.135 4.355 ;
      RECT 37.12 3.881 37.125 4.37 ;
      RECT 37.1 3.889 37.12 4.375 ;
      RECT 37.07 3.905 37.1 4.375 ;
      RECT 37.06 3.917 37.065 4.375 ;
      RECT 37.025 3.932 37.06 4.375 ;
      RECT 36.995 3.952 37.025 4.375 ;
      RECT 36.985 3.977 36.995 4.375 ;
      RECT 36.98 4.005 36.985 4.375 ;
      RECT 36.975 4.035 36.98 4.375 ;
      RECT 36.97 4.052 36.975 4.375 ;
      RECT 36.96 4.08 36.97 4.375 ;
      RECT 36.95 4.115 36.96 4.375 ;
      RECT 36.945 4.15 36.95 4.375 ;
      RECT 37.065 3.915 37.07 4.375 ;
      RECT 36.58 4.017 36.765 4.19 ;
      RECT 36.54 3.935 36.725 4.188 ;
      RECT 36.501 3.94 36.725 4.184 ;
      RECT 36.415 3.949 36.725 4.179 ;
      RECT 36.331 3.965 36.73 4.174 ;
      RECT 36.245 3.985 36.755 4.168 ;
      RECT 36.245 4.005 36.76 4.168 ;
      RECT 36.331 3.975 36.755 4.174 ;
      RECT 36.415 3.95 36.73 4.179 ;
      RECT 36.58 3.932 36.725 4.19 ;
      RECT 36.58 3.927 36.68 4.19 ;
      RECT 36.666 3.921 36.68 4.19 ;
      RECT 36.055 3.245 36.06 3.644 ;
      RECT 35.8 3.245 35.835 3.642 ;
      RECT 35.395 3.28 35.4 3.636 ;
      RECT 36.14 3.283 36.145 3.538 ;
      RECT 36.135 3.281 36.14 3.544 ;
      RECT 36.13 3.28 36.135 3.551 ;
      RECT 36.105 3.273 36.13 3.575 ;
      RECT 36.1 3.266 36.105 3.599 ;
      RECT 36.095 3.262 36.1 3.608 ;
      RECT 36.085 3.257 36.095 3.621 ;
      RECT 36.08 3.254 36.085 3.63 ;
      RECT 36.075 3.252 36.08 3.635 ;
      RECT 36.06 3.248 36.075 3.645 ;
      RECT 36.045 3.242 36.055 3.644 ;
      RECT 36.007 3.24 36.045 3.644 ;
      RECT 35.921 3.242 36.007 3.644 ;
      RECT 35.835 3.244 35.921 3.643 ;
      RECT 35.764 3.245 35.8 3.642 ;
      RECT 35.678 3.247 35.764 3.642 ;
      RECT 35.592 3.249 35.678 3.641 ;
      RECT 35.506 3.251 35.592 3.641 ;
      RECT 35.42 3.254 35.506 3.64 ;
      RECT 35.41 3.26 35.42 3.639 ;
      RECT 35.4 3.272 35.41 3.637 ;
      RECT 35.34 3.307 35.395 3.633 ;
      RECT 35.335 3.337 35.34 3.395 ;
      RECT 36.08 4.417 36.095 4.61 ;
      RECT 36.075 4.385 36.08 4.61 ;
      RECT 36.065 4.36 36.075 4.61 ;
      RECT 36.06 4.332 36.065 4.61 ;
      RECT 36.03 4.255 36.06 4.61 ;
      RECT 36.005 4.137 36.03 4.61 ;
      RECT 36 4.075 36.005 4.61 ;
      RECT 35.99 4.062 36 4.61 ;
      RECT 35.97 4.052 35.99 4.61 ;
      RECT 35.955 4.035 35.97 4.61 ;
      RECT 35.925 4.023 35.955 4.61 ;
      RECT 35.92 4.022 35.925 4.555 ;
      RECT 35.915 4.022 35.92 4.513 ;
      RECT 35.9 4.021 35.915 4.465 ;
      RECT 35.885 4.021 35.9 4.403 ;
      RECT 35.865 4.021 35.885 4.363 ;
      RECT 35.86 4.021 35.865 4.348 ;
      RECT 35.835 4.02 35.86 4.343 ;
      RECT 35.765 4.019 35.835 4.33 ;
      RECT 35.75 4.018 35.765 4.315 ;
      RECT 35.72 4.017 35.75 4.298 ;
      RECT 35.715 4.017 35.72 4.283 ;
      RECT 35.665 4.016 35.715 4.263 ;
      RECT 35.6 4.015 35.665 4.218 ;
      RECT 35.595 4.015 35.6 4.19 ;
      RECT 35.68 4.552 35.685 4.809 ;
      RECT 35.66 4.471 35.68 4.826 ;
      RECT 35.64 4.465 35.66 4.855 ;
      RECT 35.58 4.452 35.64 4.875 ;
      RECT 35.535 4.436 35.58 4.876 ;
      RECT 35.451 4.424 35.535 4.864 ;
      RECT 35.365 4.411 35.451 4.848 ;
      RECT 35.355 4.404 35.365 4.84 ;
      RECT 35.31 4.401 35.355 4.78 ;
      RECT 35.29 4.397 35.31 4.695 ;
      RECT 35.275 4.395 35.29 4.648 ;
      RECT 35.245 4.392 35.275 4.618 ;
      RECT 35.21 4.388 35.245 4.595 ;
      RECT 35.167 4.383 35.21 4.583 ;
      RECT 35.081 4.374 35.167 4.592 ;
      RECT 34.995 4.363 35.081 4.604 ;
      RECT 34.93 4.354 34.995 4.613 ;
      RECT 34.91 4.345 34.93 4.618 ;
      RECT 34.905 4.338 34.91 4.62 ;
      RECT 34.865 4.323 34.905 4.617 ;
      RECT 34.845 4.302 34.865 4.612 ;
      RECT 34.83 4.29 34.845 4.605 ;
      RECT 34.825 4.282 34.83 4.598 ;
      RECT 34.81 4.262 34.825 4.591 ;
      RECT 34.805 4.125 34.81 4.585 ;
      RECT 34.725 4.014 34.805 4.557 ;
      RECT 34.716 4.007 34.725 4.523 ;
      RECT 34.63 4.001 34.716 4.448 ;
      RECT 34.605 3.992 34.63 4.36 ;
      RECT 34.575 3.987 34.605 4.335 ;
      RECT 34.51 3.996 34.575 4.32 ;
      RECT 34.49 4.012 34.51 4.295 ;
      RECT 34.48 4.018 34.49 4.243 ;
      RECT 34.46 4.04 34.48 4.125 ;
      RECT 35.115 4.005 35.285 4.19 ;
      RECT 35.115 4.005 35.32 4.188 ;
      RECT 35.165 3.915 35.335 4.179 ;
      RECT 35.115 4.072 35.34 4.172 ;
      RECT 35.13 3.95 35.335 4.179 ;
      RECT 34.33 4.683 34.395 5.126 ;
      RECT 34.27 4.708 34.395 5.124 ;
      RECT 34.27 4.708 34.45 5.118 ;
      RECT 34.255 4.733 34.45 5.117 ;
      RECT 34.395 4.67 34.47 5.114 ;
      RECT 34.33 4.695 34.55 5.108 ;
      RECT 34.255 4.734 34.595 5.102 ;
      RECT 34.24 4.761 34.595 5.093 ;
      RECT 34.255 4.754 34.615 5.085 ;
      RECT 34.24 4.763 34.62 5.068 ;
      RECT 34.235 4.78 34.62 4.895 ;
      RECT 34.24 3.502 34.275 3.74 ;
      RECT 34.24 3.502 34.305 3.739 ;
      RECT 34.24 3.502 34.42 3.735 ;
      RECT 34.24 3.502 34.475 3.713 ;
      RECT 34.25 3.445 34.53 3.613 ;
      RECT 34.355 3.285 34.385 3.736 ;
      RECT 34.385 3.28 34.565 3.493 ;
      RECT 34.255 3.421 34.565 3.493 ;
      RECT 34.305 3.317 34.355 3.737 ;
      RECT 34.275 3.373 34.565 3.493 ;
      RECT 32.775 3.035 32.945 4.225 ;
      RECT 32.775 3.035 33.245 3.205 ;
      RECT 32.775 9.405 33.245 9.575 ;
      RECT 32.775 8.385 32.945 9.575 ;
      RECT 31.785 3.035 31.955 4.225 ;
      RECT 31.785 3.035 32.255 3.205 ;
      RECT 31.785 9.405 32.255 9.575 ;
      RECT 31.785 8.385 31.955 9.575 ;
      RECT 29.935 3.93 30.105 5.16 ;
      RECT 29.99 2.15 30.16 4.1 ;
      RECT 29.935 1.87 30.105 2.32 ;
      RECT 29.935 10.29 30.105 10.74 ;
      RECT 29.99 8.51 30.16 10.46 ;
      RECT 29.935 7.45 30.105 8.68 ;
      RECT 29.415 1.87 29.585 5.16 ;
      RECT 29.415 3.37 29.82 3.7 ;
      RECT 29.415 2.53 29.82 2.86 ;
      RECT 29.415 7.45 29.585 10.74 ;
      RECT 29.415 9.75 29.82 10.08 ;
      RECT 29.415 8.91 29.82 9.24 ;
      RECT 27.515 4.687 27.53 4.738 ;
      RECT 27.51 4.667 27.515 4.785 ;
      RECT 27.495 4.657 27.51 4.853 ;
      RECT 27.47 4.637 27.495 4.908 ;
      RECT 27.43 4.622 27.47 4.928 ;
      RECT 27.385 4.616 27.43 4.956 ;
      RECT 27.315 4.606 27.385 4.973 ;
      RECT 27.295 4.598 27.315 4.973 ;
      RECT 27.235 4.592 27.295 4.965 ;
      RECT 27.176 4.583 27.235 4.953 ;
      RECT 27.09 4.572 27.176 4.936 ;
      RECT 27.068 4.563 27.09 4.924 ;
      RECT 26.982 4.556 27.068 4.911 ;
      RECT 26.896 4.543 26.982 4.892 ;
      RECT 26.81 4.531 26.896 4.872 ;
      RECT 26.78 4.52 26.81 4.859 ;
      RECT 26.73 4.506 26.78 4.851 ;
      RECT 26.71 4.495 26.73 4.843 ;
      RECT 26.661 4.484 26.71 4.835 ;
      RECT 26.575 4.463 26.661 4.82 ;
      RECT 26.53 4.45 26.575 4.805 ;
      RECT 26.485 4.45 26.53 4.785 ;
      RECT 26.43 4.45 26.485 4.72 ;
      RECT 26.405 4.45 26.43 4.643 ;
      RECT 26.93 4.187 27.1 4.37 ;
      RECT 26.93 4.187 27.115 4.328 ;
      RECT 26.93 4.187 27.12 4.27 ;
      RECT 26.99 3.955 27.125 4.246 ;
      RECT 26.99 3.959 27.13 4.229 ;
      RECT 26.935 4.122 27.13 4.229 ;
      RECT 26.96 3.967 27.1 4.37 ;
      RECT 26.96 3.971 27.14 4.17 ;
      RECT 26.945 4.057 27.14 4.17 ;
      RECT 26.955 3.987 27.1 4.37 ;
      RECT 26.955 3.99 27.15 4.083 ;
      RECT 26.95 4.007 27.15 4.083 ;
      RECT 26.72 3.227 26.89 3.71 ;
      RECT 26.715 3.222 26.865 3.7 ;
      RECT 26.715 3.229 26.895 3.694 ;
      RECT 26.705 3.223 26.865 3.673 ;
      RECT 26.705 3.239 26.91 3.632 ;
      RECT 26.675 3.224 26.865 3.595 ;
      RECT 26.675 3.254 26.92 3.535 ;
      RECT 26.67 3.226 26.865 3.533 ;
      RECT 26.65 3.235 26.895 3.49 ;
      RECT 26.625 3.251 26.91 3.402 ;
      RECT 26.625 3.27 26.935 3.393 ;
      RECT 26.62 3.307 26.935 3.345 ;
      RECT 26.625 3.287 26.94 3.313 ;
      RECT 26.72 3.221 26.83 3.71 ;
      RECT 26.806 3.22 26.83 3.71 ;
      RECT 26.04 4.005 26.045 4.216 ;
      RECT 26.64 4.005 26.645 4.19 ;
      RECT 26.705 4.045 26.71 4.158 ;
      RECT 26.7 4.037 26.705 4.164 ;
      RECT 26.695 4.027 26.7 4.172 ;
      RECT 26.69 4.017 26.695 4.181 ;
      RECT 26.685 4.007 26.69 4.185 ;
      RECT 26.645 4.005 26.685 4.188 ;
      RECT 26.617 4.004 26.64 4.192 ;
      RECT 26.531 4.001 26.617 4.199 ;
      RECT 26.445 3.997 26.531 4.21 ;
      RECT 26.425 3.995 26.445 4.216 ;
      RECT 26.407 3.994 26.425 4.219 ;
      RECT 26.321 3.992 26.407 4.226 ;
      RECT 26.235 3.987 26.321 4.239 ;
      RECT 26.216 3.984 26.235 4.244 ;
      RECT 26.13 3.982 26.216 4.235 ;
      RECT 26.12 3.982 26.13 4.228 ;
      RECT 26.045 3.995 26.12 4.222 ;
      RECT 26.03 4.006 26.04 4.216 ;
      RECT 26.02 4.008 26.03 4.215 ;
      RECT 26.01 4.012 26.02 4.211 ;
      RECT 26.005 4.015 26.01 4.205 ;
      RECT 25.995 4.017 26.005 4.199 ;
      RECT 25.99 4.02 25.995 4.193 ;
      RECT 25.97 4.606 25.975 4.81 ;
      RECT 25.955 4.593 25.97 4.903 ;
      RECT 25.94 4.574 25.955 5.18 ;
      RECT 25.905 4.54 25.94 5.18 ;
      RECT 25.901 4.51 25.905 5.18 ;
      RECT 25.815 4.392 25.901 5.18 ;
      RECT 25.805 4.267 25.815 5.18 ;
      RECT 25.79 4.235 25.805 5.18 ;
      RECT 25.785 4.21 25.79 5.18 ;
      RECT 25.78 4.2 25.785 5.136 ;
      RECT 25.765 4.172 25.78 5.041 ;
      RECT 25.75 4.138 25.765 4.94 ;
      RECT 25.745 4.116 25.75 4.893 ;
      RECT 25.74 4.105 25.745 4.863 ;
      RECT 25.735 4.095 25.74 4.829 ;
      RECT 25.725 4.082 25.735 4.797 ;
      RECT 25.7 4.058 25.725 4.723 ;
      RECT 25.695 4.038 25.7 4.648 ;
      RECT 25.69 4.032 25.695 4.623 ;
      RECT 25.685 4.027 25.69 4.588 ;
      RECT 25.68 4.022 25.685 4.563 ;
      RECT 25.675 4.02 25.68 4.543 ;
      RECT 25.67 4.02 25.675 4.528 ;
      RECT 25.665 4.02 25.67 4.488 ;
      RECT 25.655 4.02 25.665 4.46 ;
      RECT 25.645 4.02 25.655 4.405 ;
      RECT 25.63 4.02 25.645 4.343 ;
      RECT 25.625 4.019 25.63 4.288 ;
      RECT 25.61 4.018 25.625 4.268 ;
      RECT 25.55 4.016 25.61 4.242 ;
      RECT 25.515 4.017 25.55 4.222 ;
      RECT 25.51 4.019 25.515 4.212 ;
      RECT 25.5 4.038 25.51 4.202 ;
      RECT 25.495 4.065 25.5 4.133 ;
      RECT 25.61 3.49 25.78 3.735 ;
      RECT 25.645 3.261 25.78 3.735 ;
      RECT 25.645 3.263 25.79 3.73 ;
      RECT 25.645 3.265 25.815 3.718 ;
      RECT 25.645 3.268 25.84 3.7 ;
      RECT 25.645 3.273 25.89 3.673 ;
      RECT 25.645 3.278 25.91 3.638 ;
      RECT 25.625 3.28 25.92 3.613 ;
      RECT 25.615 3.375 25.92 3.613 ;
      RECT 25.645 3.26 25.755 3.735 ;
      RECT 25.655 3.257 25.75 3.735 ;
      RECT 25.175 4.522 25.365 4.88 ;
      RECT 25.175 4.534 25.4 4.879 ;
      RECT 25.175 4.562 25.42 4.877 ;
      RECT 25.175 4.587 25.425 4.876 ;
      RECT 25.175 4.645 25.44 4.875 ;
      RECT 25.16 4.518 25.32 4.86 ;
      RECT 25.14 4.527 25.365 4.813 ;
      RECT 25.115 4.538 25.4 4.75 ;
      RECT 25.115 4.622 25.435 4.75 ;
      RECT 25.115 4.597 25.43 4.75 ;
      RECT 25.175 4.513 25.32 4.88 ;
      RECT 25.261 4.512 25.32 4.88 ;
      RECT 25.261 4.511 25.305 4.88 ;
      RECT 24.655 7.45 24.825 10.74 ;
      RECT 24.655 9.75 25.06 10.08 ;
      RECT 24.655 8.91 25.06 9.24 ;
      RECT 24.96 4.027 24.965 4.405 ;
      RECT 24.955 3.995 24.96 4.405 ;
      RECT 24.95 3.967 24.955 4.405 ;
      RECT 24.945 3.947 24.95 4.405 ;
      RECT 24.89 3.93 24.945 4.405 ;
      RECT 24.85 3.915 24.89 4.405 ;
      RECT 24.795 3.902 24.85 4.405 ;
      RECT 24.76 3.893 24.795 4.405 ;
      RECT 24.756 3.891 24.76 4.404 ;
      RECT 24.67 3.887 24.756 4.387 ;
      RECT 24.585 3.879 24.67 4.35 ;
      RECT 24.575 3.875 24.585 4.323 ;
      RECT 24.565 3.875 24.575 4.305 ;
      RECT 24.555 3.877 24.565 4.288 ;
      RECT 24.55 3.882 24.555 4.274 ;
      RECT 24.545 3.886 24.55 4.261 ;
      RECT 24.535 3.891 24.545 4.245 ;
      RECT 24.52 3.905 24.535 4.22 ;
      RECT 24.515 3.911 24.52 4.2 ;
      RECT 24.51 3.913 24.515 4.193 ;
      RECT 24.505 3.917 24.51 4.068 ;
      RECT 24.685 4.717 24.93 5.18 ;
      RECT 24.605 4.69 24.925 5.176 ;
      RECT 24.535 4.725 24.93 5.169 ;
      RECT 24.325 4.98 24.93 5.165 ;
      RECT 24.505 4.748 24.93 5.165 ;
      RECT 24.345 4.94 24.93 5.165 ;
      RECT 24.495 4.76 24.93 5.165 ;
      RECT 24.38 4.877 24.93 5.165 ;
      RECT 24.435 4.802 24.93 5.165 ;
      RECT 24.685 4.667 24.925 5.18 ;
      RECT 24.715 4.66 24.925 5.18 ;
      RECT 24.705 4.662 24.925 5.18 ;
      RECT 24.715 4.657 24.845 5.18 ;
      RECT 24.27 3.22 24.356 3.659 ;
      RECT 24.265 3.22 24.356 3.657 ;
      RECT 24.265 3.22 24.425 3.656 ;
      RECT 24.265 3.22 24.455 3.653 ;
      RECT 24.25 3.227 24.455 3.644 ;
      RECT 24.25 3.227 24.46 3.64 ;
      RECT 24.245 3.237 24.46 3.633 ;
      RECT 24.24 3.242 24.46 3.608 ;
      RECT 24.24 3.242 24.475 3.59 ;
      RECT 24.265 3.22 24.495 3.505 ;
      RECT 24.235 3.247 24.495 3.503 ;
      RECT 24.245 3.24 24.5 3.441 ;
      RECT 24.235 3.362 24.505 3.424 ;
      RECT 24.22 3.257 24.5 3.375 ;
      RECT 24.215 3.267 24.5 3.275 ;
      RECT 24.295 4.038 24.3 4.115 ;
      RECT 24.285 4.032 24.295 4.305 ;
      RECT 24.275 4.024 24.285 4.326 ;
      RECT 24.265 4.015 24.275 4.348 ;
      RECT 24.26 4.01 24.265 4.365 ;
      RECT 24.22 4.01 24.26 4.405 ;
      RECT 24.2 4.01 24.22 4.46 ;
      RECT 24.195 4.01 24.2 4.488 ;
      RECT 24.185 4.01 24.195 4.503 ;
      RECT 24.15 4.01 24.185 4.545 ;
      RECT 24.145 4.01 24.15 4.588 ;
      RECT 24.135 4.01 24.145 4.603 ;
      RECT 24.12 4.01 24.135 4.623 ;
      RECT 24.105 4.01 24.12 4.65 ;
      RECT 24.1 4.011 24.105 4.668 ;
      RECT 24.08 4.012 24.1 4.675 ;
      RECT 24.025 4.013 24.08 4.695 ;
      RECT 24.015 4.014 24.025 4.709 ;
      RECT 24.01 4.017 24.015 4.708 ;
      RECT 23.97 4.09 24.01 4.706 ;
      RECT 23.955 4.17 23.97 4.704 ;
      RECT 23.93 4.225 23.955 4.702 ;
      RECT 23.915 4.29 23.93 4.701 ;
      RECT 23.87 4.322 23.915 4.698 ;
      RECT 23.785 4.345 23.87 4.693 ;
      RECT 23.76 4.365 23.785 4.688 ;
      RECT 23.69 4.37 23.76 4.684 ;
      RECT 23.67 4.372 23.69 4.681 ;
      RECT 23.585 4.383 23.67 4.675 ;
      RECT 23.58 4.394 23.585 4.67 ;
      RECT 23.57 4.396 23.58 4.67 ;
      RECT 23.535 4.4 23.57 4.668 ;
      RECT 23.485 4.41 23.535 4.655 ;
      RECT 23.465 4.418 23.485 4.64 ;
      RECT 23.385 4.43 23.465 4.623 ;
      RECT 23.55 3.98 23.72 4.19 ;
      RECT 23.666 3.976 23.72 4.19 ;
      RECT 23.471 3.98 23.72 4.181 ;
      RECT 23.471 3.98 23.725 4.17 ;
      RECT 23.385 3.98 23.725 4.161 ;
      RECT 23.385 3.988 23.735 4.105 ;
      RECT 23.385 4 23.74 4.018 ;
      RECT 23.385 4.007 23.745 4.01 ;
      RECT 23.58 3.978 23.72 4.19 ;
      RECT 23.335 4.923 23.58 5.255 ;
      RECT 23.33 4.915 23.335 5.252 ;
      RECT 23.3 4.935 23.58 5.233 ;
      RECT 23.28 4.967 23.58 5.206 ;
      RECT 23.33 4.92 23.507 5.252 ;
      RECT 23.33 4.917 23.421 5.252 ;
      RECT 23.27 3.265 23.44 3.685 ;
      RECT 23.265 3.265 23.44 3.683 ;
      RECT 23.265 3.265 23.465 3.673 ;
      RECT 23.265 3.265 23.485 3.648 ;
      RECT 23.26 3.265 23.485 3.643 ;
      RECT 23.26 3.265 23.495 3.633 ;
      RECT 23.26 3.265 23.5 3.628 ;
      RECT 23.26 3.27 23.505 3.623 ;
      RECT 23.26 3.302 23.52 3.613 ;
      RECT 23.26 3.372 23.545 3.596 ;
      RECT 23.24 3.372 23.545 3.588 ;
      RECT 23.24 3.432 23.555 3.565 ;
      RECT 23.24 3.472 23.565 3.51 ;
      RECT 23.225 3.265 23.5 3.49 ;
      RECT 23.215 3.28 23.505 3.388 ;
      RECT 22.805 4.67 22.975 5.195 ;
      RECT 22.8 4.67 22.975 5.188 ;
      RECT 22.79 4.67 22.98 5.153 ;
      RECT 22.785 4.68 22.98 5.125 ;
      RECT 22.78 4.7 22.98 5.108 ;
      RECT 22.79 4.675 22.985 5.098 ;
      RECT 22.775 4.72 22.985 5.09 ;
      RECT 22.77 4.74 22.985 5.075 ;
      RECT 22.765 4.77 22.985 5.065 ;
      RECT 22.755 4.815 22.985 5.04 ;
      RECT 22.785 4.685 22.99 5.023 ;
      RECT 22.75 4.867 22.99 5.018 ;
      RECT 22.785 4.695 22.995 4.988 ;
      RECT 22.745 4.9 22.995 4.985 ;
      RECT 22.74 4.925 22.995 4.965 ;
      RECT 22.78 4.712 23.005 4.905 ;
      RECT 22.775 4.734 23.015 4.798 ;
      RECT 22.725 3.981 22.74 4.25 ;
      RECT 22.68 3.965 22.725 4.295 ;
      RECT 22.675 3.953 22.68 4.345 ;
      RECT 22.665 3.949 22.675 4.378 ;
      RECT 22.66 3.946 22.665 4.406 ;
      RECT 22.645 3.948 22.66 4.448 ;
      RECT 22.64 3.952 22.645 4.488 ;
      RECT 22.62 3.957 22.64 4.54 ;
      RECT 22.616 3.962 22.62 4.597 ;
      RECT 22.53 3.981 22.616 4.634 ;
      RECT 22.52 4.002 22.53 4.67 ;
      RECT 22.515 4.01 22.52 4.671 ;
      RECT 22.51 4.052 22.515 4.672 ;
      RECT 22.495 4.14 22.51 4.673 ;
      RECT 22.485 4.29 22.495 4.675 ;
      RECT 22.48 4.335 22.485 4.677 ;
      RECT 22.445 4.377 22.48 4.68 ;
      RECT 22.44 4.395 22.445 4.683 ;
      RECT 22.363 4.401 22.44 4.689 ;
      RECT 22.277 4.415 22.363 4.702 ;
      RECT 22.191 4.429 22.277 4.716 ;
      RECT 22.105 4.443 22.191 4.729 ;
      RECT 22.045 4.455 22.105 4.741 ;
      RECT 22.02 4.462 22.045 4.748 ;
      RECT 22.006 4.465 22.02 4.753 ;
      RECT 21.92 4.473 22.006 4.769 ;
      RECT 21.915 4.48 21.92 4.784 ;
      RECT 21.891 4.48 21.915 4.791 ;
      RECT 21.805 4.483 21.891 4.819 ;
      RECT 21.72 4.487 21.805 4.863 ;
      RECT 21.655 4.491 21.72 4.9 ;
      RECT 21.63 4.494 21.655 4.916 ;
      RECT 21.555 4.507 21.63 4.92 ;
      RECT 21.53 4.525 21.555 4.924 ;
      RECT 21.52 4.532 21.53 4.926 ;
      RECT 21.505 4.535 21.52 4.927 ;
      RECT 21.445 4.547 21.505 4.931 ;
      RECT 21.435 4.561 21.445 4.935 ;
      RECT 21.38 4.571 21.435 4.923 ;
      RECT 21.355 4.592 21.38 4.906 ;
      RECT 21.335 4.612 21.355 4.897 ;
      RECT 21.33 4.625 21.335 4.892 ;
      RECT 21.315 4.637 21.33 4.888 ;
      RECT 22.55 3.292 22.555 3.315 ;
      RECT 22.545 3.283 22.55 3.355 ;
      RECT 22.54 3.281 22.545 3.398 ;
      RECT 22.535 3.272 22.54 3.433 ;
      RECT 22.53 3.262 22.535 3.505 ;
      RECT 22.525 3.252 22.53 3.57 ;
      RECT 22.52 3.249 22.525 3.61 ;
      RECT 22.495 3.243 22.52 3.7 ;
      RECT 22.46 3.231 22.495 3.725 ;
      RECT 22.45 3.222 22.46 3.725 ;
      RECT 22.315 3.22 22.325 3.708 ;
      RECT 22.305 3.22 22.315 3.675 ;
      RECT 22.3 3.22 22.305 3.65 ;
      RECT 22.295 3.22 22.3 3.638 ;
      RECT 22.29 3.22 22.295 3.62 ;
      RECT 22.28 3.22 22.29 3.585 ;
      RECT 22.275 3.222 22.28 3.563 ;
      RECT 22.27 3.228 22.275 3.548 ;
      RECT 22.265 3.234 22.27 3.533 ;
      RECT 22.25 3.246 22.265 3.506 ;
      RECT 22.245 3.257 22.25 3.474 ;
      RECT 22.24 3.267 22.245 3.458 ;
      RECT 22.23 3.275 22.24 3.427 ;
      RECT 22.225 3.285 22.23 3.401 ;
      RECT 22.22 3.342 22.225 3.384 ;
      RECT 22.325 3.22 22.45 3.725 ;
      RECT 22.04 3.907 22.3 4.205 ;
      RECT 22.035 3.914 22.3 4.203 ;
      RECT 22.04 3.909 22.315 4.198 ;
      RECT 22.03 3.922 22.315 4.195 ;
      RECT 22.03 3.927 22.32 4.188 ;
      RECT 22.025 3.935 22.32 4.185 ;
      RECT 22.025 3.952 22.325 3.983 ;
      RECT 22.04 3.904 22.271 4.205 ;
      RECT 22.095 3.903 22.271 4.205 ;
      RECT 22.095 3.9 22.185 4.205 ;
      RECT 22.095 3.897 22.181 4.205 ;
      RECT 21.785 4.17 21.79 4.183 ;
      RECT 21.78 4.137 21.785 4.188 ;
      RECT 21.775 4.092 21.78 4.195 ;
      RECT 21.77 4.047 21.775 4.203 ;
      RECT 21.765 4.015 21.77 4.211 ;
      RECT 21.76 3.975 21.765 4.212 ;
      RECT 21.745 3.955 21.76 4.214 ;
      RECT 21.67 3.937 21.745 4.226 ;
      RECT 21.66 3.93 21.67 4.237 ;
      RECT 21.655 3.93 21.66 4.239 ;
      RECT 21.625 3.936 21.655 4.243 ;
      RECT 21.585 3.949 21.625 4.243 ;
      RECT 21.56 3.96 21.585 4.229 ;
      RECT 21.545 3.966 21.56 4.212 ;
      RECT 21.535 3.968 21.545 4.203 ;
      RECT 21.53 3.969 21.535 4.198 ;
      RECT 21.525 3.97 21.53 4.193 ;
      RECT 21.52 3.971 21.525 4.19 ;
      RECT 21.495 3.976 21.52 4.18 ;
      RECT 21.485 3.992 21.495 4.167 ;
      RECT 21.48 4.012 21.485 4.162 ;
      RECT 21.49 3.405 21.495 3.601 ;
      RECT 21.475 3.369 21.49 3.603 ;
      RECT 21.465 3.351 21.475 3.608 ;
      RECT 21.455 3.337 21.465 3.612 ;
      RECT 21.41 3.321 21.455 3.622 ;
      RECT 21.405 3.311 21.41 3.631 ;
      RECT 21.36 3.3 21.405 3.637 ;
      RECT 21.355 3.288 21.36 3.644 ;
      RECT 21.34 3.283 21.355 3.648 ;
      RECT 21.325 3.275 21.34 3.653 ;
      RECT 21.315 3.268 21.325 3.658 ;
      RECT 21.305 3.265 21.315 3.663 ;
      RECT 21.295 3.265 21.305 3.664 ;
      RECT 21.29 3.262 21.295 3.663 ;
      RECT 21.255 3.257 21.28 3.662 ;
      RECT 21.231 3.253 21.255 3.661 ;
      RECT 21.145 3.244 21.231 3.658 ;
      RECT 21.13 3.236 21.145 3.655 ;
      RECT 21.108 3.235 21.13 3.654 ;
      RECT 21.022 3.235 21.108 3.652 ;
      RECT 20.936 3.235 21.022 3.65 ;
      RECT 20.85 3.235 20.936 3.647 ;
      RECT 20.84 3.235 20.85 3.638 ;
      RECT 20.81 3.235 20.84 3.598 ;
      RECT 20.8 3.245 20.81 3.553 ;
      RECT 20.795 3.285 20.8 3.538 ;
      RECT 20.79 3.3 20.795 3.525 ;
      RECT 20.76 3.38 20.79 3.487 ;
      RECT 21.28 3.26 21.29 3.663 ;
      RECT 21.105 4.025 21.12 4.63 ;
      RECT 21.11 4.02 21.12 4.63 ;
      RECT 21.275 4.02 21.28 4.203 ;
      RECT 21.265 4.02 21.275 4.233 ;
      RECT 21.25 4.02 21.265 4.293 ;
      RECT 21.245 4.02 21.25 4.338 ;
      RECT 21.24 4.02 21.245 4.368 ;
      RECT 21.235 4.02 21.24 4.388 ;
      RECT 21.225 4.02 21.235 4.423 ;
      RECT 21.21 4.02 21.225 4.455 ;
      RECT 21.165 4.02 21.21 4.483 ;
      RECT 21.16 4.02 21.165 4.513 ;
      RECT 21.155 4.02 21.16 4.525 ;
      RECT 21.15 4.02 21.155 4.533 ;
      RECT 21.14 4.02 21.15 4.548 ;
      RECT 21.135 4.02 21.14 4.57 ;
      RECT 21.125 4.02 21.135 4.593 ;
      RECT 21.12 4.02 21.125 4.613 ;
      RECT 21.085 4.035 21.105 4.63 ;
      RECT 21.06 4.052 21.085 4.63 ;
      RECT 21.055 4.062 21.06 4.63 ;
      RECT 21.025 4.077 21.055 4.63 ;
      RECT 20.95 4.119 21.025 4.63 ;
      RECT 20.945 4.15 20.95 4.613 ;
      RECT 20.94 4.154 20.945 4.595 ;
      RECT 20.935 4.158 20.94 4.558 ;
      RECT 20.93 4.342 20.935 4.525 ;
      RECT 20.415 4.531 20.501 5.096 ;
      RECT 20.37 4.533 20.535 5.09 ;
      RECT 20.501 4.53 20.535 5.09 ;
      RECT 20.415 4.532 20.62 5.084 ;
      RECT 20.37 4.542 20.63 5.08 ;
      RECT 20.345 4.534 20.62 5.076 ;
      RECT 20.34 4.537 20.62 5.071 ;
      RECT 20.315 4.552 20.63 5.065 ;
      RECT 20.315 4.577 20.67 5.06 ;
      RECT 20.275 4.585 20.67 5.035 ;
      RECT 20.275 4.612 20.685 5.033 ;
      RECT 20.275 4.642 20.695 5.02 ;
      RECT 20.27 4.787 20.695 5.008 ;
      RECT 20.275 4.716 20.715 5.005 ;
      RECT 20.275 4.773 20.72 4.813 ;
      RECT 20.465 4.052 20.635 4.23 ;
      RECT 20.415 3.991 20.465 4.215 ;
      RECT 20.15 3.971 20.415 4.2 ;
      RECT 20.11 4.035 20.585 4.2 ;
      RECT 20.11 4.025 20.54 4.2 ;
      RECT 20.11 4.022 20.53 4.2 ;
      RECT 20.11 4.01 20.52 4.2 ;
      RECT 20.11 3.995 20.465 4.2 ;
      RECT 20.15 3.967 20.351 4.2 ;
      RECT 20.16 3.945 20.351 4.2 ;
      RECT 20.185 3.93 20.265 4.2 ;
      RECT 19.94 4.46 20.06 4.905 ;
      RECT 19.925 4.46 20.06 4.904 ;
      RECT 19.88 4.482 20.06 4.899 ;
      RECT 19.84 4.531 20.06 4.893 ;
      RECT 19.84 4.531 20.065 4.868 ;
      RECT 19.84 4.531 20.085 4.758 ;
      RECT 19.835 4.561 20.085 4.755 ;
      RECT 19.925 4.46 20.095 4.65 ;
      RECT 19.585 3.245 19.59 3.69 ;
      RECT 19.395 3.245 19.415 3.655 ;
      RECT 19.365 3.245 19.37 3.63 ;
      RECT 20.045 3.552 20.06 3.74 ;
      RECT 20.04 3.537 20.045 3.746 ;
      RECT 20.02 3.51 20.04 3.749 ;
      RECT 19.97 3.477 20.02 3.758 ;
      RECT 19.94 3.457 19.97 3.762 ;
      RECT 19.921 3.445 19.94 3.758 ;
      RECT 19.835 3.417 19.921 3.748 ;
      RECT 19.825 3.392 19.835 3.738 ;
      RECT 19.755 3.36 19.825 3.73 ;
      RECT 19.73 3.32 19.755 3.722 ;
      RECT 19.71 3.302 19.73 3.716 ;
      RECT 19.7 3.292 19.71 3.713 ;
      RECT 19.69 3.285 19.7 3.711 ;
      RECT 19.67 3.272 19.69 3.708 ;
      RECT 19.66 3.262 19.67 3.705 ;
      RECT 19.65 3.255 19.66 3.703 ;
      RECT 19.6 3.247 19.65 3.697 ;
      RECT 19.59 3.245 19.6 3.691 ;
      RECT 19.56 3.245 19.585 3.688 ;
      RECT 19.531 3.245 19.56 3.683 ;
      RECT 19.445 3.245 19.531 3.673 ;
      RECT 19.415 3.245 19.445 3.66 ;
      RECT 19.37 3.245 19.395 3.643 ;
      RECT 19.355 3.245 19.365 3.625 ;
      RECT 19.335 3.252 19.355 3.61 ;
      RECT 19.33 3.267 19.335 3.598 ;
      RECT 19.325 3.272 19.33 3.538 ;
      RECT 19.32 3.277 19.325 3.38 ;
      RECT 19.315 3.28 19.32 3.298 ;
      RECT 19.58 3.965 19.666 4.286 ;
      RECT 19.58 3.965 19.7 4.279 ;
      RECT 19.53 3.965 19.7 4.275 ;
      RECT 19.53 3.967 19.786 4.273 ;
      RECT 19.53 3.969 19.81 4.267 ;
      RECT 19.53 3.976 19.82 4.266 ;
      RECT 19.53 3.985 19.825 4.263 ;
      RECT 19.53 3.991 19.83 4.258 ;
      RECT 19.53 4.035 19.835 4.255 ;
      RECT 19.53 4.127 19.84 4.252 ;
      RECT 19.055 4.57 19.09 4.89 ;
      RECT 19.64 4.755 19.645 4.937 ;
      RECT 19.595 4.637 19.64 4.956 ;
      RECT 19.58 4.614 19.595 4.979 ;
      RECT 19.57 4.604 19.58 4.989 ;
      RECT 19.55 4.599 19.57 5.002 ;
      RECT 19.525 4.597 19.55 5.023 ;
      RECT 19.506 4.596 19.525 5.035 ;
      RECT 19.42 4.593 19.506 5.035 ;
      RECT 19.35 4.588 19.42 5.023 ;
      RECT 19.275 4.584 19.35 4.998 ;
      RECT 19.21 4.58 19.275 4.965 ;
      RECT 19.14 4.577 19.21 4.925 ;
      RECT 19.11 4.573 19.14 4.9 ;
      RECT 19.09 4.571 19.11 4.893 ;
      RECT 19.006 4.569 19.055 4.891 ;
      RECT 18.92 4.566 19.006 4.892 ;
      RECT 18.845 4.565 18.92 4.894 ;
      RECT 18.76 4.565 18.845 4.92 ;
      RECT 18.683 4.566 18.76 4.945 ;
      RECT 18.597 4.567 18.683 4.945 ;
      RECT 18.511 4.567 18.597 4.945 ;
      RECT 18.425 4.568 18.511 4.945 ;
      RECT 18.405 4.569 18.425 4.937 ;
      RECT 18.39 4.575 18.405 4.922 ;
      RECT 18.355 4.595 18.39 4.902 ;
      RECT 18.345 4.615 18.355 4.884 ;
      RECT 19.315 3.92 19.32 4.19 ;
      RECT 19.31 3.911 19.315 4.195 ;
      RECT 19.3 3.901 19.31 4.207 ;
      RECT 19.295 3.89 19.3 4.218 ;
      RECT 19.275 3.884 19.295 4.236 ;
      RECT 19.23 3.881 19.275 4.285 ;
      RECT 19.215 3.88 19.23 4.33 ;
      RECT 19.21 3.88 19.215 4.343 ;
      RECT 19.2 3.88 19.21 4.355 ;
      RECT 19.195 3.881 19.2 4.37 ;
      RECT 19.175 3.889 19.195 4.375 ;
      RECT 19.145 3.905 19.175 4.375 ;
      RECT 19.135 3.917 19.14 4.375 ;
      RECT 19.1 3.932 19.135 4.375 ;
      RECT 19.07 3.952 19.1 4.375 ;
      RECT 19.06 3.977 19.07 4.375 ;
      RECT 19.055 4.005 19.06 4.375 ;
      RECT 19.05 4.035 19.055 4.375 ;
      RECT 19.045 4.052 19.05 4.375 ;
      RECT 19.035 4.08 19.045 4.375 ;
      RECT 19.025 4.115 19.035 4.375 ;
      RECT 19.02 4.15 19.025 4.375 ;
      RECT 19.14 3.915 19.145 4.375 ;
      RECT 18.655 4.017 18.84 4.19 ;
      RECT 18.615 3.935 18.8 4.188 ;
      RECT 18.576 3.94 18.8 4.184 ;
      RECT 18.49 3.949 18.8 4.179 ;
      RECT 18.406 3.965 18.805 4.174 ;
      RECT 18.32 3.985 18.83 4.168 ;
      RECT 18.32 4.005 18.835 4.168 ;
      RECT 18.406 3.975 18.83 4.174 ;
      RECT 18.49 3.95 18.805 4.179 ;
      RECT 18.655 3.932 18.8 4.19 ;
      RECT 18.655 3.927 18.755 4.19 ;
      RECT 18.741 3.921 18.755 4.19 ;
      RECT 18.13 3.245 18.135 3.644 ;
      RECT 17.875 3.245 17.91 3.642 ;
      RECT 17.47 3.28 17.475 3.636 ;
      RECT 18.215 3.283 18.22 3.538 ;
      RECT 18.21 3.281 18.215 3.544 ;
      RECT 18.205 3.28 18.21 3.551 ;
      RECT 18.18 3.273 18.205 3.575 ;
      RECT 18.175 3.266 18.18 3.599 ;
      RECT 18.17 3.262 18.175 3.608 ;
      RECT 18.16 3.257 18.17 3.621 ;
      RECT 18.155 3.254 18.16 3.63 ;
      RECT 18.15 3.252 18.155 3.635 ;
      RECT 18.135 3.248 18.15 3.645 ;
      RECT 18.12 3.242 18.13 3.644 ;
      RECT 18.082 3.24 18.12 3.644 ;
      RECT 17.996 3.242 18.082 3.644 ;
      RECT 17.91 3.244 17.996 3.643 ;
      RECT 17.839 3.245 17.875 3.642 ;
      RECT 17.753 3.247 17.839 3.642 ;
      RECT 17.667 3.249 17.753 3.641 ;
      RECT 17.581 3.251 17.667 3.641 ;
      RECT 17.495 3.254 17.581 3.64 ;
      RECT 17.485 3.26 17.495 3.639 ;
      RECT 17.475 3.272 17.485 3.637 ;
      RECT 17.415 3.307 17.47 3.633 ;
      RECT 17.41 3.337 17.415 3.395 ;
      RECT 18.155 4.417 18.17 4.61 ;
      RECT 18.15 4.385 18.155 4.61 ;
      RECT 18.14 4.36 18.15 4.61 ;
      RECT 18.135 4.332 18.14 4.61 ;
      RECT 18.105 4.255 18.135 4.61 ;
      RECT 18.08 4.137 18.105 4.61 ;
      RECT 18.075 4.075 18.08 4.61 ;
      RECT 18.065 4.062 18.075 4.61 ;
      RECT 18.045 4.052 18.065 4.61 ;
      RECT 18.03 4.035 18.045 4.61 ;
      RECT 18 4.023 18.03 4.61 ;
      RECT 17.995 4.022 18 4.555 ;
      RECT 17.99 4.022 17.995 4.513 ;
      RECT 17.975 4.021 17.99 4.465 ;
      RECT 17.96 4.021 17.975 4.403 ;
      RECT 17.94 4.021 17.96 4.363 ;
      RECT 17.935 4.021 17.94 4.348 ;
      RECT 17.91 4.02 17.935 4.343 ;
      RECT 17.84 4.019 17.91 4.33 ;
      RECT 17.825 4.018 17.84 4.315 ;
      RECT 17.795 4.017 17.825 4.298 ;
      RECT 17.79 4.017 17.795 4.283 ;
      RECT 17.74 4.016 17.79 4.263 ;
      RECT 17.675 4.015 17.74 4.218 ;
      RECT 17.67 4.015 17.675 4.19 ;
      RECT 17.755 4.552 17.76 4.809 ;
      RECT 17.735 4.471 17.755 4.826 ;
      RECT 17.715 4.465 17.735 4.855 ;
      RECT 17.655 4.452 17.715 4.875 ;
      RECT 17.61 4.436 17.655 4.876 ;
      RECT 17.526 4.424 17.61 4.864 ;
      RECT 17.44 4.411 17.526 4.848 ;
      RECT 17.43 4.404 17.44 4.84 ;
      RECT 17.385 4.401 17.43 4.78 ;
      RECT 17.365 4.397 17.385 4.695 ;
      RECT 17.35 4.395 17.365 4.648 ;
      RECT 17.32 4.392 17.35 4.618 ;
      RECT 17.285 4.388 17.32 4.595 ;
      RECT 17.242 4.383 17.285 4.583 ;
      RECT 17.156 4.374 17.242 4.592 ;
      RECT 17.07 4.363 17.156 4.604 ;
      RECT 17.005 4.354 17.07 4.613 ;
      RECT 16.985 4.345 17.005 4.618 ;
      RECT 16.98 4.338 16.985 4.62 ;
      RECT 16.94 4.323 16.98 4.617 ;
      RECT 16.92 4.302 16.94 4.612 ;
      RECT 16.905 4.29 16.92 4.605 ;
      RECT 16.9 4.282 16.905 4.598 ;
      RECT 16.885 4.262 16.9 4.591 ;
      RECT 16.88 4.125 16.885 4.585 ;
      RECT 16.8 4.014 16.88 4.557 ;
      RECT 16.791 4.007 16.8 4.523 ;
      RECT 16.705 4.001 16.791 4.448 ;
      RECT 16.68 3.992 16.705 4.36 ;
      RECT 16.65 3.987 16.68 4.335 ;
      RECT 16.585 3.996 16.65 4.32 ;
      RECT 16.565 4.012 16.585 4.295 ;
      RECT 16.555 4.018 16.565 4.243 ;
      RECT 16.535 4.04 16.555 4.125 ;
      RECT 17.19 4.005 17.36 4.19 ;
      RECT 17.19 4.005 17.395 4.188 ;
      RECT 17.24 3.915 17.41 4.179 ;
      RECT 17.19 4.072 17.415 4.172 ;
      RECT 17.205 3.95 17.41 4.179 ;
      RECT 16.405 4.683 16.47 5.126 ;
      RECT 16.345 4.708 16.47 5.124 ;
      RECT 16.345 4.708 16.525 5.118 ;
      RECT 16.33 4.733 16.525 5.117 ;
      RECT 16.47 4.67 16.545 5.114 ;
      RECT 16.405 4.695 16.625 5.108 ;
      RECT 16.33 4.734 16.67 5.102 ;
      RECT 16.315 4.761 16.67 5.093 ;
      RECT 16.33 4.754 16.69 5.085 ;
      RECT 16.315 4.763 16.695 5.068 ;
      RECT 16.31 4.78 16.695 4.895 ;
      RECT 16.315 3.502 16.35 3.74 ;
      RECT 16.315 3.502 16.38 3.739 ;
      RECT 16.315 3.502 16.495 3.735 ;
      RECT 16.315 3.502 16.55 3.713 ;
      RECT 16.325 3.445 16.605 3.613 ;
      RECT 16.43 3.285 16.46 3.736 ;
      RECT 16.46 3.28 16.64 3.493 ;
      RECT 16.33 3.421 16.64 3.493 ;
      RECT 16.38 3.317 16.43 3.737 ;
      RECT 16.35 3.373 16.64 3.493 ;
      RECT 14.145 10.29 14.315 10.74 ;
      RECT 14.2 8.51 14.37 10.46 ;
      RECT 14.145 7.45 14.315 8.68 ;
      RECT 13.625 7.45 13.795 10.74 ;
      RECT 13.625 9.75 14.03 10.08 ;
      RECT 13.625 8.91 14.03 9.24 ;
      RECT 104.845 7.455 105.015 8.925 ;
      RECT 104.845 10.235 105.015 10.745 ;
      RECT 103.855 1.865 104.025 2.375 ;
      RECT 103.855 3.685 104.025 5.155 ;
      RECT 103.855 7.455 104.025 8.925 ;
      RECT 103.855 10.235 104.025 10.745 ;
      RECT 102.495 1.87 102.665 5.16 ;
      RECT 102.495 7.45 102.665 10.74 ;
      RECT 102.065 1.87 102.235 2.38 ;
      RECT 102.065 2.95 102.235 5.16 ;
      RECT 102.065 7.45 102.235 9.66 ;
      RECT 102.065 10.23 102.235 10.74 ;
      RECT 97.735 7.45 97.905 10.74 ;
      RECT 97.305 7.45 97.475 9.66 ;
      RECT 97.305 10.23 97.475 10.74 ;
      RECT 86.92 7.455 87.09 8.925 ;
      RECT 86.92 10.235 87.09 10.745 ;
      RECT 85.93 1.865 86.1 2.375 ;
      RECT 85.93 3.685 86.1 5.155 ;
      RECT 85.93 7.455 86.1 8.925 ;
      RECT 85.93 10.235 86.1 10.745 ;
      RECT 84.57 1.87 84.74 5.16 ;
      RECT 84.57 7.45 84.74 10.74 ;
      RECT 84.14 1.87 84.31 2.38 ;
      RECT 84.14 2.95 84.31 5.16 ;
      RECT 84.14 7.45 84.31 9.66 ;
      RECT 84.14 10.23 84.31 10.74 ;
      RECT 79.81 7.45 79.98 10.74 ;
      RECT 79.38 7.45 79.55 9.66 ;
      RECT 79.38 10.23 79.55 10.74 ;
      RECT 68.995 7.455 69.165 8.925 ;
      RECT 68.995 10.235 69.165 10.745 ;
      RECT 68.005 1.865 68.175 2.375 ;
      RECT 68.005 3.685 68.175 5.155 ;
      RECT 68.005 7.455 68.175 8.925 ;
      RECT 68.005 10.235 68.175 10.745 ;
      RECT 66.645 1.87 66.815 5.16 ;
      RECT 66.645 7.45 66.815 10.74 ;
      RECT 66.215 1.87 66.385 2.38 ;
      RECT 66.215 2.95 66.385 5.16 ;
      RECT 66.215 7.45 66.385 9.66 ;
      RECT 66.215 10.23 66.385 10.74 ;
      RECT 61.885 7.45 62.055 10.74 ;
      RECT 61.455 7.45 61.625 9.66 ;
      RECT 61.455 10.23 61.625 10.74 ;
      RECT 51.07 7.455 51.24 8.925 ;
      RECT 51.07 10.235 51.24 10.745 ;
      RECT 50.08 1.865 50.25 2.375 ;
      RECT 50.08 3.685 50.25 5.155 ;
      RECT 50.08 7.455 50.25 8.925 ;
      RECT 50.08 10.235 50.25 10.745 ;
      RECT 48.72 1.87 48.89 5.16 ;
      RECT 48.72 7.45 48.89 10.74 ;
      RECT 48.29 1.87 48.46 2.38 ;
      RECT 48.29 2.95 48.46 5.16 ;
      RECT 48.29 7.45 48.46 9.66 ;
      RECT 48.29 10.23 48.46 10.74 ;
      RECT 43.96 7.45 44.13 10.74 ;
      RECT 43.53 7.45 43.7 9.66 ;
      RECT 43.53 10.23 43.7 10.74 ;
      RECT 33.145 7.455 33.315 8.925 ;
      RECT 33.145 10.235 33.315 10.745 ;
      RECT 32.155 1.865 32.325 2.375 ;
      RECT 32.155 3.685 32.325 5.155 ;
      RECT 32.155 7.455 32.325 8.925 ;
      RECT 32.155 10.235 32.325 10.745 ;
      RECT 30.795 1.87 30.965 5.16 ;
      RECT 30.795 7.45 30.965 10.74 ;
      RECT 30.365 1.87 30.535 2.38 ;
      RECT 30.365 2.95 30.535 5.16 ;
      RECT 30.365 7.45 30.535 9.66 ;
      RECT 30.365 10.23 30.535 10.74 ;
      RECT 26.035 7.45 26.205 10.74 ;
      RECT 25.605 7.45 25.775 9.66 ;
      RECT 25.605 10.23 25.775 10.74 ;
      RECT 14.575 7.45 14.745 9.66 ;
      RECT 14.575 10.23 14.745 10.74 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r2 ;
  SIZE 92.605 BY 12.61 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 20.355 1.865 20.525 2.375 ;
        RECT 20.355 3.685 20.525 5.155 ;
      LAYER met1 ;
        RECT 20.295 3.655 20.585 3.885 ;
        RECT 20.295 2.175 20.585 2.405 ;
        RECT 20.355 2.175 20.525 3.885 ;
      LAYER mcon ;
        RECT 20.355 3.685 20.525 3.855 ;
        RECT 20.355 2.205 20.525 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 38.28 1.865 38.45 2.375 ;
        RECT 38.28 3.685 38.45 5.155 ;
      LAYER met1 ;
        RECT 38.22 3.655 38.51 3.885 ;
        RECT 38.22 2.175 38.51 2.405 ;
        RECT 38.28 2.175 38.45 3.885 ;
      LAYER mcon ;
        RECT 38.28 3.685 38.45 3.855 ;
        RECT 38.28 2.205 38.45 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 56.205 1.865 56.375 2.375 ;
        RECT 56.205 3.685 56.375 5.155 ;
      LAYER met1 ;
        RECT 56.145 3.655 56.435 3.885 ;
        RECT 56.145 2.175 56.435 2.405 ;
        RECT 56.205 2.175 56.375 3.885 ;
      LAYER mcon ;
        RECT 56.205 3.685 56.375 3.855 ;
        RECT 56.205 2.205 56.375 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 74.13 1.865 74.3 2.375 ;
        RECT 74.13 3.685 74.3 5.155 ;
      LAYER met1 ;
        RECT 74.07 3.655 74.36 3.885 ;
        RECT 74.07 2.175 74.36 2.405 ;
        RECT 74.13 2.175 74.3 3.885 ;
      LAYER mcon ;
        RECT 74.13 3.685 74.3 3.855 ;
        RECT 74.13 2.205 74.3 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 92.055 1.865 92.225 2.375 ;
        RECT 92.055 3.685 92.225 5.155 ;
      LAYER met1 ;
        RECT 91.995 3.655 92.285 3.885 ;
        RECT 91.995 2.175 92.285 2.405 ;
        RECT 92.055 2.175 92.225 3.885 ;
      LAYER mcon ;
        RECT 92.055 3.685 92.225 3.855 ;
        RECT 92.055 2.205 92.225 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 16.205 2.955 16.375 4.23 ;
        RECT 16.205 8.38 16.375 9.655 ;
        RECT 11.445 8.38 11.615 9.655 ;
      LAYER met2 ;
        RECT 16.125 4 16.475 4.35 ;
        RECT 16.115 8.275 16.465 8.625 ;
        RECT 16.19 4 16.365 8.625 ;
      LAYER met1 ;
        RECT 16.125 4.06 16.605 4.23 ;
        RECT 16.125 4 16.475 4.35 ;
        RECT 11.385 8.38 16.605 8.55 ;
        RECT 16.115 8.275 16.465 8.625 ;
        RECT 11.385 8.35 11.675 8.58 ;
      LAYER via1 ;
        RECT 16.215 8.375 16.365 8.525 ;
        RECT 16.225 4.1 16.375 4.25 ;
      LAYER mcon ;
        RECT 11.445 8.38 11.615 8.55 ;
        RECT 16.205 8.38 16.375 8.55 ;
        RECT 16.205 4.06 16.375 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 34.13 2.955 34.3 4.23 ;
        RECT 34.13 8.38 34.3 9.655 ;
        RECT 29.37 8.38 29.54 9.655 ;
      LAYER met2 ;
        RECT 34.05 4 34.4 4.35 ;
        RECT 34.04 8.275 34.39 8.625 ;
        RECT 34.115 4 34.29 8.625 ;
      LAYER met1 ;
        RECT 34.05 4.06 34.53 4.23 ;
        RECT 34.05 4 34.4 4.35 ;
        RECT 29.31 8.38 34.53 8.55 ;
        RECT 34.04 8.275 34.39 8.625 ;
        RECT 29.31 8.35 29.6 8.58 ;
      LAYER via1 ;
        RECT 34.14 8.375 34.29 8.525 ;
        RECT 34.15 4.1 34.3 4.25 ;
      LAYER mcon ;
        RECT 29.37 8.38 29.54 8.55 ;
        RECT 34.13 8.38 34.3 8.55 ;
        RECT 34.13 4.06 34.3 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 52.055 2.955 52.225 4.23 ;
        RECT 52.055 8.38 52.225 9.655 ;
        RECT 47.295 8.38 47.465 9.655 ;
      LAYER met2 ;
        RECT 51.975 4 52.325 4.35 ;
        RECT 51.965 8.275 52.315 8.625 ;
        RECT 52.04 4 52.215 8.625 ;
      LAYER met1 ;
        RECT 51.975 4.06 52.455 4.23 ;
        RECT 51.975 4 52.325 4.35 ;
        RECT 47.235 8.38 52.455 8.55 ;
        RECT 51.965 8.275 52.315 8.625 ;
        RECT 47.235 8.35 47.525 8.58 ;
      LAYER via1 ;
        RECT 52.065 8.375 52.215 8.525 ;
        RECT 52.075 4.1 52.225 4.25 ;
      LAYER mcon ;
        RECT 47.295 8.38 47.465 8.55 ;
        RECT 52.055 8.38 52.225 8.55 ;
        RECT 52.055 4.06 52.225 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 69.98 2.955 70.15 4.23 ;
        RECT 69.98 8.38 70.15 9.655 ;
        RECT 65.22 8.38 65.39 9.655 ;
      LAYER met2 ;
        RECT 69.9 4 70.25 4.35 ;
        RECT 69.89 8.275 70.24 8.625 ;
        RECT 69.965 4 70.14 8.625 ;
      LAYER met1 ;
        RECT 69.9 4.06 70.38 4.23 ;
        RECT 69.9 4 70.25 4.35 ;
        RECT 65.16 8.38 70.38 8.55 ;
        RECT 69.89 8.275 70.24 8.625 ;
        RECT 65.16 8.35 65.45 8.58 ;
      LAYER via1 ;
        RECT 69.99 8.375 70.14 8.525 ;
        RECT 70 4.1 70.15 4.25 ;
      LAYER mcon ;
        RECT 65.22 8.38 65.39 8.55 ;
        RECT 69.98 8.38 70.15 8.55 ;
        RECT 69.98 4.06 70.15 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 87.905 2.955 88.075 4.23 ;
        RECT 87.905 8.38 88.075 9.655 ;
        RECT 83.145 8.38 83.315 9.655 ;
      LAYER met2 ;
        RECT 87.825 4 88.175 4.35 ;
        RECT 87.815 8.275 88.165 8.625 ;
        RECT 87.89 4 88.065 8.625 ;
      LAYER met1 ;
        RECT 87.825 4.06 88.305 4.23 ;
        RECT 87.825 4 88.175 4.35 ;
        RECT 83.085 8.38 88.305 8.55 ;
        RECT 87.815 8.275 88.165 8.625 ;
        RECT 83.085 8.35 83.375 8.58 ;
      LAYER via1 ;
        RECT 87.915 8.375 88.065 8.525 ;
        RECT 87.925 4.1 88.075 4.25 ;
      LAYER mcon ;
        RECT 83.145 8.38 83.315 8.55 ;
        RECT 87.905 8.38 88.075 8.55 ;
        RECT 87.905 4.06 88.075 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.415 8.38 0.585 9.655 ;
      LAYER met1 ;
        RECT 0.355 8.38 0.815 8.55 ;
        RECT 0.355 8.35 0.645 8.58 ;
      LAYER mcon ;
        RECT 0.415 8.38 0.585 8.55 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.025 5.58 92.6 7.18 ;
        RECT 86.64 5.43 92.6 7.18 ;
        RECT 90.465 5.425 92.445 7.185 ;
        RECT 91.625 4.695 91.795 7.915 ;
        RECT 90.635 4.695 90.805 7.915 ;
        RECT 87.895 4.7 88.065 7.91 ;
        RECT 85.14 5.08 85.31 7.18 ;
        RECT 83.135 5.58 83.305 7.91 ;
        RECT 82.7 5.08 82.87 7.18 ;
        RECT 80.74 5.08 80.91 7.18 ;
        RECT 79.78 5.08 79.95 7.18 ;
        RECT 77.82 5.08 77.99 7.18 ;
        RECT 76.82 5.08 76.99 7.18 ;
        RECT 75.86 5.08 76.03 7.18 ;
        RECT 68.715 5.43 74.675 7.18 ;
        RECT 72.54 5.425 74.52 7.185 ;
        RECT 73.7 4.695 73.87 7.915 ;
        RECT 72.71 4.695 72.88 7.915 ;
        RECT 69.97 4.7 70.14 7.91 ;
        RECT 67.215 5.08 67.385 7.18 ;
        RECT 65.21 5.58 65.38 7.91 ;
        RECT 64.775 5.08 64.945 7.18 ;
        RECT 62.815 5.08 62.985 7.18 ;
        RECT 61.855 5.08 62.025 7.18 ;
        RECT 59.895 5.08 60.065 7.18 ;
        RECT 58.895 5.08 59.065 7.18 ;
        RECT 57.935 5.08 58.105 7.18 ;
        RECT 50.79 5.43 56.75 7.18 ;
        RECT 54.615 5.425 56.595 7.185 ;
        RECT 55.775 4.695 55.945 7.915 ;
        RECT 54.785 4.695 54.955 7.915 ;
        RECT 52.045 4.7 52.215 7.91 ;
        RECT 49.29 5.08 49.46 7.18 ;
        RECT 47.285 5.58 47.455 7.91 ;
        RECT 46.85 5.08 47.02 7.18 ;
        RECT 44.89 5.08 45.06 7.18 ;
        RECT 43.93 5.08 44.1 7.18 ;
        RECT 41.97 5.08 42.14 7.18 ;
        RECT 40.97 5.08 41.14 7.18 ;
        RECT 40.01 5.08 40.18 7.18 ;
        RECT 32.865 5.43 38.825 7.18 ;
        RECT 36.69 5.425 38.67 7.185 ;
        RECT 37.85 4.695 38.02 7.915 ;
        RECT 36.86 4.695 37.03 7.915 ;
        RECT 34.12 4.7 34.29 7.91 ;
        RECT 31.365 5.08 31.535 7.18 ;
        RECT 29.36 5.58 29.53 7.91 ;
        RECT 28.925 5.08 29.095 7.18 ;
        RECT 26.965 5.08 27.135 7.18 ;
        RECT 26.005 5.08 26.175 7.18 ;
        RECT 24.045 5.08 24.215 7.18 ;
        RECT 23.045 5.08 23.215 7.18 ;
        RECT 22.085 5.08 22.255 7.18 ;
        RECT 14.94 5.43 20.9 7.18 ;
        RECT 18.765 5.425 20.745 7.185 ;
        RECT 19.925 4.695 20.095 7.915 ;
        RECT 18.935 4.695 19.105 7.915 ;
        RECT 16.195 4.7 16.365 7.91 ;
        RECT 13.44 5.08 13.61 7.18 ;
        RECT 11.435 5.58 11.605 7.91 ;
        RECT 11 5.08 11.17 7.18 ;
        RECT 9.04 5.08 9.21 7.18 ;
        RECT 8.08 5.08 8.25 7.18 ;
        RECT 6.12 5.08 6.29 7.18 ;
        RECT 5.12 5.08 5.29 7.18 ;
        RECT 4.16 5.08 4.33 7.18 ;
        RECT 2.215 5.58 2.385 10.74 ;
        RECT 0.405 5.58 0.575 7.91 ;
      LAYER met1 ;
        RECT 0.025 5.58 92.6 7.18 ;
        RECT 75.05 5.43 92.6 7.18 ;
        RECT 90.465 5.425 92.445 7.185 ;
        RECT 75.05 5.425 87.01 7.18 ;
        RECT 57.125 5.43 74.675 7.18 ;
        RECT 72.54 5.425 74.52 7.185 ;
        RECT 57.125 5.425 69.085 7.18 ;
        RECT 39.2 5.43 56.75 7.18 ;
        RECT 54.615 5.425 56.595 7.185 ;
        RECT 39.2 5.425 51.16 7.18 ;
        RECT 21.275 5.43 38.825 7.18 ;
        RECT 36.69 5.425 38.67 7.185 ;
        RECT 21.275 5.425 33.235 7.18 ;
        RECT 3.35 5.43 20.9 7.18 ;
        RECT 18.765 5.425 20.745 7.185 ;
        RECT 3.35 5.425 15.31 7.18 ;
        RECT 2.155 9.09 2.445 9.32 ;
        RECT 1.985 9.12 2.445 9.29 ;
      LAYER mcon ;
        RECT 2.215 9.12 2.385 9.29 ;
        RECT 2.525 6.98 2.695 7.15 ;
        RECT 3.495 5.58 3.665 5.75 ;
        RECT 3.955 5.58 4.125 5.75 ;
        RECT 4.415 5.58 4.585 5.75 ;
        RECT 4.875 5.58 5.045 5.75 ;
        RECT 5.335 5.58 5.505 5.75 ;
        RECT 5.795 5.58 5.965 5.75 ;
        RECT 6.255 5.58 6.425 5.75 ;
        RECT 6.715 5.58 6.885 5.75 ;
        RECT 7.175 5.58 7.345 5.75 ;
        RECT 7.635 5.58 7.805 5.75 ;
        RECT 8.095 5.58 8.265 5.75 ;
        RECT 8.555 5.58 8.725 5.75 ;
        RECT 9.015 5.58 9.185 5.75 ;
        RECT 9.475 5.58 9.645 5.75 ;
        RECT 9.935 5.58 10.105 5.75 ;
        RECT 10.395 5.58 10.565 5.75 ;
        RECT 10.855 5.58 11.025 5.75 ;
        RECT 11.315 5.58 11.485 5.75 ;
        RECT 11.775 5.58 11.945 5.75 ;
        RECT 12.235 5.58 12.405 5.75 ;
        RECT 12.695 5.58 12.865 5.75 ;
        RECT 13.155 5.58 13.325 5.75 ;
        RECT 13.555 6.98 13.725 7.15 ;
        RECT 13.615 5.58 13.785 5.75 ;
        RECT 14.075 5.58 14.245 5.75 ;
        RECT 14.535 5.58 14.705 5.75 ;
        RECT 14.995 5.58 15.165 5.75 ;
        RECT 18.315 6.98 18.485 7.15 ;
        RECT 18.315 5.46 18.485 5.63 ;
        RECT 19.015 6.985 19.185 7.155 ;
        RECT 19.015 5.455 19.185 5.625 ;
        RECT 20.005 6.985 20.175 7.155 ;
        RECT 20.005 5.455 20.175 5.625 ;
        RECT 21.42 5.58 21.59 5.75 ;
        RECT 21.88 5.58 22.05 5.75 ;
        RECT 22.34 5.58 22.51 5.75 ;
        RECT 22.8 5.58 22.97 5.75 ;
        RECT 23.26 5.58 23.43 5.75 ;
        RECT 23.72 5.58 23.89 5.75 ;
        RECT 24.18 5.58 24.35 5.75 ;
        RECT 24.64 5.58 24.81 5.75 ;
        RECT 25.1 5.58 25.27 5.75 ;
        RECT 25.56 5.58 25.73 5.75 ;
        RECT 26.02 5.58 26.19 5.75 ;
        RECT 26.48 5.58 26.65 5.75 ;
        RECT 26.94 5.58 27.11 5.75 ;
        RECT 27.4 5.58 27.57 5.75 ;
        RECT 27.86 5.58 28.03 5.75 ;
        RECT 28.32 5.58 28.49 5.75 ;
        RECT 28.78 5.58 28.95 5.75 ;
        RECT 29.24 5.58 29.41 5.75 ;
        RECT 29.7 5.58 29.87 5.75 ;
        RECT 30.16 5.58 30.33 5.75 ;
        RECT 30.62 5.58 30.79 5.75 ;
        RECT 31.08 5.58 31.25 5.75 ;
        RECT 31.48 6.98 31.65 7.15 ;
        RECT 31.54 5.58 31.71 5.75 ;
        RECT 32 5.58 32.17 5.75 ;
        RECT 32.46 5.58 32.63 5.75 ;
        RECT 32.92 5.58 33.09 5.75 ;
        RECT 36.24 6.98 36.41 7.15 ;
        RECT 36.24 5.46 36.41 5.63 ;
        RECT 36.94 6.985 37.11 7.155 ;
        RECT 36.94 5.455 37.11 5.625 ;
        RECT 37.93 6.985 38.1 7.155 ;
        RECT 37.93 5.455 38.1 5.625 ;
        RECT 39.345 5.58 39.515 5.75 ;
        RECT 39.805 5.58 39.975 5.75 ;
        RECT 40.265 5.58 40.435 5.75 ;
        RECT 40.725 5.58 40.895 5.75 ;
        RECT 41.185 5.58 41.355 5.75 ;
        RECT 41.645 5.58 41.815 5.75 ;
        RECT 42.105 5.58 42.275 5.75 ;
        RECT 42.565 5.58 42.735 5.75 ;
        RECT 43.025 5.58 43.195 5.75 ;
        RECT 43.485 5.58 43.655 5.75 ;
        RECT 43.945 5.58 44.115 5.75 ;
        RECT 44.405 5.58 44.575 5.75 ;
        RECT 44.865 5.58 45.035 5.75 ;
        RECT 45.325 5.58 45.495 5.75 ;
        RECT 45.785 5.58 45.955 5.75 ;
        RECT 46.245 5.58 46.415 5.75 ;
        RECT 46.705 5.58 46.875 5.75 ;
        RECT 47.165 5.58 47.335 5.75 ;
        RECT 47.625 5.58 47.795 5.75 ;
        RECT 48.085 5.58 48.255 5.75 ;
        RECT 48.545 5.58 48.715 5.75 ;
        RECT 49.005 5.58 49.175 5.75 ;
        RECT 49.405 6.98 49.575 7.15 ;
        RECT 49.465 5.58 49.635 5.75 ;
        RECT 49.925 5.58 50.095 5.75 ;
        RECT 50.385 5.58 50.555 5.75 ;
        RECT 50.845 5.58 51.015 5.75 ;
        RECT 54.165 6.98 54.335 7.15 ;
        RECT 54.165 5.46 54.335 5.63 ;
        RECT 54.865 6.985 55.035 7.155 ;
        RECT 54.865 5.455 55.035 5.625 ;
        RECT 55.855 6.985 56.025 7.155 ;
        RECT 55.855 5.455 56.025 5.625 ;
        RECT 57.27 5.58 57.44 5.75 ;
        RECT 57.73 5.58 57.9 5.75 ;
        RECT 58.19 5.58 58.36 5.75 ;
        RECT 58.65 5.58 58.82 5.75 ;
        RECT 59.11 5.58 59.28 5.75 ;
        RECT 59.57 5.58 59.74 5.75 ;
        RECT 60.03 5.58 60.2 5.75 ;
        RECT 60.49 5.58 60.66 5.75 ;
        RECT 60.95 5.58 61.12 5.75 ;
        RECT 61.41 5.58 61.58 5.75 ;
        RECT 61.87 5.58 62.04 5.75 ;
        RECT 62.33 5.58 62.5 5.75 ;
        RECT 62.79 5.58 62.96 5.75 ;
        RECT 63.25 5.58 63.42 5.75 ;
        RECT 63.71 5.58 63.88 5.75 ;
        RECT 64.17 5.58 64.34 5.75 ;
        RECT 64.63 5.58 64.8 5.75 ;
        RECT 65.09 5.58 65.26 5.75 ;
        RECT 65.55 5.58 65.72 5.75 ;
        RECT 66.01 5.58 66.18 5.75 ;
        RECT 66.47 5.58 66.64 5.75 ;
        RECT 66.93 5.58 67.1 5.75 ;
        RECT 67.33 6.98 67.5 7.15 ;
        RECT 67.39 5.58 67.56 5.75 ;
        RECT 67.85 5.58 68.02 5.75 ;
        RECT 68.31 5.58 68.48 5.75 ;
        RECT 68.77 5.58 68.94 5.75 ;
        RECT 72.09 6.98 72.26 7.15 ;
        RECT 72.09 5.46 72.26 5.63 ;
        RECT 72.79 6.985 72.96 7.155 ;
        RECT 72.79 5.455 72.96 5.625 ;
        RECT 73.78 6.985 73.95 7.155 ;
        RECT 73.78 5.455 73.95 5.625 ;
        RECT 75.195 5.58 75.365 5.75 ;
        RECT 75.655 5.58 75.825 5.75 ;
        RECT 76.115 5.58 76.285 5.75 ;
        RECT 76.575 5.58 76.745 5.75 ;
        RECT 77.035 5.58 77.205 5.75 ;
        RECT 77.495 5.58 77.665 5.75 ;
        RECT 77.955 5.58 78.125 5.75 ;
        RECT 78.415 5.58 78.585 5.75 ;
        RECT 78.875 5.58 79.045 5.75 ;
        RECT 79.335 5.58 79.505 5.75 ;
        RECT 79.795 5.58 79.965 5.75 ;
        RECT 80.255 5.58 80.425 5.75 ;
        RECT 80.715 5.58 80.885 5.75 ;
        RECT 81.175 5.58 81.345 5.75 ;
        RECT 81.635 5.58 81.805 5.75 ;
        RECT 82.095 5.58 82.265 5.75 ;
        RECT 82.555 5.58 82.725 5.75 ;
        RECT 83.015 5.58 83.185 5.75 ;
        RECT 83.475 5.58 83.645 5.75 ;
        RECT 83.935 5.58 84.105 5.75 ;
        RECT 84.395 5.58 84.565 5.75 ;
        RECT 84.855 5.58 85.025 5.75 ;
        RECT 85.255 6.98 85.425 7.15 ;
        RECT 85.315 5.58 85.485 5.75 ;
        RECT 85.775 5.58 85.945 5.75 ;
        RECT 86.235 5.58 86.405 5.75 ;
        RECT 86.695 5.58 86.865 5.75 ;
        RECT 90.015 6.98 90.185 7.15 ;
        RECT 90.015 5.46 90.185 5.63 ;
        RECT 90.715 6.985 90.885 7.155 ;
        RECT 90.715 5.455 90.885 5.625 ;
        RECT 91.705 6.985 91.875 7.155 ;
        RECT 91.705 5.455 91.875 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.05 11.445 92.605 12.61 ;
        RECT 0.055 11.01 92.605 12.61 ;
        RECT 91.625 10.385 91.795 12.61 ;
        RECT 90.635 10.385 90.805 12.61 ;
        RECT 87.895 10.38 88.065 12.61 ;
        RECT 83.135 10.38 83.305 12.61 ;
        RECT 73.7 10.385 73.87 12.61 ;
        RECT 72.71 10.385 72.88 12.61 ;
        RECT 69.97 10.38 70.14 12.61 ;
        RECT 65.21 10.38 65.38 12.61 ;
        RECT 55.775 10.385 55.945 12.61 ;
        RECT 54.785 10.385 54.955 12.61 ;
        RECT 52.045 10.38 52.215 12.61 ;
        RECT 47.285 10.38 47.455 12.61 ;
        RECT 37.85 10.385 38.02 12.61 ;
        RECT 36.86 10.385 37.03 12.61 ;
        RECT 34.12 10.38 34.29 12.61 ;
        RECT 29.36 10.38 29.53 12.61 ;
        RECT 19.925 10.385 20.095 12.61 ;
        RECT 18.935 10.385 19.105 12.61 ;
        RECT 16.195 10.38 16.365 12.61 ;
        RECT 11.435 10.38 11.605 12.61 ;
        RECT 0.405 10.38 0.575 12.61 ;
        RECT 84.14 8.51 84.31 10.46 ;
        RECT 84.085 10.29 84.255 10.74 ;
        RECT 84.085 7.45 84.255 8.68 ;
        RECT 66.215 8.51 66.385 10.46 ;
        RECT 66.16 10.29 66.33 10.74 ;
        RECT 66.16 7.45 66.33 8.68 ;
        RECT 48.29 8.51 48.46 10.46 ;
        RECT 48.235 10.29 48.405 10.74 ;
        RECT 48.235 7.45 48.405 8.68 ;
        RECT 30.365 8.51 30.535 10.46 ;
        RECT 30.31 10.29 30.48 10.74 ;
        RECT 30.31 7.45 30.48 8.68 ;
        RECT 12.44 8.51 12.61 10.46 ;
        RECT 12.385 10.29 12.555 10.74 ;
        RECT 12.385 7.45 12.555 8.68 ;
      LAYER met1 ;
        RECT 0.05 11.445 92.605 12.61 ;
        RECT 0.055 11.01 92.605 12.61 ;
        RECT 84.08 8.72 84.37 8.95 ;
        RECT 83.745 8.75 84.37 8.92 ;
        RECT 83.745 8.75 83.915 12.61 ;
        RECT 66.155 8.72 66.445 8.95 ;
        RECT 65.82 8.75 66.445 8.92 ;
        RECT 65.82 8.75 65.99 12.61 ;
        RECT 48.23 8.72 48.52 8.95 ;
        RECT 47.895 8.75 48.52 8.92 ;
        RECT 47.895 8.75 48.065 12.61 ;
        RECT 30.305 8.72 30.595 8.95 ;
        RECT 29.97 8.75 30.595 8.92 ;
        RECT 29.97 8.75 30.14 12.61 ;
        RECT 12.38 8.72 12.67 8.95 ;
        RECT 12.045 8.75 12.67 8.92 ;
        RECT 12.045 8.75 12.215 12.61 ;
      LAYER mcon ;
        RECT 0.485 11.04 0.655 11.21 ;
        RECT 1.165 11.04 1.335 11.21 ;
        RECT 1.845 11.04 2.015 11.21 ;
        RECT 2.525 11.04 2.695 11.21 ;
        RECT 11.515 11.04 11.685 11.21 ;
        RECT 12.195 11.04 12.365 11.21 ;
        RECT 12.44 8.75 12.61 8.92 ;
        RECT 12.875 11.04 13.045 11.21 ;
        RECT 13.555 11.04 13.725 11.21 ;
        RECT 16.275 11.04 16.445 11.21 ;
        RECT 16.955 11.04 17.125 11.21 ;
        RECT 17.635 11.04 17.805 11.21 ;
        RECT 18.315 11.04 18.485 11.21 ;
        RECT 19.015 11.045 19.185 11.215 ;
        RECT 20.005 11.045 20.175 11.215 ;
        RECT 29.44 11.04 29.61 11.21 ;
        RECT 30.12 11.04 30.29 11.21 ;
        RECT 30.365 8.75 30.535 8.92 ;
        RECT 30.8 11.04 30.97 11.21 ;
        RECT 31.48 11.04 31.65 11.21 ;
        RECT 34.2 11.04 34.37 11.21 ;
        RECT 34.88 11.04 35.05 11.21 ;
        RECT 35.56 11.04 35.73 11.21 ;
        RECT 36.24 11.04 36.41 11.21 ;
        RECT 36.94 11.045 37.11 11.215 ;
        RECT 37.93 11.045 38.1 11.215 ;
        RECT 47.365 11.04 47.535 11.21 ;
        RECT 48.045 11.04 48.215 11.21 ;
        RECT 48.29 8.75 48.46 8.92 ;
        RECT 48.725 11.04 48.895 11.21 ;
        RECT 49.405 11.04 49.575 11.21 ;
        RECT 52.125 11.04 52.295 11.21 ;
        RECT 52.805 11.04 52.975 11.21 ;
        RECT 53.485 11.04 53.655 11.21 ;
        RECT 54.165 11.04 54.335 11.21 ;
        RECT 54.865 11.045 55.035 11.215 ;
        RECT 55.855 11.045 56.025 11.215 ;
        RECT 65.29 11.04 65.46 11.21 ;
        RECT 65.97 11.04 66.14 11.21 ;
        RECT 66.215 8.75 66.385 8.92 ;
        RECT 66.65 11.04 66.82 11.21 ;
        RECT 67.33 11.04 67.5 11.21 ;
        RECT 70.05 11.04 70.22 11.21 ;
        RECT 70.73 11.04 70.9 11.21 ;
        RECT 71.41 11.04 71.58 11.21 ;
        RECT 72.09 11.04 72.26 11.21 ;
        RECT 72.79 11.045 72.96 11.215 ;
        RECT 73.78 11.045 73.95 11.215 ;
        RECT 83.215 11.04 83.385 11.21 ;
        RECT 83.895 11.04 84.065 11.21 ;
        RECT 84.14 8.75 84.31 8.92 ;
        RECT 84.575 11.04 84.745 11.21 ;
        RECT 85.255 11.04 85.425 11.21 ;
        RECT 87.975 11.04 88.145 11.21 ;
        RECT 88.655 11.04 88.825 11.21 ;
        RECT 89.335 11.04 89.505 11.21 ;
        RECT 90.015 11.04 90.185 11.21 ;
        RECT 90.715 11.045 90.885 11.215 ;
        RECT 91.705 11.045 91.875 11.215 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 84.405 9.49 84.78 9.86 ;
      RECT 84.44 7.36 84.75 9.86 ;
      RECT 84.44 7.36 87.535 7.67 ;
      RECT 87.225 2.42 87.535 7.67 ;
      RECT 87.225 2.435 87.6 2.805 ;
      RECT 84.355 4.98 84.91 5.31 ;
      RECT 84.355 3.315 84.655 5.31 ;
      RECT 80.42 4.42 80.975 4.75 ;
      RECT 80.675 3.315 80.975 4.75 ;
      RECT 81.47 3.18 81.62 3.83 ;
      RECT 80.675 3.315 84.655 3.615 ;
      RECT 79.19 2.255 79.49 5.205 ;
      RECT 79.18 3.86 79.91 4.19 ;
      RECT 79.145 2.255 79.52 2.625 ;
      RECT 77.74 4.42 78.47 4.75 ;
      RECT 77.755 2.255 78.055 4.75 ;
      RECT 75.63 3.86 76.36 4.19 ;
      RECT 75.785 2.225 76.085 4.19 ;
      RECT 77.71 2.255 78.085 2.625 ;
      RECT 75.74 2.225 76.115 2.595 ;
      RECT 75.74 2.265 78.085 2.565 ;
      RECT 66.48 9.49 66.855 9.86 ;
      RECT 66.515 7.36 66.825 9.86 ;
      RECT 66.515 7.36 69.61 7.67 ;
      RECT 69.3 2.42 69.61 7.67 ;
      RECT 69.3 2.435 69.675 2.805 ;
      RECT 66.43 4.98 66.985 5.31 ;
      RECT 66.43 3.315 66.73 5.31 ;
      RECT 62.495 4.42 63.05 4.75 ;
      RECT 62.75 3.315 63.05 4.75 ;
      RECT 63.545 3.18 63.695 3.83 ;
      RECT 62.75 3.315 66.73 3.615 ;
      RECT 61.265 2.255 61.565 5.205 ;
      RECT 61.255 3.86 61.985 4.19 ;
      RECT 61.22 2.255 61.595 2.625 ;
      RECT 59.815 4.42 60.545 4.75 ;
      RECT 59.83 2.255 60.13 4.75 ;
      RECT 57.705 3.86 58.435 4.19 ;
      RECT 57.86 2.225 58.16 4.19 ;
      RECT 59.785 2.255 60.16 2.625 ;
      RECT 57.815 2.225 58.19 2.595 ;
      RECT 57.815 2.265 60.16 2.565 ;
      RECT 48.555 9.49 48.93 9.86 ;
      RECT 48.59 7.36 48.9 9.86 ;
      RECT 48.59 7.36 51.685 7.67 ;
      RECT 51.375 2.42 51.685 7.67 ;
      RECT 51.375 2.435 51.75 2.805 ;
      RECT 48.505 4.98 49.06 5.31 ;
      RECT 48.505 3.315 48.805 5.31 ;
      RECT 44.57 4.42 45.125 4.75 ;
      RECT 44.825 3.315 45.125 4.75 ;
      RECT 45.62 3.18 45.77 3.83 ;
      RECT 44.825 3.315 48.805 3.615 ;
      RECT 43.34 2.255 43.64 5.205 ;
      RECT 43.33 3.86 44.06 4.19 ;
      RECT 43.295 2.255 43.67 2.625 ;
      RECT 41.89 4.42 42.62 4.75 ;
      RECT 41.905 2.255 42.205 4.75 ;
      RECT 39.78 3.86 40.51 4.19 ;
      RECT 39.935 2.225 40.235 4.19 ;
      RECT 41.86 2.255 42.235 2.625 ;
      RECT 39.89 2.225 40.265 2.595 ;
      RECT 39.89 2.265 42.235 2.565 ;
      RECT 30.63 9.49 31.005 9.86 ;
      RECT 30.665 7.36 30.975 9.86 ;
      RECT 30.665 7.36 33.76 7.67 ;
      RECT 33.45 2.42 33.76 7.67 ;
      RECT 33.45 2.435 33.825 2.805 ;
      RECT 30.58 4.98 31.135 5.31 ;
      RECT 30.58 3.315 30.88 5.31 ;
      RECT 26.645 4.42 27.2 4.75 ;
      RECT 26.9 3.315 27.2 4.75 ;
      RECT 27.695 3.18 27.845 3.83 ;
      RECT 26.9 3.315 30.88 3.615 ;
      RECT 25.415 2.255 25.715 5.205 ;
      RECT 25.405 3.86 26.135 4.19 ;
      RECT 25.37 2.255 25.745 2.625 ;
      RECT 23.965 4.42 24.695 4.75 ;
      RECT 23.98 2.255 24.28 4.75 ;
      RECT 21.855 3.86 22.585 4.19 ;
      RECT 22.01 2.225 22.31 4.19 ;
      RECT 23.935 2.255 24.31 2.625 ;
      RECT 21.965 2.225 22.34 2.595 ;
      RECT 21.965 2.265 24.31 2.565 ;
      RECT 12.705 9.49 13.08 9.86 ;
      RECT 12.74 7.36 13.05 9.86 ;
      RECT 12.74 7.36 15.835 7.67 ;
      RECT 15.525 2.42 15.835 7.67 ;
      RECT 15.525 2.435 15.9 2.805 ;
      RECT 12.655 4.98 13.21 5.31 ;
      RECT 12.655 3.315 12.955 5.31 ;
      RECT 8.72 4.42 9.275 4.75 ;
      RECT 8.975 3.315 9.275 4.75 ;
      RECT 9.77 3.18 9.92 3.83 ;
      RECT 8.975 3.315 12.955 3.615 ;
      RECT 7.49 2.255 7.79 5.205 ;
      RECT 7.48 3.86 8.21 4.19 ;
      RECT 7.445 2.255 7.82 2.625 ;
      RECT 6.04 4.42 6.77 4.75 ;
      RECT 6.055 2.255 6.355 4.75 ;
      RECT 3.93 3.86 4.66 4.19 ;
      RECT 4.085 2.225 4.385 4.19 ;
      RECT 6.01 2.255 6.385 2.625 ;
      RECT 4.04 2.225 4.415 2.595 ;
      RECT 4.04 2.265 6.385 2.565 ;
      RECT 85.54 3.3 86.27 3.63 ;
      RECT 83.32 4.98 84.05 5.31 ;
      RECT 81.62 4.98 82.35 5.31 ;
      RECT 76.665 3.86 77.395 4.19 ;
      RECT 75.3 4.98 76.03 5.31 ;
      RECT 67.615 3.3 68.345 3.63 ;
      RECT 65.395 4.98 66.125 5.31 ;
      RECT 63.695 4.98 64.425 5.31 ;
      RECT 58.74 3.86 59.47 4.19 ;
      RECT 57.375 4.98 58.105 5.31 ;
      RECT 49.69 3.3 50.42 3.63 ;
      RECT 47.47 4.98 48.2 5.31 ;
      RECT 45.77 4.98 46.5 5.31 ;
      RECT 40.815 3.86 41.545 4.19 ;
      RECT 39.45 4.98 40.18 5.31 ;
      RECT 31.765 3.3 32.495 3.63 ;
      RECT 29.545 4.98 30.275 5.31 ;
      RECT 27.845 4.98 28.575 5.31 ;
      RECT 22.89 3.86 23.62 4.19 ;
      RECT 21.525 4.98 22.255 5.31 ;
      RECT 13.84 3.3 14.57 3.63 ;
      RECT 11.62 4.98 12.35 5.31 ;
      RECT 9.92 4.98 10.65 5.31 ;
      RECT 4.965 3.86 5.695 4.19 ;
      RECT 3.6 4.98 4.33 5.31 ;
    LAYER via2 ;
      RECT 87.315 2.52 87.515 2.72 ;
      RECT 85.605 3.365 85.805 3.565 ;
      RECT 84.645 5.045 84.845 5.245 ;
      RECT 84.495 9.575 84.695 9.775 ;
      RECT 83.645 5.045 83.845 5.245 ;
      RECT 81.685 5.045 81.885 5.245 ;
      RECT 80.485 4.485 80.685 4.685 ;
      RECT 79.245 3.925 79.445 4.125 ;
      RECT 79.235 2.34 79.435 2.54 ;
      RECT 77.805 4.485 78.005 4.685 ;
      RECT 77.8 2.335 78 2.535 ;
      RECT 77.065 3.925 77.265 4.125 ;
      RECT 75.845 3.925 76.045 4.125 ;
      RECT 75.83 2.31 76.03 2.51 ;
      RECT 75.365 5.045 75.565 5.245 ;
      RECT 69.39 2.52 69.59 2.72 ;
      RECT 67.68 3.365 67.88 3.565 ;
      RECT 66.72 5.045 66.92 5.245 ;
      RECT 66.57 9.575 66.77 9.775 ;
      RECT 65.72 5.045 65.92 5.245 ;
      RECT 63.76 5.045 63.96 5.245 ;
      RECT 62.56 4.485 62.76 4.685 ;
      RECT 61.32 3.925 61.52 4.125 ;
      RECT 61.31 2.34 61.51 2.54 ;
      RECT 59.88 4.485 60.08 4.685 ;
      RECT 59.875 2.335 60.075 2.535 ;
      RECT 59.14 3.925 59.34 4.125 ;
      RECT 57.92 3.925 58.12 4.125 ;
      RECT 57.905 2.31 58.105 2.51 ;
      RECT 57.44 5.045 57.64 5.245 ;
      RECT 51.465 2.52 51.665 2.72 ;
      RECT 49.755 3.365 49.955 3.565 ;
      RECT 48.795 5.045 48.995 5.245 ;
      RECT 48.645 9.575 48.845 9.775 ;
      RECT 47.795 5.045 47.995 5.245 ;
      RECT 45.835 5.045 46.035 5.245 ;
      RECT 44.635 4.485 44.835 4.685 ;
      RECT 43.395 3.925 43.595 4.125 ;
      RECT 43.385 2.34 43.585 2.54 ;
      RECT 41.955 4.485 42.155 4.685 ;
      RECT 41.95 2.335 42.15 2.535 ;
      RECT 41.215 3.925 41.415 4.125 ;
      RECT 39.995 3.925 40.195 4.125 ;
      RECT 39.98 2.31 40.18 2.51 ;
      RECT 39.515 5.045 39.715 5.245 ;
      RECT 33.54 2.52 33.74 2.72 ;
      RECT 31.83 3.365 32.03 3.565 ;
      RECT 30.87 5.045 31.07 5.245 ;
      RECT 30.72 9.575 30.92 9.775 ;
      RECT 29.87 5.045 30.07 5.245 ;
      RECT 27.91 5.045 28.11 5.245 ;
      RECT 26.71 4.485 26.91 4.685 ;
      RECT 25.47 3.925 25.67 4.125 ;
      RECT 25.46 2.34 25.66 2.54 ;
      RECT 24.03 4.485 24.23 4.685 ;
      RECT 24.025 2.335 24.225 2.535 ;
      RECT 23.29 3.925 23.49 4.125 ;
      RECT 22.07 3.925 22.27 4.125 ;
      RECT 22.055 2.31 22.255 2.51 ;
      RECT 21.59 5.045 21.79 5.245 ;
      RECT 15.615 2.52 15.815 2.72 ;
      RECT 13.905 3.365 14.105 3.565 ;
      RECT 12.945 5.045 13.145 5.245 ;
      RECT 12.795 9.575 12.995 9.775 ;
      RECT 11.945 5.045 12.145 5.245 ;
      RECT 9.985 5.045 10.185 5.245 ;
      RECT 8.785 4.485 8.985 4.685 ;
      RECT 7.545 3.925 7.745 4.125 ;
      RECT 7.535 2.34 7.735 2.54 ;
      RECT 6.105 4.485 6.305 4.685 ;
      RECT 6.1 2.335 6.3 2.535 ;
      RECT 5.365 3.925 5.565 4.125 ;
      RECT 4.145 3.925 4.345 4.125 ;
      RECT 4.13 2.31 4.33 2.51 ;
      RECT 3.665 5.045 3.865 5.245 ;
    LAYER met2 ;
      RECT 1.41 10.835 92.225 11.005 ;
      RECT 92.055 9.71 92.225 11.005 ;
      RECT 1.41 8.69 1.58 11.005 ;
      RECT 92.025 9.71 92.375 10.06 ;
      RECT 1.35 8.69 1.64 9.04 ;
      RECT 88.87 8.66 89.19 8.98 ;
      RECT 88.9 8.13 89.07 8.98 ;
      RECT 88.9 8.13 89.075 8.48 ;
      RECT 88.9 8.13 89.875 8.305 ;
      RECT 89.7 3.26 89.875 8.305 ;
      RECT 89.645 3.26 89.995 3.61 ;
      RECT 89.67 9.09 89.995 9.415 ;
      RECT 88.555 9.18 89.995 9.35 ;
      RECT 88.555 3.69 88.715 9.35 ;
      RECT 88.87 3.66 89.19 3.98 ;
      RECT 88.555 3.69 89.19 3.86 ;
      RECT 87.225 2.435 87.6 2.805 ;
      RECT 79.145 2.255 79.52 2.625 ;
      RECT 77.71 2.255 78.085 2.625 ;
      RECT 77.71 2.375 87.53 2.545 ;
      RECT 81.83 5.655 87.51 5.825 ;
      RECT 87.34 4.72 87.51 5.825 ;
      RECT 81.64 4.895 81.665 5.825 ;
      RECT 81.895 5.005 81.925 5.285 ;
      RECT 81.6 4.895 81.665 5.155 ;
      RECT 87.25 4.725 87.6 5.075 ;
      RECT 81.43 3.52 81.465 3.78 ;
      RECT 81.205 3.52 81.265 3.78 ;
      RECT 81.885 4.985 81.895 5.285 ;
      RECT 81.88 4.945 81.885 5.285 ;
      RECT 81.865 4.9 81.88 5.285 ;
      RECT 81.86 4.865 81.865 5.285 ;
      RECT 81.855 4.845 81.86 5.285 ;
      RECT 81.83 4.782 81.855 5.285 ;
      RECT 81.825 4.72 81.83 5.825 ;
      RECT 81.805 4.67 81.825 5.825 ;
      RECT 81.795 4.6 81.805 5.825 ;
      RECT 81.75 4.54 81.795 5.825 ;
      RECT 81.665 4.501 81.75 5.825 ;
      RECT 81.66 4.492 81.665 4.865 ;
      RECT 81.65 4.491 81.66 4.848 ;
      RECT 81.625 4.472 81.65 4.818 ;
      RECT 81.62 4.447 81.625 4.797 ;
      RECT 81.61 4.425 81.62 4.788 ;
      RECT 81.605 4.396 81.61 4.778 ;
      RECT 81.565 4.322 81.605 4.75 ;
      RECT 81.545 4.223 81.565 4.715 ;
      RECT 81.53 4.159 81.545 4.698 ;
      RECT 81.5 4.083 81.53 4.67 ;
      RECT 81.48 3.998 81.5 4.643 ;
      RECT 81.44 3.894 81.48 4.55 ;
      RECT 81.435 3.815 81.44 4.458 ;
      RECT 81.43 3.798 81.435 4.435 ;
      RECT 81.425 3.52 81.43 4.415 ;
      RECT 81.395 3.52 81.425 4.353 ;
      RECT 81.39 3.52 81.395 4.285 ;
      RECT 81.38 3.52 81.39 4.25 ;
      RECT 81.37 3.52 81.38 4.215 ;
      RECT 81.305 3.52 81.37 4.07 ;
      RECT 81.3 3.52 81.305 3.94 ;
      RECT 81.27 3.52 81.3 3.873 ;
      RECT 81.265 3.52 81.27 3.798 ;
      RECT 85.6 3.455 85.86 3.715 ;
      RECT 85.595 3.455 85.86 3.663 ;
      RECT 85.59 3.455 85.86 3.633 ;
      RECT 85.565 3.325 85.845 3.605 ;
      RECT 74.08 9.09 74.43 9.44 ;
      RECT 85.325 9.045 85.675 9.395 ;
      RECT 74.08 9.12 85.675 9.32 ;
      RECT 84.605 5.005 84.885 5.285 ;
      RECT 84.645 4.96 84.91 5.22 ;
      RECT 84.635 4.995 84.91 5.22 ;
      RECT 84.64 4.98 84.885 5.285 ;
      RECT 84.645 4.957 84.855 5.285 ;
      RECT 84.645 4.955 84.84 5.285 ;
      RECT 84.685 4.945 84.84 5.285 ;
      RECT 84.655 4.95 84.84 5.285 ;
      RECT 84.685 4.942 84.785 5.285 ;
      RECT 84.71 4.935 84.785 5.285 ;
      RECT 84.69 4.937 84.785 5.285 ;
      RECT 84.02 4.45 84.28 4.71 ;
      RECT 84.07 4.442 84.26 4.71 ;
      RECT 84.075 4.362 84.26 4.71 ;
      RECT 84.195 3.75 84.26 4.71 ;
      RECT 84.1 4.147 84.26 4.71 ;
      RECT 84.175 3.835 84.26 4.71 ;
      RECT 84.21 3.46 84.346 4.188 ;
      RECT 84.155 3.957 84.346 4.188 ;
      RECT 84.17 3.897 84.26 4.71 ;
      RECT 84.21 3.46 84.37 3.853 ;
      RECT 84.21 3.46 84.38 3.75 ;
      RECT 84.2 3.46 84.46 3.72 ;
      RECT 83.605 5.005 83.885 5.285 ;
      RECT 83.625 4.965 83.885 5.285 ;
      RECT 83.265 4.92 83.37 5.18 ;
      RECT 83.12 3.41 83.21 3.67 ;
      RECT 83.66 4.475 83.665 4.515 ;
      RECT 83.655 4.465 83.66 4.6 ;
      RECT 83.65 4.455 83.655 4.693 ;
      RECT 83.64 4.435 83.65 4.749 ;
      RECT 83.56 4.363 83.64 4.829 ;
      RECT 83.595 5.007 83.605 5.232 ;
      RECT 83.59 5.004 83.595 5.227 ;
      RECT 83.575 5.001 83.59 5.22 ;
      RECT 83.54 4.995 83.575 5.202 ;
      RECT 83.555 4.298 83.56 4.903 ;
      RECT 83.535 4.249 83.555 4.918 ;
      RECT 83.525 4.982 83.54 5.185 ;
      RECT 83.53 4.191 83.535 4.933 ;
      RECT 83.525 4.169 83.53 4.943 ;
      RECT 83.49 4.079 83.525 5.18 ;
      RECT 83.475 3.957 83.49 5.18 ;
      RECT 83.47 3.91 83.475 5.18 ;
      RECT 83.445 3.835 83.47 5.18 ;
      RECT 83.43 3.75 83.445 5.18 ;
      RECT 83.425 3.697 83.43 5.18 ;
      RECT 83.42 3.677 83.425 5.18 ;
      RECT 83.415 3.652 83.42 4.414 ;
      RECT 83.4 4.612 83.42 5.18 ;
      RECT 83.41 3.63 83.415 4.391 ;
      RECT 83.4 3.582 83.41 4.356 ;
      RECT 83.395 3.545 83.4 4.322 ;
      RECT 83.395 4.692 83.4 5.18 ;
      RECT 83.38 3.522 83.395 4.277 ;
      RECT 83.375 4.79 83.395 5.18 ;
      RECT 83.325 3.41 83.38 4.119 ;
      RECT 83.37 4.912 83.375 5.18 ;
      RECT 83.31 3.41 83.325 3.958 ;
      RECT 83.305 3.41 83.31 3.91 ;
      RECT 83.3 3.41 83.305 3.898 ;
      RECT 83.255 3.41 83.3 3.835 ;
      RECT 83.23 3.41 83.255 3.753 ;
      RECT 83.215 3.41 83.23 3.705 ;
      RECT 83.21 3.41 83.215 3.675 ;
      RECT 82.535 4.86 82.58 5.12 ;
      RECT 82.44 3.395 82.585 3.655 ;
      RECT 82.945 4.017 82.955 4.108 ;
      RECT 82.93 3.955 82.945 4.164 ;
      RECT 82.925 3.902 82.93 4.21 ;
      RECT 82.875 3.849 82.925 4.336 ;
      RECT 82.87 3.804 82.875 4.483 ;
      RECT 82.86 3.792 82.87 4.525 ;
      RECT 82.825 3.756 82.86 4.63 ;
      RECT 82.82 3.724 82.825 4.736 ;
      RECT 82.805 3.706 82.82 4.781 ;
      RECT 82.8 3.689 82.805 4.015 ;
      RECT 82.795 4.07 82.805 4.838 ;
      RECT 82.79 3.675 82.8 3.988 ;
      RECT 82.785 4.125 82.795 5.12 ;
      RECT 82.78 3.661 82.79 3.973 ;
      RECT 82.78 4.175 82.785 5.12 ;
      RECT 82.765 3.638 82.78 3.953 ;
      RECT 82.745 4.297 82.78 5.12 ;
      RECT 82.76 3.62 82.765 3.935 ;
      RECT 82.755 3.612 82.76 3.925 ;
      RECT 82.725 3.58 82.755 3.889 ;
      RECT 82.735 4.425 82.745 5.12 ;
      RECT 82.73 4.452 82.735 5.12 ;
      RECT 82.725 4.502 82.73 5.12 ;
      RECT 82.715 3.546 82.725 3.854 ;
      RECT 82.675 4.57 82.725 5.12 ;
      RECT 82.7 3.523 82.715 3.83 ;
      RECT 82.675 3.395 82.7 3.793 ;
      RECT 82.67 3.395 82.675 3.765 ;
      RECT 82.64 4.67 82.675 5.12 ;
      RECT 82.665 3.395 82.67 3.758 ;
      RECT 82.66 3.395 82.665 3.748 ;
      RECT 82.645 3.395 82.66 3.733 ;
      RECT 82.63 3.395 82.645 3.705 ;
      RECT 82.595 4.775 82.64 5.12 ;
      RECT 82.615 3.395 82.63 3.678 ;
      RECT 82.585 3.395 82.615 3.663 ;
      RECT 82.58 4.847 82.595 5.12 ;
      RECT 82.505 3.93 82.545 4.19 ;
      RECT 82.28 3.877 82.285 4.135 ;
      RECT 78.235 3.355 78.495 3.615 ;
      RECT 78.235 3.38 78.51 3.595 ;
      RECT 80.625 3.205 80.63 3.35 ;
      RECT 82.495 3.925 82.505 4.19 ;
      RECT 82.475 3.917 82.495 4.19 ;
      RECT 82.457 3.913 82.475 4.19 ;
      RECT 82.371 3.902 82.457 4.19 ;
      RECT 82.285 3.885 82.371 4.19 ;
      RECT 82.23 3.872 82.28 4.12 ;
      RECT 82.196 3.864 82.23 4.095 ;
      RECT 82.11 3.853 82.196 4.06 ;
      RECT 82.075 3.83 82.11 4.025 ;
      RECT 82.065 3.792 82.075 4.011 ;
      RECT 82.06 3.765 82.065 4.007 ;
      RECT 82.055 3.752 82.06 4.004 ;
      RECT 82.045 3.732 82.055 4 ;
      RECT 82.04 3.707 82.045 3.996 ;
      RECT 82.015 3.662 82.04 3.99 ;
      RECT 82.005 3.603 82.015 3.982 ;
      RECT 81.995 3.571 82.005 3.973 ;
      RECT 81.975 3.523 81.995 3.953 ;
      RECT 81.97 3.483 81.975 3.923 ;
      RECT 81.955 3.457 81.97 3.897 ;
      RECT 81.95 3.435 81.955 3.873 ;
      RECT 81.935 3.407 81.95 3.849 ;
      RECT 81.92 3.38 81.935 3.813 ;
      RECT 81.905 3.357 81.92 3.775 ;
      RECT 81.9 3.347 81.905 3.75 ;
      RECT 81.89 3.34 81.9 3.733 ;
      RECT 81.875 3.327 81.89 3.703 ;
      RECT 81.87 3.317 81.875 3.678 ;
      RECT 81.865 3.312 81.87 3.665 ;
      RECT 81.855 3.305 81.865 3.645 ;
      RECT 81.85 3.298 81.855 3.63 ;
      RECT 81.825 3.291 81.85 3.588 ;
      RECT 81.81 3.281 81.825 3.538 ;
      RECT 81.8 3.276 81.81 3.508 ;
      RECT 81.79 3.272 81.8 3.483 ;
      RECT 81.775 3.269 81.79 3.473 ;
      RECT 81.725 3.266 81.775 3.458 ;
      RECT 81.705 3.264 81.725 3.443 ;
      RECT 81.656 3.262 81.705 3.438 ;
      RECT 81.57 3.258 81.656 3.433 ;
      RECT 81.531 3.255 81.57 3.429 ;
      RECT 81.445 3.251 81.531 3.424 ;
      RECT 81.395 3.248 81.445 3.418 ;
      RECT 81.346 3.245 81.395 3.413 ;
      RECT 81.26 3.242 81.346 3.408 ;
      RECT 81.256 3.24 81.26 3.405 ;
      RECT 81.17 3.237 81.256 3.4 ;
      RECT 81.121 3.233 81.17 3.393 ;
      RECT 81.035 3.23 81.121 3.388 ;
      RECT 81.011 3.227 81.035 3.384 ;
      RECT 80.925 3.225 81.011 3.379 ;
      RECT 80.86 3.221 80.925 3.372 ;
      RECT 80.857 3.22 80.86 3.369 ;
      RECT 80.771 3.217 80.857 3.366 ;
      RECT 80.685 3.211 80.771 3.359 ;
      RECT 80.655 3.207 80.685 3.355 ;
      RECT 80.63 3.205 80.655 3.353 ;
      RECT 80.575 3.202 80.625 3.35 ;
      RECT 80.495 3.201 80.575 3.35 ;
      RECT 80.44 3.203 80.495 3.353 ;
      RECT 80.425 3.204 80.44 3.357 ;
      RECT 80.37 3.212 80.425 3.367 ;
      RECT 80.34 3.22 80.37 3.38 ;
      RECT 80.321 3.221 80.34 3.386 ;
      RECT 80.235 3.224 80.321 3.391 ;
      RECT 80.165 3.229 80.235 3.4 ;
      RECT 80.146 3.232 80.165 3.406 ;
      RECT 80.06 3.236 80.146 3.411 ;
      RECT 80.02 3.24 80.06 3.418 ;
      RECT 80.011 3.242 80.02 3.421 ;
      RECT 79.925 3.246 80.011 3.426 ;
      RECT 79.922 3.249 79.925 3.43 ;
      RECT 79.836 3.252 79.922 3.434 ;
      RECT 79.75 3.258 79.836 3.442 ;
      RECT 79.726 3.262 79.75 3.446 ;
      RECT 79.64 3.266 79.726 3.451 ;
      RECT 79.595 3.271 79.64 3.458 ;
      RECT 79.515 3.276 79.595 3.465 ;
      RECT 79.435 3.282 79.515 3.48 ;
      RECT 79.41 3.286 79.435 3.493 ;
      RECT 79.345 3.289 79.41 3.505 ;
      RECT 79.29 3.294 79.345 3.52 ;
      RECT 79.26 3.297 79.29 3.538 ;
      RECT 79.25 3.299 79.26 3.551 ;
      RECT 79.19 3.314 79.25 3.561 ;
      RECT 79.175 3.331 79.19 3.57 ;
      RECT 79.17 3.34 79.175 3.57 ;
      RECT 79.16 3.35 79.17 3.57 ;
      RECT 79.15 3.367 79.16 3.57 ;
      RECT 79.13 3.377 79.15 3.571 ;
      RECT 79.085 3.387 79.13 3.572 ;
      RECT 79.05 3.396 79.085 3.574 ;
      RECT 78.985 3.401 79.05 3.576 ;
      RECT 78.905 3.402 78.985 3.579 ;
      RECT 78.901 3.4 78.905 3.58 ;
      RECT 78.815 3.397 78.901 3.582 ;
      RECT 78.768 3.394 78.815 3.584 ;
      RECT 78.682 3.39 78.768 3.587 ;
      RECT 78.596 3.386 78.682 3.59 ;
      RECT 78.51 3.382 78.596 3.594 ;
      RECT 80.445 4.445 80.725 4.725 ;
      RECT 80.485 4.425 80.745 4.685 ;
      RECT 80.475 4.435 80.745 4.685 ;
      RECT 80.485 4.362 80.7 4.725 ;
      RECT 80.54 4.285 80.695 4.725 ;
      RECT 80.545 4.07 80.695 4.725 ;
      RECT 80.535 3.872 80.685 4.123 ;
      RECT 80.525 3.872 80.685 3.99 ;
      RECT 80.52 3.75 80.68 3.893 ;
      RECT 80.505 3.75 80.68 3.798 ;
      RECT 80.5 3.46 80.675 3.775 ;
      RECT 80.485 3.46 80.675 3.745 ;
      RECT 80.445 3.46 80.705 3.72 ;
      RECT 80.355 4.93 80.435 5.19 ;
      RECT 79.76 3.65 79.765 3.915 ;
      RECT 79.64 3.65 79.765 3.91 ;
      RECT 80.315 4.895 80.355 5.19 ;
      RECT 80.27 4.817 80.315 5.19 ;
      RECT 80.25 4.745 80.27 5.19 ;
      RECT 80.24 4.697 80.25 5.19 ;
      RECT 80.205 4.63 80.24 5.19 ;
      RECT 80.175 4.53 80.205 5.19 ;
      RECT 80.155 4.455 80.175 4.99 ;
      RECT 80.145 4.405 80.155 4.945 ;
      RECT 80.14 4.382 80.145 4.918 ;
      RECT 80.135 4.367 80.14 4.905 ;
      RECT 80.13 4.352 80.135 4.883 ;
      RECT 80.125 4.337 80.13 4.865 ;
      RECT 80.1 4.292 80.125 4.82 ;
      RECT 80.09 4.24 80.1 4.763 ;
      RECT 80.08 4.21 80.09 4.73 ;
      RECT 80.07 4.175 80.08 4.698 ;
      RECT 80.035 4.107 80.07 4.63 ;
      RECT 80.03 4.046 80.035 4.565 ;
      RECT 80.02 4.034 80.03 4.545 ;
      RECT 80.015 4.022 80.02 4.525 ;
      RECT 80.01 4.014 80.015 4.513 ;
      RECT 80.005 4.006 80.01 4.493 ;
      RECT 79.995 3.994 80.005 4.465 ;
      RECT 79.985 3.978 79.995 4.435 ;
      RECT 79.96 3.95 79.985 4.373 ;
      RECT 79.95 3.921 79.96 4.318 ;
      RECT 79.935 3.9 79.95 4.278 ;
      RECT 79.93 3.884 79.935 4.25 ;
      RECT 79.925 3.872 79.93 4.24 ;
      RECT 79.92 3.867 79.925 4.213 ;
      RECT 79.915 3.86 79.92 4.2 ;
      RECT 79.9 3.843 79.915 4.173 ;
      RECT 79.89 3.65 79.9 4.133 ;
      RECT 79.88 3.65 79.89 4.1 ;
      RECT 79.87 3.65 79.88 4.075 ;
      RECT 79.8 3.65 79.87 4.01 ;
      RECT 79.79 3.65 79.8 3.958 ;
      RECT 79.775 3.65 79.79 3.94 ;
      RECT 79.765 3.65 79.775 3.925 ;
      RECT 79.595 4.52 79.855 4.78 ;
      RECT 78.13 4.555 78.135 4.762 ;
      RECT 77.765 4.445 77.84 4.76 ;
      RECT 77.58 4.5 77.735 4.76 ;
      RECT 77.765 4.445 77.87 4.725 ;
      RECT 79.58 4.617 79.595 4.778 ;
      RECT 79.555 4.625 79.58 4.783 ;
      RECT 79.53 4.632 79.555 4.788 ;
      RECT 79.467 4.643 79.53 4.797 ;
      RECT 79.381 4.662 79.467 4.814 ;
      RECT 79.295 4.684 79.381 4.833 ;
      RECT 79.28 4.697 79.295 4.844 ;
      RECT 79.24 4.705 79.28 4.851 ;
      RECT 79.22 4.71 79.24 4.858 ;
      RECT 79.182 4.711 79.22 4.861 ;
      RECT 79.096 4.714 79.182 4.862 ;
      RECT 79.01 4.718 79.096 4.863 ;
      RECT 78.961 4.72 79.01 4.865 ;
      RECT 78.875 4.72 78.961 4.867 ;
      RECT 78.835 4.715 78.875 4.869 ;
      RECT 78.825 4.709 78.835 4.87 ;
      RECT 78.785 4.704 78.825 4.867 ;
      RECT 78.775 4.697 78.785 4.863 ;
      RECT 78.76 4.693 78.775 4.861 ;
      RECT 78.743 4.689 78.76 4.859 ;
      RECT 78.657 4.679 78.743 4.851 ;
      RECT 78.571 4.661 78.657 4.837 ;
      RECT 78.485 4.644 78.571 4.823 ;
      RECT 78.46 4.632 78.485 4.814 ;
      RECT 78.39 4.622 78.46 4.807 ;
      RECT 78.345 4.61 78.39 4.798 ;
      RECT 78.285 4.597 78.345 4.79 ;
      RECT 78.28 4.589 78.285 4.785 ;
      RECT 78.245 4.584 78.28 4.783 ;
      RECT 78.19 4.575 78.245 4.776 ;
      RECT 78.15 4.564 78.19 4.768 ;
      RECT 78.135 4.557 78.15 4.764 ;
      RECT 78.115 4.55 78.13 4.761 ;
      RECT 78.1 4.54 78.115 4.759 ;
      RECT 78.085 4.527 78.1 4.756 ;
      RECT 78.06 4.51 78.085 4.752 ;
      RECT 78.045 4.492 78.06 4.749 ;
      RECT 78.02 4.445 78.045 4.747 ;
      RECT 77.996 4.445 78.02 4.744 ;
      RECT 77.91 4.445 77.996 4.736 ;
      RECT 77.87 4.445 77.91 4.728 ;
      RECT 77.735 4.492 77.765 4.76 ;
      RECT 79.415 4.075 79.675 4.335 ;
      RECT 79.375 4.075 79.675 4.213 ;
      RECT 79.34 4.075 79.675 4.198 ;
      RECT 79.285 4.075 79.675 4.178 ;
      RECT 79.205 3.885 79.485 4.165 ;
      RECT 79.205 4.067 79.555 4.165 ;
      RECT 79.205 4.01 79.54 4.165 ;
      RECT 79.205 3.957 79.49 4.165 ;
      RECT 77.035 3.885 77.23 4.67 ;
      RECT 77.115 2.5 77.23 4.67 ;
      RECT 76.97 4.41 77.03 4.67 ;
      RECT 78.34 3.93 78.6 4.19 ;
      RECT 77.025 3.885 77.23 4.165 ;
      RECT 78.335 3.94 78.6 4.125 ;
      RECT 78.05 3.915 78.06 4.065 ;
      RECT 77.285 2.5 77.365 2.845 ;
      RECT 77.02 2.5 77.23 2.845 ;
      RECT 78.325 3.94 78.335 4.124 ;
      RECT 78.315 3.939 78.325 4.121 ;
      RECT 78.306 3.938 78.315 4.119 ;
      RECT 78.22 3.934 78.306 4.109 ;
      RECT 78.146 3.926 78.22 4.091 ;
      RECT 78.06 3.919 78.146 4.074 ;
      RECT 78 3.915 78.05 4.064 ;
      RECT 77.965 3.914 78 4.061 ;
      RECT 77.91 3.914 77.965 4.063 ;
      RECT 77.875 3.914 77.91 4.067 ;
      RECT 77.789 3.913 77.875 4.074 ;
      RECT 77.703 3.912 77.789 4.084 ;
      RECT 77.617 3.911 77.703 4.095 ;
      RECT 77.531 3.911 77.617 4.105 ;
      RECT 77.445 3.91 77.531 4.115 ;
      RECT 77.41 3.91 77.445 4.155 ;
      RECT 77.405 3.91 77.41 4.198 ;
      RECT 77.38 3.91 77.405 4.215 ;
      RECT 77.305 3.91 77.38 4.23 ;
      RECT 77.285 3.885 77.305 4.243 ;
      RECT 77.28 2.5 77.285 4.253 ;
      RECT 77.255 2.5 77.28 4.295 ;
      RECT 77.23 2.5 77.255 4.373 ;
      RECT 77.03 4.292 77.035 4.67 ;
      RECT 76.365 4.244 76.38 4.7 ;
      RECT 76.36 4.316 76.466 4.698 ;
      RECT 76.38 3.41 76.515 4.696 ;
      RECT 76.365 4.26 76.52 4.695 ;
      RECT 76.365 4.31 76.525 4.693 ;
      RECT 76.35 4.375 76.525 4.692 ;
      RECT 76.36 4.367 76.53 4.689 ;
      RECT 76.34 4.415 76.53 4.684 ;
      RECT 76.34 4.415 76.545 4.681 ;
      RECT 76.335 4.415 76.545 4.678 ;
      RECT 76.31 4.415 76.57 4.675 ;
      RECT 76.38 3.41 76.54 4.063 ;
      RECT 76.375 3.41 76.54 4.035 ;
      RECT 76.37 3.41 76.54 3.863 ;
      RECT 76.37 3.41 76.56 3.803 ;
      RECT 76.325 3.41 76.585 3.67 ;
      RECT 75.805 3.885 76.085 4.165 ;
      RECT 75.795 3.9 76.085 4.16 ;
      RECT 75.75 3.962 76.085 4.158 ;
      RECT 75.825 3.877 75.99 4.165 ;
      RECT 75.825 3.862 75.946 4.165 ;
      RECT 75.86 3.855 75.946 4.165 ;
      RECT 75.325 5.005 75.605 5.285 ;
      RECT 75.285 4.967 75.58 5.078 ;
      RECT 75.27 4.917 75.56 4.973 ;
      RECT 75.215 4.68 75.475 4.94 ;
      RECT 75.215 4.882 75.555 4.94 ;
      RECT 75.215 4.822 75.55 4.94 ;
      RECT 75.215 4.772 75.53 4.94 ;
      RECT 75.215 4.752 75.525 4.94 ;
      RECT 75.215 4.73 75.52 4.94 ;
      RECT 75.215 4.715 75.49 4.94 ;
      RECT 70.945 8.66 71.265 8.98 ;
      RECT 70.975 8.13 71.145 8.98 ;
      RECT 70.975 8.13 71.15 8.48 ;
      RECT 70.975 8.13 71.95 8.305 ;
      RECT 71.775 3.26 71.95 8.305 ;
      RECT 71.72 3.26 72.07 3.61 ;
      RECT 71.745 9.09 72.07 9.415 ;
      RECT 70.63 9.18 72.07 9.35 ;
      RECT 70.63 3.69 70.79 9.35 ;
      RECT 70.945 3.66 71.265 3.98 ;
      RECT 70.63 3.69 71.265 3.86 ;
      RECT 69.3 2.435 69.675 2.805 ;
      RECT 61.22 2.255 61.595 2.625 ;
      RECT 59.785 2.255 60.16 2.625 ;
      RECT 59.785 2.375 69.605 2.545 ;
      RECT 63.905 5.655 69.585 5.825 ;
      RECT 69.415 4.72 69.585 5.825 ;
      RECT 63.715 4.895 63.74 5.825 ;
      RECT 63.97 5.005 64 5.285 ;
      RECT 63.675 4.895 63.74 5.155 ;
      RECT 69.325 4.725 69.675 5.075 ;
      RECT 63.505 3.52 63.54 3.78 ;
      RECT 63.28 3.52 63.34 3.78 ;
      RECT 63.96 4.985 63.97 5.285 ;
      RECT 63.955 4.945 63.96 5.285 ;
      RECT 63.94 4.9 63.955 5.285 ;
      RECT 63.935 4.865 63.94 5.285 ;
      RECT 63.93 4.845 63.935 5.285 ;
      RECT 63.905 4.782 63.93 5.285 ;
      RECT 63.9 4.72 63.905 5.825 ;
      RECT 63.88 4.67 63.9 5.825 ;
      RECT 63.87 4.6 63.88 5.825 ;
      RECT 63.825 4.54 63.87 5.825 ;
      RECT 63.74 4.501 63.825 5.825 ;
      RECT 63.735 4.492 63.74 4.865 ;
      RECT 63.725 4.491 63.735 4.848 ;
      RECT 63.7 4.472 63.725 4.818 ;
      RECT 63.695 4.447 63.7 4.797 ;
      RECT 63.685 4.425 63.695 4.788 ;
      RECT 63.68 4.396 63.685 4.778 ;
      RECT 63.64 4.322 63.68 4.75 ;
      RECT 63.62 4.223 63.64 4.715 ;
      RECT 63.605 4.159 63.62 4.698 ;
      RECT 63.575 4.083 63.605 4.67 ;
      RECT 63.555 3.998 63.575 4.643 ;
      RECT 63.515 3.894 63.555 4.55 ;
      RECT 63.51 3.815 63.515 4.458 ;
      RECT 63.505 3.798 63.51 4.435 ;
      RECT 63.5 3.52 63.505 4.415 ;
      RECT 63.47 3.52 63.5 4.353 ;
      RECT 63.465 3.52 63.47 4.285 ;
      RECT 63.455 3.52 63.465 4.25 ;
      RECT 63.445 3.52 63.455 4.215 ;
      RECT 63.38 3.52 63.445 4.07 ;
      RECT 63.375 3.52 63.38 3.94 ;
      RECT 63.345 3.52 63.375 3.873 ;
      RECT 63.34 3.52 63.345 3.798 ;
      RECT 67.675 3.455 67.935 3.715 ;
      RECT 67.67 3.455 67.935 3.663 ;
      RECT 67.665 3.455 67.935 3.633 ;
      RECT 67.64 3.325 67.92 3.605 ;
      RECT 56.155 9.09 56.505 9.44 ;
      RECT 67.12 9.045 67.47 9.395 ;
      RECT 56.155 9.12 67.47 9.32 ;
      RECT 66.68 5.005 66.96 5.285 ;
      RECT 66.72 4.96 66.985 5.22 ;
      RECT 66.71 4.995 66.985 5.22 ;
      RECT 66.715 4.98 66.96 5.285 ;
      RECT 66.72 4.957 66.93 5.285 ;
      RECT 66.72 4.955 66.915 5.285 ;
      RECT 66.76 4.945 66.915 5.285 ;
      RECT 66.73 4.95 66.915 5.285 ;
      RECT 66.76 4.942 66.86 5.285 ;
      RECT 66.785 4.935 66.86 5.285 ;
      RECT 66.765 4.937 66.86 5.285 ;
      RECT 66.095 4.45 66.355 4.71 ;
      RECT 66.145 4.442 66.335 4.71 ;
      RECT 66.15 4.362 66.335 4.71 ;
      RECT 66.27 3.75 66.335 4.71 ;
      RECT 66.175 4.147 66.335 4.71 ;
      RECT 66.25 3.835 66.335 4.71 ;
      RECT 66.285 3.46 66.421 4.188 ;
      RECT 66.23 3.957 66.421 4.188 ;
      RECT 66.245 3.897 66.335 4.71 ;
      RECT 66.285 3.46 66.445 3.853 ;
      RECT 66.285 3.46 66.455 3.75 ;
      RECT 66.275 3.46 66.535 3.72 ;
      RECT 65.68 5.005 65.96 5.285 ;
      RECT 65.7 4.965 65.96 5.285 ;
      RECT 65.34 4.92 65.445 5.18 ;
      RECT 65.195 3.41 65.285 3.67 ;
      RECT 65.735 4.475 65.74 4.515 ;
      RECT 65.73 4.465 65.735 4.6 ;
      RECT 65.725 4.455 65.73 4.693 ;
      RECT 65.715 4.435 65.725 4.749 ;
      RECT 65.635 4.363 65.715 4.829 ;
      RECT 65.67 5.007 65.68 5.232 ;
      RECT 65.665 5.004 65.67 5.227 ;
      RECT 65.65 5.001 65.665 5.22 ;
      RECT 65.615 4.995 65.65 5.202 ;
      RECT 65.63 4.298 65.635 4.903 ;
      RECT 65.61 4.249 65.63 4.918 ;
      RECT 65.6 4.982 65.615 5.185 ;
      RECT 65.605 4.191 65.61 4.933 ;
      RECT 65.6 4.169 65.605 4.943 ;
      RECT 65.565 4.079 65.6 5.18 ;
      RECT 65.55 3.957 65.565 5.18 ;
      RECT 65.545 3.91 65.55 5.18 ;
      RECT 65.52 3.835 65.545 5.18 ;
      RECT 65.505 3.75 65.52 5.18 ;
      RECT 65.5 3.697 65.505 5.18 ;
      RECT 65.495 3.677 65.5 5.18 ;
      RECT 65.49 3.652 65.495 4.414 ;
      RECT 65.475 4.612 65.495 5.18 ;
      RECT 65.485 3.63 65.49 4.391 ;
      RECT 65.475 3.582 65.485 4.356 ;
      RECT 65.47 3.545 65.475 4.322 ;
      RECT 65.47 4.692 65.475 5.18 ;
      RECT 65.455 3.522 65.47 4.277 ;
      RECT 65.45 4.79 65.47 5.18 ;
      RECT 65.4 3.41 65.455 4.119 ;
      RECT 65.445 4.912 65.45 5.18 ;
      RECT 65.385 3.41 65.4 3.958 ;
      RECT 65.38 3.41 65.385 3.91 ;
      RECT 65.375 3.41 65.38 3.898 ;
      RECT 65.33 3.41 65.375 3.835 ;
      RECT 65.305 3.41 65.33 3.753 ;
      RECT 65.29 3.41 65.305 3.705 ;
      RECT 65.285 3.41 65.29 3.675 ;
      RECT 64.61 4.86 64.655 5.12 ;
      RECT 64.515 3.395 64.66 3.655 ;
      RECT 65.02 4.017 65.03 4.108 ;
      RECT 65.005 3.955 65.02 4.164 ;
      RECT 65 3.902 65.005 4.21 ;
      RECT 64.95 3.849 65 4.336 ;
      RECT 64.945 3.804 64.95 4.483 ;
      RECT 64.935 3.792 64.945 4.525 ;
      RECT 64.9 3.756 64.935 4.63 ;
      RECT 64.895 3.724 64.9 4.736 ;
      RECT 64.88 3.706 64.895 4.781 ;
      RECT 64.875 3.689 64.88 4.015 ;
      RECT 64.87 4.07 64.88 4.838 ;
      RECT 64.865 3.675 64.875 3.988 ;
      RECT 64.86 4.125 64.87 5.12 ;
      RECT 64.855 3.661 64.865 3.973 ;
      RECT 64.855 4.175 64.86 5.12 ;
      RECT 64.84 3.638 64.855 3.953 ;
      RECT 64.82 4.297 64.855 5.12 ;
      RECT 64.835 3.62 64.84 3.935 ;
      RECT 64.83 3.612 64.835 3.925 ;
      RECT 64.8 3.58 64.83 3.889 ;
      RECT 64.81 4.425 64.82 5.12 ;
      RECT 64.805 4.452 64.81 5.12 ;
      RECT 64.8 4.502 64.805 5.12 ;
      RECT 64.79 3.546 64.8 3.854 ;
      RECT 64.75 4.57 64.8 5.12 ;
      RECT 64.775 3.523 64.79 3.83 ;
      RECT 64.75 3.395 64.775 3.793 ;
      RECT 64.745 3.395 64.75 3.765 ;
      RECT 64.715 4.67 64.75 5.12 ;
      RECT 64.74 3.395 64.745 3.758 ;
      RECT 64.735 3.395 64.74 3.748 ;
      RECT 64.72 3.395 64.735 3.733 ;
      RECT 64.705 3.395 64.72 3.705 ;
      RECT 64.67 4.775 64.715 5.12 ;
      RECT 64.69 3.395 64.705 3.678 ;
      RECT 64.66 3.395 64.69 3.663 ;
      RECT 64.655 4.847 64.67 5.12 ;
      RECT 64.58 3.93 64.62 4.19 ;
      RECT 64.355 3.877 64.36 4.135 ;
      RECT 60.31 3.355 60.57 3.615 ;
      RECT 60.31 3.38 60.585 3.595 ;
      RECT 62.7 3.205 62.705 3.35 ;
      RECT 64.57 3.925 64.58 4.19 ;
      RECT 64.55 3.917 64.57 4.19 ;
      RECT 64.532 3.913 64.55 4.19 ;
      RECT 64.446 3.902 64.532 4.19 ;
      RECT 64.36 3.885 64.446 4.19 ;
      RECT 64.305 3.872 64.355 4.12 ;
      RECT 64.271 3.864 64.305 4.095 ;
      RECT 64.185 3.853 64.271 4.06 ;
      RECT 64.15 3.83 64.185 4.025 ;
      RECT 64.14 3.792 64.15 4.011 ;
      RECT 64.135 3.765 64.14 4.007 ;
      RECT 64.13 3.752 64.135 4.004 ;
      RECT 64.12 3.732 64.13 4 ;
      RECT 64.115 3.707 64.12 3.996 ;
      RECT 64.09 3.662 64.115 3.99 ;
      RECT 64.08 3.603 64.09 3.982 ;
      RECT 64.07 3.571 64.08 3.973 ;
      RECT 64.05 3.523 64.07 3.953 ;
      RECT 64.045 3.483 64.05 3.923 ;
      RECT 64.03 3.457 64.045 3.897 ;
      RECT 64.025 3.435 64.03 3.873 ;
      RECT 64.01 3.407 64.025 3.849 ;
      RECT 63.995 3.38 64.01 3.813 ;
      RECT 63.98 3.357 63.995 3.775 ;
      RECT 63.975 3.347 63.98 3.75 ;
      RECT 63.965 3.34 63.975 3.733 ;
      RECT 63.95 3.327 63.965 3.703 ;
      RECT 63.945 3.317 63.95 3.678 ;
      RECT 63.94 3.312 63.945 3.665 ;
      RECT 63.93 3.305 63.94 3.645 ;
      RECT 63.925 3.298 63.93 3.63 ;
      RECT 63.9 3.291 63.925 3.588 ;
      RECT 63.885 3.281 63.9 3.538 ;
      RECT 63.875 3.276 63.885 3.508 ;
      RECT 63.865 3.272 63.875 3.483 ;
      RECT 63.85 3.269 63.865 3.473 ;
      RECT 63.8 3.266 63.85 3.458 ;
      RECT 63.78 3.264 63.8 3.443 ;
      RECT 63.731 3.262 63.78 3.438 ;
      RECT 63.645 3.258 63.731 3.433 ;
      RECT 63.606 3.255 63.645 3.429 ;
      RECT 63.52 3.251 63.606 3.424 ;
      RECT 63.47 3.248 63.52 3.418 ;
      RECT 63.421 3.245 63.47 3.413 ;
      RECT 63.335 3.242 63.421 3.408 ;
      RECT 63.331 3.24 63.335 3.405 ;
      RECT 63.245 3.237 63.331 3.4 ;
      RECT 63.196 3.233 63.245 3.393 ;
      RECT 63.11 3.23 63.196 3.388 ;
      RECT 63.086 3.227 63.11 3.384 ;
      RECT 63 3.225 63.086 3.379 ;
      RECT 62.935 3.221 63 3.372 ;
      RECT 62.932 3.22 62.935 3.369 ;
      RECT 62.846 3.217 62.932 3.366 ;
      RECT 62.76 3.211 62.846 3.359 ;
      RECT 62.73 3.207 62.76 3.355 ;
      RECT 62.705 3.205 62.73 3.353 ;
      RECT 62.65 3.202 62.7 3.35 ;
      RECT 62.57 3.201 62.65 3.35 ;
      RECT 62.515 3.203 62.57 3.353 ;
      RECT 62.5 3.204 62.515 3.357 ;
      RECT 62.445 3.212 62.5 3.367 ;
      RECT 62.415 3.22 62.445 3.38 ;
      RECT 62.396 3.221 62.415 3.386 ;
      RECT 62.31 3.224 62.396 3.391 ;
      RECT 62.24 3.229 62.31 3.4 ;
      RECT 62.221 3.232 62.24 3.406 ;
      RECT 62.135 3.236 62.221 3.411 ;
      RECT 62.095 3.24 62.135 3.418 ;
      RECT 62.086 3.242 62.095 3.421 ;
      RECT 62 3.246 62.086 3.426 ;
      RECT 61.997 3.249 62 3.43 ;
      RECT 61.911 3.252 61.997 3.434 ;
      RECT 61.825 3.258 61.911 3.442 ;
      RECT 61.801 3.262 61.825 3.446 ;
      RECT 61.715 3.266 61.801 3.451 ;
      RECT 61.67 3.271 61.715 3.458 ;
      RECT 61.59 3.276 61.67 3.465 ;
      RECT 61.51 3.282 61.59 3.48 ;
      RECT 61.485 3.286 61.51 3.493 ;
      RECT 61.42 3.289 61.485 3.505 ;
      RECT 61.365 3.294 61.42 3.52 ;
      RECT 61.335 3.297 61.365 3.538 ;
      RECT 61.325 3.299 61.335 3.551 ;
      RECT 61.265 3.314 61.325 3.561 ;
      RECT 61.25 3.331 61.265 3.57 ;
      RECT 61.245 3.34 61.25 3.57 ;
      RECT 61.235 3.35 61.245 3.57 ;
      RECT 61.225 3.367 61.235 3.57 ;
      RECT 61.205 3.377 61.225 3.571 ;
      RECT 61.16 3.387 61.205 3.572 ;
      RECT 61.125 3.396 61.16 3.574 ;
      RECT 61.06 3.401 61.125 3.576 ;
      RECT 60.98 3.402 61.06 3.579 ;
      RECT 60.976 3.4 60.98 3.58 ;
      RECT 60.89 3.397 60.976 3.582 ;
      RECT 60.843 3.394 60.89 3.584 ;
      RECT 60.757 3.39 60.843 3.587 ;
      RECT 60.671 3.386 60.757 3.59 ;
      RECT 60.585 3.382 60.671 3.594 ;
      RECT 62.52 4.445 62.8 4.725 ;
      RECT 62.56 4.425 62.82 4.685 ;
      RECT 62.55 4.435 62.82 4.685 ;
      RECT 62.56 4.362 62.775 4.725 ;
      RECT 62.615 4.285 62.77 4.725 ;
      RECT 62.62 4.07 62.77 4.725 ;
      RECT 62.61 3.872 62.76 4.123 ;
      RECT 62.6 3.872 62.76 3.99 ;
      RECT 62.595 3.75 62.755 3.893 ;
      RECT 62.58 3.75 62.755 3.798 ;
      RECT 62.575 3.46 62.75 3.775 ;
      RECT 62.56 3.46 62.75 3.745 ;
      RECT 62.52 3.46 62.78 3.72 ;
      RECT 62.43 4.93 62.51 5.19 ;
      RECT 61.835 3.65 61.84 3.915 ;
      RECT 61.715 3.65 61.84 3.91 ;
      RECT 62.39 4.895 62.43 5.19 ;
      RECT 62.345 4.817 62.39 5.19 ;
      RECT 62.325 4.745 62.345 5.19 ;
      RECT 62.315 4.697 62.325 5.19 ;
      RECT 62.28 4.63 62.315 5.19 ;
      RECT 62.25 4.53 62.28 5.19 ;
      RECT 62.23 4.455 62.25 4.99 ;
      RECT 62.22 4.405 62.23 4.945 ;
      RECT 62.215 4.382 62.22 4.918 ;
      RECT 62.21 4.367 62.215 4.905 ;
      RECT 62.205 4.352 62.21 4.883 ;
      RECT 62.2 4.337 62.205 4.865 ;
      RECT 62.175 4.292 62.2 4.82 ;
      RECT 62.165 4.24 62.175 4.763 ;
      RECT 62.155 4.21 62.165 4.73 ;
      RECT 62.145 4.175 62.155 4.698 ;
      RECT 62.11 4.107 62.145 4.63 ;
      RECT 62.105 4.046 62.11 4.565 ;
      RECT 62.095 4.034 62.105 4.545 ;
      RECT 62.09 4.022 62.095 4.525 ;
      RECT 62.085 4.014 62.09 4.513 ;
      RECT 62.08 4.006 62.085 4.493 ;
      RECT 62.07 3.994 62.08 4.465 ;
      RECT 62.06 3.978 62.07 4.435 ;
      RECT 62.035 3.95 62.06 4.373 ;
      RECT 62.025 3.921 62.035 4.318 ;
      RECT 62.01 3.9 62.025 4.278 ;
      RECT 62.005 3.884 62.01 4.25 ;
      RECT 62 3.872 62.005 4.24 ;
      RECT 61.995 3.867 62 4.213 ;
      RECT 61.99 3.86 61.995 4.2 ;
      RECT 61.975 3.843 61.99 4.173 ;
      RECT 61.965 3.65 61.975 4.133 ;
      RECT 61.955 3.65 61.965 4.1 ;
      RECT 61.945 3.65 61.955 4.075 ;
      RECT 61.875 3.65 61.945 4.01 ;
      RECT 61.865 3.65 61.875 3.958 ;
      RECT 61.85 3.65 61.865 3.94 ;
      RECT 61.84 3.65 61.85 3.925 ;
      RECT 61.67 4.52 61.93 4.78 ;
      RECT 60.205 4.555 60.21 4.762 ;
      RECT 59.84 4.445 59.915 4.76 ;
      RECT 59.655 4.5 59.81 4.76 ;
      RECT 59.84 4.445 59.945 4.725 ;
      RECT 61.655 4.617 61.67 4.778 ;
      RECT 61.63 4.625 61.655 4.783 ;
      RECT 61.605 4.632 61.63 4.788 ;
      RECT 61.542 4.643 61.605 4.797 ;
      RECT 61.456 4.662 61.542 4.814 ;
      RECT 61.37 4.684 61.456 4.833 ;
      RECT 61.355 4.697 61.37 4.844 ;
      RECT 61.315 4.705 61.355 4.851 ;
      RECT 61.295 4.71 61.315 4.858 ;
      RECT 61.257 4.711 61.295 4.861 ;
      RECT 61.171 4.714 61.257 4.862 ;
      RECT 61.085 4.718 61.171 4.863 ;
      RECT 61.036 4.72 61.085 4.865 ;
      RECT 60.95 4.72 61.036 4.867 ;
      RECT 60.91 4.715 60.95 4.869 ;
      RECT 60.9 4.709 60.91 4.87 ;
      RECT 60.86 4.704 60.9 4.867 ;
      RECT 60.85 4.697 60.86 4.863 ;
      RECT 60.835 4.693 60.85 4.861 ;
      RECT 60.818 4.689 60.835 4.859 ;
      RECT 60.732 4.679 60.818 4.851 ;
      RECT 60.646 4.661 60.732 4.837 ;
      RECT 60.56 4.644 60.646 4.823 ;
      RECT 60.535 4.632 60.56 4.814 ;
      RECT 60.465 4.622 60.535 4.807 ;
      RECT 60.42 4.61 60.465 4.798 ;
      RECT 60.36 4.597 60.42 4.79 ;
      RECT 60.355 4.589 60.36 4.785 ;
      RECT 60.32 4.584 60.355 4.783 ;
      RECT 60.265 4.575 60.32 4.776 ;
      RECT 60.225 4.564 60.265 4.768 ;
      RECT 60.21 4.557 60.225 4.764 ;
      RECT 60.19 4.55 60.205 4.761 ;
      RECT 60.175 4.54 60.19 4.759 ;
      RECT 60.16 4.527 60.175 4.756 ;
      RECT 60.135 4.51 60.16 4.752 ;
      RECT 60.12 4.492 60.135 4.749 ;
      RECT 60.095 4.445 60.12 4.747 ;
      RECT 60.071 4.445 60.095 4.744 ;
      RECT 59.985 4.445 60.071 4.736 ;
      RECT 59.945 4.445 59.985 4.728 ;
      RECT 59.81 4.492 59.84 4.76 ;
      RECT 61.49 4.075 61.75 4.335 ;
      RECT 61.45 4.075 61.75 4.213 ;
      RECT 61.415 4.075 61.75 4.198 ;
      RECT 61.36 4.075 61.75 4.178 ;
      RECT 61.28 3.885 61.56 4.165 ;
      RECT 61.28 4.067 61.63 4.165 ;
      RECT 61.28 4.01 61.615 4.165 ;
      RECT 61.28 3.957 61.565 4.165 ;
      RECT 59.11 3.885 59.305 4.67 ;
      RECT 59.19 2.5 59.305 4.67 ;
      RECT 59.045 4.41 59.105 4.67 ;
      RECT 60.415 3.93 60.675 4.19 ;
      RECT 59.1 3.885 59.305 4.165 ;
      RECT 60.41 3.94 60.675 4.125 ;
      RECT 60.125 3.915 60.135 4.065 ;
      RECT 59.36 2.5 59.44 2.845 ;
      RECT 59.095 2.5 59.305 2.845 ;
      RECT 60.4 3.94 60.41 4.124 ;
      RECT 60.39 3.939 60.4 4.121 ;
      RECT 60.381 3.938 60.39 4.119 ;
      RECT 60.295 3.934 60.381 4.109 ;
      RECT 60.221 3.926 60.295 4.091 ;
      RECT 60.135 3.919 60.221 4.074 ;
      RECT 60.075 3.915 60.125 4.064 ;
      RECT 60.04 3.914 60.075 4.061 ;
      RECT 59.985 3.914 60.04 4.063 ;
      RECT 59.95 3.914 59.985 4.067 ;
      RECT 59.864 3.913 59.95 4.074 ;
      RECT 59.778 3.912 59.864 4.084 ;
      RECT 59.692 3.911 59.778 4.095 ;
      RECT 59.606 3.911 59.692 4.105 ;
      RECT 59.52 3.91 59.606 4.115 ;
      RECT 59.485 3.91 59.52 4.155 ;
      RECT 59.48 3.91 59.485 4.198 ;
      RECT 59.455 3.91 59.48 4.215 ;
      RECT 59.38 3.91 59.455 4.23 ;
      RECT 59.36 3.885 59.38 4.243 ;
      RECT 59.355 2.5 59.36 4.253 ;
      RECT 59.33 2.5 59.355 4.295 ;
      RECT 59.305 2.5 59.33 4.373 ;
      RECT 59.105 4.292 59.11 4.67 ;
      RECT 58.44 4.244 58.455 4.7 ;
      RECT 58.435 4.316 58.541 4.698 ;
      RECT 58.455 3.41 58.59 4.696 ;
      RECT 58.44 4.26 58.595 4.695 ;
      RECT 58.44 4.31 58.6 4.693 ;
      RECT 58.425 4.375 58.6 4.692 ;
      RECT 58.435 4.367 58.605 4.689 ;
      RECT 58.415 4.415 58.605 4.684 ;
      RECT 58.415 4.415 58.62 4.681 ;
      RECT 58.41 4.415 58.62 4.678 ;
      RECT 58.385 4.415 58.645 4.675 ;
      RECT 58.455 3.41 58.615 4.063 ;
      RECT 58.45 3.41 58.615 4.035 ;
      RECT 58.445 3.41 58.615 3.863 ;
      RECT 58.445 3.41 58.635 3.803 ;
      RECT 58.4 3.41 58.66 3.67 ;
      RECT 57.88 3.885 58.16 4.165 ;
      RECT 57.87 3.9 58.16 4.16 ;
      RECT 57.825 3.962 58.16 4.158 ;
      RECT 57.9 3.877 58.065 4.165 ;
      RECT 57.9 3.862 58.021 4.165 ;
      RECT 57.935 3.855 58.021 4.165 ;
      RECT 57.4 5.005 57.68 5.285 ;
      RECT 57.36 4.967 57.655 5.078 ;
      RECT 57.345 4.917 57.635 4.973 ;
      RECT 57.29 4.68 57.55 4.94 ;
      RECT 57.29 4.882 57.63 4.94 ;
      RECT 57.29 4.822 57.625 4.94 ;
      RECT 57.29 4.772 57.605 4.94 ;
      RECT 57.29 4.752 57.6 4.94 ;
      RECT 57.29 4.73 57.595 4.94 ;
      RECT 57.29 4.715 57.565 4.94 ;
      RECT 53.02 8.66 53.34 8.98 ;
      RECT 53.05 8.13 53.22 8.98 ;
      RECT 53.05 8.13 53.225 8.48 ;
      RECT 53.05 8.13 54.025 8.305 ;
      RECT 53.85 3.26 54.025 8.305 ;
      RECT 53.795 3.26 54.145 3.61 ;
      RECT 53.82 9.09 54.145 9.415 ;
      RECT 52.705 9.18 54.145 9.35 ;
      RECT 52.705 3.69 52.865 9.35 ;
      RECT 53.02 3.66 53.34 3.98 ;
      RECT 52.705 3.69 53.34 3.86 ;
      RECT 51.375 2.435 51.75 2.805 ;
      RECT 43.295 2.255 43.67 2.625 ;
      RECT 41.86 2.255 42.235 2.625 ;
      RECT 41.86 2.375 51.68 2.545 ;
      RECT 45.98 5.655 51.66 5.825 ;
      RECT 51.49 4.72 51.66 5.825 ;
      RECT 45.79 4.895 45.815 5.825 ;
      RECT 46.045 5.005 46.075 5.285 ;
      RECT 45.75 4.895 45.815 5.155 ;
      RECT 51.4 4.725 51.75 5.075 ;
      RECT 45.58 3.52 45.615 3.78 ;
      RECT 45.355 3.52 45.415 3.78 ;
      RECT 46.035 4.985 46.045 5.285 ;
      RECT 46.03 4.945 46.035 5.285 ;
      RECT 46.015 4.9 46.03 5.285 ;
      RECT 46.01 4.865 46.015 5.285 ;
      RECT 46.005 4.845 46.01 5.285 ;
      RECT 45.98 4.782 46.005 5.285 ;
      RECT 45.975 4.72 45.98 5.825 ;
      RECT 45.955 4.67 45.975 5.825 ;
      RECT 45.945 4.6 45.955 5.825 ;
      RECT 45.9 4.54 45.945 5.825 ;
      RECT 45.815 4.501 45.9 5.825 ;
      RECT 45.81 4.492 45.815 4.865 ;
      RECT 45.8 4.491 45.81 4.848 ;
      RECT 45.775 4.472 45.8 4.818 ;
      RECT 45.77 4.447 45.775 4.797 ;
      RECT 45.76 4.425 45.77 4.788 ;
      RECT 45.755 4.396 45.76 4.778 ;
      RECT 45.715 4.322 45.755 4.75 ;
      RECT 45.695 4.223 45.715 4.715 ;
      RECT 45.68 4.159 45.695 4.698 ;
      RECT 45.65 4.083 45.68 4.67 ;
      RECT 45.63 3.998 45.65 4.643 ;
      RECT 45.59 3.894 45.63 4.55 ;
      RECT 45.585 3.815 45.59 4.458 ;
      RECT 45.58 3.798 45.585 4.435 ;
      RECT 45.575 3.52 45.58 4.415 ;
      RECT 45.545 3.52 45.575 4.353 ;
      RECT 45.54 3.52 45.545 4.285 ;
      RECT 45.53 3.52 45.54 4.25 ;
      RECT 45.52 3.52 45.53 4.215 ;
      RECT 45.455 3.52 45.52 4.07 ;
      RECT 45.45 3.52 45.455 3.94 ;
      RECT 45.42 3.52 45.45 3.873 ;
      RECT 45.415 3.52 45.42 3.798 ;
      RECT 49.75 3.455 50.01 3.715 ;
      RECT 49.745 3.455 50.01 3.663 ;
      RECT 49.74 3.455 50.01 3.633 ;
      RECT 49.715 3.325 49.995 3.605 ;
      RECT 38.275 9.095 38.625 9.445 ;
      RECT 49.25 9.05 49.6 9.4 ;
      RECT 38.275 9.125 49.6 9.325 ;
      RECT 48.755 5.005 49.035 5.285 ;
      RECT 48.795 4.96 49.06 5.22 ;
      RECT 48.785 4.995 49.06 5.22 ;
      RECT 48.79 4.98 49.035 5.285 ;
      RECT 48.795 4.957 49.005 5.285 ;
      RECT 48.795 4.955 48.99 5.285 ;
      RECT 48.835 4.945 48.99 5.285 ;
      RECT 48.805 4.95 48.99 5.285 ;
      RECT 48.835 4.942 48.935 5.285 ;
      RECT 48.86 4.935 48.935 5.285 ;
      RECT 48.84 4.937 48.935 5.285 ;
      RECT 48.17 4.45 48.43 4.71 ;
      RECT 48.22 4.442 48.41 4.71 ;
      RECT 48.225 4.362 48.41 4.71 ;
      RECT 48.345 3.75 48.41 4.71 ;
      RECT 48.25 4.147 48.41 4.71 ;
      RECT 48.325 3.835 48.41 4.71 ;
      RECT 48.36 3.46 48.496 4.188 ;
      RECT 48.305 3.957 48.496 4.188 ;
      RECT 48.32 3.897 48.41 4.71 ;
      RECT 48.36 3.46 48.52 3.853 ;
      RECT 48.36 3.46 48.53 3.75 ;
      RECT 48.35 3.46 48.61 3.72 ;
      RECT 47.755 5.005 48.035 5.285 ;
      RECT 47.775 4.965 48.035 5.285 ;
      RECT 47.415 4.92 47.52 5.18 ;
      RECT 47.27 3.41 47.36 3.67 ;
      RECT 47.81 4.475 47.815 4.515 ;
      RECT 47.805 4.465 47.81 4.6 ;
      RECT 47.8 4.455 47.805 4.693 ;
      RECT 47.79 4.435 47.8 4.749 ;
      RECT 47.71 4.363 47.79 4.829 ;
      RECT 47.745 5.007 47.755 5.232 ;
      RECT 47.74 5.004 47.745 5.227 ;
      RECT 47.725 5.001 47.74 5.22 ;
      RECT 47.69 4.995 47.725 5.202 ;
      RECT 47.705 4.298 47.71 4.903 ;
      RECT 47.685 4.249 47.705 4.918 ;
      RECT 47.675 4.982 47.69 5.185 ;
      RECT 47.68 4.191 47.685 4.933 ;
      RECT 47.675 4.169 47.68 4.943 ;
      RECT 47.64 4.079 47.675 5.18 ;
      RECT 47.625 3.957 47.64 5.18 ;
      RECT 47.62 3.91 47.625 5.18 ;
      RECT 47.595 3.835 47.62 5.18 ;
      RECT 47.58 3.75 47.595 5.18 ;
      RECT 47.575 3.697 47.58 5.18 ;
      RECT 47.57 3.677 47.575 5.18 ;
      RECT 47.565 3.652 47.57 4.414 ;
      RECT 47.55 4.612 47.57 5.18 ;
      RECT 47.56 3.63 47.565 4.391 ;
      RECT 47.55 3.582 47.56 4.356 ;
      RECT 47.545 3.545 47.55 4.322 ;
      RECT 47.545 4.692 47.55 5.18 ;
      RECT 47.53 3.522 47.545 4.277 ;
      RECT 47.525 4.79 47.545 5.18 ;
      RECT 47.475 3.41 47.53 4.119 ;
      RECT 47.52 4.912 47.525 5.18 ;
      RECT 47.46 3.41 47.475 3.958 ;
      RECT 47.455 3.41 47.46 3.91 ;
      RECT 47.45 3.41 47.455 3.898 ;
      RECT 47.405 3.41 47.45 3.835 ;
      RECT 47.38 3.41 47.405 3.753 ;
      RECT 47.365 3.41 47.38 3.705 ;
      RECT 47.36 3.41 47.365 3.675 ;
      RECT 46.685 4.86 46.73 5.12 ;
      RECT 46.59 3.395 46.735 3.655 ;
      RECT 47.095 4.017 47.105 4.108 ;
      RECT 47.08 3.955 47.095 4.164 ;
      RECT 47.075 3.902 47.08 4.21 ;
      RECT 47.025 3.849 47.075 4.336 ;
      RECT 47.02 3.804 47.025 4.483 ;
      RECT 47.01 3.792 47.02 4.525 ;
      RECT 46.975 3.756 47.01 4.63 ;
      RECT 46.97 3.724 46.975 4.736 ;
      RECT 46.955 3.706 46.97 4.781 ;
      RECT 46.95 3.689 46.955 4.015 ;
      RECT 46.945 4.07 46.955 4.838 ;
      RECT 46.94 3.675 46.95 3.988 ;
      RECT 46.935 4.125 46.945 5.12 ;
      RECT 46.93 3.661 46.94 3.973 ;
      RECT 46.93 4.175 46.935 5.12 ;
      RECT 46.915 3.638 46.93 3.953 ;
      RECT 46.895 4.297 46.93 5.12 ;
      RECT 46.91 3.62 46.915 3.935 ;
      RECT 46.905 3.612 46.91 3.925 ;
      RECT 46.875 3.58 46.905 3.889 ;
      RECT 46.885 4.425 46.895 5.12 ;
      RECT 46.88 4.452 46.885 5.12 ;
      RECT 46.875 4.502 46.88 5.12 ;
      RECT 46.865 3.546 46.875 3.854 ;
      RECT 46.825 4.57 46.875 5.12 ;
      RECT 46.85 3.523 46.865 3.83 ;
      RECT 46.825 3.395 46.85 3.793 ;
      RECT 46.82 3.395 46.825 3.765 ;
      RECT 46.79 4.67 46.825 5.12 ;
      RECT 46.815 3.395 46.82 3.758 ;
      RECT 46.81 3.395 46.815 3.748 ;
      RECT 46.795 3.395 46.81 3.733 ;
      RECT 46.78 3.395 46.795 3.705 ;
      RECT 46.745 4.775 46.79 5.12 ;
      RECT 46.765 3.395 46.78 3.678 ;
      RECT 46.735 3.395 46.765 3.663 ;
      RECT 46.73 4.847 46.745 5.12 ;
      RECT 46.655 3.93 46.695 4.19 ;
      RECT 46.43 3.877 46.435 4.135 ;
      RECT 42.385 3.355 42.645 3.615 ;
      RECT 42.385 3.38 42.66 3.595 ;
      RECT 44.775 3.205 44.78 3.35 ;
      RECT 46.645 3.925 46.655 4.19 ;
      RECT 46.625 3.917 46.645 4.19 ;
      RECT 46.607 3.913 46.625 4.19 ;
      RECT 46.521 3.902 46.607 4.19 ;
      RECT 46.435 3.885 46.521 4.19 ;
      RECT 46.38 3.872 46.43 4.12 ;
      RECT 46.346 3.864 46.38 4.095 ;
      RECT 46.26 3.853 46.346 4.06 ;
      RECT 46.225 3.83 46.26 4.025 ;
      RECT 46.215 3.792 46.225 4.011 ;
      RECT 46.21 3.765 46.215 4.007 ;
      RECT 46.205 3.752 46.21 4.004 ;
      RECT 46.195 3.732 46.205 4 ;
      RECT 46.19 3.707 46.195 3.996 ;
      RECT 46.165 3.662 46.19 3.99 ;
      RECT 46.155 3.603 46.165 3.982 ;
      RECT 46.145 3.571 46.155 3.973 ;
      RECT 46.125 3.523 46.145 3.953 ;
      RECT 46.12 3.483 46.125 3.923 ;
      RECT 46.105 3.457 46.12 3.897 ;
      RECT 46.1 3.435 46.105 3.873 ;
      RECT 46.085 3.407 46.1 3.849 ;
      RECT 46.07 3.38 46.085 3.813 ;
      RECT 46.055 3.357 46.07 3.775 ;
      RECT 46.05 3.347 46.055 3.75 ;
      RECT 46.04 3.34 46.05 3.733 ;
      RECT 46.025 3.327 46.04 3.703 ;
      RECT 46.02 3.317 46.025 3.678 ;
      RECT 46.015 3.312 46.02 3.665 ;
      RECT 46.005 3.305 46.015 3.645 ;
      RECT 46 3.298 46.005 3.63 ;
      RECT 45.975 3.291 46 3.588 ;
      RECT 45.96 3.281 45.975 3.538 ;
      RECT 45.95 3.276 45.96 3.508 ;
      RECT 45.94 3.272 45.95 3.483 ;
      RECT 45.925 3.269 45.94 3.473 ;
      RECT 45.875 3.266 45.925 3.458 ;
      RECT 45.855 3.264 45.875 3.443 ;
      RECT 45.806 3.262 45.855 3.438 ;
      RECT 45.72 3.258 45.806 3.433 ;
      RECT 45.681 3.255 45.72 3.429 ;
      RECT 45.595 3.251 45.681 3.424 ;
      RECT 45.545 3.248 45.595 3.418 ;
      RECT 45.496 3.245 45.545 3.413 ;
      RECT 45.41 3.242 45.496 3.408 ;
      RECT 45.406 3.24 45.41 3.405 ;
      RECT 45.32 3.237 45.406 3.4 ;
      RECT 45.271 3.233 45.32 3.393 ;
      RECT 45.185 3.23 45.271 3.388 ;
      RECT 45.161 3.227 45.185 3.384 ;
      RECT 45.075 3.225 45.161 3.379 ;
      RECT 45.01 3.221 45.075 3.372 ;
      RECT 45.007 3.22 45.01 3.369 ;
      RECT 44.921 3.217 45.007 3.366 ;
      RECT 44.835 3.211 44.921 3.359 ;
      RECT 44.805 3.207 44.835 3.355 ;
      RECT 44.78 3.205 44.805 3.353 ;
      RECT 44.725 3.202 44.775 3.35 ;
      RECT 44.645 3.201 44.725 3.35 ;
      RECT 44.59 3.203 44.645 3.353 ;
      RECT 44.575 3.204 44.59 3.357 ;
      RECT 44.52 3.212 44.575 3.367 ;
      RECT 44.49 3.22 44.52 3.38 ;
      RECT 44.471 3.221 44.49 3.386 ;
      RECT 44.385 3.224 44.471 3.391 ;
      RECT 44.315 3.229 44.385 3.4 ;
      RECT 44.296 3.232 44.315 3.406 ;
      RECT 44.21 3.236 44.296 3.411 ;
      RECT 44.17 3.24 44.21 3.418 ;
      RECT 44.161 3.242 44.17 3.421 ;
      RECT 44.075 3.246 44.161 3.426 ;
      RECT 44.072 3.249 44.075 3.43 ;
      RECT 43.986 3.252 44.072 3.434 ;
      RECT 43.9 3.258 43.986 3.442 ;
      RECT 43.876 3.262 43.9 3.446 ;
      RECT 43.79 3.266 43.876 3.451 ;
      RECT 43.745 3.271 43.79 3.458 ;
      RECT 43.665 3.276 43.745 3.465 ;
      RECT 43.585 3.282 43.665 3.48 ;
      RECT 43.56 3.286 43.585 3.493 ;
      RECT 43.495 3.289 43.56 3.505 ;
      RECT 43.44 3.294 43.495 3.52 ;
      RECT 43.41 3.297 43.44 3.538 ;
      RECT 43.4 3.299 43.41 3.551 ;
      RECT 43.34 3.314 43.4 3.561 ;
      RECT 43.325 3.331 43.34 3.57 ;
      RECT 43.32 3.34 43.325 3.57 ;
      RECT 43.31 3.35 43.32 3.57 ;
      RECT 43.3 3.367 43.31 3.57 ;
      RECT 43.28 3.377 43.3 3.571 ;
      RECT 43.235 3.387 43.28 3.572 ;
      RECT 43.2 3.396 43.235 3.574 ;
      RECT 43.135 3.401 43.2 3.576 ;
      RECT 43.055 3.402 43.135 3.579 ;
      RECT 43.051 3.4 43.055 3.58 ;
      RECT 42.965 3.397 43.051 3.582 ;
      RECT 42.918 3.394 42.965 3.584 ;
      RECT 42.832 3.39 42.918 3.587 ;
      RECT 42.746 3.386 42.832 3.59 ;
      RECT 42.66 3.382 42.746 3.594 ;
      RECT 44.595 4.445 44.875 4.725 ;
      RECT 44.635 4.425 44.895 4.685 ;
      RECT 44.625 4.435 44.895 4.685 ;
      RECT 44.635 4.362 44.85 4.725 ;
      RECT 44.69 4.285 44.845 4.725 ;
      RECT 44.695 4.07 44.845 4.725 ;
      RECT 44.685 3.872 44.835 4.123 ;
      RECT 44.675 3.872 44.835 3.99 ;
      RECT 44.67 3.75 44.83 3.893 ;
      RECT 44.655 3.75 44.83 3.798 ;
      RECT 44.65 3.46 44.825 3.775 ;
      RECT 44.635 3.46 44.825 3.745 ;
      RECT 44.595 3.46 44.855 3.72 ;
      RECT 44.505 4.93 44.585 5.19 ;
      RECT 43.91 3.65 43.915 3.915 ;
      RECT 43.79 3.65 43.915 3.91 ;
      RECT 44.465 4.895 44.505 5.19 ;
      RECT 44.42 4.817 44.465 5.19 ;
      RECT 44.4 4.745 44.42 5.19 ;
      RECT 44.39 4.697 44.4 5.19 ;
      RECT 44.355 4.63 44.39 5.19 ;
      RECT 44.325 4.53 44.355 5.19 ;
      RECT 44.305 4.455 44.325 4.99 ;
      RECT 44.295 4.405 44.305 4.945 ;
      RECT 44.29 4.382 44.295 4.918 ;
      RECT 44.285 4.367 44.29 4.905 ;
      RECT 44.28 4.352 44.285 4.883 ;
      RECT 44.275 4.337 44.28 4.865 ;
      RECT 44.25 4.292 44.275 4.82 ;
      RECT 44.24 4.24 44.25 4.763 ;
      RECT 44.23 4.21 44.24 4.73 ;
      RECT 44.22 4.175 44.23 4.698 ;
      RECT 44.185 4.107 44.22 4.63 ;
      RECT 44.18 4.046 44.185 4.565 ;
      RECT 44.17 4.034 44.18 4.545 ;
      RECT 44.165 4.022 44.17 4.525 ;
      RECT 44.16 4.014 44.165 4.513 ;
      RECT 44.155 4.006 44.16 4.493 ;
      RECT 44.145 3.994 44.155 4.465 ;
      RECT 44.135 3.978 44.145 4.435 ;
      RECT 44.11 3.95 44.135 4.373 ;
      RECT 44.1 3.921 44.11 4.318 ;
      RECT 44.085 3.9 44.1 4.278 ;
      RECT 44.08 3.884 44.085 4.25 ;
      RECT 44.075 3.872 44.08 4.24 ;
      RECT 44.07 3.867 44.075 4.213 ;
      RECT 44.065 3.86 44.07 4.2 ;
      RECT 44.05 3.843 44.065 4.173 ;
      RECT 44.04 3.65 44.05 4.133 ;
      RECT 44.03 3.65 44.04 4.1 ;
      RECT 44.02 3.65 44.03 4.075 ;
      RECT 43.95 3.65 44.02 4.01 ;
      RECT 43.94 3.65 43.95 3.958 ;
      RECT 43.925 3.65 43.94 3.94 ;
      RECT 43.915 3.65 43.925 3.925 ;
      RECT 43.745 4.52 44.005 4.78 ;
      RECT 42.28 4.555 42.285 4.762 ;
      RECT 41.915 4.445 41.99 4.76 ;
      RECT 41.73 4.5 41.885 4.76 ;
      RECT 41.915 4.445 42.02 4.725 ;
      RECT 43.73 4.617 43.745 4.778 ;
      RECT 43.705 4.625 43.73 4.783 ;
      RECT 43.68 4.632 43.705 4.788 ;
      RECT 43.617 4.643 43.68 4.797 ;
      RECT 43.531 4.662 43.617 4.814 ;
      RECT 43.445 4.684 43.531 4.833 ;
      RECT 43.43 4.697 43.445 4.844 ;
      RECT 43.39 4.705 43.43 4.851 ;
      RECT 43.37 4.71 43.39 4.858 ;
      RECT 43.332 4.711 43.37 4.861 ;
      RECT 43.246 4.714 43.332 4.862 ;
      RECT 43.16 4.718 43.246 4.863 ;
      RECT 43.111 4.72 43.16 4.865 ;
      RECT 43.025 4.72 43.111 4.867 ;
      RECT 42.985 4.715 43.025 4.869 ;
      RECT 42.975 4.709 42.985 4.87 ;
      RECT 42.935 4.704 42.975 4.867 ;
      RECT 42.925 4.697 42.935 4.863 ;
      RECT 42.91 4.693 42.925 4.861 ;
      RECT 42.893 4.689 42.91 4.859 ;
      RECT 42.807 4.679 42.893 4.851 ;
      RECT 42.721 4.661 42.807 4.837 ;
      RECT 42.635 4.644 42.721 4.823 ;
      RECT 42.61 4.632 42.635 4.814 ;
      RECT 42.54 4.622 42.61 4.807 ;
      RECT 42.495 4.61 42.54 4.798 ;
      RECT 42.435 4.597 42.495 4.79 ;
      RECT 42.43 4.589 42.435 4.785 ;
      RECT 42.395 4.584 42.43 4.783 ;
      RECT 42.34 4.575 42.395 4.776 ;
      RECT 42.3 4.564 42.34 4.768 ;
      RECT 42.285 4.557 42.3 4.764 ;
      RECT 42.265 4.55 42.28 4.761 ;
      RECT 42.25 4.54 42.265 4.759 ;
      RECT 42.235 4.527 42.25 4.756 ;
      RECT 42.21 4.51 42.235 4.752 ;
      RECT 42.195 4.492 42.21 4.749 ;
      RECT 42.17 4.445 42.195 4.747 ;
      RECT 42.146 4.445 42.17 4.744 ;
      RECT 42.06 4.445 42.146 4.736 ;
      RECT 42.02 4.445 42.06 4.728 ;
      RECT 41.885 4.492 41.915 4.76 ;
      RECT 43.565 4.075 43.825 4.335 ;
      RECT 43.525 4.075 43.825 4.213 ;
      RECT 43.49 4.075 43.825 4.198 ;
      RECT 43.435 4.075 43.825 4.178 ;
      RECT 43.355 3.885 43.635 4.165 ;
      RECT 43.355 4.067 43.705 4.165 ;
      RECT 43.355 4.01 43.69 4.165 ;
      RECT 43.355 3.957 43.64 4.165 ;
      RECT 41.185 3.885 41.38 4.67 ;
      RECT 41.265 2.5 41.38 4.67 ;
      RECT 41.12 4.41 41.18 4.67 ;
      RECT 42.49 3.93 42.75 4.19 ;
      RECT 41.175 3.885 41.38 4.165 ;
      RECT 42.485 3.94 42.75 4.125 ;
      RECT 42.2 3.915 42.21 4.065 ;
      RECT 41.435 2.5 41.515 2.845 ;
      RECT 41.17 2.5 41.38 2.845 ;
      RECT 42.475 3.94 42.485 4.124 ;
      RECT 42.465 3.939 42.475 4.121 ;
      RECT 42.456 3.938 42.465 4.119 ;
      RECT 42.37 3.934 42.456 4.109 ;
      RECT 42.296 3.926 42.37 4.091 ;
      RECT 42.21 3.919 42.296 4.074 ;
      RECT 42.15 3.915 42.2 4.064 ;
      RECT 42.115 3.914 42.15 4.061 ;
      RECT 42.06 3.914 42.115 4.063 ;
      RECT 42.025 3.914 42.06 4.067 ;
      RECT 41.939 3.913 42.025 4.074 ;
      RECT 41.853 3.912 41.939 4.084 ;
      RECT 41.767 3.911 41.853 4.095 ;
      RECT 41.681 3.911 41.767 4.105 ;
      RECT 41.595 3.91 41.681 4.115 ;
      RECT 41.56 3.91 41.595 4.155 ;
      RECT 41.555 3.91 41.56 4.198 ;
      RECT 41.53 3.91 41.555 4.215 ;
      RECT 41.455 3.91 41.53 4.23 ;
      RECT 41.435 3.885 41.455 4.243 ;
      RECT 41.43 2.5 41.435 4.253 ;
      RECT 41.405 2.5 41.43 4.295 ;
      RECT 41.38 2.5 41.405 4.373 ;
      RECT 41.18 4.292 41.185 4.67 ;
      RECT 40.515 4.244 40.53 4.7 ;
      RECT 40.51 4.316 40.616 4.698 ;
      RECT 40.53 3.41 40.665 4.696 ;
      RECT 40.515 4.26 40.67 4.695 ;
      RECT 40.515 4.31 40.675 4.693 ;
      RECT 40.5 4.375 40.675 4.692 ;
      RECT 40.51 4.367 40.68 4.689 ;
      RECT 40.49 4.415 40.68 4.684 ;
      RECT 40.49 4.415 40.695 4.681 ;
      RECT 40.485 4.415 40.695 4.678 ;
      RECT 40.46 4.415 40.72 4.675 ;
      RECT 40.53 3.41 40.69 4.063 ;
      RECT 40.525 3.41 40.69 4.035 ;
      RECT 40.52 3.41 40.69 3.863 ;
      RECT 40.52 3.41 40.71 3.803 ;
      RECT 40.475 3.41 40.735 3.67 ;
      RECT 39.955 3.885 40.235 4.165 ;
      RECT 39.945 3.9 40.235 4.16 ;
      RECT 39.9 3.962 40.235 4.158 ;
      RECT 39.975 3.877 40.14 4.165 ;
      RECT 39.975 3.862 40.096 4.165 ;
      RECT 40.01 3.855 40.096 4.165 ;
      RECT 39.475 5.005 39.755 5.285 ;
      RECT 39.435 4.967 39.73 5.078 ;
      RECT 39.42 4.917 39.71 4.973 ;
      RECT 39.365 4.68 39.625 4.94 ;
      RECT 39.365 4.882 39.705 4.94 ;
      RECT 39.365 4.822 39.7 4.94 ;
      RECT 39.365 4.772 39.68 4.94 ;
      RECT 39.365 4.752 39.675 4.94 ;
      RECT 39.365 4.73 39.67 4.94 ;
      RECT 39.365 4.715 39.64 4.94 ;
      RECT 35.095 8.66 35.415 8.98 ;
      RECT 35.125 8.13 35.295 8.98 ;
      RECT 35.125 8.13 35.3 8.48 ;
      RECT 35.125 8.13 36.1 8.305 ;
      RECT 35.925 3.26 36.1 8.305 ;
      RECT 35.87 3.26 36.22 3.61 ;
      RECT 35.895 9.09 36.22 9.415 ;
      RECT 34.78 9.18 36.22 9.35 ;
      RECT 34.78 3.69 34.94 9.35 ;
      RECT 35.095 3.66 35.415 3.98 ;
      RECT 34.78 3.69 35.415 3.86 ;
      RECT 33.45 2.435 33.825 2.805 ;
      RECT 25.37 2.255 25.745 2.625 ;
      RECT 23.935 2.255 24.31 2.625 ;
      RECT 23.935 2.375 33.755 2.545 ;
      RECT 28.055 5.655 33.735 5.825 ;
      RECT 33.565 4.72 33.735 5.825 ;
      RECT 27.865 4.895 27.89 5.825 ;
      RECT 28.12 5.005 28.15 5.285 ;
      RECT 27.825 4.895 27.89 5.155 ;
      RECT 33.475 4.725 33.825 5.075 ;
      RECT 27.655 3.52 27.69 3.78 ;
      RECT 27.43 3.52 27.49 3.78 ;
      RECT 28.11 4.985 28.12 5.285 ;
      RECT 28.105 4.945 28.11 5.285 ;
      RECT 28.09 4.9 28.105 5.285 ;
      RECT 28.085 4.865 28.09 5.285 ;
      RECT 28.08 4.845 28.085 5.285 ;
      RECT 28.055 4.782 28.08 5.285 ;
      RECT 28.05 4.72 28.055 5.825 ;
      RECT 28.03 4.67 28.05 5.825 ;
      RECT 28.02 4.6 28.03 5.825 ;
      RECT 27.975 4.54 28.02 5.825 ;
      RECT 27.89 4.501 27.975 5.825 ;
      RECT 27.885 4.492 27.89 4.865 ;
      RECT 27.875 4.491 27.885 4.848 ;
      RECT 27.85 4.472 27.875 4.818 ;
      RECT 27.845 4.447 27.85 4.797 ;
      RECT 27.835 4.425 27.845 4.788 ;
      RECT 27.83 4.396 27.835 4.778 ;
      RECT 27.79 4.322 27.83 4.75 ;
      RECT 27.77 4.223 27.79 4.715 ;
      RECT 27.755 4.159 27.77 4.698 ;
      RECT 27.725 4.083 27.755 4.67 ;
      RECT 27.705 3.998 27.725 4.643 ;
      RECT 27.665 3.894 27.705 4.55 ;
      RECT 27.66 3.815 27.665 4.458 ;
      RECT 27.655 3.798 27.66 4.435 ;
      RECT 27.65 3.52 27.655 4.415 ;
      RECT 27.62 3.52 27.65 4.353 ;
      RECT 27.615 3.52 27.62 4.285 ;
      RECT 27.605 3.52 27.615 4.25 ;
      RECT 27.595 3.52 27.605 4.215 ;
      RECT 27.53 3.52 27.595 4.07 ;
      RECT 27.525 3.52 27.53 3.94 ;
      RECT 27.495 3.52 27.525 3.873 ;
      RECT 27.49 3.52 27.495 3.798 ;
      RECT 31.825 3.455 32.085 3.715 ;
      RECT 31.82 3.455 32.085 3.663 ;
      RECT 31.815 3.455 32.085 3.633 ;
      RECT 31.79 3.325 32.07 3.605 ;
      RECT 20.35 9.09 20.7 9.44 ;
      RECT 31.32 9.045 31.67 9.395 ;
      RECT 20.35 9.12 31.67 9.32 ;
      RECT 30.83 5.005 31.11 5.285 ;
      RECT 30.87 4.96 31.135 5.22 ;
      RECT 30.86 4.995 31.135 5.22 ;
      RECT 30.865 4.98 31.11 5.285 ;
      RECT 30.87 4.957 31.08 5.285 ;
      RECT 30.87 4.955 31.065 5.285 ;
      RECT 30.91 4.945 31.065 5.285 ;
      RECT 30.88 4.95 31.065 5.285 ;
      RECT 30.91 4.942 31.01 5.285 ;
      RECT 30.935 4.935 31.01 5.285 ;
      RECT 30.915 4.937 31.01 5.285 ;
      RECT 30.245 4.45 30.505 4.71 ;
      RECT 30.295 4.442 30.485 4.71 ;
      RECT 30.3 4.362 30.485 4.71 ;
      RECT 30.42 3.75 30.485 4.71 ;
      RECT 30.325 4.147 30.485 4.71 ;
      RECT 30.4 3.835 30.485 4.71 ;
      RECT 30.435 3.46 30.571 4.188 ;
      RECT 30.38 3.957 30.571 4.188 ;
      RECT 30.395 3.897 30.485 4.71 ;
      RECT 30.435 3.46 30.595 3.853 ;
      RECT 30.435 3.46 30.605 3.75 ;
      RECT 30.425 3.46 30.685 3.72 ;
      RECT 29.83 5.005 30.11 5.285 ;
      RECT 29.85 4.965 30.11 5.285 ;
      RECT 29.49 4.92 29.595 5.18 ;
      RECT 29.345 3.41 29.435 3.67 ;
      RECT 29.885 4.475 29.89 4.515 ;
      RECT 29.88 4.465 29.885 4.6 ;
      RECT 29.875 4.455 29.88 4.693 ;
      RECT 29.865 4.435 29.875 4.749 ;
      RECT 29.785 4.363 29.865 4.829 ;
      RECT 29.82 5.007 29.83 5.232 ;
      RECT 29.815 5.004 29.82 5.227 ;
      RECT 29.8 5.001 29.815 5.22 ;
      RECT 29.765 4.995 29.8 5.202 ;
      RECT 29.78 4.298 29.785 4.903 ;
      RECT 29.76 4.249 29.78 4.918 ;
      RECT 29.75 4.982 29.765 5.185 ;
      RECT 29.755 4.191 29.76 4.933 ;
      RECT 29.75 4.169 29.755 4.943 ;
      RECT 29.715 4.079 29.75 5.18 ;
      RECT 29.7 3.957 29.715 5.18 ;
      RECT 29.695 3.91 29.7 5.18 ;
      RECT 29.67 3.835 29.695 5.18 ;
      RECT 29.655 3.75 29.67 5.18 ;
      RECT 29.65 3.697 29.655 5.18 ;
      RECT 29.645 3.677 29.65 5.18 ;
      RECT 29.64 3.652 29.645 4.414 ;
      RECT 29.625 4.612 29.645 5.18 ;
      RECT 29.635 3.63 29.64 4.391 ;
      RECT 29.625 3.582 29.635 4.356 ;
      RECT 29.62 3.545 29.625 4.322 ;
      RECT 29.62 4.692 29.625 5.18 ;
      RECT 29.605 3.522 29.62 4.277 ;
      RECT 29.6 4.79 29.62 5.18 ;
      RECT 29.55 3.41 29.605 4.119 ;
      RECT 29.595 4.912 29.6 5.18 ;
      RECT 29.535 3.41 29.55 3.958 ;
      RECT 29.53 3.41 29.535 3.91 ;
      RECT 29.525 3.41 29.53 3.898 ;
      RECT 29.48 3.41 29.525 3.835 ;
      RECT 29.455 3.41 29.48 3.753 ;
      RECT 29.44 3.41 29.455 3.705 ;
      RECT 29.435 3.41 29.44 3.675 ;
      RECT 28.76 4.86 28.805 5.12 ;
      RECT 28.665 3.395 28.81 3.655 ;
      RECT 29.17 4.017 29.18 4.108 ;
      RECT 29.155 3.955 29.17 4.164 ;
      RECT 29.15 3.902 29.155 4.21 ;
      RECT 29.1 3.849 29.15 4.336 ;
      RECT 29.095 3.804 29.1 4.483 ;
      RECT 29.085 3.792 29.095 4.525 ;
      RECT 29.05 3.756 29.085 4.63 ;
      RECT 29.045 3.724 29.05 4.736 ;
      RECT 29.03 3.706 29.045 4.781 ;
      RECT 29.025 3.689 29.03 4.015 ;
      RECT 29.02 4.07 29.03 4.838 ;
      RECT 29.015 3.675 29.025 3.988 ;
      RECT 29.01 4.125 29.02 5.12 ;
      RECT 29.005 3.661 29.015 3.973 ;
      RECT 29.005 4.175 29.01 5.12 ;
      RECT 28.99 3.638 29.005 3.953 ;
      RECT 28.97 4.297 29.005 5.12 ;
      RECT 28.985 3.62 28.99 3.935 ;
      RECT 28.98 3.612 28.985 3.925 ;
      RECT 28.95 3.58 28.98 3.889 ;
      RECT 28.96 4.425 28.97 5.12 ;
      RECT 28.955 4.452 28.96 5.12 ;
      RECT 28.95 4.502 28.955 5.12 ;
      RECT 28.94 3.546 28.95 3.854 ;
      RECT 28.9 4.57 28.95 5.12 ;
      RECT 28.925 3.523 28.94 3.83 ;
      RECT 28.9 3.395 28.925 3.793 ;
      RECT 28.895 3.395 28.9 3.765 ;
      RECT 28.865 4.67 28.9 5.12 ;
      RECT 28.89 3.395 28.895 3.758 ;
      RECT 28.885 3.395 28.89 3.748 ;
      RECT 28.87 3.395 28.885 3.733 ;
      RECT 28.855 3.395 28.87 3.705 ;
      RECT 28.82 4.775 28.865 5.12 ;
      RECT 28.84 3.395 28.855 3.678 ;
      RECT 28.81 3.395 28.84 3.663 ;
      RECT 28.805 4.847 28.82 5.12 ;
      RECT 28.73 3.93 28.77 4.19 ;
      RECT 28.505 3.877 28.51 4.135 ;
      RECT 24.46 3.355 24.72 3.615 ;
      RECT 24.46 3.38 24.735 3.595 ;
      RECT 26.85 3.205 26.855 3.35 ;
      RECT 28.72 3.925 28.73 4.19 ;
      RECT 28.7 3.917 28.72 4.19 ;
      RECT 28.682 3.913 28.7 4.19 ;
      RECT 28.596 3.902 28.682 4.19 ;
      RECT 28.51 3.885 28.596 4.19 ;
      RECT 28.455 3.872 28.505 4.12 ;
      RECT 28.421 3.864 28.455 4.095 ;
      RECT 28.335 3.853 28.421 4.06 ;
      RECT 28.3 3.83 28.335 4.025 ;
      RECT 28.29 3.792 28.3 4.011 ;
      RECT 28.285 3.765 28.29 4.007 ;
      RECT 28.28 3.752 28.285 4.004 ;
      RECT 28.27 3.732 28.28 4 ;
      RECT 28.265 3.707 28.27 3.996 ;
      RECT 28.24 3.662 28.265 3.99 ;
      RECT 28.23 3.603 28.24 3.982 ;
      RECT 28.22 3.571 28.23 3.973 ;
      RECT 28.2 3.523 28.22 3.953 ;
      RECT 28.195 3.483 28.2 3.923 ;
      RECT 28.18 3.457 28.195 3.897 ;
      RECT 28.175 3.435 28.18 3.873 ;
      RECT 28.16 3.407 28.175 3.849 ;
      RECT 28.145 3.38 28.16 3.813 ;
      RECT 28.13 3.357 28.145 3.775 ;
      RECT 28.125 3.347 28.13 3.75 ;
      RECT 28.115 3.34 28.125 3.733 ;
      RECT 28.1 3.327 28.115 3.703 ;
      RECT 28.095 3.317 28.1 3.678 ;
      RECT 28.09 3.312 28.095 3.665 ;
      RECT 28.08 3.305 28.09 3.645 ;
      RECT 28.075 3.298 28.08 3.63 ;
      RECT 28.05 3.291 28.075 3.588 ;
      RECT 28.035 3.281 28.05 3.538 ;
      RECT 28.025 3.276 28.035 3.508 ;
      RECT 28.015 3.272 28.025 3.483 ;
      RECT 28 3.269 28.015 3.473 ;
      RECT 27.95 3.266 28 3.458 ;
      RECT 27.93 3.264 27.95 3.443 ;
      RECT 27.881 3.262 27.93 3.438 ;
      RECT 27.795 3.258 27.881 3.433 ;
      RECT 27.756 3.255 27.795 3.429 ;
      RECT 27.67 3.251 27.756 3.424 ;
      RECT 27.62 3.248 27.67 3.418 ;
      RECT 27.571 3.245 27.62 3.413 ;
      RECT 27.485 3.242 27.571 3.408 ;
      RECT 27.481 3.24 27.485 3.405 ;
      RECT 27.395 3.237 27.481 3.4 ;
      RECT 27.346 3.233 27.395 3.393 ;
      RECT 27.26 3.23 27.346 3.388 ;
      RECT 27.236 3.227 27.26 3.384 ;
      RECT 27.15 3.225 27.236 3.379 ;
      RECT 27.085 3.221 27.15 3.372 ;
      RECT 27.082 3.22 27.085 3.369 ;
      RECT 26.996 3.217 27.082 3.366 ;
      RECT 26.91 3.211 26.996 3.359 ;
      RECT 26.88 3.207 26.91 3.355 ;
      RECT 26.855 3.205 26.88 3.353 ;
      RECT 26.8 3.202 26.85 3.35 ;
      RECT 26.72 3.201 26.8 3.35 ;
      RECT 26.665 3.203 26.72 3.353 ;
      RECT 26.65 3.204 26.665 3.357 ;
      RECT 26.595 3.212 26.65 3.367 ;
      RECT 26.565 3.22 26.595 3.38 ;
      RECT 26.546 3.221 26.565 3.386 ;
      RECT 26.46 3.224 26.546 3.391 ;
      RECT 26.39 3.229 26.46 3.4 ;
      RECT 26.371 3.232 26.39 3.406 ;
      RECT 26.285 3.236 26.371 3.411 ;
      RECT 26.245 3.24 26.285 3.418 ;
      RECT 26.236 3.242 26.245 3.421 ;
      RECT 26.15 3.246 26.236 3.426 ;
      RECT 26.147 3.249 26.15 3.43 ;
      RECT 26.061 3.252 26.147 3.434 ;
      RECT 25.975 3.258 26.061 3.442 ;
      RECT 25.951 3.262 25.975 3.446 ;
      RECT 25.865 3.266 25.951 3.451 ;
      RECT 25.82 3.271 25.865 3.458 ;
      RECT 25.74 3.276 25.82 3.465 ;
      RECT 25.66 3.282 25.74 3.48 ;
      RECT 25.635 3.286 25.66 3.493 ;
      RECT 25.57 3.289 25.635 3.505 ;
      RECT 25.515 3.294 25.57 3.52 ;
      RECT 25.485 3.297 25.515 3.538 ;
      RECT 25.475 3.299 25.485 3.551 ;
      RECT 25.415 3.314 25.475 3.561 ;
      RECT 25.4 3.331 25.415 3.57 ;
      RECT 25.395 3.34 25.4 3.57 ;
      RECT 25.385 3.35 25.395 3.57 ;
      RECT 25.375 3.367 25.385 3.57 ;
      RECT 25.355 3.377 25.375 3.571 ;
      RECT 25.31 3.387 25.355 3.572 ;
      RECT 25.275 3.396 25.31 3.574 ;
      RECT 25.21 3.401 25.275 3.576 ;
      RECT 25.13 3.402 25.21 3.579 ;
      RECT 25.126 3.4 25.13 3.58 ;
      RECT 25.04 3.397 25.126 3.582 ;
      RECT 24.993 3.394 25.04 3.584 ;
      RECT 24.907 3.39 24.993 3.587 ;
      RECT 24.821 3.386 24.907 3.59 ;
      RECT 24.735 3.382 24.821 3.594 ;
      RECT 26.67 4.445 26.95 4.725 ;
      RECT 26.71 4.425 26.97 4.685 ;
      RECT 26.7 4.435 26.97 4.685 ;
      RECT 26.71 4.362 26.925 4.725 ;
      RECT 26.765 4.285 26.92 4.725 ;
      RECT 26.77 4.07 26.92 4.725 ;
      RECT 26.76 3.872 26.91 4.123 ;
      RECT 26.75 3.872 26.91 3.99 ;
      RECT 26.745 3.75 26.905 3.893 ;
      RECT 26.73 3.75 26.905 3.798 ;
      RECT 26.725 3.46 26.9 3.775 ;
      RECT 26.71 3.46 26.9 3.745 ;
      RECT 26.67 3.46 26.93 3.72 ;
      RECT 26.58 4.93 26.66 5.19 ;
      RECT 25.985 3.65 25.99 3.915 ;
      RECT 25.865 3.65 25.99 3.91 ;
      RECT 26.54 4.895 26.58 5.19 ;
      RECT 26.495 4.817 26.54 5.19 ;
      RECT 26.475 4.745 26.495 5.19 ;
      RECT 26.465 4.697 26.475 5.19 ;
      RECT 26.43 4.63 26.465 5.19 ;
      RECT 26.4 4.53 26.43 5.19 ;
      RECT 26.38 4.455 26.4 4.99 ;
      RECT 26.37 4.405 26.38 4.945 ;
      RECT 26.365 4.382 26.37 4.918 ;
      RECT 26.36 4.367 26.365 4.905 ;
      RECT 26.355 4.352 26.36 4.883 ;
      RECT 26.35 4.337 26.355 4.865 ;
      RECT 26.325 4.292 26.35 4.82 ;
      RECT 26.315 4.24 26.325 4.763 ;
      RECT 26.305 4.21 26.315 4.73 ;
      RECT 26.295 4.175 26.305 4.698 ;
      RECT 26.26 4.107 26.295 4.63 ;
      RECT 26.255 4.046 26.26 4.565 ;
      RECT 26.245 4.034 26.255 4.545 ;
      RECT 26.24 4.022 26.245 4.525 ;
      RECT 26.235 4.014 26.24 4.513 ;
      RECT 26.23 4.006 26.235 4.493 ;
      RECT 26.22 3.994 26.23 4.465 ;
      RECT 26.21 3.978 26.22 4.435 ;
      RECT 26.185 3.95 26.21 4.373 ;
      RECT 26.175 3.921 26.185 4.318 ;
      RECT 26.16 3.9 26.175 4.278 ;
      RECT 26.155 3.884 26.16 4.25 ;
      RECT 26.15 3.872 26.155 4.24 ;
      RECT 26.145 3.867 26.15 4.213 ;
      RECT 26.14 3.86 26.145 4.2 ;
      RECT 26.125 3.843 26.14 4.173 ;
      RECT 26.115 3.65 26.125 4.133 ;
      RECT 26.105 3.65 26.115 4.1 ;
      RECT 26.095 3.65 26.105 4.075 ;
      RECT 26.025 3.65 26.095 4.01 ;
      RECT 26.015 3.65 26.025 3.958 ;
      RECT 26 3.65 26.015 3.94 ;
      RECT 25.99 3.65 26 3.925 ;
      RECT 25.82 4.52 26.08 4.78 ;
      RECT 24.355 4.555 24.36 4.762 ;
      RECT 23.99 4.445 24.065 4.76 ;
      RECT 23.805 4.5 23.96 4.76 ;
      RECT 23.99 4.445 24.095 4.725 ;
      RECT 25.805 4.617 25.82 4.778 ;
      RECT 25.78 4.625 25.805 4.783 ;
      RECT 25.755 4.632 25.78 4.788 ;
      RECT 25.692 4.643 25.755 4.797 ;
      RECT 25.606 4.662 25.692 4.814 ;
      RECT 25.52 4.684 25.606 4.833 ;
      RECT 25.505 4.697 25.52 4.844 ;
      RECT 25.465 4.705 25.505 4.851 ;
      RECT 25.445 4.71 25.465 4.858 ;
      RECT 25.407 4.711 25.445 4.861 ;
      RECT 25.321 4.714 25.407 4.862 ;
      RECT 25.235 4.718 25.321 4.863 ;
      RECT 25.186 4.72 25.235 4.865 ;
      RECT 25.1 4.72 25.186 4.867 ;
      RECT 25.06 4.715 25.1 4.869 ;
      RECT 25.05 4.709 25.06 4.87 ;
      RECT 25.01 4.704 25.05 4.867 ;
      RECT 25 4.697 25.01 4.863 ;
      RECT 24.985 4.693 25 4.861 ;
      RECT 24.968 4.689 24.985 4.859 ;
      RECT 24.882 4.679 24.968 4.851 ;
      RECT 24.796 4.661 24.882 4.837 ;
      RECT 24.71 4.644 24.796 4.823 ;
      RECT 24.685 4.632 24.71 4.814 ;
      RECT 24.615 4.622 24.685 4.807 ;
      RECT 24.57 4.61 24.615 4.798 ;
      RECT 24.51 4.597 24.57 4.79 ;
      RECT 24.505 4.589 24.51 4.785 ;
      RECT 24.47 4.584 24.505 4.783 ;
      RECT 24.415 4.575 24.47 4.776 ;
      RECT 24.375 4.564 24.415 4.768 ;
      RECT 24.36 4.557 24.375 4.764 ;
      RECT 24.34 4.55 24.355 4.761 ;
      RECT 24.325 4.54 24.34 4.759 ;
      RECT 24.31 4.527 24.325 4.756 ;
      RECT 24.285 4.51 24.31 4.752 ;
      RECT 24.27 4.492 24.285 4.749 ;
      RECT 24.245 4.445 24.27 4.747 ;
      RECT 24.221 4.445 24.245 4.744 ;
      RECT 24.135 4.445 24.221 4.736 ;
      RECT 24.095 4.445 24.135 4.728 ;
      RECT 23.96 4.492 23.99 4.76 ;
      RECT 25.64 4.075 25.9 4.335 ;
      RECT 25.6 4.075 25.9 4.213 ;
      RECT 25.565 4.075 25.9 4.198 ;
      RECT 25.51 4.075 25.9 4.178 ;
      RECT 25.43 3.885 25.71 4.165 ;
      RECT 25.43 4.067 25.78 4.165 ;
      RECT 25.43 4.01 25.765 4.165 ;
      RECT 25.43 3.957 25.715 4.165 ;
      RECT 23.26 3.885 23.455 4.67 ;
      RECT 23.34 2.5 23.455 4.67 ;
      RECT 23.195 4.41 23.255 4.67 ;
      RECT 24.565 3.93 24.825 4.19 ;
      RECT 23.25 3.885 23.455 4.165 ;
      RECT 24.56 3.94 24.825 4.125 ;
      RECT 24.275 3.915 24.285 4.065 ;
      RECT 23.51 2.5 23.59 2.845 ;
      RECT 23.245 2.5 23.455 2.845 ;
      RECT 24.55 3.94 24.56 4.124 ;
      RECT 24.54 3.939 24.55 4.121 ;
      RECT 24.531 3.938 24.54 4.119 ;
      RECT 24.445 3.934 24.531 4.109 ;
      RECT 24.371 3.926 24.445 4.091 ;
      RECT 24.285 3.919 24.371 4.074 ;
      RECT 24.225 3.915 24.275 4.064 ;
      RECT 24.19 3.914 24.225 4.061 ;
      RECT 24.135 3.914 24.19 4.063 ;
      RECT 24.1 3.914 24.135 4.067 ;
      RECT 24.014 3.913 24.1 4.074 ;
      RECT 23.928 3.912 24.014 4.084 ;
      RECT 23.842 3.911 23.928 4.095 ;
      RECT 23.756 3.911 23.842 4.105 ;
      RECT 23.67 3.91 23.756 4.115 ;
      RECT 23.635 3.91 23.67 4.155 ;
      RECT 23.63 3.91 23.635 4.198 ;
      RECT 23.605 3.91 23.63 4.215 ;
      RECT 23.53 3.91 23.605 4.23 ;
      RECT 23.51 3.885 23.53 4.243 ;
      RECT 23.505 2.5 23.51 4.253 ;
      RECT 23.48 2.5 23.505 4.295 ;
      RECT 23.455 2.5 23.48 4.373 ;
      RECT 23.255 4.292 23.26 4.67 ;
      RECT 22.59 4.244 22.605 4.7 ;
      RECT 22.585 4.316 22.691 4.698 ;
      RECT 22.605 3.41 22.74 4.696 ;
      RECT 22.59 4.26 22.745 4.695 ;
      RECT 22.59 4.31 22.75 4.693 ;
      RECT 22.575 4.375 22.75 4.692 ;
      RECT 22.585 4.367 22.755 4.689 ;
      RECT 22.565 4.415 22.755 4.684 ;
      RECT 22.565 4.415 22.77 4.681 ;
      RECT 22.56 4.415 22.77 4.678 ;
      RECT 22.535 4.415 22.795 4.675 ;
      RECT 22.605 3.41 22.765 4.063 ;
      RECT 22.6 3.41 22.765 4.035 ;
      RECT 22.595 3.41 22.765 3.863 ;
      RECT 22.595 3.41 22.785 3.803 ;
      RECT 22.55 3.41 22.81 3.67 ;
      RECT 22.03 3.885 22.31 4.165 ;
      RECT 22.02 3.9 22.31 4.16 ;
      RECT 21.975 3.962 22.31 4.158 ;
      RECT 22.05 3.877 22.215 4.165 ;
      RECT 22.05 3.862 22.171 4.165 ;
      RECT 22.085 3.855 22.171 4.165 ;
      RECT 21.55 5.005 21.83 5.285 ;
      RECT 21.51 4.967 21.805 5.078 ;
      RECT 21.495 4.917 21.785 4.973 ;
      RECT 21.44 4.68 21.7 4.94 ;
      RECT 21.44 4.882 21.78 4.94 ;
      RECT 21.44 4.822 21.775 4.94 ;
      RECT 21.44 4.772 21.755 4.94 ;
      RECT 21.44 4.752 21.75 4.94 ;
      RECT 21.44 4.73 21.745 4.94 ;
      RECT 21.44 4.715 21.715 4.94 ;
      RECT 17.17 8.66 17.49 8.98 ;
      RECT 17.2 8.13 17.37 8.98 ;
      RECT 17.2 8.13 17.375 8.48 ;
      RECT 17.2 8.13 18.175 8.305 ;
      RECT 18 3.26 18.175 8.305 ;
      RECT 17.945 3.26 18.295 3.61 ;
      RECT 17.97 9.09 18.295 9.415 ;
      RECT 16.855 9.18 18.295 9.35 ;
      RECT 16.855 3.69 17.015 9.35 ;
      RECT 17.17 3.66 17.49 3.98 ;
      RECT 16.855 3.69 17.49 3.86 ;
      RECT 15.525 2.435 15.9 2.805 ;
      RECT 7.445 2.255 7.82 2.625 ;
      RECT 6.01 2.255 6.385 2.625 ;
      RECT 6.01 2.375 15.83 2.545 ;
      RECT 10.13 5.655 15.81 5.825 ;
      RECT 15.64 4.72 15.81 5.825 ;
      RECT 9.94 4.895 9.965 5.825 ;
      RECT 10.195 5.005 10.225 5.285 ;
      RECT 9.9 4.895 9.965 5.155 ;
      RECT 15.55 4.725 15.9 5.075 ;
      RECT 9.73 3.52 9.765 3.78 ;
      RECT 9.505 3.52 9.565 3.78 ;
      RECT 10.185 4.985 10.195 5.285 ;
      RECT 10.18 4.945 10.185 5.285 ;
      RECT 10.165 4.9 10.18 5.285 ;
      RECT 10.16 4.865 10.165 5.285 ;
      RECT 10.155 4.845 10.16 5.285 ;
      RECT 10.13 4.782 10.155 5.285 ;
      RECT 10.125 4.72 10.13 5.825 ;
      RECT 10.105 4.67 10.125 5.825 ;
      RECT 10.095 4.6 10.105 5.825 ;
      RECT 10.05 4.54 10.095 5.825 ;
      RECT 9.965 4.501 10.05 5.825 ;
      RECT 9.96 4.492 9.965 4.865 ;
      RECT 9.95 4.491 9.96 4.848 ;
      RECT 9.925 4.472 9.95 4.818 ;
      RECT 9.92 4.447 9.925 4.797 ;
      RECT 9.91 4.425 9.92 4.788 ;
      RECT 9.905 4.396 9.91 4.778 ;
      RECT 9.865 4.322 9.905 4.75 ;
      RECT 9.845 4.223 9.865 4.715 ;
      RECT 9.83 4.159 9.845 4.698 ;
      RECT 9.8 4.083 9.83 4.67 ;
      RECT 9.78 3.998 9.8 4.643 ;
      RECT 9.74 3.894 9.78 4.55 ;
      RECT 9.735 3.815 9.74 4.458 ;
      RECT 9.73 3.798 9.735 4.435 ;
      RECT 9.725 3.52 9.73 4.415 ;
      RECT 9.695 3.52 9.725 4.353 ;
      RECT 9.69 3.52 9.695 4.285 ;
      RECT 9.68 3.52 9.69 4.25 ;
      RECT 9.67 3.52 9.68 4.215 ;
      RECT 9.605 3.52 9.67 4.07 ;
      RECT 9.6 3.52 9.605 3.94 ;
      RECT 9.57 3.52 9.6 3.873 ;
      RECT 9.565 3.52 9.57 3.798 ;
      RECT 13.9 3.455 14.16 3.715 ;
      RECT 13.895 3.455 14.16 3.663 ;
      RECT 13.89 3.455 14.16 3.633 ;
      RECT 13.865 3.325 14.145 3.605 ;
      RECT 1.725 9.43 2.015 9.78 ;
      RECT 1.725 9.49 3.035 9.66 ;
      RECT 2.865 9.12 3.035 9.66 ;
      RECT 13.365 9.04 13.715 9.39 ;
      RECT 2.865 9.12 13.715 9.29 ;
      RECT 12.905 5.005 13.185 5.285 ;
      RECT 12.945 4.96 13.21 5.22 ;
      RECT 12.935 4.995 13.21 5.22 ;
      RECT 12.94 4.98 13.185 5.285 ;
      RECT 12.945 4.957 13.155 5.285 ;
      RECT 12.945 4.955 13.14 5.285 ;
      RECT 12.985 4.945 13.14 5.285 ;
      RECT 12.955 4.95 13.14 5.285 ;
      RECT 12.985 4.942 13.085 5.285 ;
      RECT 13.01 4.935 13.085 5.285 ;
      RECT 12.99 4.937 13.085 5.285 ;
      RECT 12.32 4.45 12.58 4.71 ;
      RECT 12.37 4.442 12.56 4.71 ;
      RECT 12.375 4.362 12.56 4.71 ;
      RECT 12.495 3.75 12.56 4.71 ;
      RECT 12.4 4.147 12.56 4.71 ;
      RECT 12.475 3.835 12.56 4.71 ;
      RECT 12.51 3.46 12.646 4.188 ;
      RECT 12.455 3.957 12.646 4.188 ;
      RECT 12.47 3.897 12.56 4.71 ;
      RECT 12.51 3.46 12.67 3.853 ;
      RECT 12.51 3.46 12.68 3.75 ;
      RECT 12.5 3.46 12.76 3.72 ;
      RECT 11.905 5.005 12.185 5.285 ;
      RECT 11.925 4.965 12.185 5.285 ;
      RECT 11.565 4.92 11.67 5.18 ;
      RECT 11.42 3.41 11.51 3.67 ;
      RECT 11.96 4.475 11.965 4.515 ;
      RECT 11.955 4.465 11.96 4.6 ;
      RECT 11.95 4.455 11.955 4.693 ;
      RECT 11.94 4.435 11.95 4.749 ;
      RECT 11.86 4.363 11.94 4.829 ;
      RECT 11.895 5.007 11.905 5.232 ;
      RECT 11.89 5.004 11.895 5.227 ;
      RECT 11.875 5.001 11.89 5.22 ;
      RECT 11.84 4.995 11.875 5.202 ;
      RECT 11.855 4.298 11.86 4.903 ;
      RECT 11.835 4.249 11.855 4.918 ;
      RECT 11.825 4.982 11.84 5.185 ;
      RECT 11.83 4.191 11.835 4.933 ;
      RECT 11.825 4.169 11.83 4.943 ;
      RECT 11.79 4.079 11.825 5.18 ;
      RECT 11.775 3.957 11.79 5.18 ;
      RECT 11.77 3.91 11.775 5.18 ;
      RECT 11.745 3.835 11.77 5.18 ;
      RECT 11.73 3.75 11.745 5.18 ;
      RECT 11.725 3.697 11.73 5.18 ;
      RECT 11.72 3.677 11.725 5.18 ;
      RECT 11.715 3.652 11.72 4.414 ;
      RECT 11.7 4.612 11.72 5.18 ;
      RECT 11.71 3.63 11.715 4.391 ;
      RECT 11.7 3.582 11.71 4.356 ;
      RECT 11.695 3.545 11.7 4.322 ;
      RECT 11.695 4.692 11.7 5.18 ;
      RECT 11.68 3.522 11.695 4.277 ;
      RECT 11.675 4.79 11.695 5.18 ;
      RECT 11.625 3.41 11.68 4.119 ;
      RECT 11.67 4.912 11.675 5.18 ;
      RECT 11.61 3.41 11.625 3.958 ;
      RECT 11.605 3.41 11.61 3.91 ;
      RECT 11.6 3.41 11.605 3.898 ;
      RECT 11.555 3.41 11.6 3.835 ;
      RECT 11.53 3.41 11.555 3.753 ;
      RECT 11.515 3.41 11.53 3.705 ;
      RECT 11.51 3.41 11.515 3.675 ;
      RECT 10.835 4.86 10.88 5.12 ;
      RECT 10.74 3.395 10.885 3.655 ;
      RECT 11.245 4.017 11.255 4.108 ;
      RECT 11.23 3.955 11.245 4.164 ;
      RECT 11.225 3.902 11.23 4.21 ;
      RECT 11.175 3.849 11.225 4.336 ;
      RECT 11.17 3.804 11.175 4.483 ;
      RECT 11.16 3.792 11.17 4.525 ;
      RECT 11.125 3.756 11.16 4.63 ;
      RECT 11.12 3.724 11.125 4.736 ;
      RECT 11.105 3.706 11.12 4.781 ;
      RECT 11.1 3.689 11.105 4.015 ;
      RECT 11.095 4.07 11.105 4.838 ;
      RECT 11.09 3.675 11.1 3.988 ;
      RECT 11.085 4.125 11.095 5.12 ;
      RECT 11.08 3.661 11.09 3.973 ;
      RECT 11.08 4.175 11.085 5.12 ;
      RECT 11.065 3.638 11.08 3.953 ;
      RECT 11.045 4.297 11.08 5.12 ;
      RECT 11.06 3.62 11.065 3.935 ;
      RECT 11.055 3.612 11.06 3.925 ;
      RECT 11.025 3.58 11.055 3.889 ;
      RECT 11.035 4.425 11.045 5.12 ;
      RECT 11.03 4.452 11.035 5.12 ;
      RECT 11.025 4.502 11.03 5.12 ;
      RECT 11.015 3.546 11.025 3.854 ;
      RECT 10.975 4.57 11.025 5.12 ;
      RECT 11 3.523 11.015 3.83 ;
      RECT 10.975 3.395 11 3.793 ;
      RECT 10.97 3.395 10.975 3.765 ;
      RECT 10.94 4.67 10.975 5.12 ;
      RECT 10.965 3.395 10.97 3.758 ;
      RECT 10.96 3.395 10.965 3.748 ;
      RECT 10.945 3.395 10.96 3.733 ;
      RECT 10.93 3.395 10.945 3.705 ;
      RECT 10.895 4.775 10.94 5.12 ;
      RECT 10.915 3.395 10.93 3.678 ;
      RECT 10.885 3.395 10.915 3.663 ;
      RECT 10.88 4.847 10.895 5.12 ;
      RECT 10.805 3.93 10.845 4.19 ;
      RECT 10.58 3.877 10.585 4.135 ;
      RECT 6.535 3.355 6.795 3.615 ;
      RECT 6.535 3.38 6.81 3.595 ;
      RECT 8.925 3.205 8.93 3.35 ;
      RECT 10.795 3.925 10.805 4.19 ;
      RECT 10.775 3.917 10.795 4.19 ;
      RECT 10.757 3.913 10.775 4.19 ;
      RECT 10.671 3.902 10.757 4.19 ;
      RECT 10.585 3.885 10.671 4.19 ;
      RECT 10.53 3.872 10.58 4.12 ;
      RECT 10.496 3.864 10.53 4.095 ;
      RECT 10.41 3.853 10.496 4.06 ;
      RECT 10.375 3.83 10.41 4.025 ;
      RECT 10.365 3.792 10.375 4.011 ;
      RECT 10.36 3.765 10.365 4.007 ;
      RECT 10.355 3.752 10.36 4.004 ;
      RECT 10.345 3.732 10.355 4 ;
      RECT 10.34 3.707 10.345 3.996 ;
      RECT 10.315 3.662 10.34 3.99 ;
      RECT 10.305 3.603 10.315 3.982 ;
      RECT 10.295 3.571 10.305 3.973 ;
      RECT 10.275 3.523 10.295 3.953 ;
      RECT 10.27 3.483 10.275 3.923 ;
      RECT 10.255 3.457 10.27 3.897 ;
      RECT 10.25 3.435 10.255 3.873 ;
      RECT 10.235 3.407 10.25 3.849 ;
      RECT 10.22 3.38 10.235 3.813 ;
      RECT 10.205 3.357 10.22 3.775 ;
      RECT 10.2 3.347 10.205 3.75 ;
      RECT 10.19 3.34 10.2 3.733 ;
      RECT 10.175 3.327 10.19 3.703 ;
      RECT 10.17 3.317 10.175 3.678 ;
      RECT 10.165 3.312 10.17 3.665 ;
      RECT 10.155 3.305 10.165 3.645 ;
      RECT 10.15 3.298 10.155 3.63 ;
      RECT 10.125 3.291 10.15 3.588 ;
      RECT 10.11 3.281 10.125 3.538 ;
      RECT 10.1 3.276 10.11 3.508 ;
      RECT 10.09 3.272 10.1 3.483 ;
      RECT 10.075 3.269 10.09 3.473 ;
      RECT 10.025 3.266 10.075 3.458 ;
      RECT 10.005 3.264 10.025 3.443 ;
      RECT 9.956 3.262 10.005 3.438 ;
      RECT 9.87 3.258 9.956 3.433 ;
      RECT 9.831 3.255 9.87 3.429 ;
      RECT 9.745 3.251 9.831 3.424 ;
      RECT 9.695 3.248 9.745 3.418 ;
      RECT 9.646 3.245 9.695 3.413 ;
      RECT 9.56 3.242 9.646 3.408 ;
      RECT 9.556 3.24 9.56 3.405 ;
      RECT 9.47 3.237 9.556 3.4 ;
      RECT 9.421 3.233 9.47 3.393 ;
      RECT 9.335 3.23 9.421 3.388 ;
      RECT 9.311 3.227 9.335 3.384 ;
      RECT 9.225 3.225 9.311 3.379 ;
      RECT 9.16 3.221 9.225 3.372 ;
      RECT 9.157 3.22 9.16 3.369 ;
      RECT 9.071 3.217 9.157 3.366 ;
      RECT 8.985 3.211 9.071 3.359 ;
      RECT 8.955 3.207 8.985 3.355 ;
      RECT 8.93 3.205 8.955 3.353 ;
      RECT 8.875 3.202 8.925 3.35 ;
      RECT 8.795 3.201 8.875 3.35 ;
      RECT 8.74 3.203 8.795 3.353 ;
      RECT 8.725 3.204 8.74 3.357 ;
      RECT 8.67 3.212 8.725 3.367 ;
      RECT 8.64 3.22 8.67 3.38 ;
      RECT 8.621 3.221 8.64 3.386 ;
      RECT 8.535 3.224 8.621 3.391 ;
      RECT 8.465 3.229 8.535 3.4 ;
      RECT 8.446 3.232 8.465 3.406 ;
      RECT 8.36 3.236 8.446 3.411 ;
      RECT 8.32 3.24 8.36 3.418 ;
      RECT 8.311 3.242 8.32 3.421 ;
      RECT 8.225 3.246 8.311 3.426 ;
      RECT 8.222 3.249 8.225 3.43 ;
      RECT 8.136 3.252 8.222 3.434 ;
      RECT 8.05 3.258 8.136 3.442 ;
      RECT 8.026 3.262 8.05 3.446 ;
      RECT 7.94 3.266 8.026 3.451 ;
      RECT 7.895 3.271 7.94 3.458 ;
      RECT 7.815 3.276 7.895 3.465 ;
      RECT 7.735 3.282 7.815 3.48 ;
      RECT 7.71 3.286 7.735 3.493 ;
      RECT 7.645 3.289 7.71 3.505 ;
      RECT 7.59 3.294 7.645 3.52 ;
      RECT 7.56 3.297 7.59 3.538 ;
      RECT 7.55 3.299 7.56 3.551 ;
      RECT 7.49 3.314 7.55 3.561 ;
      RECT 7.475 3.331 7.49 3.57 ;
      RECT 7.47 3.34 7.475 3.57 ;
      RECT 7.46 3.35 7.47 3.57 ;
      RECT 7.45 3.367 7.46 3.57 ;
      RECT 7.43 3.377 7.45 3.571 ;
      RECT 7.385 3.387 7.43 3.572 ;
      RECT 7.35 3.396 7.385 3.574 ;
      RECT 7.285 3.401 7.35 3.576 ;
      RECT 7.205 3.402 7.285 3.579 ;
      RECT 7.201 3.4 7.205 3.58 ;
      RECT 7.115 3.397 7.201 3.582 ;
      RECT 7.068 3.394 7.115 3.584 ;
      RECT 6.982 3.39 7.068 3.587 ;
      RECT 6.896 3.386 6.982 3.59 ;
      RECT 6.81 3.382 6.896 3.594 ;
      RECT 8.745 4.445 9.025 4.725 ;
      RECT 8.785 4.425 9.045 4.685 ;
      RECT 8.775 4.435 9.045 4.685 ;
      RECT 8.785 4.362 9 4.725 ;
      RECT 8.84 4.285 8.995 4.725 ;
      RECT 8.845 4.07 8.995 4.725 ;
      RECT 8.835 3.872 8.985 4.123 ;
      RECT 8.825 3.872 8.985 3.99 ;
      RECT 8.82 3.75 8.98 3.893 ;
      RECT 8.805 3.75 8.98 3.798 ;
      RECT 8.8 3.46 8.975 3.775 ;
      RECT 8.785 3.46 8.975 3.745 ;
      RECT 8.745 3.46 9.005 3.72 ;
      RECT 8.655 4.93 8.735 5.19 ;
      RECT 8.06 3.65 8.065 3.915 ;
      RECT 7.94 3.65 8.065 3.91 ;
      RECT 8.615 4.895 8.655 5.19 ;
      RECT 8.57 4.817 8.615 5.19 ;
      RECT 8.55 4.745 8.57 5.19 ;
      RECT 8.54 4.697 8.55 5.19 ;
      RECT 8.505 4.63 8.54 5.19 ;
      RECT 8.475 4.53 8.505 5.19 ;
      RECT 8.455 4.455 8.475 4.99 ;
      RECT 8.445 4.405 8.455 4.945 ;
      RECT 8.44 4.382 8.445 4.918 ;
      RECT 8.435 4.367 8.44 4.905 ;
      RECT 8.43 4.352 8.435 4.883 ;
      RECT 8.425 4.337 8.43 4.865 ;
      RECT 8.4 4.292 8.425 4.82 ;
      RECT 8.39 4.24 8.4 4.763 ;
      RECT 8.38 4.21 8.39 4.73 ;
      RECT 8.37 4.175 8.38 4.698 ;
      RECT 8.335 4.107 8.37 4.63 ;
      RECT 8.33 4.046 8.335 4.565 ;
      RECT 8.32 4.034 8.33 4.545 ;
      RECT 8.315 4.022 8.32 4.525 ;
      RECT 8.31 4.014 8.315 4.513 ;
      RECT 8.305 4.006 8.31 4.493 ;
      RECT 8.295 3.994 8.305 4.465 ;
      RECT 8.285 3.978 8.295 4.435 ;
      RECT 8.26 3.95 8.285 4.373 ;
      RECT 8.25 3.921 8.26 4.318 ;
      RECT 8.235 3.9 8.25 4.278 ;
      RECT 8.23 3.884 8.235 4.25 ;
      RECT 8.225 3.872 8.23 4.24 ;
      RECT 8.22 3.867 8.225 4.213 ;
      RECT 8.215 3.86 8.22 4.2 ;
      RECT 8.2 3.843 8.215 4.173 ;
      RECT 8.19 3.65 8.2 4.133 ;
      RECT 8.18 3.65 8.19 4.1 ;
      RECT 8.17 3.65 8.18 4.075 ;
      RECT 8.1 3.65 8.17 4.01 ;
      RECT 8.09 3.65 8.1 3.958 ;
      RECT 8.075 3.65 8.09 3.94 ;
      RECT 8.065 3.65 8.075 3.925 ;
      RECT 7.895 4.52 8.155 4.78 ;
      RECT 6.43 4.555 6.435 4.762 ;
      RECT 6.065 4.445 6.14 4.76 ;
      RECT 5.88 4.5 6.035 4.76 ;
      RECT 6.065 4.445 6.17 4.725 ;
      RECT 7.88 4.617 7.895 4.778 ;
      RECT 7.855 4.625 7.88 4.783 ;
      RECT 7.83 4.632 7.855 4.788 ;
      RECT 7.767 4.643 7.83 4.797 ;
      RECT 7.681 4.662 7.767 4.814 ;
      RECT 7.595 4.684 7.681 4.833 ;
      RECT 7.58 4.697 7.595 4.844 ;
      RECT 7.54 4.705 7.58 4.851 ;
      RECT 7.52 4.71 7.54 4.858 ;
      RECT 7.482 4.711 7.52 4.861 ;
      RECT 7.396 4.714 7.482 4.862 ;
      RECT 7.31 4.718 7.396 4.863 ;
      RECT 7.261 4.72 7.31 4.865 ;
      RECT 7.175 4.72 7.261 4.867 ;
      RECT 7.135 4.715 7.175 4.869 ;
      RECT 7.125 4.709 7.135 4.87 ;
      RECT 7.085 4.704 7.125 4.867 ;
      RECT 7.075 4.697 7.085 4.863 ;
      RECT 7.06 4.693 7.075 4.861 ;
      RECT 7.043 4.689 7.06 4.859 ;
      RECT 6.957 4.679 7.043 4.851 ;
      RECT 6.871 4.661 6.957 4.837 ;
      RECT 6.785 4.644 6.871 4.823 ;
      RECT 6.76 4.632 6.785 4.814 ;
      RECT 6.69 4.622 6.76 4.807 ;
      RECT 6.645 4.61 6.69 4.798 ;
      RECT 6.585 4.597 6.645 4.79 ;
      RECT 6.58 4.589 6.585 4.785 ;
      RECT 6.545 4.584 6.58 4.783 ;
      RECT 6.49 4.575 6.545 4.776 ;
      RECT 6.45 4.564 6.49 4.768 ;
      RECT 6.435 4.557 6.45 4.764 ;
      RECT 6.415 4.55 6.43 4.761 ;
      RECT 6.4 4.54 6.415 4.759 ;
      RECT 6.385 4.527 6.4 4.756 ;
      RECT 6.36 4.51 6.385 4.752 ;
      RECT 6.345 4.492 6.36 4.749 ;
      RECT 6.32 4.445 6.345 4.747 ;
      RECT 6.296 4.445 6.32 4.744 ;
      RECT 6.21 4.445 6.296 4.736 ;
      RECT 6.17 4.445 6.21 4.728 ;
      RECT 6.035 4.492 6.065 4.76 ;
      RECT 7.715 4.075 7.975 4.335 ;
      RECT 7.675 4.075 7.975 4.213 ;
      RECT 7.64 4.075 7.975 4.198 ;
      RECT 7.585 4.075 7.975 4.178 ;
      RECT 7.505 3.885 7.785 4.165 ;
      RECT 7.505 4.067 7.855 4.165 ;
      RECT 7.505 4.01 7.84 4.165 ;
      RECT 7.505 3.957 7.79 4.165 ;
      RECT 5.335 3.885 5.53 4.67 ;
      RECT 5.415 2.5 5.53 4.67 ;
      RECT 5.27 4.41 5.33 4.67 ;
      RECT 6.64 3.93 6.9 4.19 ;
      RECT 5.325 3.885 5.53 4.165 ;
      RECT 6.635 3.94 6.9 4.125 ;
      RECT 6.35 3.915 6.36 4.065 ;
      RECT 5.585 2.5 5.665 2.845 ;
      RECT 5.32 2.5 5.53 2.845 ;
      RECT 6.625 3.94 6.635 4.124 ;
      RECT 6.615 3.939 6.625 4.121 ;
      RECT 6.606 3.938 6.615 4.119 ;
      RECT 6.52 3.934 6.606 4.109 ;
      RECT 6.446 3.926 6.52 4.091 ;
      RECT 6.36 3.919 6.446 4.074 ;
      RECT 6.3 3.915 6.35 4.064 ;
      RECT 6.265 3.914 6.3 4.061 ;
      RECT 6.21 3.914 6.265 4.063 ;
      RECT 6.175 3.914 6.21 4.067 ;
      RECT 6.089 3.913 6.175 4.074 ;
      RECT 6.003 3.912 6.089 4.084 ;
      RECT 5.917 3.911 6.003 4.095 ;
      RECT 5.831 3.911 5.917 4.105 ;
      RECT 5.745 3.91 5.831 4.115 ;
      RECT 5.71 3.91 5.745 4.155 ;
      RECT 5.705 3.91 5.71 4.198 ;
      RECT 5.68 3.91 5.705 4.215 ;
      RECT 5.605 3.91 5.68 4.23 ;
      RECT 5.585 3.885 5.605 4.243 ;
      RECT 5.58 2.5 5.585 4.253 ;
      RECT 5.555 2.5 5.58 4.295 ;
      RECT 5.53 2.5 5.555 4.373 ;
      RECT 5.33 4.292 5.335 4.67 ;
      RECT 4.665 4.244 4.68 4.7 ;
      RECT 4.66 4.316 4.766 4.698 ;
      RECT 4.68 3.41 4.815 4.696 ;
      RECT 4.665 4.26 4.82 4.695 ;
      RECT 4.665 4.31 4.825 4.693 ;
      RECT 4.65 4.375 4.825 4.692 ;
      RECT 4.66 4.367 4.83 4.689 ;
      RECT 4.64 4.415 4.83 4.684 ;
      RECT 4.64 4.415 4.845 4.681 ;
      RECT 4.635 4.415 4.845 4.678 ;
      RECT 4.61 4.415 4.87 4.675 ;
      RECT 4.68 3.41 4.84 4.063 ;
      RECT 4.675 3.41 4.84 4.035 ;
      RECT 4.67 3.41 4.84 3.863 ;
      RECT 4.67 3.41 4.86 3.803 ;
      RECT 4.625 3.41 4.885 3.67 ;
      RECT 4.105 3.885 4.385 4.165 ;
      RECT 4.095 3.9 4.385 4.16 ;
      RECT 4.05 3.962 4.385 4.158 ;
      RECT 4.125 3.877 4.29 4.165 ;
      RECT 4.125 3.862 4.246 4.165 ;
      RECT 4.16 3.855 4.246 4.165 ;
      RECT 3.625 5.005 3.905 5.285 ;
      RECT 3.585 4.967 3.88 5.078 ;
      RECT 3.57 4.917 3.86 4.973 ;
      RECT 3.515 4.68 3.775 4.94 ;
      RECT 3.515 4.882 3.855 4.94 ;
      RECT 3.515 4.822 3.85 4.94 ;
      RECT 3.515 4.772 3.83 4.94 ;
      RECT 3.515 4.752 3.825 4.94 ;
      RECT 3.515 4.73 3.82 4.94 ;
      RECT 3.515 4.715 3.79 4.94 ;
      RECT 84.405 9.49 84.78 9.86 ;
      RECT 75.74 2.225 76.115 2.595 ;
      RECT 66.48 9.49 66.855 9.86 ;
      RECT 57.815 2.225 58.19 2.595 ;
      RECT 48.555 9.49 48.93 9.86 ;
      RECT 39.89 2.225 40.265 2.595 ;
      RECT 30.63 9.49 31.005 9.86 ;
      RECT 21.965 2.225 22.34 2.595 ;
      RECT 12.705 9.49 13.08 9.86 ;
      RECT 4.04 2.225 4.415 2.595 ;
    LAYER via1 ;
      RECT 92.125 9.81 92.275 9.96 ;
      RECT 89.76 9.175 89.91 9.325 ;
      RECT 89.745 3.36 89.895 3.51 ;
      RECT 88.955 3.745 89.105 3.895 ;
      RECT 88.955 8.76 89.105 8.91 ;
      RECT 87.35 4.825 87.5 4.975 ;
      RECT 87.34 2.545 87.49 2.695 ;
      RECT 85.655 3.51 85.805 3.66 ;
      RECT 85.425 9.145 85.575 9.295 ;
      RECT 84.705 5.015 84.855 5.165 ;
      RECT 84.52 9.6 84.67 9.75 ;
      RECT 84.255 3.515 84.405 3.665 ;
      RECT 84.075 4.505 84.225 4.655 ;
      RECT 83.68 5.02 83.83 5.17 ;
      RECT 83.32 4.975 83.47 5.125 ;
      RECT 83.175 3.465 83.325 3.615 ;
      RECT 82.59 4.915 82.74 5.065 ;
      RECT 82.495 3.45 82.645 3.6 ;
      RECT 82.34 3.985 82.49 4.135 ;
      RECT 81.655 4.95 81.805 5.1 ;
      RECT 81.26 3.575 81.41 3.725 ;
      RECT 80.54 4.48 80.69 4.63 ;
      RECT 80.5 3.515 80.65 3.665 ;
      RECT 80.23 4.985 80.38 5.135 ;
      RECT 79.695 3.705 79.845 3.855 ;
      RECT 79.65 4.575 79.8 4.725 ;
      RECT 79.47 4.13 79.62 4.28 ;
      RECT 78.395 3.985 78.545 4.135 ;
      RECT 78.29 3.41 78.44 3.56 ;
      RECT 77.635 4.555 77.785 4.705 ;
      RECT 77.115 2.595 77.265 2.745 ;
      RECT 77.025 4.465 77.175 4.615 ;
      RECT 76.38 3.465 76.53 3.615 ;
      RECT 76.365 4.47 76.515 4.62 ;
      RECT 75.85 3.955 76 4.105 ;
      RECT 75.27 4.735 75.42 4.885 ;
      RECT 74.18 9.19 74.33 9.34 ;
      RECT 71.835 9.175 71.985 9.325 ;
      RECT 71.82 3.36 71.97 3.51 ;
      RECT 71.03 3.745 71.18 3.895 ;
      RECT 71.03 8.76 71.18 8.91 ;
      RECT 69.425 4.825 69.575 4.975 ;
      RECT 69.415 2.545 69.565 2.695 ;
      RECT 67.73 3.51 67.88 3.66 ;
      RECT 67.22 9.145 67.37 9.295 ;
      RECT 66.78 5.015 66.93 5.165 ;
      RECT 66.595 9.6 66.745 9.75 ;
      RECT 66.33 3.515 66.48 3.665 ;
      RECT 66.15 4.505 66.3 4.655 ;
      RECT 65.755 5.02 65.905 5.17 ;
      RECT 65.395 4.975 65.545 5.125 ;
      RECT 65.25 3.465 65.4 3.615 ;
      RECT 64.665 4.915 64.815 5.065 ;
      RECT 64.57 3.45 64.72 3.6 ;
      RECT 64.415 3.985 64.565 4.135 ;
      RECT 63.73 4.95 63.88 5.1 ;
      RECT 63.335 3.575 63.485 3.725 ;
      RECT 62.615 4.48 62.765 4.63 ;
      RECT 62.575 3.515 62.725 3.665 ;
      RECT 62.305 4.985 62.455 5.135 ;
      RECT 61.77 3.705 61.92 3.855 ;
      RECT 61.725 4.575 61.875 4.725 ;
      RECT 61.545 4.13 61.695 4.28 ;
      RECT 60.47 3.985 60.62 4.135 ;
      RECT 60.365 3.41 60.515 3.56 ;
      RECT 59.71 4.555 59.86 4.705 ;
      RECT 59.19 2.595 59.34 2.745 ;
      RECT 59.1 4.465 59.25 4.615 ;
      RECT 58.455 3.465 58.605 3.615 ;
      RECT 58.44 4.47 58.59 4.62 ;
      RECT 57.925 3.955 58.075 4.105 ;
      RECT 57.345 4.735 57.495 4.885 ;
      RECT 56.255 9.19 56.405 9.34 ;
      RECT 53.91 9.175 54.06 9.325 ;
      RECT 53.895 3.36 54.045 3.51 ;
      RECT 53.105 3.745 53.255 3.895 ;
      RECT 53.105 8.76 53.255 8.91 ;
      RECT 51.5 4.825 51.65 4.975 ;
      RECT 51.49 2.545 51.64 2.695 ;
      RECT 49.805 3.51 49.955 3.66 ;
      RECT 49.35 9.15 49.5 9.3 ;
      RECT 48.855 5.015 49.005 5.165 ;
      RECT 48.67 9.6 48.82 9.75 ;
      RECT 48.405 3.515 48.555 3.665 ;
      RECT 48.225 4.505 48.375 4.655 ;
      RECT 47.83 5.02 47.98 5.17 ;
      RECT 47.47 4.975 47.62 5.125 ;
      RECT 47.325 3.465 47.475 3.615 ;
      RECT 46.74 4.915 46.89 5.065 ;
      RECT 46.645 3.45 46.795 3.6 ;
      RECT 46.49 3.985 46.64 4.135 ;
      RECT 45.805 4.95 45.955 5.1 ;
      RECT 45.41 3.575 45.56 3.725 ;
      RECT 44.69 4.48 44.84 4.63 ;
      RECT 44.65 3.515 44.8 3.665 ;
      RECT 44.38 4.985 44.53 5.135 ;
      RECT 43.845 3.705 43.995 3.855 ;
      RECT 43.8 4.575 43.95 4.725 ;
      RECT 43.62 4.13 43.77 4.28 ;
      RECT 42.545 3.985 42.695 4.135 ;
      RECT 42.44 3.41 42.59 3.56 ;
      RECT 41.785 4.555 41.935 4.705 ;
      RECT 41.265 2.595 41.415 2.745 ;
      RECT 41.175 4.465 41.325 4.615 ;
      RECT 40.53 3.465 40.68 3.615 ;
      RECT 40.515 4.47 40.665 4.62 ;
      RECT 40 3.955 40.15 4.105 ;
      RECT 39.42 4.735 39.57 4.885 ;
      RECT 38.375 9.195 38.525 9.345 ;
      RECT 35.985 9.175 36.135 9.325 ;
      RECT 35.97 3.36 36.12 3.51 ;
      RECT 35.18 3.745 35.33 3.895 ;
      RECT 35.18 8.76 35.33 8.91 ;
      RECT 33.575 4.825 33.725 4.975 ;
      RECT 33.565 2.545 33.715 2.695 ;
      RECT 31.88 3.51 32.03 3.66 ;
      RECT 31.42 9.145 31.57 9.295 ;
      RECT 30.93 5.015 31.08 5.165 ;
      RECT 30.745 9.6 30.895 9.75 ;
      RECT 30.48 3.515 30.63 3.665 ;
      RECT 30.3 4.505 30.45 4.655 ;
      RECT 29.905 5.02 30.055 5.17 ;
      RECT 29.545 4.975 29.695 5.125 ;
      RECT 29.4 3.465 29.55 3.615 ;
      RECT 28.815 4.915 28.965 5.065 ;
      RECT 28.72 3.45 28.87 3.6 ;
      RECT 28.565 3.985 28.715 4.135 ;
      RECT 27.88 4.95 28.03 5.1 ;
      RECT 27.485 3.575 27.635 3.725 ;
      RECT 26.765 4.48 26.915 4.63 ;
      RECT 26.725 3.515 26.875 3.665 ;
      RECT 26.455 4.985 26.605 5.135 ;
      RECT 25.92 3.705 26.07 3.855 ;
      RECT 25.875 4.575 26.025 4.725 ;
      RECT 25.695 4.13 25.845 4.28 ;
      RECT 24.62 3.985 24.77 4.135 ;
      RECT 24.515 3.41 24.665 3.56 ;
      RECT 23.86 4.555 24.01 4.705 ;
      RECT 23.34 2.595 23.49 2.745 ;
      RECT 23.25 4.465 23.4 4.615 ;
      RECT 22.605 3.465 22.755 3.615 ;
      RECT 22.59 4.47 22.74 4.62 ;
      RECT 22.075 3.955 22.225 4.105 ;
      RECT 21.495 4.735 21.645 4.885 ;
      RECT 20.45 9.19 20.6 9.34 ;
      RECT 18.06 9.175 18.21 9.325 ;
      RECT 18.045 3.36 18.195 3.51 ;
      RECT 17.255 3.745 17.405 3.895 ;
      RECT 17.255 8.76 17.405 8.91 ;
      RECT 15.65 4.825 15.8 4.975 ;
      RECT 15.64 2.545 15.79 2.695 ;
      RECT 13.955 3.51 14.105 3.66 ;
      RECT 13.465 9.14 13.615 9.29 ;
      RECT 13.005 5.015 13.155 5.165 ;
      RECT 12.82 9.6 12.97 9.75 ;
      RECT 12.555 3.515 12.705 3.665 ;
      RECT 12.375 4.505 12.525 4.655 ;
      RECT 11.98 5.02 12.13 5.17 ;
      RECT 11.62 4.975 11.77 5.125 ;
      RECT 11.475 3.465 11.625 3.615 ;
      RECT 10.89 4.915 11.04 5.065 ;
      RECT 10.795 3.45 10.945 3.6 ;
      RECT 10.64 3.985 10.79 4.135 ;
      RECT 9.955 4.95 10.105 5.1 ;
      RECT 9.56 3.575 9.71 3.725 ;
      RECT 8.84 4.48 8.99 4.63 ;
      RECT 8.8 3.515 8.95 3.665 ;
      RECT 8.53 4.985 8.68 5.135 ;
      RECT 7.995 3.705 8.145 3.855 ;
      RECT 7.95 4.575 8.1 4.725 ;
      RECT 7.77 4.13 7.92 4.28 ;
      RECT 6.695 3.985 6.845 4.135 ;
      RECT 6.59 3.41 6.74 3.56 ;
      RECT 5.935 4.555 6.085 4.705 ;
      RECT 5.415 2.595 5.565 2.745 ;
      RECT 5.325 4.465 5.475 4.615 ;
      RECT 4.68 3.465 4.83 3.615 ;
      RECT 4.665 4.47 4.815 4.62 ;
      RECT 4.15 3.955 4.3 4.105 ;
      RECT 3.57 4.735 3.72 4.885 ;
      RECT 1.795 9.53 1.945 9.68 ;
      RECT 1.42 8.79 1.57 8.94 ;
    LAYER met1 ;
      RECT 75.05 2.58 87.01 3.185 ;
      RECT 79.475 0 87.01 3.185 ;
      RECT 57.125 2.58 69.085 3.185 ;
      RECT 61.55 0 69.085 3.185 ;
      RECT 39.2 2.58 51.16 3.185 ;
      RECT 43.625 0 51.16 3.185 ;
      RECT 21.275 2.58 33.235 3.185 ;
      RECT 25.7 0 33.235 3.185 ;
      RECT 3.35 2.435 15.31 3.185 ;
      RECT 7.775 0 15.31 3.185 ;
      RECT 75.045 0 75.79 2.975 ;
      RECT 57.12 0 57.865 2.975 ;
      RECT 39.195 0 39.94 2.975 ;
      RECT 21.27 0 22.015 2.975 ;
      RECT 3.345 0 4.09 2.975 ;
      RECT 15.525 2.435 15.9 2.805 ;
      RECT 3.345 2.435 16.275 2.74 ;
      RECT 78.04 0 79.195 3.185 ;
      RECT 75.045 2.55 77.76 2.975 ;
      RECT 76.07 0 77.76 3.185 ;
      RECT 60.115 0 61.27 3.185 ;
      RECT 57.12 2.55 59.835 2.975 ;
      RECT 58.145 0 59.835 3.185 ;
      RECT 42.19 0 43.345 3.185 ;
      RECT 39.195 2.55 41.91 2.975 ;
      RECT 40.22 0 41.91 3.185 ;
      RECT 24.265 0 25.42 3.185 ;
      RECT 21.27 2.55 23.985 2.975 ;
      RECT 22.295 0 23.985 3.185 ;
      RECT 6.34 0 7.495 3.185 ;
      RECT 4.37 0 6.06 3.185 ;
      RECT 76.07 0 87.01 2.3 ;
      RECT 58.145 0 69.085 2.3 ;
      RECT 40.22 0 51.16 2.3 ;
      RECT 22.295 0 33.235 2.3 ;
      RECT 4.37 0 15.31 2.3 ;
      RECT 75.045 0 87.01 2.27 ;
      RECT 57.12 0 69.085 2.27 ;
      RECT 39.195 0 51.16 2.27 ;
      RECT 21.27 0 33.235 2.27 ;
      RECT 3.345 0 15.31 2.27 ;
      RECT 0.02 0 92.6 1.6 ;
      RECT 91.995 10.205 92.285 10.435 ;
      RECT 92.055 8.725 92.225 10.435 ;
      RECT 92.025 9.71 92.375 10.06 ;
      RECT 91.995 8.725 92.285 8.955 ;
      RECT 91.59 3.69 91.695 4.26 ;
      RECT 91.59 4.025 91.915 4.255 ;
      RECT 91.59 4.055 92.085 4.225 ;
      RECT 91.59 3.69 91.78 4.255 ;
      RECT 91.005 3.655 91.295 3.885 ;
      RECT 91.005 3.69 91.78 3.86 ;
      RECT 91.065 2.175 91.235 3.885 ;
      RECT 91.005 2.175 91.295 2.405 ;
      RECT 91.005 10.205 91.295 10.435 ;
      RECT 91.065 8.725 91.235 10.435 ;
      RECT 91.005 8.725 91.295 8.955 ;
      RECT 91.005 8.76 91.86 8.92 ;
      RECT 91.69 8.355 91.86 8.92 ;
      RECT 91.005 8.755 91.4 8.92 ;
      RECT 91.625 8.355 91.915 8.585 ;
      RECT 91.625 8.385 92.085 8.555 ;
      RECT 90.635 4.025 90.925 4.255 ;
      RECT 90.635 4.055 91.095 4.225 ;
      RECT 90.7 2.95 90.865 4.255 ;
      RECT 89.215 2.92 89.505 3.15 ;
      RECT 89.215 2.95 90.865 3.12 ;
      RECT 89.275 2.18 89.445 3.15 ;
      RECT 89.215 2.18 89.505 2.41 ;
      RECT 89.215 10.2 89.505 10.43 ;
      RECT 89.275 9.46 89.445 10.43 ;
      RECT 89.275 9.555 90.865 9.725 ;
      RECT 90.695 8.355 90.865 9.725 ;
      RECT 89.215 9.46 89.505 9.69 ;
      RECT 90.635 8.355 90.925 8.585 ;
      RECT 90.635 8.385 91.095 8.555 ;
      RECT 87.25 4.725 87.6 5.075 ;
      RECT 87.34 3.32 87.51 5.075 ;
      RECT 89.645 3.26 89.995 3.61 ;
      RECT 87.34 3.32 88.96 3.495 ;
      RECT 87.34 3.32 89.995 3.49 ;
      RECT 89.67 9.09 89.995 9.415 ;
      RECT 85.325 9.045 85.675 9.395 ;
      RECT 89.645 9.09 89.995 9.32 ;
      RECT 84.885 9.09 85.175 9.32 ;
      RECT 84.715 9.12 89.995 9.29 ;
      RECT 88.87 3.66 89.19 3.98 ;
      RECT 88.84 3.66 89.19 3.89 ;
      RECT 88.67 3.69 89.19 3.86 ;
      RECT 88.87 8.66 89.19 8.98 ;
      RECT 88.84 8.72 89.19 8.95 ;
      RECT 88.67 8.75 89.19 8.92 ;
      RECT 84.65 4.96 84.69 5.22 ;
      RECT 84.69 4.94 84.695 4.95 ;
      RECT 86.02 4.185 86.03 4.406 ;
      RECT 85.95 4.18 86.02 4.531 ;
      RECT 85.94 4.18 85.95 4.658 ;
      RECT 85.915 4.18 85.94 4.705 ;
      RECT 85.89 4.18 85.915 4.783 ;
      RECT 85.87 4.18 85.89 4.853 ;
      RECT 85.845 4.18 85.87 4.893 ;
      RECT 85.835 4.18 85.845 4.913 ;
      RECT 85.825 4.182 85.835 4.921 ;
      RECT 85.82 4.187 85.825 4.378 ;
      RECT 85.82 4.387 85.825 4.922 ;
      RECT 85.815 4.432 85.82 4.923 ;
      RECT 85.805 4.497 85.815 4.924 ;
      RECT 85.795 4.592 85.805 4.926 ;
      RECT 85.79 4.645 85.795 4.928 ;
      RECT 85.785 4.665 85.79 4.929 ;
      RECT 85.73 4.69 85.785 4.935 ;
      RECT 85.69 4.725 85.73 4.944 ;
      RECT 85.68 4.742 85.69 4.949 ;
      RECT 85.671 4.748 85.68 4.951 ;
      RECT 85.585 4.786 85.671 4.962 ;
      RECT 85.58 4.825 85.585 4.972 ;
      RECT 85.505 4.832 85.58 4.982 ;
      RECT 85.485 4.842 85.505 4.993 ;
      RECT 85.455 4.849 85.485 5.001 ;
      RECT 85.43 4.856 85.455 5.008 ;
      RECT 85.406 4.862 85.43 5.013 ;
      RECT 85.32 4.875 85.406 5.025 ;
      RECT 85.242 4.882 85.32 5.043 ;
      RECT 85.156 4.877 85.242 5.061 ;
      RECT 85.07 4.872 85.156 5.081 ;
      RECT 84.99 4.866 85.07 5.098 ;
      RECT 84.925 4.862 84.99 5.127 ;
      RECT 84.92 4.576 84.925 4.6 ;
      RECT 84.91 4.852 84.925 5.155 ;
      RECT 84.915 4.57 84.92 4.64 ;
      RECT 84.91 4.564 84.915 4.71 ;
      RECT 84.905 4.558 84.91 4.788 ;
      RECT 84.905 4.835 84.91 5.22 ;
      RECT 84.897 4.555 84.905 5.22 ;
      RECT 84.811 4.553 84.897 5.22 ;
      RECT 84.725 4.551 84.811 5.22 ;
      RECT 84.715 4.552 84.725 5.22 ;
      RECT 84.71 4.557 84.715 5.22 ;
      RECT 84.7 4.57 84.71 5.22 ;
      RECT 84.695 4.592 84.7 5.22 ;
      RECT 84.69 4.952 84.695 5.22 ;
      RECT 85.32 4.42 85.325 4.64 ;
      RECT 85.825 3.455 85.86 3.715 ;
      RECT 85.81 3.455 85.825 3.723 ;
      RECT 85.781 3.455 85.81 3.745 ;
      RECT 85.695 3.455 85.781 3.805 ;
      RECT 85.675 3.455 85.695 3.87 ;
      RECT 85.615 3.455 85.675 4.035 ;
      RECT 85.61 3.455 85.615 4.183 ;
      RECT 85.605 3.455 85.61 4.195 ;
      RECT 85.6 3.455 85.605 4.221 ;
      RECT 85.57 3.641 85.6 4.301 ;
      RECT 85.565 3.689 85.57 4.39 ;
      RECT 85.56 3.703 85.565 4.405 ;
      RECT 85.555 3.722 85.56 4.435 ;
      RECT 85.55 3.737 85.555 4.451 ;
      RECT 85.545 3.752 85.55 4.473 ;
      RECT 85.54 3.772 85.545 4.495 ;
      RECT 85.53 3.792 85.54 4.528 ;
      RECT 85.515 3.834 85.53 4.59 ;
      RECT 85.51 3.865 85.515 4.63 ;
      RECT 85.505 3.877 85.51 4.635 ;
      RECT 85.5 3.889 85.505 4.64 ;
      RECT 85.495 3.902 85.5 4.64 ;
      RECT 85.49 3.92 85.495 4.64 ;
      RECT 85.485 3.94 85.49 4.64 ;
      RECT 85.48 3.952 85.485 4.64 ;
      RECT 85.475 3.965 85.48 4.64 ;
      RECT 85.455 4 85.475 4.64 ;
      RECT 85.405 4.102 85.455 4.64 ;
      RECT 85.4 4.187 85.405 4.64 ;
      RECT 85.395 4.195 85.4 4.64 ;
      RECT 85.39 4.212 85.395 4.64 ;
      RECT 85.385 4.227 85.39 4.64 ;
      RECT 85.35 4.292 85.385 4.64 ;
      RECT 85.335 4.357 85.35 4.64 ;
      RECT 85.33 4.387 85.335 4.64 ;
      RECT 85.325 4.412 85.33 4.64 ;
      RECT 85.31 4.422 85.32 4.64 ;
      RECT 85.295 4.435 85.31 4.633 ;
      RECT 85.04 4.025 85.11 4.235 ;
      RECT 84.83 4.002 84.835 4.195 ;
      RECT 82.285 3.93 82.545 4.19 ;
      RECT 85.12 4.212 85.125 4.215 ;
      RECT 85.11 4.03 85.12 4.23 ;
      RECT 85.011 4.023 85.04 4.235 ;
      RECT 84.925 4.015 85.011 4.235 ;
      RECT 84.91 4.009 84.925 4.233 ;
      RECT 84.89 4.008 84.91 4.22 ;
      RECT 84.885 4.007 84.89 4.203 ;
      RECT 84.835 4.004 84.885 4.198 ;
      RECT 84.805 4.001 84.83 4.193 ;
      RECT 84.785 3.999 84.805 4.188 ;
      RECT 84.77 3.997 84.785 4.185 ;
      RECT 84.74 3.995 84.77 4.183 ;
      RECT 84.675 3.991 84.74 4.175 ;
      RECT 84.645 3.986 84.675 4.17 ;
      RECT 84.625 3.984 84.645 4.168 ;
      RECT 84.595 3.981 84.625 4.163 ;
      RECT 84.535 3.977 84.595 4.155 ;
      RECT 84.53 3.974 84.535 4.15 ;
      RECT 84.46 3.972 84.53 4.145 ;
      RECT 84.431 3.968 84.46 4.138 ;
      RECT 84.345 3.963 84.431 4.13 ;
      RECT 84.311 3.958 84.345 4.122 ;
      RECT 84.225 3.95 84.311 4.114 ;
      RECT 84.186 3.943 84.225 4.106 ;
      RECT 84.1 3.938 84.186 4.098 ;
      RECT 84.035 3.932 84.1 4.088 ;
      RECT 84.015 3.927 84.035 4.083 ;
      RECT 84.006 3.924 84.015 4.082 ;
      RECT 83.92 3.92 84.006 4.076 ;
      RECT 83.88 3.916 83.92 4.068 ;
      RECT 83.86 3.912 83.88 4.066 ;
      RECT 83.8 3.912 83.86 4.063 ;
      RECT 83.78 3.915 83.8 4.061 ;
      RECT 83.759 3.915 83.78 4.061 ;
      RECT 83.673 3.917 83.759 4.065 ;
      RECT 83.587 3.919 83.673 4.071 ;
      RECT 83.501 3.921 83.587 4.078 ;
      RECT 83.415 3.924 83.501 4.084 ;
      RECT 83.381 3.925 83.415 4.089 ;
      RECT 83.295 3.928 83.381 4.094 ;
      RECT 83.266 3.935 83.295 4.099 ;
      RECT 83.18 3.935 83.266 4.104 ;
      RECT 83.147 3.935 83.18 4.109 ;
      RECT 83.061 3.937 83.147 4.114 ;
      RECT 82.975 3.939 83.061 4.121 ;
      RECT 82.911 3.941 82.975 4.127 ;
      RECT 82.825 3.943 82.911 4.133 ;
      RECT 82.822 3.945 82.825 4.136 ;
      RECT 82.736 3.946 82.822 4.14 ;
      RECT 82.65 3.949 82.736 4.147 ;
      RECT 82.631 3.951 82.65 4.151 ;
      RECT 82.545 3.953 82.631 4.156 ;
      RECT 82.275 3.965 82.285 4.16 ;
      RECT 84.455 10.2 84.745 10.43 ;
      RECT 84.515 9.46 84.685 10.43 ;
      RECT 84.405 9.49 84.78 9.86 ;
      RECT 84.455 9.46 84.745 9.86 ;
      RECT 84.51 3.545 84.695 3.755 ;
      RECT 84.505 3.546 84.7 3.753 ;
      RECT 84.5 3.551 84.71 3.748 ;
      RECT 84.495 3.527 84.5 3.745 ;
      RECT 84.465 3.524 84.495 3.738 ;
      RECT 84.46 3.52 84.465 3.729 ;
      RECT 84.425 3.551 84.71 3.724 ;
      RECT 84.2 3.46 84.46 3.72 ;
      RECT 84.5 3.529 84.505 3.748 ;
      RECT 84.505 3.53 84.51 3.753 ;
      RECT 84.2 3.542 84.58 3.72 ;
      RECT 84.2 3.54 84.565 3.72 ;
      RECT 84.2 3.535 84.555 3.72 ;
      RECT 84.155 4.45 84.205 4.735 ;
      RECT 84.1 4.42 84.105 4.735 ;
      RECT 84.07 4.4 84.075 4.735 ;
      RECT 84.22 4.45 84.28 4.71 ;
      RECT 84.215 4.45 84.22 4.718 ;
      RECT 84.205 4.45 84.215 4.73 ;
      RECT 84.12 4.44 84.155 4.735 ;
      RECT 84.115 4.427 84.12 4.735 ;
      RECT 84.105 4.422 84.115 4.735 ;
      RECT 84.085 4.412 84.1 4.735 ;
      RECT 84.075 4.405 84.085 4.735 ;
      RECT 84.065 4.397 84.07 4.735 ;
      RECT 84.035 4.387 84.065 4.735 ;
      RECT 84.02 4.375 84.035 4.735 ;
      RECT 84.005 4.365 84.02 4.73 ;
      RECT 83.985 4.355 84.005 4.705 ;
      RECT 83.975 4.347 83.985 4.682 ;
      RECT 83.945 4.33 83.975 4.672 ;
      RECT 83.94 4.307 83.945 4.663 ;
      RECT 83.935 4.294 83.94 4.661 ;
      RECT 83.92 4.27 83.935 4.655 ;
      RECT 83.915 4.246 83.92 4.649 ;
      RECT 83.905 4.235 83.915 4.644 ;
      RECT 83.9 4.225 83.905 4.64 ;
      RECT 83.895 4.217 83.9 4.637 ;
      RECT 83.885 4.212 83.895 4.633 ;
      RECT 83.88 4.207 83.885 4.629 ;
      RECT 83.795 4.205 83.88 4.604 ;
      RECT 83.765 4.205 83.795 4.57 ;
      RECT 83.75 4.205 83.765 4.553 ;
      RECT 83.695 4.205 83.75 4.498 ;
      RECT 83.69 4.21 83.695 4.447 ;
      RECT 83.68 4.215 83.69 4.437 ;
      RECT 83.675 4.225 83.68 4.423 ;
      RECT 83.625 4.965 83.885 5.225 ;
      RECT 83.545 4.98 83.885 5.201 ;
      RECT 83.525 4.98 83.885 5.196 ;
      RECT 83.501 4.98 83.885 5.194 ;
      RECT 83.415 4.98 83.885 5.189 ;
      RECT 83.265 4.92 83.525 5.185 ;
      RECT 83.22 4.98 83.885 5.18 ;
      RECT 83.215 4.987 83.885 5.175 ;
      RECT 83.23 4.975 83.545 5.185 ;
      RECT 83.12 3.41 83.38 3.67 ;
      RECT 83.12 3.467 83.385 3.663 ;
      RECT 83.12 3.497 83.39 3.595 ;
      RECT 83.18 3.928 83.295 3.93 ;
      RECT 83.266 3.925 83.295 3.93 ;
      RECT 82.29 4.929 82.315 5.169 ;
      RECT 82.275 4.932 82.365 5.163 ;
      RECT 82.27 4.937 82.451 5.158 ;
      RECT 82.265 4.945 82.515 5.156 ;
      RECT 82.265 4.945 82.525 5.155 ;
      RECT 82.26 4.952 82.535 5.148 ;
      RECT 82.26 4.952 82.621 5.137 ;
      RECT 82.255 4.987 82.621 5.133 ;
      RECT 82.255 4.987 82.63 5.122 ;
      RECT 82.535 4.86 82.795 5.12 ;
      RECT 82.245 5.037 82.795 5.118 ;
      RECT 82.515 4.905 82.535 5.153 ;
      RECT 82.451 4.908 82.515 5.157 ;
      RECT 82.365 4.913 82.451 5.162 ;
      RECT 82.295 4.924 82.795 5.12 ;
      RECT 82.315 4.918 82.365 5.167 ;
      RECT 82.44 3.395 82.45 3.657 ;
      RECT 82.43 3.452 82.44 3.66 ;
      RECT 82.405 3.457 82.43 3.666 ;
      RECT 82.38 3.461 82.405 3.678 ;
      RECT 82.37 3.464 82.38 3.688 ;
      RECT 82.365 3.465 82.37 3.693 ;
      RECT 82.36 3.466 82.365 3.698 ;
      RECT 82.355 3.467 82.36 3.7 ;
      RECT 82.33 3.47 82.355 3.703 ;
      RECT 82.3 3.476 82.33 3.706 ;
      RECT 82.235 3.487 82.3 3.709 ;
      RECT 82.19 3.495 82.235 3.713 ;
      RECT 82.175 3.495 82.19 3.721 ;
      RECT 82.17 3.496 82.175 3.728 ;
      RECT 82.165 3.498 82.17 3.731 ;
      RECT 82.16 3.502 82.165 3.734 ;
      RECT 82.15 3.51 82.16 3.738 ;
      RECT 82.145 3.523 82.15 3.743 ;
      RECT 82.14 3.531 82.145 3.745 ;
      RECT 82.135 3.537 82.14 3.745 ;
      RECT 82.13 3.541 82.135 3.748 ;
      RECT 82.125 3.543 82.13 3.751 ;
      RECT 82.12 3.546 82.125 3.754 ;
      RECT 82.11 3.551 82.12 3.758 ;
      RECT 82.105 3.557 82.11 3.763 ;
      RECT 82.095 3.563 82.105 3.767 ;
      RECT 82.08 3.57 82.095 3.773 ;
      RECT 82.051 3.584 82.08 3.783 ;
      RECT 81.965 3.619 82.051 3.815 ;
      RECT 81.945 3.652 81.965 3.844 ;
      RECT 81.925 3.665 81.945 3.855 ;
      RECT 81.905 3.677 81.925 3.866 ;
      RECT 81.855 3.699 81.905 3.886 ;
      RECT 81.84 3.717 81.855 3.903 ;
      RECT 81.835 3.723 81.84 3.906 ;
      RECT 81.83 3.727 81.835 3.909 ;
      RECT 81.825 3.731 81.83 3.913 ;
      RECT 81.82 3.733 81.825 3.916 ;
      RECT 81.81 3.74 81.82 3.919 ;
      RECT 81.805 3.745 81.81 3.923 ;
      RECT 81.8 3.747 81.805 3.926 ;
      RECT 81.795 3.751 81.8 3.929 ;
      RECT 81.79 3.753 81.795 3.933 ;
      RECT 81.775 3.758 81.79 3.938 ;
      RECT 81.77 3.763 81.775 3.941 ;
      RECT 81.765 3.771 81.77 3.944 ;
      RECT 81.76 3.773 81.765 3.947 ;
      RECT 81.755 3.775 81.76 3.95 ;
      RECT 81.745 3.777 81.755 3.956 ;
      RECT 81.71 3.791 81.745 3.968 ;
      RECT 81.7 3.806 81.71 3.978 ;
      RECT 81.625 3.835 81.7 4.002 ;
      RECT 81.62 3.86 81.625 4.025 ;
      RECT 81.605 3.864 81.62 4.031 ;
      RECT 81.595 3.872 81.605 4.036 ;
      RECT 81.565 3.885 81.595 4.04 ;
      RECT 81.555 3.9 81.565 4.045 ;
      RECT 81.545 3.905 81.555 4.048 ;
      RECT 81.54 3.907 81.545 4.05 ;
      RECT 81.525 3.91 81.54 4.053 ;
      RECT 81.52 3.912 81.525 4.056 ;
      RECT 81.5 3.917 81.52 4.06 ;
      RECT 81.47 3.922 81.5 4.068 ;
      RECT 81.445 3.929 81.47 4.076 ;
      RECT 81.44 3.934 81.445 4.081 ;
      RECT 81.41 3.937 81.44 4.085 ;
      RECT 81.37 3.94 81.41 4.095 ;
      RECT 81.335 3.937 81.37 4.107 ;
      RECT 81.325 3.933 81.335 4.114 ;
      RECT 81.3 3.929 81.325 4.12 ;
      RECT 81.295 3.925 81.3 4.125 ;
      RECT 81.255 3.922 81.295 4.125 ;
      RECT 81.24 3.907 81.255 4.126 ;
      RECT 81.217 3.895 81.24 4.126 ;
      RECT 81.131 3.895 81.217 4.127 ;
      RECT 81.045 3.895 81.131 4.129 ;
      RECT 81.025 3.895 81.045 4.126 ;
      RECT 81.02 3.9 81.025 4.121 ;
      RECT 81.015 3.905 81.02 4.119 ;
      RECT 81.005 3.915 81.015 4.117 ;
      RECT 81 3.921 81.005 4.11 ;
      RECT 80.995 3.923 81 4.095 ;
      RECT 80.99 3.927 80.995 4.085 ;
      RECT 82.45 3.395 82.7 3.655 ;
      RECT 80.175 4.93 80.435 5.19 ;
      RECT 82.47 4.42 82.475 4.63 ;
      RECT 82.475 4.425 82.485 4.625 ;
      RECT 82.425 4.42 82.47 4.645 ;
      RECT 82.415 4.42 82.425 4.665 ;
      RECT 82.396 4.42 82.415 4.67 ;
      RECT 82.31 4.42 82.396 4.667 ;
      RECT 82.28 4.422 82.31 4.665 ;
      RECT 82.225 4.432 82.28 4.663 ;
      RECT 82.16 4.446 82.225 4.661 ;
      RECT 82.155 4.454 82.16 4.66 ;
      RECT 82.14 4.457 82.155 4.658 ;
      RECT 82.075 4.467 82.14 4.654 ;
      RECT 82.027 4.481 82.075 4.655 ;
      RECT 81.941 4.498 82.027 4.669 ;
      RECT 81.855 4.519 81.941 4.686 ;
      RECT 81.835 4.532 81.855 4.696 ;
      RECT 81.79 4.54 81.835 4.703 ;
      RECT 81.755 4.548 81.79 4.711 ;
      RECT 81.721 4.556 81.755 4.719 ;
      RECT 81.635 4.57 81.721 4.731 ;
      RECT 81.6 4.587 81.635 4.743 ;
      RECT 81.591 4.596 81.6 4.747 ;
      RECT 81.505 4.614 81.591 4.764 ;
      RECT 81.446 4.641 81.505 4.791 ;
      RECT 81.36 4.668 81.446 4.819 ;
      RECT 81.34 4.69 81.36 4.839 ;
      RECT 81.28 4.705 81.34 4.855 ;
      RECT 81.27 4.717 81.28 4.868 ;
      RECT 81.265 4.722 81.27 4.871 ;
      RECT 81.255 4.725 81.265 4.874 ;
      RECT 81.25 4.727 81.255 4.877 ;
      RECT 81.22 4.735 81.25 4.884 ;
      RECT 81.205 4.742 81.22 4.892 ;
      RECT 81.195 4.747 81.205 4.896 ;
      RECT 81.19 4.75 81.195 4.899 ;
      RECT 81.18 4.752 81.19 4.902 ;
      RECT 81.145 4.762 81.18 4.911 ;
      RECT 81.07 4.785 81.145 4.933 ;
      RECT 81.05 4.803 81.07 4.951 ;
      RECT 81.02 4.81 81.05 4.961 ;
      RECT 81 4.818 81.02 4.971 ;
      RECT 80.99 4.824 81 4.978 ;
      RECT 80.971 4.829 80.99 4.984 ;
      RECT 80.885 4.849 80.971 5.004 ;
      RECT 80.87 4.869 80.885 5.023 ;
      RECT 80.825 4.881 80.87 5.034 ;
      RECT 80.76 4.902 80.825 5.057 ;
      RECT 80.72 4.922 80.76 5.078 ;
      RECT 80.71 4.932 80.72 5.088 ;
      RECT 80.66 4.944 80.71 5.099 ;
      RECT 80.64 4.96 80.66 5.111 ;
      RECT 80.61 4.97 80.64 5.117 ;
      RECT 80.6 4.975 80.61 5.119 ;
      RECT 80.531 4.976 80.6 5.125 ;
      RECT 80.445 4.978 80.531 5.135 ;
      RECT 80.435 4.979 80.445 5.14 ;
      RECT 81.705 5.005 81.895 5.215 ;
      RECT 81.695 5.01 81.905 5.208 ;
      RECT 81.68 5.01 81.905 5.173 ;
      RECT 81.6 4.895 81.86 5.155 ;
      RECT 80.515 4.425 80.7 4.72 ;
      RECT 80.505 4.425 80.7 4.718 ;
      RECT 80.49 4.425 80.705 4.713 ;
      RECT 80.49 4.425 80.71 4.71 ;
      RECT 80.485 4.425 80.71 4.708 ;
      RECT 80.48 4.68 80.71 4.698 ;
      RECT 80.485 4.425 80.745 4.685 ;
      RECT 80.445 3.46 80.705 3.72 ;
      RECT 80.255 3.385 80.341 3.718 ;
      RECT 80.23 3.389 80.385 3.714 ;
      RECT 80.341 3.381 80.385 3.714 ;
      RECT 80.341 3.382 80.39 3.713 ;
      RECT 80.255 3.387 80.405 3.712 ;
      RECT 80.23 3.395 80.445 3.711 ;
      RECT 80.225 3.39 80.405 3.706 ;
      RECT 80.215 3.405 80.445 3.613 ;
      RECT 80.215 3.457 80.645 3.613 ;
      RECT 80.215 3.45 80.625 3.613 ;
      RECT 80.215 3.437 80.595 3.613 ;
      RECT 80.215 3.425 80.535 3.613 ;
      RECT 80.215 3.41 80.51 3.613 ;
      RECT 79.415 4.04 79.55 4.335 ;
      RECT 79.675 4.063 79.68 4.25 ;
      RECT 80.395 3.96 80.54 4.195 ;
      RECT 80.555 3.96 80.56 4.185 ;
      RECT 80.59 3.971 80.595 4.165 ;
      RECT 80.585 3.963 80.59 4.17 ;
      RECT 80.565 3.96 80.585 4.175 ;
      RECT 80.56 3.96 80.565 4.183 ;
      RECT 80.55 3.96 80.555 4.188 ;
      RECT 80.54 3.96 80.55 4.193 ;
      RECT 80.37 3.962 80.395 4.195 ;
      RECT 80.32 3.969 80.37 4.195 ;
      RECT 80.315 3.974 80.32 4.195 ;
      RECT 80.276 3.979 80.315 4.196 ;
      RECT 80.19 3.991 80.276 4.197 ;
      RECT 80.181 4.001 80.19 4.197 ;
      RECT 80.095 4.01 80.181 4.199 ;
      RECT 80.071 4.02 80.095 4.201 ;
      RECT 79.985 4.031 80.071 4.202 ;
      RECT 79.955 4.042 79.985 4.204 ;
      RECT 79.925 4.047 79.955 4.206 ;
      RECT 79.9 4.053 79.925 4.209 ;
      RECT 79.885 4.058 79.9 4.21 ;
      RECT 79.84 4.064 79.885 4.21 ;
      RECT 79.835 4.069 79.84 4.211 ;
      RECT 79.815 4.069 79.835 4.213 ;
      RECT 79.795 4.067 79.815 4.218 ;
      RECT 79.76 4.066 79.795 4.225 ;
      RECT 79.73 4.065 79.76 4.235 ;
      RECT 79.68 4.064 79.73 4.245 ;
      RECT 79.59 4.061 79.675 4.335 ;
      RECT 79.565 4.055 79.59 4.335 ;
      RECT 79.55 4.045 79.565 4.335 ;
      RECT 79.365 4.04 79.415 4.255 ;
      RECT 79.355 4.045 79.365 4.245 ;
      RECT 79.595 4.52 79.855 4.78 ;
      RECT 79.595 4.52 79.885 4.673 ;
      RECT 79.595 4.52 79.92 4.658 ;
      RECT 79.85 4.44 80.04 4.65 ;
      RECT 79.84 4.445 80.05 4.643 ;
      RECT 79.805 4.515 80.05 4.643 ;
      RECT 79.835 4.457 79.855 4.78 ;
      RECT 79.82 4.505 80.05 4.643 ;
      RECT 79.825 4.477 79.855 4.78 ;
      RECT 78.905 3.545 78.975 4.65 ;
      RECT 79.64 3.65 79.9 3.91 ;
      RECT 79.22 3.696 79.235 3.905 ;
      RECT 79.556 3.709 79.64 3.86 ;
      RECT 79.47 3.706 79.556 3.86 ;
      RECT 79.431 3.704 79.47 3.86 ;
      RECT 79.345 3.702 79.431 3.86 ;
      RECT 79.285 3.7 79.345 3.871 ;
      RECT 79.25 3.698 79.285 3.889 ;
      RECT 79.235 3.696 79.25 3.9 ;
      RECT 79.205 3.696 79.22 3.913 ;
      RECT 79.195 3.696 79.205 3.918 ;
      RECT 79.17 3.695 79.195 3.923 ;
      RECT 79.155 3.69 79.17 3.929 ;
      RECT 79.15 3.683 79.155 3.934 ;
      RECT 79.125 3.674 79.15 3.94 ;
      RECT 79.08 3.653 79.125 3.953 ;
      RECT 79.07 3.637 79.08 3.963 ;
      RECT 79.055 3.63 79.07 3.973 ;
      RECT 79.045 3.623 79.055 3.99 ;
      RECT 79.04 3.62 79.045 4.02 ;
      RECT 79.035 3.618 79.04 4.05 ;
      RECT 79.03 3.616 79.035 4.087 ;
      RECT 79.015 3.612 79.03 4.154 ;
      RECT 79.015 4.445 79.025 4.645 ;
      RECT 79.01 3.608 79.015 4.28 ;
      RECT 79.01 4.432 79.015 4.65 ;
      RECT 79.005 3.606 79.01 4.365 ;
      RECT 79.005 4.422 79.01 4.65 ;
      RECT 78.99 3.577 79.005 4.65 ;
      RECT 78.975 3.55 78.99 4.65 ;
      RECT 78.9 3.545 78.905 3.9 ;
      RECT 78.9 3.955 78.905 4.65 ;
      RECT 78.885 3.545 78.9 3.878 ;
      RECT 78.895 3.977 78.9 4.65 ;
      RECT 78.885 4.017 78.895 4.65 ;
      RECT 78.85 3.545 78.885 3.82 ;
      RECT 78.88 4.052 78.885 4.65 ;
      RECT 78.865 4.107 78.88 4.65 ;
      RECT 78.86 4.172 78.865 4.65 ;
      RECT 78.845 4.22 78.86 4.65 ;
      RECT 78.82 3.545 78.85 3.775 ;
      RECT 78.84 4.275 78.845 4.65 ;
      RECT 78.825 4.335 78.84 4.65 ;
      RECT 78.82 4.383 78.825 4.648 ;
      RECT 78.815 3.545 78.82 3.768 ;
      RECT 78.815 4.415 78.82 4.643 ;
      RECT 78.79 3.545 78.815 3.76 ;
      RECT 78.78 3.55 78.79 3.75 ;
      RECT 78.995 4.825 79.015 5.065 ;
      RECT 78.225 4.755 78.23 4.965 ;
      RECT 79.505 4.828 79.515 5.023 ;
      RECT 79.5 4.818 79.505 5.026 ;
      RECT 79.42 4.815 79.5 5.049 ;
      RECT 79.416 4.815 79.42 5.071 ;
      RECT 79.33 4.815 79.416 5.081 ;
      RECT 79.315 4.815 79.33 5.089 ;
      RECT 79.286 4.816 79.315 5.087 ;
      RECT 79.2 4.821 79.286 5.083 ;
      RECT 79.187 4.825 79.2 5.079 ;
      RECT 79.101 4.825 79.187 5.075 ;
      RECT 79.015 4.825 79.101 5.069 ;
      RECT 78.931 4.825 78.995 5.063 ;
      RECT 78.845 4.825 78.931 5.058 ;
      RECT 78.825 4.825 78.845 5.054 ;
      RECT 78.765 4.82 78.825 5.051 ;
      RECT 78.737 4.814 78.765 5.048 ;
      RECT 78.651 4.809 78.737 5.044 ;
      RECT 78.565 4.803 78.651 5.038 ;
      RECT 78.49 4.785 78.565 5.033 ;
      RECT 78.455 4.762 78.49 5.029 ;
      RECT 78.445 4.752 78.455 5.028 ;
      RECT 78.39 4.75 78.445 5.027 ;
      RECT 78.315 4.75 78.39 5.023 ;
      RECT 78.305 4.75 78.315 5.018 ;
      RECT 78.29 4.75 78.305 5.01 ;
      RECT 78.24 4.752 78.29 4.988 ;
      RECT 78.23 4.755 78.24 4.968 ;
      RECT 78.22 4.76 78.225 4.963 ;
      RECT 78.215 4.765 78.22 4.958 ;
      RECT 78.34 3.93 78.6 4.19 ;
      RECT 78.34 3.945 78.62 4.155 ;
      RECT 78.34 3.95 78.63 4.15 ;
      RECT 76.325 3.41 76.585 3.67 ;
      RECT 76.315 3.44 76.585 3.65 ;
      RECT 78.235 3.355 78.495 3.615 ;
      RECT 78.23 3.43 78.235 3.616 ;
      RECT 78.205 3.435 78.23 3.618 ;
      RECT 78.19 3.442 78.205 3.621 ;
      RECT 78.13 3.46 78.19 3.626 ;
      RECT 78.1 3.48 78.13 3.633 ;
      RECT 78.075 3.488 78.1 3.638 ;
      RECT 78.05 3.496 78.075 3.64 ;
      RECT 78.032 3.5 78.05 3.639 ;
      RECT 77.946 3.498 78.032 3.639 ;
      RECT 77.86 3.496 77.946 3.639 ;
      RECT 77.774 3.494 77.86 3.638 ;
      RECT 77.688 3.492 77.774 3.638 ;
      RECT 77.602 3.49 77.688 3.638 ;
      RECT 77.516 3.488 77.602 3.638 ;
      RECT 77.43 3.486 77.516 3.637 ;
      RECT 77.412 3.485 77.43 3.637 ;
      RECT 77.326 3.484 77.412 3.637 ;
      RECT 77.24 3.482 77.326 3.637 ;
      RECT 77.154 3.481 77.24 3.636 ;
      RECT 77.068 3.48 77.154 3.636 ;
      RECT 76.982 3.478 77.068 3.636 ;
      RECT 76.896 3.477 76.982 3.636 ;
      RECT 76.81 3.475 76.896 3.635 ;
      RECT 76.786 3.473 76.81 3.635 ;
      RECT 76.7 3.466 76.786 3.635 ;
      RECT 76.671 3.458 76.7 3.635 ;
      RECT 76.585 3.45 76.671 3.635 ;
      RECT 76.305 3.447 76.315 3.645 ;
      RECT 77.81 4.41 77.815 4.76 ;
      RECT 77.58 4.5 77.72 4.76 ;
      RECT 78.055 4.185 78.1 4.395 ;
      RECT 78.11 4.196 78.12 4.39 ;
      RECT 78.1 4.188 78.11 4.395 ;
      RECT 78.035 4.185 78.055 4.4 ;
      RECT 78.005 4.185 78.035 4.423 ;
      RECT 77.995 4.185 78.005 4.448 ;
      RECT 77.99 4.185 77.995 4.458 ;
      RECT 77.935 4.185 77.99 4.498 ;
      RECT 77.93 4.185 77.935 4.538 ;
      RECT 77.925 4.187 77.93 4.543 ;
      RECT 77.91 4.197 77.925 4.554 ;
      RECT 77.865 4.255 77.91 4.59 ;
      RECT 77.855 4.31 77.865 4.624 ;
      RECT 77.84 4.337 77.855 4.64 ;
      RECT 77.83 4.364 77.84 4.76 ;
      RECT 77.815 4.387 77.83 4.76 ;
      RECT 77.805 4.427 77.81 4.76 ;
      RECT 77.8 4.437 77.805 4.76 ;
      RECT 77.795 4.452 77.8 4.76 ;
      RECT 77.785 4.457 77.795 4.76 ;
      RECT 77.72 4.48 77.785 4.76 ;
      RECT 77.22 3.975 77.41 4.185 ;
      RECT 75.795 3.9 76.055 4.16 ;
      RECT 76.145 3.895 76.24 4.105 ;
      RECT 76.12 3.91 76.13 4.105 ;
      RECT 77.41 3.982 77.42 4.18 ;
      RECT 77.21 3.982 77.22 4.18 ;
      RECT 77.195 3.997 77.21 4.17 ;
      RECT 77.19 4.005 77.195 4.163 ;
      RECT 77.18 4.008 77.19 4.16 ;
      RECT 77.145 4.007 77.18 4.158 ;
      RECT 77.116 4.003 77.145 4.155 ;
      RECT 77.03 3.998 77.116 4.152 ;
      RECT 76.97 3.992 77.03 4.148 ;
      RECT 76.941 3.988 76.97 4.145 ;
      RECT 76.855 3.98 76.941 4.142 ;
      RECT 76.846 3.974 76.855 4.14 ;
      RECT 76.76 3.969 76.846 4.138 ;
      RECT 76.737 3.964 76.76 4.135 ;
      RECT 76.651 3.958 76.737 4.132 ;
      RECT 76.565 3.949 76.651 4.127 ;
      RECT 76.555 3.944 76.565 4.125 ;
      RECT 76.536 3.943 76.555 4.124 ;
      RECT 76.45 3.938 76.536 4.12 ;
      RECT 76.43 3.933 76.45 4.116 ;
      RECT 76.37 3.928 76.43 4.113 ;
      RECT 76.345 3.918 76.37 4.111 ;
      RECT 76.34 3.911 76.345 4.11 ;
      RECT 76.33 3.902 76.34 4.109 ;
      RECT 76.326 3.895 76.33 4.109 ;
      RECT 76.24 3.895 76.326 4.107 ;
      RECT 76.13 3.902 76.145 4.105 ;
      RECT 76.115 3.912 76.12 4.105 ;
      RECT 76.095 3.915 76.115 4.102 ;
      RECT 76.065 3.915 76.095 4.098 ;
      RECT 76.055 3.915 76.065 4.098 ;
      RECT 76.97 4.41 77.23 4.67 ;
      RECT 76.9 4.42 77.23 4.63 ;
      RECT 76.89 4.427 77.23 4.625 ;
      RECT 76.31 4.415 76.57 4.675 ;
      RECT 76.31 4.455 76.675 4.665 ;
      RECT 76.31 4.457 76.68 4.664 ;
      RECT 76.31 4.465 76.685 4.661 ;
      RECT 75.235 3.54 75.335 5.065 ;
      RECT 75.425 4.68 75.475 4.94 ;
      RECT 75.42 3.553 75.425 3.74 ;
      RECT 75.415 4.661 75.425 4.94 ;
      RECT 75.415 3.55 75.42 3.748 ;
      RECT 75.4 3.544 75.415 3.755 ;
      RECT 75.41 4.649 75.415 5.023 ;
      RECT 75.4 4.637 75.41 5.06 ;
      RECT 75.39 3.54 75.4 3.762 ;
      RECT 75.39 4.622 75.4 5.065 ;
      RECT 75.385 3.54 75.39 3.77 ;
      RECT 75.365 4.592 75.39 5.065 ;
      RECT 75.345 3.54 75.385 3.818 ;
      RECT 75.355 4.552 75.365 5.065 ;
      RECT 75.345 4.507 75.355 5.065 ;
      RECT 75.34 3.54 75.345 3.888 ;
      RECT 75.34 4.465 75.345 5.065 ;
      RECT 75.335 3.54 75.34 4.365 ;
      RECT 75.335 4.447 75.34 5.065 ;
      RECT 75.225 3.543 75.235 5.065 ;
      RECT 75.21 3.55 75.225 5.061 ;
      RECT 75.205 3.56 75.21 5.056 ;
      RECT 75.2 3.76 75.205 4.948 ;
      RECT 75.195 3.845 75.2 4.5 ;
      RECT 74.07 10.205 74.36 10.435 ;
      RECT 74.13 8.725 74.3 10.435 ;
      RECT 74.08 9.09 74.43 9.44 ;
      RECT 74.07 8.725 74.36 8.955 ;
      RECT 73.665 3.69 73.77 4.26 ;
      RECT 73.665 4.025 73.99 4.255 ;
      RECT 73.665 4.055 74.16 4.225 ;
      RECT 73.665 3.69 73.855 4.255 ;
      RECT 73.08 3.655 73.37 3.885 ;
      RECT 73.08 3.69 73.855 3.86 ;
      RECT 73.14 2.175 73.31 3.885 ;
      RECT 73.08 2.175 73.37 2.405 ;
      RECT 73.08 10.205 73.37 10.435 ;
      RECT 73.14 8.725 73.31 10.435 ;
      RECT 73.08 8.725 73.37 8.955 ;
      RECT 73.08 8.76 73.935 8.92 ;
      RECT 73.765 8.355 73.935 8.92 ;
      RECT 73.08 8.755 73.475 8.92 ;
      RECT 73.7 8.355 73.99 8.585 ;
      RECT 73.7 8.385 74.16 8.555 ;
      RECT 72.71 4.025 73 4.255 ;
      RECT 72.71 4.055 73.17 4.225 ;
      RECT 72.775 2.95 72.94 4.255 ;
      RECT 71.29 2.92 71.58 3.15 ;
      RECT 71.29 2.95 72.94 3.12 ;
      RECT 71.35 2.18 71.52 3.15 ;
      RECT 71.29 2.18 71.58 2.41 ;
      RECT 71.29 10.2 71.58 10.43 ;
      RECT 71.35 9.46 71.52 10.43 ;
      RECT 71.35 9.555 72.94 9.725 ;
      RECT 72.77 8.355 72.94 9.725 ;
      RECT 71.29 9.46 71.58 9.69 ;
      RECT 72.71 8.355 73 8.585 ;
      RECT 72.71 8.385 73.17 8.555 ;
      RECT 69.325 4.725 69.675 5.075 ;
      RECT 69.415 3.32 69.585 5.075 ;
      RECT 71.72 3.26 72.07 3.61 ;
      RECT 69.415 3.32 71.035 3.495 ;
      RECT 69.415 3.32 72.07 3.49 ;
      RECT 71.745 9.09 72.07 9.415 ;
      RECT 67.12 9.045 67.47 9.395 ;
      RECT 71.72 9.09 72.07 9.32 ;
      RECT 66.96 9.09 67.47 9.32 ;
      RECT 66.79 9.12 72.07 9.29 ;
      RECT 70.945 3.66 71.265 3.98 ;
      RECT 70.915 3.66 71.265 3.89 ;
      RECT 70.745 3.69 71.265 3.86 ;
      RECT 70.945 8.66 71.265 8.98 ;
      RECT 70.915 8.72 71.265 8.95 ;
      RECT 70.745 8.75 71.265 8.92 ;
      RECT 66.725 4.96 66.765 5.22 ;
      RECT 66.765 4.94 66.77 4.95 ;
      RECT 68.095 4.185 68.105 4.406 ;
      RECT 68.025 4.18 68.095 4.531 ;
      RECT 68.015 4.18 68.025 4.658 ;
      RECT 67.99 4.18 68.015 4.705 ;
      RECT 67.965 4.18 67.99 4.783 ;
      RECT 67.945 4.18 67.965 4.853 ;
      RECT 67.92 4.18 67.945 4.893 ;
      RECT 67.91 4.18 67.92 4.913 ;
      RECT 67.9 4.182 67.91 4.921 ;
      RECT 67.895 4.187 67.9 4.378 ;
      RECT 67.895 4.387 67.9 4.922 ;
      RECT 67.89 4.432 67.895 4.923 ;
      RECT 67.88 4.497 67.89 4.924 ;
      RECT 67.87 4.592 67.88 4.926 ;
      RECT 67.865 4.645 67.87 4.928 ;
      RECT 67.86 4.665 67.865 4.929 ;
      RECT 67.805 4.69 67.86 4.935 ;
      RECT 67.765 4.725 67.805 4.944 ;
      RECT 67.755 4.742 67.765 4.949 ;
      RECT 67.746 4.748 67.755 4.951 ;
      RECT 67.66 4.786 67.746 4.962 ;
      RECT 67.655 4.825 67.66 4.972 ;
      RECT 67.58 4.832 67.655 4.982 ;
      RECT 67.56 4.842 67.58 4.993 ;
      RECT 67.53 4.849 67.56 5.001 ;
      RECT 67.505 4.856 67.53 5.008 ;
      RECT 67.481 4.862 67.505 5.013 ;
      RECT 67.395 4.875 67.481 5.025 ;
      RECT 67.317 4.882 67.395 5.043 ;
      RECT 67.231 4.877 67.317 5.061 ;
      RECT 67.145 4.872 67.231 5.081 ;
      RECT 67.065 4.866 67.145 5.098 ;
      RECT 67 4.862 67.065 5.127 ;
      RECT 66.995 4.576 67 4.6 ;
      RECT 66.985 4.852 67 5.155 ;
      RECT 66.99 4.57 66.995 4.64 ;
      RECT 66.985 4.564 66.99 4.71 ;
      RECT 66.98 4.558 66.985 4.788 ;
      RECT 66.98 4.835 66.985 5.22 ;
      RECT 66.972 4.555 66.98 5.22 ;
      RECT 66.886 4.553 66.972 5.22 ;
      RECT 66.8 4.551 66.886 5.22 ;
      RECT 66.79 4.552 66.8 5.22 ;
      RECT 66.785 4.557 66.79 5.22 ;
      RECT 66.775 4.57 66.785 5.22 ;
      RECT 66.77 4.592 66.775 5.22 ;
      RECT 66.765 4.952 66.77 5.22 ;
      RECT 67.395 4.42 67.4 4.64 ;
      RECT 67.9 3.455 67.935 3.715 ;
      RECT 67.885 3.455 67.9 3.723 ;
      RECT 67.856 3.455 67.885 3.745 ;
      RECT 67.77 3.455 67.856 3.805 ;
      RECT 67.75 3.455 67.77 3.87 ;
      RECT 67.69 3.455 67.75 4.035 ;
      RECT 67.685 3.455 67.69 4.183 ;
      RECT 67.68 3.455 67.685 4.195 ;
      RECT 67.675 3.455 67.68 4.221 ;
      RECT 67.645 3.641 67.675 4.301 ;
      RECT 67.64 3.689 67.645 4.39 ;
      RECT 67.635 3.703 67.64 4.405 ;
      RECT 67.63 3.722 67.635 4.435 ;
      RECT 67.625 3.737 67.63 4.451 ;
      RECT 67.62 3.752 67.625 4.473 ;
      RECT 67.615 3.772 67.62 4.495 ;
      RECT 67.605 3.792 67.615 4.528 ;
      RECT 67.59 3.834 67.605 4.59 ;
      RECT 67.585 3.865 67.59 4.63 ;
      RECT 67.58 3.877 67.585 4.635 ;
      RECT 67.575 3.889 67.58 4.64 ;
      RECT 67.57 3.902 67.575 4.64 ;
      RECT 67.565 3.92 67.57 4.64 ;
      RECT 67.56 3.94 67.565 4.64 ;
      RECT 67.555 3.952 67.56 4.64 ;
      RECT 67.55 3.965 67.555 4.64 ;
      RECT 67.53 4 67.55 4.64 ;
      RECT 67.48 4.102 67.53 4.64 ;
      RECT 67.475 4.187 67.48 4.64 ;
      RECT 67.47 4.195 67.475 4.64 ;
      RECT 67.465 4.212 67.47 4.64 ;
      RECT 67.46 4.227 67.465 4.64 ;
      RECT 67.425 4.292 67.46 4.64 ;
      RECT 67.41 4.357 67.425 4.64 ;
      RECT 67.405 4.387 67.41 4.64 ;
      RECT 67.4 4.412 67.405 4.64 ;
      RECT 67.385 4.422 67.395 4.64 ;
      RECT 67.37 4.435 67.385 4.633 ;
      RECT 67.115 4.025 67.185 4.235 ;
      RECT 66.905 4.002 66.91 4.195 ;
      RECT 64.36 3.93 64.62 4.19 ;
      RECT 67.195 4.212 67.2 4.215 ;
      RECT 67.185 4.03 67.195 4.23 ;
      RECT 67.086 4.023 67.115 4.235 ;
      RECT 67 4.015 67.086 4.235 ;
      RECT 66.985 4.009 67 4.233 ;
      RECT 66.965 4.008 66.985 4.22 ;
      RECT 66.96 4.007 66.965 4.203 ;
      RECT 66.91 4.004 66.96 4.198 ;
      RECT 66.88 4.001 66.905 4.193 ;
      RECT 66.86 3.999 66.88 4.188 ;
      RECT 66.845 3.997 66.86 4.185 ;
      RECT 66.815 3.995 66.845 4.183 ;
      RECT 66.75 3.991 66.815 4.175 ;
      RECT 66.72 3.986 66.75 4.17 ;
      RECT 66.7 3.984 66.72 4.168 ;
      RECT 66.67 3.981 66.7 4.163 ;
      RECT 66.61 3.977 66.67 4.155 ;
      RECT 66.605 3.974 66.61 4.15 ;
      RECT 66.535 3.972 66.605 4.145 ;
      RECT 66.506 3.968 66.535 4.138 ;
      RECT 66.42 3.963 66.506 4.13 ;
      RECT 66.386 3.958 66.42 4.122 ;
      RECT 66.3 3.95 66.386 4.114 ;
      RECT 66.261 3.943 66.3 4.106 ;
      RECT 66.175 3.938 66.261 4.098 ;
      RECT 66.11 3.932 66.175 4.088 ;
      RECT 66.09 3.927 66.11 4.083 ;
      RECT 66.081 3.924 66.09 4.082 ;
      RECT 65.995 3.92 66.081 4.076 ;
      RECT 65.955 3.916 65.995 4.068 ;
      RECT 65.935 3.912 65.955 4.066 ;
      RECT 65.875 3.912 65.935 4.063 ;
      RECT 65.855 3.915 65.875 4.061 ;
      RECT 65.834 3.915 65.855 4.061 ;
      RECT 65.748 3.917 65.834 4.065 ;
      RECT 65.662 3.919 65.748 4.071 ;
      RECT 65.576 3.921 65.662 4.078 ;
      RECT 65.49 3.924 65.576 4.084 ;
      RECT 65.456 3.925 65.49 4.089 ;
      RECT 65.37 3.928 65.456 4.094 ;
      RECT 65.341 3.935 65.37 4.099 ;
      RECT 65.255 3.935 65.341 4.104 ;
      RECT 65.222 3.935 65.255 4.109 ;
      RECT 65.136 3.937 65.222 4.114 ;
      RECT 65.05 3.939 65.136 4.121 ;
      RECT 64.986 3.941 65.05 4.127 ;
      RECT 64.9 3.943 64.986 4.133 ;
      RECT 64.897 3.945 64.9 4.136 ;
      RECT 64.811 3.946 64.897 4.14 ;
      RECT 64.725 3.949 64.811 4.147 ;
      RECT 64.706 3.951 64.725 4.151 ;
      RECT 64.62 3.953 64.706 4.156 ;
      RECT 64.35 3.965 64.36 4.16 ;
      RECT 66.53 10.2 66.82 10.43 ;
      RECT 66.59 9.46 66.76 10.43 ;
      RECT 66.48 9.49 66.855 9.86 ;
      RECT 66.53 9.46 66.82 9.86 ;
      RECT 66.585 3.545 66.77 3.755 ;
      RECT 66.58 3.546 66.775 3.753 ;
      RECT 66.575 3.551 66.785 3.748 ;
      RECT 66.57 3.527 66.575 3.745 ;
      RECT 66.54 3.524 66.57 3.738 ;
      RECT 66.535 3.52 66.54 3.729 ;
      RECT 66.5 3.551 66.785 3.724 ;
      RECT 66.275 3.46 66.535 3.72 ;
      RECT 66.575 3.529 66.58 3.748 ;
      RECT 66.58 3.53 66.585 3.753 ;
      RECT 66.275 3.542 66.655 3.72 ;
      RECT 66.275 3.54 66.64 3.72 ;
      RECT 66.275 3.535 66.63 3.72 ;
      RECT 66.23 4.45 66.28 4.735 ;
      RECT 66.175 4.42 66.18 4.735 ;
      RECT 66.145 4.4 66.15 4.735 ;
      RECT 66.295 4.45 66.355 4.71 ;
      RECT 66.29 4.45 66.295 4.718 ;
      RECT 66.28 4.45 66.29 4.73 ;
      RECT 66.195 4.44 66.23 4.735 ;
      RECT 66.19 4.427 66.195 4.735 ;
      RECT 66.18 4.422 66.19 4.735 ;
      RECT 66.16 4.412 66.175 4.735 ;
      RECT 66.15 4.405 66.16 4.735 ;
      RECT 66.14 4.397 66.145 4.735 ;
      RECT 66.11 4.387 66.14 4.735 ;
      RECT 66.095 4.375 66.11 4.735 ;
      RECT 66.08 4.365 66.095 4.73 ;
      RECT 66.06 4.355 66.08 4.705 ;
      RECT 66.05 4.347 66.06 4.682 ;
      RECT 66.02 4.33 66.05 4.672 ;
      RECT 66.015 4.307 66.02 4.663 ;
      RECT 66.01 4.294 66.015 4.661 ;
      RECT 65.995 4.27 66.01 4.655 ;
      RECT 65.99 4.246 65.995 4.649 ;
      RECT 65.98 4.235 65.99 4.644 ;
      RECT 65.975 4.225 65.98 4.64 ;
      RECT 65.97 4.217 65.975 4.637 ;
      RECT 65.96 4.212 65.97 4.633 ;
      RECT 65.955 4.207 65.96 4.629 ;
      RECT 65.87 4.205 65.955 4.604 ;
      RECT 65.84 4.205 65.87 4.57 ;
      RECT 65.825 4.205 65.84 4.553 ;
      RECT 65.77 4.205 65.825 4.498 ;
      RECT 65.765 4.21 65.77 4.447 ;
      RECT 65.755 4.215 65.765 4.437 ;
      RECT 65.75 4.225 65.755 4.423 ;
      RECT 65.7 4.965 65.96 5.225 ;
      RECT 65.62 4.98 65.96 5.201 ;
      RECT 65.6 4.98 65.96 5.196 ;
      RECT 65.576 4.98 65.96 5.194 ;
      RECT 65.49 4.98 65.96 5.189 ;
      RECT 65.34 4.92 65.6 5.185 ;
      RECT 65.295 4.98 65.96 5.18 ;
      RECT 65.29 4.987 65.96 5.175 ;
      RECT 65.305 4.975 65.62 5.185 ;
      RECT 65.195 3.41 65.455 3.67 ;
      RECT 65.195 3.467 65.46 3.663 ;
      RECT 65.195 3.497 65.465 3.595 ;
      RECT 65.255 3.928 65.37 3.93 ;
      RECT 65.341 3.925 65.37 3.93 ;
      RECT 64.365 4.929 64.39 5.169 ;
      RECT 64.35 4.932 64.44 5.163 ;
      RECT 64.345 4.937 64.526 5.158 ;
      RECT 64.34 4.945 64.59 5.156 ;
      RECT 64.34 4.945 64.6 5.155 ;
      RECT 64.335 4.952 64.61 5.148 ;
      RECT 64.335 4.952 64.696 5.137 ;
      RECT 64.33 4.987 64.696 5.133 ;
      RECT 64.33 4.987 64.705 5.122 ;
      RECT 64.61 4.86 64.87 5.12 ;
      RECT 64.32 5.037 64.87 5.118 ;
      RECT 64.59 4.905 64.61 5.153 ;
      RECT 64.526 4.908 64.59 5.157 ;
      RECT 64.44 4.913 64.526 5.162 ;
      RECT 64.37 4.924 64.87 5.12 ;
      RECT 64.39 4.918 64.44 5.167 ;
      RECT 64.515 3.395 64.525 3.657 ;
      RECT 64.505 3.452 64.515 3.66 ;
      RECT 64.48 3.457 64.505 3.666 ;
      RECT 64.455 3.461 64.48 3.678 ;
      RECT 64.445 3.464 64.455 3.688 ;
      RECT 64.44 3.465 64.445 3.693 ;
      RECT 64.435 3.466 64.44 3.698 ;
      RECT 64.43 3.467 64.435 3.7 ;
      RECT 64.405 3.47 64.43 3.703 ;
      RECT 64.375 3.476 64.405 3.706 ;
      RECT 64.31 3.487 64.375 3.709 ;
      RECT 64.265 3.495 64.31 3.713 ;
      RECT 64.25 3.495 64.265 3.721 ;
      RECT 64.245 3.496 64.25 3.728 ;
      RECT 64.24 3.498 64.245 3.731 ;
      RECT 64.235 3.502 64.24 3.734 ;
      RECT 64.225 3.51 64.235 3.738 ;
      RECT 64.22 3.523 64.225 3.743 ;
      RECT 64.215 3.531 64.22 3.745 ;
      RECT 64.21 3.537 64.215 3.745 ;
      RECT 64.205 3.541 64.21 3.748 ;
      RECT 64.2 3.543 64.205 3.751 ;
      RECT 64.195 3.546 64.2 3.754 ;
      RECT 64.185 3.551 64.195 3.758 ;
      RECT 64.18 3.557 64.185 3.763 ;
      RECT 64.17 3.563 64.18 3.767 ;
      RECT 64.155 3.57 64.17 3.773 ;
      RECT 64.126 3.584 64.155 3.783 ;
      RECT 64.04 3.619 64.126 3.815 ;
      RECT 64.02 3.652 64.04 3.844 ;
      RECT 64 3.665 64.02 3.855 ;
      RECT 63.98 3.677 64 3.866 ;
      RECT 63.93 3.699 63.98 3.886 ;
      RECT 63.915 3.717 63.93 3.903 ;
      RECT 63.91 3.723 63.915 3.906 ;
      RECT 63.905 3.727 63.91 3.909 ;
      RECT 63.9 3.731 63.905 3.913 ;
      RECT 63.895 3.733 63.9 3.916 ;
      RECT 63.885 3.74 63.895 3.919 ;
      RECT 63.88 3.745 63.885 3.923 ;
      RECT 63.875 3.747 63.88 3.926 ;
      RECT 63.87 3.751 63.875 3.929 ;
      RECT 63.865 3.753 63.87 3.933 ;
      RECT 63.85 3.758 63.865 3.938 ;
      RECT 63.845 3.763 63.85 3.941 ;
      RECT 63.84 3.771 63.845 3.944 ;
      RECT 63.835 3.773 63.84 3.947 ;
      RECT 63.83 3.775 63.835 3.95 ;
      RECT 63.82 3.777 63.83 3.956 ;
      RECT 63.785 3.791 63.82 3.968 ;
      RECT 63.775 3.806 63.785 3.978 ;
      RECT 63.7 3.835 63.775 4.002 ;
      RECT 63.695 3.86 63.7 4.025 ;
      RECT 63.68 3.864 63.695 4.031 ;
      RECT 63.67 3.872 63.68 4.036 ;
      RECT 63.64 3.885 63.67 4.04 ;
      RECT 63.63 3.9 63.64 4.045 ;
      RECT 63.62 3.905 63.63 4.048 ;
      RECT 63.615 3.907 63.62 4.05 ;
      RECT 63.6 3.91 63.615 4.053 ;
      RECT 63.595 3.912 63.6 4.056 ;
      RECT 63.575 3.917 63.595 4.06 ;
      RECT 63.545 3.922 63.575 4.068 ;
      RECT 63.52 3.929 63.545 4.076 ;
      RECT 63.515 3.934 63.52 4.081 ;
      RECT 63.485 3.937 63.515 4.085 ;
      RECT 63.445 3.94 63.485 4.095 ;
      RECT 63.41 3.937 63.445 4.107 ;
      RECT 63.4 3.933 63.41 4.114 ;
      RECT 63.375 3.929 63.4 4.12 ;
      RECT 63.37 3.925 63.375 4.125 ;
      RECT 63.33 3.922 63.37 4.125 ;
      RECT 63.315 3.907 63.33 4.126 ;
      RECT 63.292 3.895 63.315 4.126 ;
      RECT 63.206 3.895 63.292 4.127 ;
      RECT 63.12 3.895 63.206 4.129 ;
      RECT 63.1 3.895 63.12 4.126 ;
      RECT 63.095 3.9 63.1 4.121 ;
      RECT 63.09 3.905 63.095 4.119 ;
      RECT 63.08 3.915 63.09 4.117 ;
      RECT 63.075 3.921 63.08 4.11 ;
      RECT 63.07 3.923 63.075 4.095 ;
      RECT 63.065 3.927 63.07 4.085 ;
      RECT 64.525 3.395 64.775 3.655 ;
      RECT 62.25 4.93 62.51 5.19 ;
      RECT 64.545 4.42 64.55 4.63 ;
      RECT 64.55 4.425 64.56 4.625 ;
      RECT 64.5 4.42 64.545 4.645 ;
      RECT 64.49 4.42 64.5 4.665 ;
      RECT 64.471 4.42 64.49 4.67 ;
      RECT 64.385 4.42 64.471 4.667 ;
      RECT 64.355 4.422 64.385 4.665 ;
      RECT 64.3 4.432 64.355 4.663 ;
      RECT 64.235 4.446 64.3 4.661 ;
      RECT 64.23 4.454 64.235 4.66 ;
      RECT 64.215 4.457 64.23 4.658 ;
      RECT 64.15 4.467 64.215 4.654 ;
      RECT 64.102 4.481 64.15 4.655 ;
      RECT 64.016 4.498 64.102 4.669 ;
      RECT 63.93 4.519 64.016 4.686 ;
      RECT 63.91 4.532 63.93 4.696 ;
      RECT 63.865 4.54 63.91 4.703 ;
      RECT 63.83 4.548 63.865 4.711 ;
      RECT 63.796 4.556 63.83 4.719 ;
      RECT 63.71 4.57 63.796 4.731 ;
      RECT 63.675 4.587 63.71 4.743 ;
      RECT 63.666 4.596 63.675 4.747 ;
      RECT 63.58 4.614 63.666 4.764 ;
      RECT 63.521 4.641 63.58 4.791 ;
      RECT 63.435 4.668 63.521 4.819 ;
      RECT 63.415 4.69 63.435 4.839 ;
      RECT 63.355 4.705 63.415 4.855 ;
      RECT 63.345 4.717 63.355 4.868 ;
      RECT 63.34 4.722 63.345 4.871 ;
      RECT 63.33 4.725 63.34 4.874 ;
      RECT 63.325 4.727 63.33 4.877 ;
      RECT 63.295 4.735 63.325 4.884 ;
      RECT 63.28 4.742 63.295 4.892 ;
      RECT 63.27 4.747 63.28 4.896 ;
      RECT 63.265 4.75 63.27 4.899 ;
      RECT 63.255 4.752 63.265 4.902 ;
      RECT 63.22 4.762 63.255 4.911 ;
      RECT 63.145 4.785 63.22 4.933 ;
      RECT 63.125 4.803 63.145 4.951 ;
      RECT 63.095 4.81 63.125 4.961 ;
      RECT 63.075 4.818 63.095 4.971 ;
      RECT 63.065 4.824 63.075 4.978 ;
      RECT 63.046 4.829 63.065 4.984 ;
      RECT 62.96 4.849 63.046 5.004 ;
      RECT 62.945 4.869 62.96 5.023 ;
      RECT 62.9 4.881 62.945 5.034 ;
      RECT 62.835 4.902 62.9 5.057 ;
      RECT 62.795 4.922 62.835 5.078 ;
      RECT 62.785 4.932 62.795 5.088 ;
      RECT 62.735 4.944 62.785 5.099 ;
      RECT 62.715 4.96 62.735 5.111 ;
      RECT 62.685 4.97 62.715 5.117 ;
      RECT 62.675 4.975 62.685 5.119 ;
      RECT 62.606 4.976 62.675 5.125 ;
      RECT 62.52 4.978 62.606 5.135 ;
      RECT 62.51 4.979 62.52 5.14 ;
      RECT 63.78 5.005 63.97 5.215 ;
      RECT 63.77 5.01 63.98 5.208 ;
      RECT 63.755 5.01 63.98 5.173 ;
      RECT 63.675 4.895 63.935 5.155 ;
      RECT 62.59 4.425 62.775 4.72 ;
      RECT 62.58 4.425 62.775 4.718 ;
      RECT 62.565 4.425 62.78 4.713 ;
      RECT 62.565 4.425 62.785 4.71 ;
      RECT 62.56 4.425 62.785 4.708 ;
      RECT 62.555 4.68 62.785 4.698 ;
      RECT 62.56 4.425 62.82 4.685 ;
      RECT 62.52 3.46 62.78 3.72 ;
      RECT 62.33 3.385 62.416 3.718 ;
      RECT 62.305 3.389 62.46 3.714 ;
      RECT 62.416 3.381 62.46 3.714 ;
      RECT 62.416 3.382 62.465 3.713 ;
      RECT 62.33 3.387 62.48 3.712 ;
      RECT 62.305 3.395 62.52 3.711 ;
      RECT 62.3 3.39 62.48 3.706 ;
      RECT 62.29 3.405 62.52 3.613 ;
      RECT 62.29 3.457 62.72 3.613 ;
      RECT 62.29 3.45 62.7 3.613 ;
      RECT 62.29 3.437 62.67 3.613 ;
      RECT 62.29 3.425 62.61 3.613 ;
      RECT 62.29 3.41 62.585 3.613 ;
      RECT 61.49 4.04 61.625 4.335 ;
      RECT 61.75 4.063 61.755 4.25 ;
      RECT 62.47 3.96 62.615 4.195 ;
      RECT 62.63 3.96 62.635 4.185 ;
      RECT 62.665 3.971 62.67 4.165 ;
      RECT 62.66 3.963 62.665 4.17 ;
      RECT 62.64 3.96 62.66 4.175 ;
      RECT 62.635 3.96 62.64 4.183 ;
      RECT 62.625 3.96 62.63 4.188 ;
      RECT 62.615 3.96 62.625 4.193 ;
      RECT 62.445 3.962 62.47 4.195 ;
      RECT 62.395 3.969 62.445 4.195 ;
      RECT 62.39 3.974 62.395 4.195 ;
      RECT 62.351 3.979 62.39 4.196 ;
      RECT 62.265 3.991 62.351 4.197 ;
      RECT 62.256 4.001 62.265 4.197 ;
      RECT 62.17 4.01 62.256 4.199 ;
      RECT 62.146 4.02 62.17 4.201 ;
      RECT 62.06 4.031 62.146 4.202 ;
      RECT 62.03 4.042 62.06 4.204 ;
      RECT 62 4.047 62.03 4.206 ;
      RECT 61.975 4.053 62 4.209 ;
      RECT 61.96 4.058 61.975 4.21 ;
      RECT 61.915 4.064 61.96 4.21 ;
      RECT 61.91 4.069 61.915 4.211 ;
      RECT 61.89 4.069 61.91 4.213 ;
      RECT 61.87 4.067 61.89 4.218 ;
      RECT 61.835 4.066 61.87 4.225 ;
      RECT 61.805 4.065 61.835 4.235 ;
      RECT 61.755 4.064 61.805 4.245 ;
      RECT 61.665 4.061 61.75 4.335 ;
      RECT 61.64 4.055 61.665 4.335 ;
      RECT 61.625 4.045 61.64 4.335 ;
      RECT 61.44 4.04 61.49 4.255 ;
      RECT 61.43 4.045 61.44 4.245 ;
      RECT 61.67 4.52 61.93 4.78 ;
      RECT 61.67 4.52 61.96 4.673 ;
      RECT 61.67 4.52 61.995 4.658 ;
      RECT 61.925 4.44 62.115 4.65 ;
      RECT 61.915 4.445 62.125 4.643 ;
      RECT 61.88 4.515 62.125 4.643 ;
      RECT 61.91 4.457 61.93 4.78 ;
      RECT 61.895 4.505 62.125 4.643 ;
      RECT 61.9 4.477 61.93 4.78 ;
      RECT 60.98 3.545 61.05 4.65 ;
      RECT 61.715 3.65 61.975 3.91 ;
      RECT 61.295 3.696 61.31 3.905 ;
      RECT 61.631 3.709 61.715 3.86 ;
      RECT 61.545 3.706 61.631 3.86 ;
      RECT 61.506 3.704 61.545 3.86 ;
      RECT 61.42 3.702 61.506 3.86 ;
      RECT 61.36 3.7 61.42 3.871 ;
      RECT 61.325 3.698 61.36 3.889 ;
      RECT 61.31 3.696 61.325 3.9 ;
      RECT 61.28 3.696 61.295 3.913 ;
      RECT 61.27 3.696 61.28 3.918 ;
      RECT 61.245 3.695 61.27 3.923 ;
      RECT 61.23 3.69 61.245 3.929 ;
      RECT 61.225 3.683 61.23 3.934 ;
      RECT 61.2 3.674 61.225 3.94 ;
      RECT 61.155 3.653 61.2 3.953 ;
      RECT 61.145 3.637 61.155 3.963 ;
      RECT 61.13 3.63 61.145 3.973 ;
      RECT 61.12 3.623 61.13 3.99 ;
      RECT 61.115 3.62 61.12 4.02 ;
      RECT 61.11 3.618 61.115 4.05 ;
      RECT 61.105 3.616 61.11 4.087 ;
      RECT 61.09 3.612 61.105 4.154 ;
      RECT 61.09 4.445 61.1 4.645 ;
      RECT 61.085 3.608 61.09 4.28 ;
      RECT 61.085 4.432 61.09 4.65 ;
      RECT 61.08 3.606 61.085 4.365 ;
      RECT 61.08 4.422 61.085 4.65 ;
      RECT 61.065 3.577 61.08 4.65 ;
      RECT 61.05 3.55 61.065 4.65 ;
      RECT 60.975 3.545 60.98 3.9 ;
      RECT 60.975 3.955 60.98 4.65 ;
      RECT 60.96 3.545 60.975 3.878 ;
      RECT 60.97 3.977 60.975 4.65 ;
      RECT 60.96 4.017 60.97 4.65 ;
      RECT 60.925 3.545 60.96 3.82 ;
      RECT 60.955 4.052 60.96 4.65 ;
      RECT 60.94 4.107 60.955 4.65 ;
      RECT 60.935 4.172 60.94 4.65 ;
      RECT 60.92 4.22 60.935 4.65 ;
      RECT 60.895 3.545 60.925 3.775 ;
      RECT 60.915 4.275 60.92 4.65 ;
      RECT 60.9 4.335 60.915 4.65 ;
      RECT 60.895 4.383 60.9 4.648 ;
      RECT 60.89 3.545 60.895 3.768 ;
      RECT 60.89 4.415 60.895 4.643 ;
      RECT 60.865 3.545 60.89 3.76 ;
      RECT 60.855 3.55 60.865 3.75 ;
      RECT 61.07 4.825 61.09 5.065 ;
      RECT 60.3 4.755 60.305 4.965 ;
      RECT 61.58 4.828 61.59 5.023 ;
      RECT 61.575 4.818 61.58 5.026 ;
      RECT 61.495 4.815 61.575 5.049 ;
      RECT 61.491 4.815 61.495 5.071 ;
      RECT 61.405 4.815 61.491 5.081 ;
      RECT 61.39 4.815 61.405 5.089 ;
      RECT 61.361 4.816 61.39 5.087 ;
      RECT 61.275 4.821 61.361 5.083 ;
      RECT 61.262 4.825 61.275 5.079 ;
      RECT 61.176 4.825 61.262 5.075 ;
      RECT 61.09 4.825 61.176 5.069 ;
      RECT 61.006 4.825 61.07 5.063 ;
      RECT 60.92 4.825 61.006 5.058 ;
      RECT 60.9 4.825 60.92 5.054 ;
      RECT 60.84 4.82 60.9 5.051 ;
      RECT 60.812 4.814 60.84 5.048 ;
      RECT 60.726 4.809 60.812 5.044 ;
      RECT 60.64 4.803 60.726 5.038 ;
      RECT 60.565 4.785 60.64 5.033 ;
      RECT 60.53 4.762 60.565 5.029 ;
      RECT 60.52 4.752 60.53 5.028 ;
      RECT 60.465 4.75 60.52 5.027 ;
      RECT 60.39 4.75 60.465 5.023 ;
      RECT 60.38 4.75 60.39 5.018 ;
      RECT 60.365 4.75 60.38 5.01 ;
      RECT 60.315 4.752 60.365 4.988 ;
      RECT 60.305 4.755 60.315 4.968 ;
      RECT 60.295 4.76 60.3 4.963 ;
      RECT 60.29 4.765 60.295 4.958 ;
      RECT 60.415 3.93 60.675 4.19 ;
      RECT 60.415 3.945 60.695 4.155 ;
      RECT 60.415 3.95 60.705 4.15 ;
      RECT 58.4 3.41 58.66 3.67 ;
      RECT 58.39 3.44 58.66 3.65 ;
      RECT 60.31 3.355 60.57 3.615 ;
      RECT 60.305 3.43 60.31 3.616 ;
      RECT 60.28 3.435 60.305 3.618 ;
      RECT 60.265 3.442 60.28 3.621 ;
      RECT 60.205 3.46 60.265 3.626 ;
      RECT 60.175 3.48 60.205 3.633 ;
      RECT 60.15 3.488 60.175 3.638 ;
      RECT 60.125 3.496 60.15 3.64 ;
      RECT 60.107 3.5 60.125 3.639 ;
      RECT 60.021 3.498 60.107 3.639 ;
      RECT 59.935 3.496 60.021 3.639 ;
      RECT 59.849 3.494 59.935 3.638 ;
      RECT 59.763 3.492 59.849 3.638 ;
      RECT 59.677 3.49 59.763 3.638 ;
      RECT 59.591 3.488 59.677 3.638 ;
      RECT 59.505 3.486 59.591 3.637 ;
      RECT 59.487 3.485 59.505 3.637 ;
      RECT 59.401 3.484 59.487 3.637 ;
      RECT 59.315 3.482 59.401 3.637 ;
      RECT 59.229 3.481 59.315 3.636 ;
      RECT 59.143 3.48 59.229 3.636 ;
      RECT 59.057 3.478 59.143 3.636 ;
      RECT 58.971 3.477 59.057 3.636 ;
      RECT 58.885 3.475 58.971 3.635 ;
      RECT 58.861 3.473 58.885 3.635 ;
      RECT 58.775 3.466 58.861 3.635 ;
      RECT 58.746 3.458 58.775 3.635 ;
      RECT 58.66 3.45 58.746 3.635 ;
      RECT 58.38 3.447 58.39 3.645 ;
      RECT 59.885 4.41 59.89 4.76 ;
      RECT 59.655 4.5 59.795 4.76 ;
      RECT 60.13 4.185 60.175 4.395 ;
      RECT 60.185 4.196 60.195 4.39 ;
      RECT 60.175 4.188 60.185 4.395 ;
      RECT 60.11 4.185 60.13 4.4 ;
      RECT 60.08 4.185 60.11 4.423 ;
      RECT 60.07 4.185 60.08 4.448 ;
      RECT 60.065 4.185 60.07 4.458 ;
      RECT 60.01 4.185 60.065 4.498 ;
      RECT 60.005 4.185 60.01 4.538 ;
      RECT 60 4.187 60.005 4.543 ;
      RECT 59.985 4.197 60 4.554 ;
      RECT 59.94 4.255 59.985 4.59 ;
      RECT 59.93 4.31 59.94 4.624 ;
      RECT 59.915 4.337 59.93 4.64 ;
      RECT 59.905 4.364 59.915 4.76 ;
      RECT 59.89 4.387 59.905 4.76 ;
      RECT 59.88 4.427 59.885 4.76 ;
      RECT 59.875 4.437 59.88 4.76 ;
      RECT 59.87 4.452 59.875 4.76 ;
      RECT 59.86 4.457 59.87 4.76 ;
      RECT 59.795 4.48 59.86 4.76 ;
      RECT 59.295 3.975 59.485 4.185 ;
      RECT 57.87 3.9 58.13 4.16 ;
      RECT 58.22 3.895 58.315 4.105 ;
      RECT 58.195 3.91 58.205 4.105 ;
      RECT 59.485 3.982 59.495 4.18 ;
      RECT 59.285 3.982 59.295 4.18 ;
      RECT 59.27 3.997 59.285 4.17 ;
      RECT 59.265 4.005 59.27 4.163 ;
      RECT 59.255 4.008 59.265 4.16 ;
      RECT 59.22 4.007 59.255 4.158 ;
      RECT 59.191 4.003 59.22 4.155 ;
      RECT 59.105 3.998 59.191 4.152 ;
      RECT 59.045 3.992 59.105 4.148 ;
      RECT 59.016 3.988 59.045 4.145 ;
      RECT 58.93 3.98 59.016 4.142 ;
      RECT 58.921 3.974 58.93 4.14 ;
      RECT 58.835 3.969 58.921 4.138 ;
      RECT 58.812 3.964 58.835 4.135 ;
      RECT 58.726 3.958 58.812 4.132 ;
      RECT 58.64 3.949 58.726 4.127 ;
      RECT 58.63 3.944 58.64 4.125 ;
      RECT 58.611 3.943 58.63 4.124 ;
      RECT 58.525 3.938 58.611 4.12 ;
      RECT 58.505 3.933 58.525 4.116 ;
      RECT 58.445 3.928 58.505 4.113 ;
      RECT 58.42 3.918 58.445 4.111 ;
      RECT 58.415 3.911 58.42 4.11 ;
      RECT 58.405 3.902 58.415 4.109 ;
      RECT 58.401 3.895 58.405 4.109 ;
      RECT 58.315 3.895 58.401 4.107 ;
      RECT 58.205 3.902 58.22 4.105 ;
      RECT 58.19 3.912 58.195 4.105 ;
      RECT 58.17 3.915 58.19 4.102 ;
      RECT 58.14 3.915 58.17 4.098 ;
      RECT 58.13 3.915 58.14 4.098 ;
      RECT 59.045 4.41 59.305 4.67 ;
      RECT 58.975 4.42 59.305 4.63 ;
      RECT 58.965 4.427 59.305 4.625 ;
      RECT 58.385 4.415 58.645 4.675 ;
      RECT 58.385 4.455 58.75 4.665 ;
      RECT 58.385 4.457 58.755 4.664 ;
      RECT 58.385 4.465 58.76 4.661 ;
      RECT 57.31 3.54 57.41 5.065 ;
      RECT 57.5 4.68 57.55 4.94 ;
      RECT 57.495 3.553 57.5 3.74 ;
      RECT 57.49 4.661 57.5 4.94 ;
      RECT 57.49 3.55 57.495 3.748 ;
      RECT 57.475 3.544 57.49 3.755 ;
      RECT 57.485 4.649 57.49 5.023 ;
      RECT 57.475 4.637 57.485 5.06 ;
      RECT 57.465 3.54 57.475 3.762 ;
      RECT 57.465 4.622 57.475 5.065 ;
      RECT 57.46 3.54 57.465 3.77 ;
      RECT 57.44 4.592 57.465 5.065 ;
      RECT 57.42 3.54 57.46 3.818 ;
      RECT 57.43 4.552 57.44 5.065 ;
      RECT 57.42 4.507 57.43 5.065 ;
      RECT 57.415 3.54 57.42 3.888 ;
      RECT 57.415 4.465 57.42 5.065 ;
      RECT 57.41 3.54 57.415 4.365 ;
      RECT 57.41 4.447 57.415 5.065 ;
      RECT 57.3 3.543 57.31 5.065 ;
      RECT 57.285 3.55 57.3 5.061 ;
      RECT 57.28 3.56 57.285 5.056 ;
      RECT 57.275 3.76 57.28 4.948 ;
      RECT 57.27 3.845 57.275 4.5 ;
      RECT 56.145 10.205 56.435 10.435 ;
      RECT 56.205 8.725 56.375 10.435 ;
      RECT 56.155 9.09 56.505 9.44 ;
      RECT 56.145 8.725 56.435 8.955 ;
      RECT 55.74 3.69 55.845 4.26 ;
      RECT 55.74 4.025 56.065 4.255 ;
      RECT 55.74 4.055 56.235 4.225 ;
      RECT 55.74 3.69 55.93 4.255 ;
      RECT 55.155 3.655 55.445 3.885 ;
      RECT 55.155 3.69 55.93 3.86 ;
      RECT 55.215 2.175 55.385 3.885 ;
      RECT 55.155 2.175 55.445 2.405 ;
      RECT 55.155 10.205 55.445 10.435 ;
      RECT 55.215 8.725 55.385 10.435 ;
      RECT 55.155 8.725 55.445 8.955 ;
      RECT 55.155 8.76 56.01 8.92 ;
      RECT 55.84 8.355 56.01 8.92 ;
      RECT 55.155 8.755 55.55 8.92 ;
      RECT 55.775 8.355 56.065 8.585 ;
      RECT 55.775 8.385 56.235 8.555 ;
      RECT 54.785 4.025 55.075 4.255 ;
      RECT 54.785 4.055 55.245 4.225 ;
      RECT 54.85 2.95 55.015 4.255 ;
      RECT 53.365 2.92 53.655 3.15 ;
      RECT 53.365 2.95 55.015 3.12 ;
      RECT 53.425 2.18 53.595 3.15 ;
      RECT 53.365 2.18 53.655 2.41 ;
      RECT 53.365 10.2 53.655 10.43 ;
      RECT 53.425 9.46 53.595 10.43 ;
      RECT 53.425 9.555 55.015 9.725 ;
      RECT 54.845 8.355 55.015 9.725 ;
      RECT 53.365 9.46 53.655 9.69 ;
      RECT 54.785 8.355 55.075 8.585 ;
      RECT 54.785 8.385 55.245 8.555 ;
      RECT 51.4 4.725 51.75 5.075 ;
      RECT 51.49 3.32 51.66 5.075 ;
      RECT 53.795 3.26 54.145 3.61 ;
      RECT 51.49 3.32 53.11 3.495 ;
      RECT 51.49 3.32 54.145 3.49 ;
      RECT 53.82 9.09 54.145 9.415 ;
      RECT 49.25 9.05 49.6 9.4 ;
      RECT 53.795 9.09 54.145 9.32 ;
      RECT 49.035 9.09 49.6 9.32 ;
      RECT 48.865 9.12 54.145 9.29 ;
      RECT 53.02 3.66 53.34 3.98 ;
      RECT 52.99 3.66 53.34 3.89 ;
      RECT 52.82 3.69 53.34 3.86 ;
      RECT 53.02 8.66 53.34 8.98 ;
      RECT 52.99 8.72 53.34 8.95 ;
      RECT 52.82 8.75 53.34 8.92 ;
      RECT 48.8 4.96 48.84 5.22 ;
      RECT 48.84 4.94 48.845 4.95 ;
      RECT 50.17 4.185 50.18 4.406 ;
      RECT 50.1 4.18 50.17 4.531 ;
      RECT 50.09 4.18 50.1 4.658 ;
      RECT 50.065 4.18 50.09 4.705 ;
      RECT 50.04 4.18 50.065 4.783 ;
      RECT 50.02 4.18 50.04 4.853 ;
      RECT 49.995 4.18 50.02 4.893 ;
      RECT 49.985 4.18 49.995 4.913 ;
      RECT 49.975 4.182 49.985 4.921 ;
      RECT 49.97 4.187 49.975 4.378 ;
      RECT 49.97 4.387 49.975 4.922 ;
      RECT 49.965 4.432 49.97 4.923 ;
      RECT 49.955 4.497 49.965 4.924 ;
      RECT 49.945 4.592 49.955 4.926 ;
      RECT 49.94 4.645 49.945 4.928 ;
      RECT 49.935 4.665 49.94 4.929 ;
      RECT 49.88 4.69 49.935 4.935 ;
      RECT 49.84 4.725 49.88 4.944 ;
      RECT 49.83 4.742 49.84 4.949 ;
      RECT 49.821 4.748 49.83 4.951 ;
      RECT 49.735 4.786 49.821 4.962 ;
      RECT 49.73 4.825 49.735 4.972 ;
      RECT 49.655 4.832 49.73 4.982 ;
      RECT 49.635 4.842 49.655 4.993 ;
      RECT 49.605 4.849 49.635 5.001 ;
      RECT 49.58 4.856 49.605 5.008 ;
      RECT 49.556 4.862 49.58 5.013 ;
      RECT 49.47 4.875 49.556 5.025 ;
      RECT 49.392 4.882 49.47 5.043 ;
      RECT 49.306 4.877 49.392 5.061 ;
      RECT 49.22 4.872 49.306 5.081 ;
      RECT 49.14 4.866 49.22 5.098 ;
      RECT 49.075 4.862 49.14 5.127 ;
      RECT 49.07 4.576 49.075 4.6 ;
      RECT 49.06 4.852 49.075 5.155 ;
      RECT 49.065 4.57 49.07 4.64 ;
      RECT 49.06 4.564 49.065 4.71 ;
      RECT 49.055 4.558 49.06 4.788 ;
      RECT 49.055 4.835 49.06 5.22 ;
      RECT 49.047 4.555 49.055 5.22 ;
      RECT 48.961 4.553 49.047 5.22 ;
      RECT 48.875 4.551 48.961 5.22 ;
      RECT 48.865 4.552 48.875 5.22 ;
      RECT 48.86 4.557 48.865 5.22 ;
      RECT 48.85 4.57 48.86 5.22 ;
      RECT 48.845 4.592 48.85 5.22 ;
      RECT 48.84 4.952 48.845 5.22 ;
      RECT 49.47 4.42 49.475 4.64 ;
      RECT 49.975 3.455 50.01 3.715 ;
      RECT 49.96 3.455 49.975 3.723 ;
      RECT 49.931 3.455 49.96 3.745 ;
      RECT 49.845 3.455 49.931 3.805 ;
      RECT 49.825 3.455 49.845 3.87 ;
      RECT 49.765 3.455 49.825 4.035 ;
      RECT 49.76 3.455 49.765 4.183 ;
      RECT 49.755 3.455 49.76 4.195 ;
      RECT 49.75 3.455 49.755 4.221 ;
      RECT 49.72 3.641 49.75 4.301 ;
      RECT 49.715 3.689 49.72 4.39 ;
      RECT 49.71 3.703 49.715 4.405 ;
      RECT 49.705 3.722 49.71 4.435 ;
      RECT 49.7 3.737 49.705 4.451 ;
      RECT 49.695 3.752 49.7 4.473 ;
      RECT 49.69 3.772 49.695 4.495 ;
      RECT 49.68 3.792 49.69 4.528 ;
      RECT 49.665 3.834 49.68 4.59 ;
      RECT 49.66 3.865 49.665 4.63 ;
      RECT 49.655 3.877 49.66 4.635 ;
      RECT 49.65 3.889 49.655 4.64 ;
      RECT 49.645 3.902 49.65 4.64 ;
      RECT 49.64 3.92 49.645 4.64 ;
      RECT 49.635 3.94 49.64 4.64 ;
      RECT 49.63 3.952 49.635 4.64 ;
      RECT 49.625 3.965 49.63 4.64 ;
      RECT 49.605 4 49.625 4.64 ;
      RECT 49.555 4.102 49.605 4.64 ;
      RECT 49.55 4.187 49.555 4.64 ;
      RECT 49.545 4.195 49.55 4.64 ;
      RECT 49.54 4.212 49.545 4.64 ;
      RECT 49.535 4.227 49.54 4.64 ;
      RECT 49.5 4.292 49.535 4.64 ;
      RECT 49.485 4.357 49.5 4.64 ;
      RECT 49.48 4.387 49.485 4.64 ;
      RECT 49.475 4.412 49.48 4.64 ;
      RECT 49.46 4.422 49.47 4.64 ;
      RECT 49.445 4.435 49.46 4.633 ;
      RECT 49.19 4.025 49.26 4.235 ;
      RECT 48.98 4.002 48.985 4.195 ;
      RECT 46.435 3.93 46.695 4.19 ;
      RECT 49.27 4.212 49.275 4.215 ;
      RECT 49.26 4.03 49.27 4.23 ;
      RECT 49.161 4.023 49.19 4.235 ;
      RECT 49.075 4.015 49.161 4.235 ;
      RECT 49.06 4.009 49.075 4.233 ;
      RECT 49.04 4.008 49.06 4.22 ;
      RECT 49.035 4.007 49.04 4.203 ;
      RECT 48.985 4.004 49.035 4.198 ;
      RECT 48.955 4.001 48.98 4.193 ;
      RECT 48.935 3.999 48.955 4.188 ;
      RECT 48.92 3.997 48.935 4.185 ;
      RECT 48.89 3.995 48.92 4.183 ;
      RECT 48.825 3.991 48.89 4.175 ;
      RECT 48.795 3.986 48.825 4.17 ;
      RECT 48.775 3.984 48.795 4.168 ;
      RECT 48.745 3.981 48.775 4.163 ;
      RECT 48.685 3.977 48.745 4.155 ;
      RECT 48.68 3.974 48.685 4.15 ;
      RECT 48.61 3.972 48.68 4.145 ;
      RECT 48.581 3.968 48.61 4.138 ;
      RECT 48.495 3.963 48.581 4.13 ;
      RECT 48.461 3.958 48.495 4.122 ;
      RECT 48.375 3.95 48.461 4.114 ;
      RECT 48.336 3.943 48.375 4.106 ;
      RECT 48.25 3.938 48.336 4.098 ;
      RECT 48.185 3.932 48.25 4.088 ;
      RECT 48.165 3.927 48.185 4.083 ;
      RECT 48.156 3.924 48.165 4.082 ;
      RECT 48.07 3.92 48.156 4.076 ;
      RECT 48.03 3.916 48.07 4.068 ;
      RECT 48.01 3.912 48.03 4.066 ;
      RECT 47.95 3.912 48.01 4.063 ;
      RECT 47.93 3.915 47.95 4.061 ;
      RECT 47.909 3.915 47.93 4.061 ;
      RECT 47.823 3.917 47.909 4.065 ;
      RECT 47.737 3.919 47.823 4.071 ;
      RECT 47.651 3.921 47.737 4.078 ;
      RECT 47.565 3.924 47.651 4.084 ;
      RECT 47.531 3.925 47.565 4.089 ;
      RECT 47.445 3.928 47.531 4.094 ;
      RECT 47.416 3.935 47.445 4.099 ;
      RECT 47.33 3.935 47.416 4.104 ;
      RECT 47.297 3.935 47.33 4.109 ;
      RECT 47.211 3.937 47.297 4.114 ;
      RECT 47.125 3.939 47.211 4.121 ;
      RECT 47.061 3.941 47.125 4.127 ;
      RECT 46.975 3.943 47.061 4.133 ;
      RECT 46.972 3.945 46.975 4.136 ;
      RECT 46.886 3.946 46.972 4.14 ;
      RECT 46.8 3.949 46.886 4.147 ;
      RECT 46.781 3.951 46.8 4.151 ;
      RECT 46.695 3.953 46.781 4.156 ;
      RECT 46.425 3.965 46.435 4.16 ;
      RECT 48.605 10.2 48.895 10.43 ;
      RECT 48.665 9.46 48.835 10.43 ;
      RECT 48.555 9.49 48.93 9.86 ;
      RECT 48.605 9.46 48.895 9.86 ;
      RECT 48.66 3.545 48.845 3.755 ;
      RECT 48.655 3.546 48.85 3.753 ;
      RECT 48.65 3.551 48.86 3.748 ;
      RECT 48.645 3.527 48.65 3.745 ;
      RECT 48.615 3.524 48.645 3.738 ;
      RECT 48.61 3.52 48.615 3.729 ;
      RECT 48.575 3.551 48.86 3.724 ;
      RECT 48.35 3.46 48.61 3.72 ;
      RECT 48.65 3.529 48.655 3.748 ;
      RECT 48.655 3.53 48.66 3.753 ;
      RECT 48.35 3.542 48.73 3.72 ;
      RECT 48.35 3.54 48.715 3.72 ;
      RECT 48.35 3.535 48.705 3.72 ;
      RECT 48.305 4.45 48.355 4.735 ;
      RECT 48.25 4.42 48.255 4.735 ;
      RECT 48.22 4.4 48.225 4.735 ;
      RECT 48.37 4.45 48.43 4.71 ;
      RECT 48.365 4.45 48.37 4.718 ;
      RECT 48.355 4.45 48.365 4.73 ;
      RECT 48.27 4.44 48.305 4.735 ;
      RECT 48.265 4.427 48.27 4.735 ;
      RECT 48.255 4.422 48.265 4.735 ;
      RECT 48.235 4.412 48.25 4.735 ;
      RECT 48.225 4.405 48.235 4.735 ;
      RECT 48.215 4.397 48.22 4.735 ;
      RECT 48.185 4.387 48.215 4.735 ;
      RECT 48.17 4.375 48.185 4.735 ;
      RECT 48.155 4.365 48.17 4.73 ;
      RECT 48.135 4.355 48.155 4.705 ;
      RECT 48.125 4.347 48.135 4.682 ;
      RECT 48.095 4.33 48.125 4.672 ;
      RECT 48.09 4.307 48.095 4.663 ;
      RECT 48.085 4.294 48.09 4.661 ;
      RECT 48.07 4.27 48.085 4.655 ;
      RECT 48.065 4.246 48.07 4.649 ;
      RECT 48.055 4.235 48.065 4.644 ;
      RECT 48.05 4.225 48.055 4.64 ;
      RECT 48.045 4.217 48.05 4.637 ;
      RECT 48.035 4.212 48.045 4.633 ;
      RECT 48.03 4.207 48.035 4.629 ;
      RECT 47.945 4.205 48.03 4.604 ;
      RECT 47.915 4.205 47.945 4.57 ;
      RECT 47.9 4.205 47.915 4.553 ;
      RECT 47.845 4.205 47.9 4.498 ;
      RECT 47.84 4.21 47.845 4.447 ;
      RECT 47.83 4.215 47.84 4.437 ;
      RECT 47.825 4.225 47.83 4.423 ;
      RECT 47.775 4.965 48.035 5.225 ;
      RECT 47.695 4.98 48.035 5.201 ;
      RECT 47.675 4.98 48.035 5.196 ;
      RECT 47.651 4.98 48.035 5.194 ;
      RECT 47.565 4.98 48.035 5.189 ;
      RECT 47.415 4.92 47.675 5.185 ;
      RECT 47.37 4.98 48.035 5.18 ;
      RECT 47.365 4.987 48.035 5.175 ;
      RECT 47.38 4.975 47.695 5.185 ;
      RECT 47.27 3.41 47.53 3.67 ;
      RECT 47.27 3.467 47.535 3.663 ;
      RECT 47.27 3.497 47.54 3.595 ;
      RECT 47.33 3.928 47.445 3.93 ;
      RECT 47.416 3.925 47.445 3.93 ;
      RECT 46.44 4.929 46.465 5.169 ;
      RECT 46.425 4.932 46.515 5.163 ;
      RECT 46.42 4.937 46.601 5.158 ;
      RECT 46.415 4.945 46.665 5.156 ;
      RECT 46.415 4.945 46.675 5.155 ;
      RECT 46.41 4.952 46.685 5.148 ;
      RECT 46.41 4.952 46.771 5.137 ;
      RECT 46.405 4.987 46.771 5.133 ;
      RECT 46.405 4.987 46.78 5.122 ;
      RECT 46.685 4.86 46.945 5.12 ;
      RECT 46.395 5.037 46.945 5.118 ;
      RECT 46.665 4.905 46.685 5.153 ;
      RECT 46.601 4.908 46.665 5.157 ;
      RECT 46.515 4.913 46.601 5.162 ;
      RECT 46.445 4.924 46.945 5.12 ;
      RECT 46.465 4.918 46.515 5.167 ;
      RECT 46.59 3.395 46.6 3.657 ;
      RECT 46.58 3.452 46.59 3.66 ;
      RECT 46.555 3.457 46.58 3.666 ;
      RECT 46.53 3.461 46.555 3.678 ;
      RECT 46.52 3.464 46.53 3.688 ;
      RECT 46.515 3.465 46.52 3.693 ;
      RECT 46.51 3.466 46.515 3.698 ;
      RECT 46.505 3.467 46.51 3.7 ;
      RECT 46.48 3.47 46.505 3.703 ;
      RECT 46.45 3.476 46.48 3.706 ;
      RECT 46.385 3.487 46.45 3.709 ;
      RECT 46.34 3.495 46.385 3.713 ;
      RECT 46.325 3.495 46.34 3.721 ;
      RECT 46.32 3.496 46.325 3.728 ;
      RECT 46.315 3.498 46.32 3.731 ;
      RECT 46.31 3.502 46.315 3.734 ;
      RECT 46.3 3.51 46.31 3.738 ;
      RECT 46.295 3.523 46.3 3.743 ;
      RECT 46.29 3.531 46.295 3.745 ;
      RECT 46.285 3.537 46.29 3.745 ;
      RECT 46.28 3.541 46.285 3.748 ;
      RECT 46.275 3.543 46.28 3.751 ;
      RECT 46.27 3.546 46.275 3.754 ;
      RECT 46.26 3.551 46.27 3.758 ;
      RECT 46.255 3.557 46.26 3.763 ;
      RECT 46.245 3.563 46.255 3.767 ;
      RECT 46.23 3.57 46.245 3.773 ;
      RECT 46.201 3.584 46.23 3.783 ;
      RECT 46.115 3.619 46.201 3.815 ;
      RECT 46.095 3.652 46.115 3.844 ;
      RECT 46.075 3.665 46.095 3.855 ;
      RECT 46.055 3.677 46.075 3.866 ;
      RECT 46.005 3.699 46.055 3.886 ;
      RECT 45.99 3.717 46.005 3.903 ;
      RECT 45.985 3.723 45.99 3.906 ;
      RECT 45.98 3.727 45.985 3.909 ;
      RECT 45.975 3.731 45.98 3.913 ;
      RECT 45.97 3.733 45.975 3.916 ;
      RECT 45.96 3.74 45.97 3.919 ;
      RECT 45.955 3.745 45.96 3.923 ;
      RECT 45.95 3.747 45.955 3.926 ;
      RECT 45.945 3.751 45.95 3.929 ;
      RECT 45.94 3.753 45.945 3.933 ;
      RECT 45.925 3.758 45.94 3.938 ;
      RECT 45.92 3.763 45.925 3.941 ;
      RECT 45.915 3.771 45.92 3.944 ;
      RECT 45.91 3.773 45.915 3.947 ;
      RECT 45.905 3.775 45.91 3.95 ;
      RECT 45.895 3.777 45.905 3.956 ;
      RECT 45.86 3.791 45.895 3.968 ;
      RECT 45.85 3.806 45.86 3.978 ;
      RECT 45.775 3.835 45.85 4.002 ;
      RECT 45.77 3.86 45.775 4.025 ;
      RECT 45.755 3.864 45.77 4.031 ;
      RECT 45.745 3.872 45.755 4.036 ;
      RECT 45.715 3.885 45.745 4.04 ;
      RECT 45.705 3.9 45.715 4.045 ;
      RECT 45.695 3.905 45.705 4.048 ;
      RECT 45.69 3.907 45.695 4.05 ;
      RECT 45.675 3.91 45.69 4.053 ;
      RECT 45.67 3.912 45.675 4.056 ;
      RECT 45.65 3.917 45.67 4.06 ;
      RECT 45.62 3.922 45.65 4.068 ;
      RECT 45.595 3.929 45.62 4.076 ;
      RECT 45.59 3.934 45.595 4.081 ;
      RECT 45.56 3.937 45.59 4.085 ;
      RECT 45.52 3.94 45.56 4.095 ;
      RECT 45.485 3.937 45.52 4.107 ;
      RECT 45.475 3.933 45.485 4.114 ;
      RECT 45.45 3.929 45.475 4.12 ;
      RECT 45.445 3.925 45.45 4.125 ;
      RECT 45.405 3.922 45.445 4.125 ;
      RECT 45.39 3.907 45.405 4.126 ;
      RECT 45.367 3.895 45.39 4.126 ;
      RECT 45.281 3.895 45.367 4.127 ;
      RECT 45.195 3.895 45.281 4.129 ;
      RECT 45.175 3.895 45.195 4.126 ;
      RECT 45.17 3.9 45.175 4.121 ;
      RECT 45.165 3.905 45.17 4.119 ;
      RECT 45.155 3.915 45.165 4.117 ;
      RECT 45.15 3.921 45.155 4.11 ;
      RECT 45.145 3.923 45.15 4.095 ;
      RECT 45.14 3.927 45.145 4.085 ;
      RECT 46.6 3.395 46.85 3.655 ;
      RECT 44.325 4.93 44.585 5.19 ;
      RECT 46.62 4.42 46.625 4.63 ;
      RECT 46.625 4.425 46.635 4.625 ;
      RECT 46.575 4.42 46.62 4.645 ;
      RECT 46.565 4.42 46.575 4.665 ;
      RECT 46.546 4.42 46.565 4.67 ;
      RECT 46.46 4.42 46.546 4.667 ;
      RECT 46.43 4.422 46.46 4.665 ;
      RECT 46.375 4.432 46.43 4.663 ;
      RECT 46.31 4.446 46.375 4.661 ;
      RECT 46.305 4.454 46.31 4.66 ;
      RECT 46.29 4.457 46.305 4.658 ;
      RECT 46.225 4.467 46.29 4.654 ;
      RECT 46.177 4.481 46.225 4.655 ;
      RECT 46.091 4.498 46.177 4.669 ;
      RECT 46.005 4.519 46.091 4.686 ;
      RECT 45.985 4.532 46.005 4.696 ;
      RECT 45.94 4.54 45.985 4.703 ;
      RECT 45.905 4.548 45.94 4.711 ;
      RECT 45.871 4.556 45.905 4.719 ;
      RECT 45.785 4.57 45.871 4.731 ;
      RECT 45.75 4.587 45.785 4.743 ;
      RECT 45.741 4.596 45.75 4.747 ;
      RECT 45.655 4.614 45.741 4.764 ;
      RECT 45.596 4.641 45.655 4.791 ;
      RECT 45.51 4.668 45.596 4.819 ;
      RECT 45.49 4.69 45.51 4.839 ;
      RECT 45.43 4.705 45.49 4.855 ;
      RECT 45.42 4.717 45.43 4.868 ;
      RECT 45.415 4.722 45.42 4.871 ;
      RECT 45.405 4.725 45.415 4.874 ;
      RECT 45.4 4.727 45.405 4.877 ;
      RECT 45.37 4.735 45.4 4.884 ;
      RECT 45.355 4.742 45.37 4.892 ;
      RECT 45.345 4.747 45.355 4.896 ;
      RECT 45.34 4.75 45.345 4.899 ;
      RECT 45.33 4.752 45.34 4.902 ;
      RECT 45.295 4.762 45.33 4.911 ;
      RECT 45.22 4.785 45.295 4.933 ;
      RECT 45.2 4.803 45.22 4.951 ;
      RECT 45.17 4.81 45.2 4.961 ;
      RECT 45.15 4.818 45.17 4.971 ;
      RECT 45.14 4.824 45.15 4.978 ;
      RECT 45.121 4.829 45.14 4.984 ;
      RECT 45.035 4.849 45.121 5.004 ;
      RECT 45.02 4.869 45.035 5.023 ;
      RECT 44.975 4.881 45.02 5.034 ;
      RECT 44.91 4.902 44.975 5.057 ;
      RECT 44.87 4.922 44.91 5.078 ;
      RECT 44.86 4.932 44.87 5.088 ;
      RECT 44.81 4.944 44.86 5.099 ;
      RECT 44.79 4.96 44.81 5.111 ;
      RECT 44.76 4.97 44.79 5.117 ;
      RECT 44.75 4.975 44.76 5.119 ;
      RECT 44.681 4.976 44.75 5.125 ;
      RECT 44.595 4.978 44.681 5.135 ;
      RECT 44.585 4.979 44.595 5.14 ;
      RECT 45.855 5.005 46.045 5.215 ;
      RECT 45.845 5.01 46.055 5.208 ;
      RECT 45.83 5.01 46.055 5.173 ;
      RECT 45.75 4.895 46.01 5.155 ;
      RECT 44.665 4.425 44.85 4.72 ;
      RECT 44.655 4.425 44.85 4.718 ;
      RECT 44.64 4.425 44.855 4.713 ;
      RECT 44.64 4.425 44.86 4.71 ;
      RECT 44.635 4.425 44.86 4.708 ;
      RECT 44.63 4.68 44.86 4.698 ;
      RECT 44.635 4.425 44.895 4.685 ;
      RECT 44.595 3.46 44.855 3.72 ;
      RECT 44.405 3.385 44.491 3.718 ;
      RECT 44.38 3.389 44.535 3.714 ;
      RECT 44.491 3.381 44.535 3.714 ;
      RECT 44.491 3.382 44.54 3.713 ;
      RECT 44.405 3.387 44.555 3.712 ;
      RECT 44.38 3.395 44.595 3.711 ;
      RECT 44.375 3.39 44.555 3.706 ;
      RECT 44.365 3.405 44.595 3.613 ;
      RECT 44.365 3.457 44.795 3.613 ;
      RECT 44.365 3.45 44.775 3.613 ;
      RECT 44.365 3.437 44.745 3.613 ;
      RECT 44.365 3.425 44.685 3.613 ;
      RECT 44.365 3.41 44.66 3.613 ;
      RECT 43.565 4.04 43.7 4.335 ;
      RECT 43.825 4.063 43.83 4.25 ;
      RECT 44.545 3.96 44.69 4.195 ;
      RECT 44.705 3.96 44.71 4.185 ;
      RECT 44.74 3.971 44.745 4.165 ;
      RECT 44.735 3.963 44.74 4.17 ;
      RECT 44.715 3.96 44.735 4.175 ;
      RECT 44.71 3.96 44.715 4.183 ;
      RECT 44.7 3.96 44.705 4.188 ;
      RECT 44.69 3.96 44.7 4.193 ;
      RECT 44.52 3.962 44.545 4.195 ;
      RECT 44.47 3.969 44.52 4.195 ;
      RECT 44.465 3.974 44.47 4.195 ;
      RECT 44.426 3.979 44.465 4.196 ;
      RECT 44.34 3.991 44.426 4.197 ;
      RECT 44.331 4.001 44.34 4.197 ;
      RECT 44.245 4.01 44.331 4.199 ;
      RECT 44.221 4.02 44.245 4.201 ;
      RECT 44.135 4.031 44.221 4.202 ;
      RECT 44.105 4.042 44.135 4.204 ;
      RECT 44.075 4.047 44.105 4.206 ;
      RECT 44.05 4.053 44.075 4.209 ;
      RECT 44.035 4.058 44.05 4.21 ;
      RECT 43.99 4.064 44.035 4.21 ;
      RECT 43.985 4.069 43.99 4.211 ;
      RECT 43.965 4.069 43.985 4.213 ;
      RECT 43.945 4.067 43.965 4.218 ;
      RECT 43.91 4.066 43.945 4.225 ;
      RECT 43.88 4.065 43.91 4.235 ;
      RECT 43.83 4.064 43.88 4.245 ;
      RECT 43.74 4.061 43.825 4.335 ;
      RECT 43.715 4.055 43.74 4.335 ;
      RECT 43.7 4.045 43.715 4.335 ;
      RECT 43.515 4.04 43.565 4.255 ;
      RECT 43.505 4.045 43.515 4.245 ;
      RECT 43.745 4.52 44.005 4.78 ;
      RECT 43.745 4.52 44.035 4.673 ;
      RECT 43.745 4.52 44.07 4.658 ;
      RECT 44 4.44 44.19 4.65 ;
      RECT 43.99 4.445 44.2 4.643 ;
      RECT 43.955 4.515 44.2 4.643 ;
      RECT 43.985 4.457 44.005 4.78 ;
      RECT 43.97 4.505 44.2 4.643 ;
      RECT 43.975 4.477 44.005 4.78 ;
      RECT 43.055 3.545 43.125 4.65 ;
      RECT 43.79 3.65 44.05 3.91 ;
      RECT 43.37 3.696 43.385 3.905 ;
      RECT 43.706 3.709 43.79 3.86 ;
      RECT 43.62 3.706 43.706 3.86 ;
      RECT 43.581 3.704 43.62 3.86 ;
      RECT 43.495 3.702 43.581 3.86 ;
      RECT 43.435 3.7 43.495 3.871 ;
      RECT 43.4 3.698 43.435 3.889 ;
      RECT 43.385 3.696 43.4 3.9 ;
      RECT 43.355 3.696 43.37 3.913 ;
      RECT 43.345 3.696 43.355 3.918 ;
      RECT 43.32 3.695 43.345 3.923 ;
      RECT 43.305 3.69 43.32 3.929 ;
      RECT 43.3 3.683 43.305 3.934 ;
      RECT 43.275 3.674 43.3 3.94 ;
      RECT 43.23 3.653 43.275 3.953 ;
      RECT 43.22 3.637 43.23 3.963 ;
      RECT 43.205 3.63 43.22 3.973 ;
      RECT 43.195 3.623 43.205 3.99 ;
      RECT 43.19 3.62 43.195 4.02 ;
      RECT 43.185 3.618 43.19 4.05 ;
      RECT 43.18 3.616 43.185 4.087 ;
      RECT 43.165 3.612 43.18 4.154 ;
      RECT 43.165 4.445 43.175 4.645 ;
      RECT 43.16 3.608 43.165 4.28 ;
      RECT 43.16 4.432 43.165 4.65 ;
      RECT 43.155 3.606 43.16 4.365 ;
      RECT 43.155 4.422 43.16 4.65 ;
      RECT 43.14 3.577 43.155 4.65 ;
      RECT 43.125 3.55 43.14 4.65 ;
      RECT 43.05 3.545 43.055 3.9 ;
      RECT 43.05 3.955 43.055 4.65 ;
      RECT 43.035 3.545 43.05 3.878 ;
      RECT 43.045 3.977 43.05 4.65 ;
      RECT 43.035 4.017 43.045 4.65 ;
      RECT 43 3.545 43.035 3.82 ;
      RECT 43.03 4.052 43.035 4.65 ;
      RECT 43.015 4.107 43.03 4.65 ;
      RECT 43.01 4.172 43.015 4.65 ;
      RECT 42.995 4.22 43.01 4.65 ;
      RECT 42.97 3.545 43 3.775 ;
      RECT 42.99 4.275 42.995 4.65 ;
      RECT 42.975 4.335 42.99 4.65 ;
      RECT 42.97 4.383 42.975 4.648 ;
      RECT 42.965 3.545 42.97 3.768 ;
      RECT 42.965 4.415 42.97 4.643 ;
      RECT 42.94 3.545 42.965 3.76 ;
      RECT 42.93 3.55 42.94 3.75 ;
      RECT 43.145 4.825 43.165 5.065 ;
      RECT 42.375 4.755 42.38 4.965 ;
      RECT 43.655 4.828 43.665 5.023 ;
      RECT 43.65 4.818 43.655 5.026 ;
      RECT 43.57 4.815 43.65 5.049 ;
      RECT 43.566 4.815 43.57 5.071 ;
      RECT 43.48 4.815 43.566 5.081 ;
      RECT 43.465 4.815 43.48 5.089 ;
      RECT 43.436 4.816 43.465 5.087 ;
      RECT 43.35 4.821 43.436 5.083 ;
      RECT 43.337 4.825 43.35 5.079 ;
      RECT 43.251 4.825 43.337 5.075 ;
      RECT 43.165 4.825 43.251 5.069 ;
      RECT 43.081 4.825 43.145 5.063 ;
      RECT 42.995 4.825 43.081 5.058 ;
      RECT 42.975 4.825 42.995 5.054 ;
      RECT 42.915 4.82 42.975 5.051 ;
      RECT 42.887 4.814 42.915 5.048 ;
      RECT 42.801 4.809 42.887 5.044 ;
      RECT 42.715 4.803 42.801 5.038 ;
      RECT 42.64 4.785 42.715 5.033 ;
      RECT 42.605 4.762 42.64 5.029 ;
      RECT 42.595 4.752 42.605 5.028 ;
      RECT 42.54 4.75 42.595 5.027 ;
      RECT 42.465 4.75 42.54 5.023 ;
      RECT 42.455 4.75 42.465 5.018 ;
      RECT 42.44 4.75 42.455 5.01 ;
      RECT 42.39 4.752 42.44 4.988 ;
      RECT 42.38 4.755 42.39 4.968 ;
      RECT 42.37 4.76 42.375 4.963 ;
      RECT 42.365 4.765 42.37 4.958 ;
      RECT 42.49 3.93 42.75 4.19 ;
      RECT 42.49 3.945 42.77 4.155 ;
      RECT 42.49 3.95 42.78 4.15 ;
      RECT 40.475 3.41 40.735 3.67 ;
      RECT 40.465 3.44 40.735 3.65 ;
      RECT 42.385 3.355 42.645 3.615 ;
      RECT 42.38 3.43 42.385 3.616 ;
      RECT 42.355 3.435 42.38 3.618 ;
      RECT 42.34 3.442 42.355 3.621 ;
      RECT 42.28 3.46 42.34 3.626 ;
      RECT 42.25 3.48 42.28 3.633 ;
      RECT 42.225 3.488 42.25 3.638 ;
      RECT 42.2 3.496 42.225 3.64 ;
      RECT 42.182 3.5 42.2 3.639 ;
      RECT 42.096 3.498 42.182 3.639 ;
      RECT 42.01 3.496 42.096 3.639 ;
      RECT 41.924 3.494 42.01 3.638 ;
      RECT 41.838 3.492 41.924 3.638 ;
      RECT 41.752 3.49 41.838 3.638 ;
      RECT 41.666 3.488 41.752 3.638 ;
      RECT 41.58 3.486 41.666 3.637 ;
      RECT 41.562 3.485 41.58 3.637 ;
      RECT 41.476 3.484 41.562 3.637 ;
      RECT 41.39 3.482 41.476 3.637 ;
      RECT 41.304 3.481 41.39 3.636 ;
      RECT 41.218 3.48 41.304 3.636 ;
      RECT 41.132 3.478 41.218 3.636 ;
      RECT 41.046 3.477 41.132 3.636 ;
      RECT 40.96 3.475 41.046 3.635 ;
      RECT 40.936 3.473 40.96 3.635 ;
      RECT 40.85 3.466 40.936 3.635 ;
      RECT 40.821 3.458 40.85 3.635 ;
      RECT 40.735 3.45 40.821 3.635 ;
      RECT 40.455 3.447 40.465 3.645 ;
      RECT 41.96 4.41 41.965 4.76 ;
      RECT 41.73 4.5 41.87 4.76 ;
      RECT 42.205 4.185 42.25 4.395 ;
      RECT 42.26 4.196 42.27 4.39 ;
      RECT 42.25 4.188 42.26 4.395 ;
      RECT 42.185 4.185 42.205 4.4 ;
      RECT 42.155 4.185 42.185 4.423 ;
      RECT 42.145 4.185 42.155 4.448 ;
      RECT 42.14 4.185 42.145 4.458 ;
      RECT 42.085 4.185 42.14 4.498 ;
      RECT 42.08 4.185 42.085 4.538 ;
      RECT 42.075 4.187 42.08 4.543 ;
      RECT 42.06 4.197 42.075 4.554 ;
      RECT 42.015 4.255 42.06 4.59 ;
      RECT 42.005 4.31 42.015 4.624 ;
      RECT 41.99 4.337 42.005 4.64 ;
      RECT 41.98 4.364 41.99 4.76 ;
      RECT 41.965 4.387 41.98 4.76 ;
      RECT 41.955 4.427 41.96 4.76 ;
      RECT 41.95 4.437 41.955 4.76 ;
      RECT 41.945 4.452 41.95 4.76 ;
      RECT 41.935 4.457 41.945 4.76 ;
      RECT 41.87 4.48 41.935 4.76 ;
      RECT 41.37 3.975 41.56 4.185 ;
      RECT 39.945 3.9 40.205 4.16 ;
      RECT 40.295 3.895 40.39 4.105 ;
      RECT 40.27 3.91 40.28 4.105 ;
      RECT 41.56 3.982 41.57 4.18 ;
      RECT 41.36 3.982 41.37 4.18 ;
      RECT 41.345 3.997 41.36 4.17 ;
      RECT 41.34 4.005 41.345 4.163 ;
      RECT 41.33 4.008 41.34 4.16 ;
      RECT 41.295 4.007 41.33 4.158 ;
      RECT 41.266 4.003 41.295 4.155 ;
      RECT 41.18 3.998 41.266 4.152 ;
      RECT 41.12 3.992 41.18 4.148 ;
      RECT 41.091 3.988 41.12 4.145 ;
      RECT 41.005 3.98 41.091 4.142 ;
      RECT 40.996 3.974 41.005 4.14 ;
      RECT 40.91 3.969 40.996 4.138 ;
      RECT 40.887 3.964 40.91 4.135 ;
      RECT 40.801 3.958 40.887 4.132 ;
      RECT 40.715 3.949 40.801 4.127 ;
      RECT 40.705 3.944 40.715 4.125 ;
      RECT 40.686 3.943 40.705 4.124 ;
      RECT 40.6 3.938 40.686 4.12 ;
      RECT 40.58 3.933 40.6 4.116 ;
      RECT 40.52 3.928 40.58 4.113 ;
      RECT 40.495 3.918 40.52 4.111 ;
      RECT 40.49 3.911 40.495 4.11 ;
      RECT 40.48 3.902 40.49 4.109 ;
      RECT 40.476 3.895 40.48 4.109 ;
      RECT 40.39 3.895 40.476 4.107 ;
      RECT 40.28 3.902 40.295 4.105 ;
      RECT 40.265 3.912 40.27 4.105 ;
      RECT 40.245 3.915 40.265 4.102 ;
      RECT 40.215 3.915 40.245 4.098 ;
      RECT 40.205 3.915 40.215 4.098 ;
      RECT 41.12 4.41 41.38 4.67 ;
      RECT 41.05 4.42 41.38 4.63 ;
      RECT 41.04 4.427 41.38 4.625 ;
      RECT 40.46 4.415 40.72 4.675 ;
      RECT 40.46 4.455 40.825 4.665 ;
      RECT 40.46 4.457 40.83 4.664 ;
      RECT 40.46 4.465 40.835 4.661 ;
      RECT 39.385 3.54 39.485 5.065 ;
      RECT 39.575 4.68 39.625 4.94 ;
      RECT 39.57 3.553 39.575 3.74 ;
      RECT 39.565 4.661 39.575 4.94 ;
      RECT 39.565 3.55 39.57 3.748 ;
      RECT 39.55 3.544 39.565 3.755 ;
      RECT 39.56 4.649 39.565 5.023 ;
      RECT 39.55 4.637 39.56 5.06 ;
      RECT 39.54 3.54 39.55 3.762 ;
      RECT 39.54 4.622 39.55 5.065 ;
      RECT 39.535 3.54 39.54 3.77 ;
      RECT 39.515 4.592 39.54 5.065 ;
      RECT 39.495 3.54 39.535 3.818 ;
      RECT 39.505 4.552 39.515 5.065 ;
      RECT 39.495 4.507 39.505 5.065 ;
      RECT 39.49 3.54 39.495 3.888 ;
      RECT 39.49 4.465 39.495 5.065 ;
      RECT 39.485 3.54 39.49 4.365 ;
      RECT 39.485 4.447 39.49 5.065 ;
      RECT 39.375 3.543 39.385 5.065 ;
      RECT 39.36 3.55 39.375 5.061 ;
      RECT 39.355 3.56 39.36 5.056 ;
      RECT 39.35 3.76 39.355 4.948 ;
      RECT 39.345 3.845 39.35 4.5 ;
      RECT 38.22 10.205 38.51 10.435 ;
      RECT 38.28 8.725 38.45 10.435 ;
      RECT 38.27 9.095 38.625 9.45 ;
      RECT 38.22 8.725 38.51 8.955 ;
      RECT 37.815 3.69 37.92 4.26 ;
      RECT 37.815 4.025 38.14 4.255 ;
      RECT 37.815 4.055 38.31 4.225 ;
      RECT 37.815 3.69 38.005 4.255 ;
      RECT 37.23 3.655 37.52 3.885 ;
      RECT 37.23 3.69 38.005 3.86 ;
      RECT 37.29 2.175 37.46 3.885 ;
      RECT 37.23 2.175 37.52 2.405 ;
      RECT 37.23 10.205 37.52 10.435 ;
      RECT 37.29 8.725 37.46 10.435 ;
      RECT 37.23 8.725 37.52 8.955 ;
      RECT 37.23 8.76 38.085 8.92 ;
      RECT 37.915 8.355 38.085 8.92 ;
      RECT 37.23 8.755 37.625 8.92 ;
      RECT 37.85 8.355 38.14 8.585 ;
      RECT 37.85 8.385 38.31 8.555 ;
      RECT 36.86 4.025 37.15 4.255 ;
      RECT 36.86 4.055 37.32 4.225 ;
      RECT 36.925 2.95 37.09 4.255 ;
      RECT 35.44 2.92 35.73 3.15 ;
      RECT 35.44 2.95 37.09 3.12 ;
      RECT 35.5 2.18 35.67 3.15 ;
      RECT 35.44 2.18 35.73 2.41 ;
      RECT 35.44 10.2 35.73 10.43 ;
      RECT 35.5 9.46 35.67 10.43 ;
      RECT 35.5 9.555 37.09 9.725 ;
      RECT 36.92 8.355 37.09 9.725 ;
      RECT 35.44 9.46 35.73 9.69 ;
      RECT 36.86 8.355 37.15 8.585 ;
      RECT 36.86 8.385 37.32 8.555 ;
      RECT 33.475 4.725 33.825 5.075 ;
      RECT 33.565 3.32 33.735 5.075 ;
      RECT 35.87 3.26 36.22 3.61 ;
      RECT 33.565 3.32 35.185 3.495 ;
      RECT 33.565 3.32 36.22 3.49 ;
      RECT 35.895 9.09 36.22 9.415 ;
      RECT 31.32 9.045 31.67 9.395 ;
      RECT 35.87 9.09 36.22 9.32 ;
      RECT 31.11 9.09 31.67 9.32 ;
      RECT 30.94 9.12 36.22 9.29 ;
      RECT 35.095 3.66 35.415 3.98 ;
      RECT 35.065 3.66 35.415 3.89 ;
      RECT 34.895 3.69 35.415 3.86 ;
      RECT 35.095 8.66 35.415 8.98 ;
      RECT 35.065 8.72 35.415 8.95 ;
      RECT 34.895 8.75 35.415 8.92 ;
      RECT 30.875 4.96 30.915 5.22 ;
      RECT 30.915 4.94 30.92 4.95 ;
      RECT 32.245 4.185 32.255 4.406 ;
      RECT 32.175 4.18 32.245 4.531 ;
      RECT 32.165 4.18 32.175 4.658 ;
      RECT 32.14 4.18 32.165 4.705 ;
      RECT 32.115 4.18 32.14 4.783 ;
      RECT 32.095 4.18 32.115 4.853 ;
      RECT 32.07 4.18 32.095 4.893 ;
      RECT 32.06 4.18 32.07 4.913 ;
      RECT 32.05 4.182 32.06 4.921 ;
      RECT 32.045 4.187 32.05 4.378 ;
      RECT 32.045 4.387 32.05 4.922 ;
      RECT 32.04 4.432 32.045 4.923 ;
      RECT 32.03 4.497 32.04 4.924 ;
      RECT 32.02 4.592 32.03 4.926 ;
      RECT 32.015 4.645 32.02 4.928 ;
      RECT 32.01 4.665 32.015 4.929 ;
      RECT 31.955 4.69 32.01 4.935 ;
      RECT 31.915 4.725 31.955 4.944 ;
      RECT 31.905 4.742 31.915 4.949 ;
      RECT 31.896 4.748 31.905 4.951 ;
      RECT 31.81 4.786 31.896 4.962 ;
      RECT 31.805 4.825 31.81 4.972 ;
      RECT 31.73 4.832 31.805 4.982 ;
      RECT 31.71 4.842 31.73 4.993 ;
      RECT 31.68 4.849 31.71 5.001 ;
      RECT 31.655 4.856 31.68 5.008 ;
      RECT 31.631 4.862 31.655 5.013 ;
      RECT 31.545 4.875 31.631 5.025 ;
      RECT 31.467 4.882 31.545 5.043 ;
      RECT 31.381 4.877 31.467 5.061 ;
      RECT 31.295 4.872 31.381 5.081 ;
      RECT 31.215 4.866 31.295 5.098 ;
      RECT 31.15 4.862 31.215 5.127 ;
      RECT 31.145 4.576 31.15 4.6 ;
      RECT 31.135 4.852 31.15 5.155 ;
      RECT 31.14 4.57 31.145 4.64 ;
      RECT 31.135 4.564 31.14 4.71 ;
      RECT 31.13 4.558 31.135 4.788 ;
      RECT 31.13 4.835 31.135 5.22 ;
      RECT 31.122 4.555 31.13 5.22 ;
      RECT 31.036 4.553 31.122 5.22 ;
      RECT 30.95 4.551 31.036 5.22 ;
      RECT 30.94 4.552 30.95 5.22 ;
      RECT 30.935 4.557 30.94 5.22 ;
      RECT 30.925 4.57 30.935 5.22 ;
      RECT 30.92 4.592 30.925 5.22 ;
      RECT 30.915 4.952 30.92 5.22 ;
      RECT 31.545 4.42 31.55 4.64 ;
      RECT 32.05 3.455 32.085 3.715 ;
      RECT 32.035 3.455 32.05 3.723 ;
      RECT 32.006 3.455 32.035 3.745 ;
      RECT 31.92 3.455 32.006 3.805 ;
      RECT 31.9 3.455 31.92 3.87 ;
      RECT 31.84 3.455 31.9 4.035 ;
      RECT 31.835 3.455 31.84 4.183 ;
      RECT 31.83 3.455 31.835 4.195 ;
      RECT 31.825 3.455 31.83 4.221 ;
      RECT 31.795 3.641 31.825 4.301 ;
      RECT 31.79 3.689 31.795 4.39 ;
      RECT 31.785 3.703 31.79 4.405 ;
      RECT 31.78 3.722 31.785 4.435 ;
      RECT 31.775 3.737 31.78 4.451 ;
      RECT 31.77 3.752 31.775 4.473 ;
      RECT 31.765 3.772 31.77 4.495 ;
      RECT 31.755 3.792 31.765 4.528 ;
      RECT 31.74 3.834 31.755 4.59 ;
      RECT 31.735 3.865 31.74 4.63 ;
      RECT 31.73 3.877 31.735 4.635 ;
      RECT 31.725 3.889 31.73 4.64 ;
      RECT 31.72 3.902 31.725 4.64 ;
      RECT 31.715 3.92 31.72 4.64 ;
      RECT 31.71 3.94 31.715 4.64 ;
      RECT 31.705 3.952 31.71 4.64 ;
      RECT 31.7 3.965 31.705 4.64 ;
      RECT 31.68 4 31.7 4.64 ;
      RECT 31.63 4.102 31.68 4.64 ;
      RECT 31.625 4.187 31.63 4.64 ;
      RECT 31.62 4.195 31.625 4.64 ;
      RECT 31.615 4.212 31.62 4.64 ;
      RECT 31.61 4.227 31.615 4.64 ;
      RECT 31.575 4.292 31.61 4.64 ;
      RECT 31.56 4.357 31.575 4.64 ;
      RECT 31.555 4.387 31.56 4.64 ;
      RECT 31.55 4.412 31.555 4.64 ;
      RECT 31.535 4.422 31.545 4.64 ;
      RECT 31.52 4.435 31.535 4.633 ;
      RECT 31.265 4.025 31.335 4.235 ;
      RECT 31.055 4.002 31.06 4.195 ;
      RECT 28.51 3.93 28.77 4.19 ;
      RECT 31.345 4.212 31.35 4.215 ;
      RECT 31.335 4.03 31.345 4.23 ;
      RECT 31.236 4.023 31.265 4.235 ;
      RECT 31.15 4.015 31.236 4.235 ;
      RECT 31.135 4.009 31.15 4.233 ;
      RECT 31.115 4.008 31.135 4.22 ;
      RECT 31.11 4.007 31.115 4.203 ;
      RECT 31.06 4.004 31.11 4.198 ;
      RECT 31.03 4.001 31.055 4.193 ;
      RECT 31.01 3.999 31.03 4.188 ;
      RECT 30.995 3.997 31.01 4.185 ;
      RECT 30.965 3.995 30.995 4.183 ;
      RECT 30.9 3.991 30.965 4.175 ;
      RECT 30.87 3.986 30.9 4.17 ;
      RECT 30.85 3.984 30.87 4.168 ;
      RECT 30.82 3.981 30.85 4.163 ;
      RECT 30.76 3.977 30.82 4.155 ;
      RECT 30.755 3.974 30.76 4.15 ;
      RECT 30.685 3.972 30.755 4.145 ;
      RECT 30.656 3.968 30.685 4.138 ;
      RECT 30.57 3.963 30.656 4.13 ;
      RECT 30.536 3.958 30.57 4.122 ;
      RECT 30.45 3.95 30.536 4.114 ;
      RECT 30.411 3.943 30.45 4.106 ;
      RECT 30.325 3.938 30.411 4.098 ;
      RECT 30.26 3.932 30.325 4.088 ;
      RECT 30.24 3.927 30.26 4.083 ;
      RECT 30.231 3.924 30.24 4.082 ;
      RECT 30.145 3.92 30.231 4.076 ;
      RECT 30.105 3.916 30.145 4.068 ;
      RECT 30.085 3.912 30.105 4.066 ;
      RECT 30.025 3.912 30.085 4.063 ;
      RECT 30.005 3.915 30.025 4.061 ;
      RECT 29.984 3.915 30.005 4.061 ;
      RECT 29.898 3.917 29.984 4.065 ;
      RECT 29.812 3.919 29.898 4.071 ;
      RECT 29.726 3.921 29.812 4.078 ;
      RECT 29.64 3.924 29.726 4.084 ;
      RECT 29.606 3.925 29.64 4.089 ;
      RECT 29.52 3.928 29.606 4.094 ;
      RECT 29.491 3.935 29.52 4.099 ;
      RECT 29.405 3.935 29.491 4.104 ;
      RECT 29.372 3.935 29.405 4.109 ;
      RECT 29.286 3.937 29.372 4.114 ;
      RECT 29.2 3.939 29.286 4.121 ;
      RECT 29.136 3.941 29.2 4.127 ;
      RECT 29.05 3.943 29.136 4.133 ;
      RECT 29.047 3.945 29.05 4.136 ;
      RECT 28.961 3.946 29.047 4.14 ;
      RECT 28.875 3.949 28.961 4.147 ;
      RECT 28.856 3.951 28.875 4.151 ;
      RECT 28.77 3.953 28.856 4.156 ;
      RECT 28.5 3.965 28.51 4.16 ;
      RECT 30.68 10.2 30.97 10.43 ;
      RECT 30.74 9.46 30.91 10.43 ;
      RECT 30.63 9.49 31.005 9.86 ;
      RECT 30.68 9.46 30.97 9.86 ;
      RECT 30.735 3.545 30.92 3.755 ;
      RECT 30.73 3.546 30.925 3.753 ;
      RECT 30.725 3.551 30.935 3.748 ;
      RECT 30.72 3.527 30.725 3.745 ;
      RECT 30.69 3.524 30.72 3.738 ;
      RECT 30.685 3.52 30.69 3.729 ;
      RECT 30.65 3.551 30.935 3.724 ;
      RECT 30.425 3.46 30.685 3.72 ;
      RECT 30.725 3.529 30.73 3.748 ;
      RECT 30.73 3.53 30.735 3.753 ;
      RECT 30.425 3.542 30.805 3.72 ;
      RECT 30.425 3.54 30.79 3.72 ;
      RECT 30.425 3.535 30.78 3.72 ;
      RECT 30.38 4.45 30.43 4.735 ;
      RECT 30.325 4.42 30.33 4.735 ;
      RECT 30.295 4.4 30.3 4.735 ;
      RECT 30.445 4.45 30.505 4.71 ;
      RECT 30.44 4.45 30.445 4.718 ;
      RECT 30.43 4.45 30.44 4.73 ;
      RECT 30.345 4.44 30.38 4.735 ;
      RECT 30.34 4.427 30.345 4.735 ;
      RECT 30.33 4.422 30.34 4.735 ;
      RECT 30.31 4.412 30.325 4.735 ;
      RECT 30.3 4.405 30.31 4.735 ;
      RECT 30.29 4.397 30.295 4.735 ;
      RECT 30.26 4.387 30.29 4.735 ;
      RECT 30.245 4.375 30.26 4.735 ;
      RECT 30.23 4.365 30.245 4.73 ;
      RECT 30.21 4.355 30.23 4.705 ;
      RECT 30.2 4.347 30.21 4.682 ;
      RECT 30.17 4.33 30.2 4.672 ;
      RECT 30.165 4.307 30.17 4.663 ;
      RECT 30.16 4.294 30.165 4.661 ;
      RECT 30.145 4.27 30.16 4.655 ;
      RECT 30.14 4.246 30.145 4.649 ;
      RECT 30.13 4.235 30.14 4.644 ;
      RECT 30.125 4.225 30.13 4.64 ;
      RECT 30.12 4.217 30.125 4.637 ;
      RECT 30.11 4.212 30.12 4.633 ;
      RECT 30.105 4.207 30.11 4.629 ;
      RECT 30.02 4.205 30.105 4.604 ;
      RECT 29.99 4.205 30.02 4.57 ;
      RECT 29.975 4.205 29.99 4.553 ;
      RECT 29.92 4.205 29.975 4.498 ;
      RECT 29.915 4.21 29.92 4.447 ;
      RECT 29.905 4.215 29.915 4.437 ;
      RECT 29.9 4.225 29.905 4.423 ;
      RECT 29.85 4.965 30.11 5.225 ;
      RECT 29.77 4.98 30.11 5.201 ;
      RECT 29.75 4.98 30.11 5.196 ;
      RECT 29.726 4.98 30.11 5.194 ;
      RECT 29.64 4.98 30.11 5.189 ;
      RECT 29.49 4.92 29.75 5.185 ;
      RECT 29.445 4.98 30.11 5.18 ;
      RECT 29.44 4.987 30.11 5.175 ;
      RECT 29.455 4.975 29.77 5.185 ;
      RECT 29.345 3.41 29.605 3.67 ;
      RECT 29.345 3.467 29.61 3.663 ;
      RECT 29.345 3.497 29.615 3.595 ;
      RECT 29.405 3.928 29.52 3.93 ;
      RECT 29.491 3.925 29.52 3.93 ;
      RECT 28.515 4.929 28.54 5.169 ;
      RECT 28.5 4.932 28.59 5.163 ;
      RECT 28.495 4.937 28.676 5.158 ;
      RECT 28.49 4.945 28.74 5.156 ;
      RECT 28.49 4.945 28.75 5.155 ;
      RECT 28.485 4.952 28.76 5.148 ;
      RECT 28.485 4.952 28.846 5.137 ;
      RECT 28.48 4.987 28.846 5.133 ;
      RECT 28.48 4.987 28.855 5.122 ;
      RECT 28.76 4.86 29.02 5.12 ;
      RECT 28.47 5.037 29.02 5.118 ;
      RECT 28.74 4.905 28.76 5.153 ;
      RECT 28.676 4.908 28.74 5.157 ;
      RECT 28.59 4.913 28.676 5.162 ;
      RECT 28.52 4.924 29.02 5.12 ;
      RECT 28.54 4.918 28.59 5.167 ;
      RECT 28.665 3.395 28.675 3.657 ;
      RECT 28.655 3.452 28.665 3.66 ;
      RECT 28.63 3.457 28.655 3.666 ;
      RECT 28.605 3.461 28.63 3.678 ;
      RECT 28.595 3.464 28.605 3.688 ;
      RECT 28.59 3.465 28.595 3.693 ;
      RECT 28.585 3.466 28.59 3.698 ;
      RECT 28.58 3.467 28.585 3.7 ;
      RECT 28.555 3.47 28.58 3.703 ;
      RECT 28.525 3.476 28.555 3.706 ;
      RECT 28.46 3.487 28.525 3.709 ;
      RECT 28.415 3.495 28.46 3.713 ;
      RECT 28.4 3.495 28.415 3.721 ;
      RECT 28.395 3.496 28.4 3.728 ;
      RECT 28.39 3.498 28.395 3.731 ;
      RECT 28.385 3.502 28.39 3.734 ;
      RECT 28.375 3.51 28.385 3.738 ;
      RECT 28.37 3.523 28.375 3.743 ;
      RECT 28.365 3.531 28.37 3.745 ;
      RECT 28.36 3.537 28.365 3.745 ;
      RECT 28.355 3.541 28.36 3.748 ;
      RECT 28.35 3.543 28.355 3.751 ;
      RECT 28.345 3.546 28.35 3.754 ;
      RECT 28.335 3.551 28.345 3.758 ;
      RECT 28.33 3.557 28.335 3.763 ;
      RECT 28.32 3.563 28.33 3.767 ;
      RECT 28.305 3.57 28.32 3.773 ;
      RECT 28.276 3.584 28.305 3.783 ;
      RECT 28.19 3.619 28.276 3.815 ;
      RECT 28.17 3.652 28.19 3.844 ;
      RECT 28.15 3.665 28.17 3.855 ;
      RECT 28.13 3.677 28.15 3.866 ;
      RECT 28.08 3.699 28.13 3.886 ;
      RECT 28.065 3.717 28.08 3.903 ;
      RECT 28.06 3.723 28.065 3.906 ;
      RECT 28.055 3.727 28.06 3.909 ;
      RECT 28.05 3.731 28.055 3.913 ;
      RECT 28.045 3.733 28.05 3.916 ;
      RECT 28.035 3.74 28.045 3.919 ;
      RECT 28.03 3.745 28.035 3.923 ;
      RECT 28.025 3.747 28.03 3.926 ;
      RECT 28.02 3.751 28.025 3.929 ;
      RECT 28.015 3.753 28.02 3.933 ;
      RECT 28 3.758 28.015 3.938 ;
      RECT 27.995 3.763 28 3.941 ;
      RECT 27.99 3.771 27.995 3.944 ;
      RECT 27.985 3.773 27.99 3.947 ;
      RECT 27.98 3.775 27.985 3.95 ;
      RECT 27.97 3.777 27.98 3.956 ;
      RECT 27.935 3.791 27.97 3.968 ;
      RECT 27.925 3.806 27.935 3.978 ;
      RECT 27.85 3.835 27.925 4.002 ;
      RECT 27.845 3.86 27.85 4.025 ;
      RECT 27.83 3.864 27.845 4.031 ;
      RECT 27.82 3.872 27.83 4.036 ;
      RECT 27.79 3.885 27.82 4.04 ;
      RECT 27.78 3.9 27.79 4.045 ;
      RECT 27.77 3.905 27.78 4.048 ;
      RECT 27.765 3.907 27.77 4.05 ;
      RECT 27.75 3.91 27.765 4.053 ;
      RECT 27.745 3.912 27.75 4.056 ;
      RECT 27.725 3.917 27.745 4.06 ;
      RECT 27.695 3.922 27.725 4.068 ;
      RECT 27.67 3.929 27.695 4.076 ;
      RECT 27.665 3.934 27.67 4.081 ;
      RECT 27.635 3.937 27.665 4.085 ;
      RECT 27.595 3.94 27.635 4.095 ;
      RECT 27.56 3.937 27.595 4.107 ;
      RECT 27.55 3.933 27.56 4.114 ;
      RECT 27.525 3.929 27.55 4.12 ;
      RECT 27.52 3.925 27.525 4.125 ;
      RECT 27.48 3.922 27.52 4.125 ;
      RECT 27.465 3.907 27.48 4.126 ;
      RECT 27.442 3.895 27.465 4.126 ;
      RECT 27.356 3.895 27.442 4.127 ;
      RECT 27.27 3.895 27.356 4.129 ;
      RECT 27.25 3.895 27.27 4.126 ;
      RECT 27.245 3.9 27.25 4.121 ;
      RECT 27.24 3.905 27.245 4.119 ;
      RECT 27.23 3.915 27.24 4.117 ;
      RECT 27.225 3.921 27.23 4.11 ;
      RECT 27.22 3.923 27.225 4.095 ;
      RECT 27.215 3.927 27.22 4.085 ;
      RECT 28.675 3.395 28.925 3.655 ;
      RECT 26.4 4.93 26.66 5.19 ;
      RECT 28.695 4.42 28.7 4.63 ;
      RECT 28.7 4.425 28.71 4.625 ;
      RECT 28.65 4.42 28.695 4.645 ;
      RECT 28.64 4.42 28.65 4.665 ;
      RECT 28.621 4.42 28.64 4.67 ;
      RECT 28.535 4.42 28.621 4.667 ;
      RECT 28.505 4.422 28.535 4.665 ;
      RECT 28.45 4.432 28.505 4.663 ;
      RECT 28.385 4.446 28.45 4.661 ;
      RECT 28.38 4.454 28.385 4.66 ;
      RECT 28.365 4.457 28.38 4.658 ;
      RECT 28.3 4.467 28.365 4.654 ;
      RECT 28.252 4.481 28.3 4.655 ;
      RECT 28.166 4.498 28.252 4.669 ;
      RECT 28.08 4.519 28.166 4.686 ;
      RECT 28.06 4.532 28.08 4.696 ;
      RECT 28.015 4.54 28.06 4.703 ;
      RECT 27.98 4.548 28.015 4.711 ;
      RECT 27.946 4.556 27.98 4.719 ;
      RECT 27.86 4.57 27.946 4.731 ;
      RECT 27.825 4.587 27.86 4.743 ;
      RECT 27.816 4.596 27.825 4.747 ;
      RECT 27.73 4.614 27.816 4.764 ;
      RECT 27.671 4.641 27.73 4.791 ;
      RECT 27.585 4.668 27.671 4.819 ;
      RECT 27.565 4.69 27.585 4.839 ;
      RECT 27.505 4.705 27.565 4.855 ;
      RECT 27.495 4.717 27.505 4.868 ;
      RECT 27.49 4.722 27.495 4.871 ;
      RECT 27.48 4.725 27.49 4.874 ;
      RECT 27.475 4.727 27.48 4.877 ;
      RECT 27.445 4.735 27.475 4.884 ;
      RECT 27.43 4.742 27.445 4.892 ;
      RECT 27.42 4.747 27.43 4.896 ;
      RECT 27.415 4.75 27.42 4.899 ;
      RECT 27.405 4.752 27.415 4.902 ;
      RECT 27.37 4.762 27.405 4.911 ;
      RECT 27.295 4.785 27.37 4.933 ;
      RECT 27.275 4.803 27.295 4.951 ;
      RECT 27.245 4.81 27.275 4.961 ;
      RECT 27.225 4.818 27.245 4.971 ;
      RECT 27.215 4.824 27.225 4.978 ;
      RECT 27.196 4.829 27.215 4.984 ;
      RECT 27.11 4.849 27.196 5.004 ;
      RECT 27.095 4.869 27.11 5.023 ;
      RECT 27.05 4.881 27.095 5.034 ;
      RECT 26.985 4.902 27.05 5.057 ;
      RECT 26.945 4.922 26.985 5.078 ;
      RECT 26.935 4.932 26.945 5.088 ;
      RECT 26.885 4.944 26.935 5.099 ;
      RECT 26.865 4.96 26.885 5.111 ;
      RECT 26.835 4.97 26.865 5.117 ;
      RECT 26.825 4.975 26.835 5.119 ;
      RECT 26.756 4.976 26.825 5.125 ;
      RECT 26.67 4.978 26.756 5.135 ;
      RECT 26.66 4.979 26.67 5.14 ;
      RECT 27.93 5.005 28.12 5.215 ;
      RECT 27.92 5.01 28.13 5.208 ;
      RECT 27.905 5.01 28.13 5.173 ;
      RECT 27.825 4.895 28.085 5.155 ;
      RECT 26.74 4.425 26.925 4.72 ;
      RECT 26.73 4.425 26.925 4.718 ;
      RECT 26.715 4.425 26.93 4.713 ;
      RECT 26.715 4.425 26.935 4.71 ;
      RECT 26.71 4.425 26.935 4.708 ;
      RECT 26.705 4.68 26.935 4.698 ;
      RECT 26.71 4.425 26.97 4.685 ;
      RECT 26.67 3.46 26.93 3.72 ;
      RECT 26.48 3.385 26.566 3.718 ;
      RECT 26.455 3.389 26.61 3.714 ;
      RECT 26.566 3.381 26.61 3.714 ;
      RECT 26.566 3.382 26.615 3.713 ;
      RECT 26.48 3.387 26.63 3.712 ;
      RECT 26.455 3.395 26.67 3.711 ;
      RECT 26.45 3.39 26.63 3.706 ;
      RECT 26.44 3.405 26.67 3.613 ;
      RECT 26.44 3.457 26.87 3.613 ;
      RECT 26.44 3.45 26.85 3.613 ;
      RECT 26.44 3.437 26.82 3.613 ;
      RECT 26.44 3.425 26.76 3.613 ;
      RECT 26.44 3.41 26.735 3.613 ;
      RECT 25.64 4.04 25.775 4.335 ;
      RECT 25.9 4.063 25.905 4.25 ;
      RECT 26.62 3.96 26.765 4.195 ;
      RECT 26.78 3.96 26.785 4.185 ;
      RECT 26.815 3.971 26.82 4.165 ;
      RECT 26.81 3.963 26.815 4.17 ;
      RECT 26.79 3.96 26.81 4.175 ;
      RECT 26.785 3.96 26.79 4.183 ;
      RECT 26.775 3.96 26.78 4.188 ;
      RECT 26.765 3.96 26.775 4.193 ;
      RECT 26.595 3.962 26.62 4.195 ;
      RECT 26.545 3.969 26.595 4.195 ;
      RECT 26.54 3.974 26.545 4.195 ;
      RECT 26.501 3.979 26.54 4.196 ;
      RECT 26.415 3.991 26.501 4.197 ;
      RECT 26.406 4.001 26.415 4.197 ;
      RECT 26.32 4.01 26.406 4.199 ;
      RECT 26.296 4.02 26.32 4.201 ;
      RECT 26.21 4.031 26.296 4.202 ;
      RECT 26.18 4.042 26.21 4.204 ;
      RECT 26.15 4.047 26.18 4.206 ;
      RECT 26.125 4.053 26.15 4.209 ;
      RECT 26.11 4.058 26.125 4.21 ;
      RECT 26.065 4.064 26.11 4.21 ;
      RECT 26.06 4.069 26.065 4.211 ;
      RECT 26.04 4.069 26.06 4.213 ;
      RECT 26.02 4.067 26.04 4.218 ;
      RECT 25.985 4.066 26.02 4.225 ;
      RECT 25.955 4.065 25.985 4.235 ;
      RECT 25.905 4.064 25.955 4.245 ;
      RECT 25.815 4.061 25.9 4.335 ;
      RECT 25.79 4.055 25.815 4.335 ;
      RECT 25.775 4.045 25.79 4.335 ;
      RECT 25.59 4.04 25.64 4.255 ;
      RECT 25.58 4.045 25.59 4.245 ;
      RECT 25.82 4.52 26.08 4.78 ;
      RECT 25.82 4.52 26.11 4.673 ;
      RECT 25.82 4.52 26.145 4.658 ;
      RECT 26.075 4.44 26.265 4.65 ;
      RECT 26.065 4.445 26.275 4.643 ;
      RECT 26.03 4.515 26.275 4.643 ;
      RECT 26.06 4.457 26.08 4.78 ;
      RECT 26.045 4.505 26.275 4.643 ;
      RECT 26.05 4.477 26.08 4.78 ;
      RECT 25.13 3.545 25.2 4.65 ;
      RECT 25.865 3.65 26.125 3.91 ;
      RECT 25.445 3.696 25.46 3.905 ;
      RECT 25.781 3.709 25.865 3.86 ;
      RECT 25.695 3.706 25.781 3.86 ;
      RECT 25.656 3.704 25.695 3.86 ;
      RECT 25.57 3.702 25.656 3.86 ;
      RECT 25.51 3.7 25.57 3.871 ;
      RECT 25.475 3.698 25.51 3.889 ;
      RECT 25.46 3.696 25.475 3.9 ;
      RECT 25.43 3.696 25.445 3.913 ;
      RECT 25.42 3.696 25.43 3.918 ;
      RECT 25.395 3.695 25.42 3.923 ;
      RECT 25.38 3.69 25.395 3.929 ;
      RECT 25.375 3.683 25.38 3.934 ;
      RECT 25.35 3.674 25.375 3.94 ;
      RECT 25.305 3.653 25.35 3.953 ;
      RECT 25.295 3.637 25.305 3.963 ;
      RECT 25.28 3.63 25.295 3.973 ;
      RECT 25.27 3.623 25.28 3.99 ;
      RECT 25.265 3.62 25.27 4.02 ;
      RECT 25.26 3.618 25.265 4.05 ;
      RECT 25.255 3.616 25.26 4.087 ;
      RECT 25.24 3.612 25.255 4.154 ;
      RECT 25.24 4.445 25.25 4.645 ;
      RECT 25.235 3.608 25.24 4.28 ;
      RECT 25.235 4.432 25.24 4.65 ;
      RECT 25.23 3.606 25.235 4.365 ;
      RECT 25.23 4.422 25.235 4.65 ;
      RECT 25.215 3.577 25.23 4.65 ;
      RECT 25.2 3.55 25.215 4.65 ;
      RECT 25.125 3.545 25.13 3.9 ;
      RECT 25.125 3.955 25.13 4.65 ;
      RECT 25.11 3.545 25.125 3.878 ;
      RECT 25.12 3.977 25.125 4.65 ;
      RECT 25.11 4.017 25.12 4.65 ;
      RECT 25.075 3.545 25.11 3.82 ;
      RECT 25.105 4.052 25.11 4.65 ;
      RECT 25.09 4.107 25.105 4.65 ;
      RECT 25.085 4.172 25.09 4.65 ;
      RECT 25.07 4.22 25.085 4.65 ;
      RECT 25.045 3.545 25.075 3.775 ;
      RECT 25.065 4.275 25.07 4.65 ;
      RECT 25.05 4.335 25.065 4.65 ;
      RECT 25.045 4.383 25.05 4.648 ;
      RECT 25.04 3.545 25.045 3.768 ;
      RECT 25.04 4.415 25.045 4.643 ;
      RECT 25.015 3.545 25.04 3.76 ;
      RECT 25.005 3.55 25.015 3.75 ;
      RECT 25.22 4.825 25.24 5.065 ;
      RECT 24.45 4.755 24.455 4.965 ;
      RECT 25.73 4.828 25.74 5.023 ;
      RECT 25.725 4.818 25.73 5.026 ;
      RECT 25.645 4.815 25.725 5.049 ;
      RECT 25.641 4.815 25.645 5.071 ;
      RECT 25.555 4.815 25.641 5.081 ;
      RECT 25.54 4.815 25.555 5.089 ;
      RECT 25.511 4.816 25.54 5.087 ;
      RECT 25.425 4.821 25.511 5.083 ;
      RECT 25.412 4.825 25.425 5.079 ;
      RECT 25.326 4.825 25.412 5.075 ;
      RECT 25.24 4.825 25.326 5.069 ;
      RECT 25.156 4.825 25.22 5.063 ;
      RECT 25.07 4.825 25.156 5.058 ;
      RECT 25.05 4.825 25.07 5.054 ;
      RECT 24.99 4.82 25.05 5.051 ;
      RECT 24.962 4.814 24.99 5.048 ;
      RECT 24.876 4.809 24.962 5.044 ;
      RECT 24.79 4.803 24.876 5.038 ;
      RECT 24.715 4.785 24.79 5.033 ;
      RECT 24.68 4.762 24.715 5.029 ;
      RECT 24.67 4.752 24.68 5.028 ;
      RECT 24.615 4.75 24.67 5.027 ;
      RECT 24.54 4.75 24.615 5.023 ;
      RECT 24.53 4.75 24.54 5.018 ;
      RECT 24.515 4.75 24.53 5.01 ;
      RECT 24.465 4.752 24.515 4.988 ;
      RECT 24.455 4.755 24.465 4.968 ;
      RECT 24.445 4.76 24.45 4.963 ;
      RECT 24.44 4.765 24.445 4.958 ;
      RECT 24.565 3.93 24.825 4.19 ;
      RECT 24.565 3.945 24.845 4.155 ;
      RECT 24.565 3.95 24.855 4.15 ;
      RECT 22.55 3.41 22.81 3.67 ;
      RECT 22.54 3.44 22.81 3.65 ;
      RECT 24.46 3.355 24.72 3.615 ;
      RECT 24.455 3.43 24.46 3.616 ;
      RECT 24.43 3.435 24.455 3.618 ;
      RECT 24.415 3.442 24.43 3.621 ;
      RECT 24.355 3.46 24.415 3.626 ;
      RECT 24.325 3.48 24.355 3.633 ;
      RECT 24.3 3.488 24.325 3.638 ;
      RECT 24.275 3.496 24.3 3.64 ;
      RECT 24.257 3.5 24.275 3.639 ;
      RECT 24.171 3.498 24.257 3.639 ;
      RECT 24.085 3.496 24.171 3.639 ;
      RECT 23.999 3.494 24.085 3.638 ;
      RECT 23.913 3.492 23.999 3.638 ;
      RECT 23.827 3.49 23.913 3.638 ;
      RECT 23.741 3.488 23.827 3.638 ;
      RECT 23.655 3.486 23.741 3.637 ;
      RECT 23.637 3.485 23.655 3.637 ;
      RECT 23.551 3.484 23.637 3.637 ;
      RECT 23.465 3.482 23.551 3.637 ;
      RECT 23.379 3.481 23.465 3.636 ;
      RECT 23.293 3.48 23.379 3.636 ;
      RECT 23.207 3.478 23.293 3.636 ;
      RECT 23.121 3.477 23.207 3.636 ;
      RECT 23.035 3.475 23.121 3.635 ;
      RECT 23.011 3.473 23.035 3.635 ;
      RECT 22.925 3.466 23.011 3.635 ;
      RECT 22.896 3.458 22.925 3.635 ;
      RECT 22.81 3.45 22.896 3.635 ;
      RECT 22.53 3.447 22.54 3.645 ;
      RECT 24.035 4.41 24.04 4.76 ;
      RECT 23.805 4.5 23.945 4.76 ;
      RECT 24.28 4.185 24.325 4.395 ;
      RECT 24.335 4.196 24.345 4.39 ;
      RECT 24.325 4.188 24.335 4.395 ;
      RECT 24.26 4.185 24.28 4.4 ;
      RECT 24.23 4.185 24.26 4.423 ;
      RECT 24.22 4.185 24.23 4.448 ;
      RECT 24.215 4.185 24.22 4.458 ;
      RECT 24.16 4.185 24.215 4.498 ;
      RECT 24.155 4.185 24.16 4.538 ;
      RECT 24.15 4.187 24.155 4.543 ;
      RECT 24.135 4.197 24.15 4.554 ;
      RECT 24.09 4.255 24.135 4.59 ;
      RECT 24.08 4.31 24.09 4.624 ;
      RECT 24.065 4.337 24.08 4.64 ;
      RECT 24.055 4.364 24.065 4.76 ;
      RECT 24.04 4.387 24.055 4.76 ;
      RECT 24.03 4.427 24.035 4.76 ;
      RECT 24.025 4.437 24.03 4.76 ;
      RECT 24.02 4.452 24.025 4.76 ;
      RECT 24.01 4.457 24.02 4.76 ;
      RECT 23.945 4.48 24.01 4.76 ;
      RECT 23.445 3.975 23.635 4.185 ;
      RECT 22.02 3.9 22.28 4.16 ;
      RECT 22.37 3.895 22.465 4.105 ;
      RECT 22.345 3.91 22.355 4.105 ;
      RECT 23.635 3.982 23.645 4.18 ;
      RECT 23.435 3.982 23.445 4.18 ;
      RECT 23.42 3.997 23.435 4.17 ;
      RECT 23.415 4.005 23.42 4.163 ;
      RECT 23.405 4.008 23.415 4.16 ;
      RECT 23.37 4.007 23.405 4.158 ;
      RECT 23.341 4.003 23.37 4.155 ;
      RECT 23.255 3.998 23.341 4.152 ;
      RECT 23.195 3.992 23.255 4.148 ;
      RECT 23.166 3.988 23.195 4.145 ;
      RECT 23.08 3.98 23.166 4.142 ;
      RECT 23.071 3.974 23.08 4.14 ;
      RECT 22.985 3.969 23.071 4.138 ;
      RECT 22.962 3.964 22.985 4.135 ;
      RECT 22.876 3.958 22.962 4.132 ;
      RECT 22.79 3.949 22.876 4.127 ;
      RECT 22.78 3.944 22.79 4.125 ;
      RECT 22.761 3.943 22.78 4.124 ;
      RECT 22.675 3.938 22.761 4.12 ;
      RECT 22.655 3.933 22.675 4.116 ;
      RECT 22.595 3.928 22.655 4.113 ;
      RECT 22.57 3.918 22.595 4.111 ;
      RECT 22.565 3.911 22.57 4.11 ;
      RECT 22.555 3.902 22.565 4.109 ;
      RECT 22.551 3.895 22.555 4.109 ;
      RECT 22.465 3.895 22.551 4.107 ;
      RECT 22.355 3.902 22.37 4.105 ;
      RECT 22.34 3.912 22.345 4.105 ;
      RECT 22.32 3.915 22.34 4.102 ;
      RECT 22.29 3.915 22.32 4.098 ;
      RECT 22.28 3.915 22.29 4.098 ;
      RECT 23.195 4.41 23.455 4.67 ;
      RECT 23.125 4.42 23.455 4.63 ;
      RECT 23.115 4.427 23.455 4.625 ;
      RECT 22.535 4.415 22.795 4.675 ;
      RECT 22.535 4.455 22.9 4.665 ;
      RECT 22.535 4.457 22.905 4.664 ;
      RECT 22.535 4.465 22.91 4.661 ;
      RECT 21.46 3.54 21.56 5.065 ;
      RECT 21.65 4.68 21.7 4.94 ;
      RECT 21.645 3.553 21.65 3.74 ;
      RECT 21.64 4.661 21.65 4.94 ;
      RECT 21.64 3.55 21.645 3.748 ;
      RECT 21.625 3.544 21.64 3.755 ;
      RECT 21.635 4.649 21.64 5.023 ;
      RECT 21.625 4.637 21.635 5.06 ;
      RECT 21.615 3.54 21.625 3.762 ;
      RECT 21.615 4.622 21.625 5.065 ;
      RECT 21.61 3.54 21.615 3.77 ;
      RECT 21.59 4.592 21.615 5.065 ;
      RECT 21.57 3.54 21.61 3.818 ;
      RECT 21.58 4.552 21.59 5.065 ;
      RECT 21.57 4.507 21.58 5.065 ;
      RECT 21.565 3.54 21.57 3.888 ;
      RECT 21.565 4.465 21.57 5.065 ;
      RECT 21.56 3.54 21.565 4.365 ;
      RECT 21.56 4.447 21.565 5.065 ;
      RECT 21.45 3.543 21.46 5.065 ;
      RECT 21.435 3.55 21.45 5.061 ;
      RECT 21.43 3.56 21.435 5.056 ;
      RECT 21.425 3.76 21.43 4.948 ;
      RECT 21.42 3.845 21.425 4.5 ;
      RECT 20.295 10.205 20.585 10.435 ;
      RECT 20.355 8.725 20.525 10.435 ;
      RECT 20.35 9.09 20.7 9.44 ;
      RECT 20.295 8.725 20.585 8.955 ;
      RECT 19.89 3.69 19.995 4.26 ;
      RECT 19.89 4.025 20.215 4.255 ;
      RECT 19.89 4.055 20.385 4.225 ;
      RECT 19.89 3.69 20.08 4.255 ;
      RECT 19.305 3.655 19.595 3.885 ;
      RECT 19.305 3.69 20.08 3.86 ;
      RECT 19.365 2.175 19.535 3.885 ;
      RECT 19.305 2.175 19.595 2.405 ;
      RECT 19.305 10.205 19.595 10.435 ;
      RECT 19.365 8.725 19.535 10.435 ;
      RECT 19.305 8.725 19.595 8.955 ;
      RECT 19.305 8.76 20.16 8.92 ;
      RECT 19.99 8.355 20.16 8.92 ;
      RECT 19.305 8.755 19.7 8.92 ;
      RECT 19.925 8.355 20.215 8.585 ;
      RECT 19.925 8.385 20.385 8.555 ;
      RECT 18.935 4.025 19.225 4.255 ;
      RECT 18.935 4.055 19.395 4.225 ;
      RECT 19 2.95 19.165 4.255 ;
      RECT 17.515 2.92 17.805 3.15 ;
      RECT 17.515 2.95 19.165 3.12 ;
      RECT 17.575 2.18 17.745 3.15 ;
      RECT 17.515 2.18 17.805 2.41 ;
      RECT 17.515 10.2 17.805 10.43 ;
      RECT 17.575 9.46 17.745 10.43 ;
      RECT 17.575 9.555 19.165 9.725 ;
      RECT 18.995 8.355 19.165 9.725 ;
      RECT 17.515 9.46 17.805 9.69 ;
      RECT 18.935 8.355 19.225 8.585 ;
      RECT 18.935 8.385 19.395 8.555 ;
      RECT 15.55 4.725 15.9 5.075 ;
      RECT 15.64 3.32 15.81 5.075 ;
      RECT 17.945 3.26 18.295 3.61 ;
      RECT 15.64 3.32 17.26 3.495 ;
      RECT 15.64 3.32 18.295 3.49 ;
      RECT 17.97 9.09 18.295 9.415 ;
      RECT 13.365 9.04 13.715 9.39 ;
      RECT 17.945 9.09 18.295 9.32 ;
      RECT 13.185 9.09 13.715 9.32 ;
      RECT 13.015 9.12 18.295 9.29 ;
      RECT 17.17 3.66 17.49 3.98 ;
      RECT 17.14 3.66 17.49 3.89 ;
      RECT 16.97 3.69 17.49 3.86 ;
      RECT 17.17 8.66 17.49 8.98 ;
      RECT 17.14 8.72 17.49 8.95 ;
      RECT 16.97 8.75 17.49 8.92 ;
      RECT 12.95 4.96 12.99 5.22 ;
      RECT 12.99 4.94 12.995 4.95 ;
      RECT 14.32 4.185 14.33 4.406 ;
      RECT 14.25 4.18 14.32 4.531 ;
      RECT 14.24 4.18 14.25 4.658 ;
      RECT 14.215 4.18 14.24 4.705 ;
      RECT 14.19 4.18 14.215 4.783 ;
      RECT 14.17 4.18 14.19 4.853 ;
      RECT 14.145 4.18 14.17 4.893 ;
      RECT 14.135 4.18 14.145 4.913 ;
      RECT 14.125 4.182 14.135 4.921 ;
      RECT 14.12 4.187 14.125 4.378 ;
      RECT 14.12 4.387 14.125 4.922 ;
      RECT 14.115 4.432 14.12 4.923 ;
      RECT 14.105 4.497 14.115 4.924 ;
      RECT 14.095 4.592 14.105 4.926 ;
      RECT 14.09 4.645 14.095 4.928 ;
      RECT 14.085 4.665 14.09 4.929 ;
      RECT 14.03 4.69 14.085 4.935 ;
      RECT 13.99 4.725 14.03 4.944 ;
      RECT 13.98 4.742 13.99 4.949 ;
      RECT 13.971 4.748 13.98 4.951 ;
      RECT 13.885 4.786 13.971 4.962 ;
      RECT 13.88 4.825 13.885 4.972 ;
      RECT 13.805 4.832 13.88 4.982 ;
      RECT 13.785 4.842 13.805 4.993 ;
      RECT 13.755 4.849 13.785 5.001 ;
      RECT 13.73 4.856 13.755 5.008 ;
      RECT 13.706 4.862 13.73 5.013 ;
      RECT 13.62 4.875 13.706 5.025 ;
      RECT 13.542 4.882 13.62 5.043 ;
      RECT 13.456 4.877 13.542 5.061 ;
      RECT 13.37 4.872 13.456 5.081 ;
      RECT 13.29 4.866 13.37 5.098 ;
      RECT 13.225 4.862 13.29 5.127 ;
      RECT 13.22 4.576 13.225 4.6 ;
      RECT 13.21 4.852 13.225 5.155 ;
      RECT 13.215 4.57 13.22 4.64 ;
      RECT 13.21 4.564 13.215 4.71 ;
      RECT 13.205 4.558 13.21 4.788 ;
      RECT 13.205 4.835 13.21 5.22 ;
      RECT 13.197 4.555 13.205 5.22 ;
      RECT 13.111 4.553 13.197 5.22 ;
      RECT 13.025 4.551 13.111 5.22 ;
      RECT 13.015 4.552 13.025 5.22 ;
      RECT 13.01 4.557 13.015 5.22 ;
      RECT 13 4.57 13.01 5.22 ;
      RECT 12.995 4.592 13 5.22 ;
      RECT 12.99 4.952 12.995 5.22 ;
      RECT 13.62 4.42 13.625 4.64 ;
      RECT 14.125 3.455 14.16 3.715 ;
      RECT 14.11 3.455 14.125 3.723 ;
      RECT 14.081 3.455 14.11 3.745 ;
      RECT 13.995 3.455 14.081 3.805 ;
      RECT 13.975 3.455 13.995 3.87 ;
      RECT 13.915 3.455 13.975 4.035 ;
      RECT 13.91 3.455 13.915 4.183 ;
      RECT 13.905 3.455 13.91 4.195 ;
      RECT 13.9 3.455 13.905 4.221 ;
      RECT 13.87 3.641 13.9 4.301 ;
      RECT 13.865 3.689 13.87 4.39 ;
      RECT 13.86 3.703 13.865 4.405 ;
      RECT 13.855 3.722 13.86 4.435 ;
      RECT 13.85 3.737 13.855 4.451 ;
      RECT 13.845 3.752 13.85 4.473 ;
      RECT 13.84 3.772 13.845 4.495 ;
      RECT 13.83 3.792 13.84 4.528 ;
      RECT 13.815 3.834 13.83 4.59 ;
      RECT 13.81 3.865 13.815 4.63 ;
      RECT 13.805 3.877 13.81 4.635 ;
      RECT 13.8 3.889 13.805 4.64 ;
      RECT 13.795 3.902 13.8 4.64 ;
      RECT 13.79 3.92 13.795 4.64 ;
      RECT 13.785 3.94 13.79 4.64 ;
      RECT 13.78 3.952 13.785 4.64 ;
      RECT 13.775 3.965 13.78 4.64 ;
      RECT 13.755 4 13.775 4.64 ;
      RECT 13.705 4.102 13.755 4.64 ;
      RECT 13.7 4.187 13.705 4.64 ;
      RECT 13.695 4.195 13.7 4.64 ;
      RECT 13.69 4.212 13.695 4.64 ;
      RECT 13.685 4.227 13.69 4.64 ;
      RECT 13.65 4.292 13.685 4.64 ;
      RECT 13.635 4.357 13.65 4.64 ;
      RECT 13.63 4.387 13.635 4.64 ;
      RECT 13.625 4.412 13.63 4.64 ;
      RECT 13.61 4.422 13.62 4.64 ;
      RECT 13.595 4.435 13.61 4.633 ;
      RECT 13.34 4.025 13.41 4.235 ;
      RECT 13.13 4.002 13.135 4.195 ;
      RECT 10.585 3.93 10.845 4.19 ;
      RECT 13.42 4.212 13.425 4.215 ;
      RECT 13.41 4.03 13.42 4.23 ;
      RECT 13.311 4.023 13.34 4.235 ;
      RECT 13.225 4.015 13.311 4.235 ;
      RECT 13.21 4.009 13.225 4.233 ;
      RECT 13.19 4.008 13.21 4.22 ;
      RECT 13.185 4.007 13.19 4.203 ;
      RECT 13.135 4.004 13.185 4.198 ;
      RECT 13.105 4.001 13.13 4.193 ;
      RECT 13.085 3.999 13.105 4.188 ;
      RECT 13.07 3.997 13.085 4.185 ;
      RECT 13.04 3.995 13.07 4.183 ;
      RECT 12.975 3.991 13.04 4.175 ;
      RECT 12.945 3.986 12.975 4.17 ;
      RECT 12.925 3.984 12.945 4.168 ;
      RECT 12.895 3.981 12.925 4.163 ;
      RECT 12.835 3.977 12.895 4.155 ;
      RECT 12.83 3.974 12.835 4.15 ;
      RECT 12.76 3.972 12.83 4.145 ;
      RECT 12.731 3.968 12.76 4.138 ;
      RECT 12.645 3.963 12.731 4.13 ;
      RECT 12.611 3.958 12.645 4.122 ;
      RECT 12.525 3.95 12.611 4.114 ;
      RECT 12.486 3.943 12.525 4.106 ;
      RECT 12.4 3.938 12.486 4.098 ;
      RECT 12.335 3.932 12.4 4.088 ;
      RECT 12.315 3.927 12.335 4.083 ;
      RECT 12.306 3.924 12.315 4.082 ;
      RECT 12.22 3.92 12.306 4.076 ;
      RECT 12.18 3.916 12.22 4.068 ;
      RECT 12.16 3.912 12.18 4.066 ;
      RECT 12.1 3.912 12.16 4.063 ;
      RECT 12.08 3.915 12.1 4.061 ;
      RECT 12.059 3.915 12.08 4.061 ;
      RECT 11.973 3.917 12.059 4.065 ;
      RECT 11.887 3.919 11.973 4.071 ;
      RECT 11.801 3.921 11.887 4.078 ;
      RECT 11.715 3.924 11.801 4.084 ;
      RECT 11.681 3.925 11.715 4.089 ;
      RECT 11.595 3.928 11.681 4.094 ;
      RECT 11.566 3.935 11.595 4.099 ;
      RECT 11.48 3.935 11.566 4.104 ;
      RECT 11.447 3.935 11.48 4.109 ;
      RECT 11.361 3.937 11.447 4.114 ;
      RECT 11.275 3.939 11.361 4.121 ;
      RECT 11.211 3.941 11.275 4.127 ;
      RECT 11.125 3.943 11.211 4.133 ;
      RECT 11.122 3.945 11.125 4.136 ;
      RECT 11.036 3.946 11.122 4.14 ;
      RECT 10.95 3.949 11.036 4.147 ;
      RECT 10.931 3.951 10.95 4.151 ;
      RECT 10.845 3.953 10.931 4.156 ;
      RECT 10.575 3.965 10.585 4.16 ;
      RECT 12.755 10.2 13.045 10.43 ;
      RECT 12.815 9.46 12.985 10.43 ;
      RECT 12.705 9.49 13.08 9.86 ;
      RECT 12.755 9.46 13.045 9.86 ;
      RECT 12.81 3.545 12.995 3.755 ;
      RECT 12.805 3.546 13 3.753 ;
      RECT 12.8 3.551 13.01 3.748 ;
      RECT 12.795 3.527 12.8 3.745 ;
      RECT 12.765 3.524 12.795 3.738 ;
      RECT 12.76 3.52 12.765 3.729 ;
      RECT 12.725 3.551 13.01 3.724 ;
      RECT 12.5 3.46 12.76 3.72 ;
      RECT 12.8 3.529 12.805 3.748 ;
      RECT 12.805 3.53 12.81 3.753 ;
      RECT 12.5 3.542 12.88 3.72 ;
      RECT 12.5 3.54 12.865 3.72 ;
      RECT 12.5 3.535 12.855 3.72 ;
      RECT 12.455 4.45 12.505 4.735 ;
      RECT 12.4 4.42 12.405 4.735 ;
      RECT 12.37 4.4 12.375 4.735 ;
      RECT 12.52 4.45 12.58 4.71 ;
      RECT 12.515 4.45 12.52 4.718 ;
      RECT 12.505 4.45 12.515 4.73 ;
      RECT 12.42 4.44 12.455 4.735 ;
      RECT 12.415 4.427 12.42 4.735 ;
      RECT 12.405 4.422 12.415 4.735 ;
      RECT 12.385 4.412 12.4 4.735 ;
      RECT 12.375 4.405 12.385 4.735 ;
      RECT 12.365 4.397 12.37 4.735 ;
      RECT 12.335 4.387 12.365 4.735 ;
      RECT 12.32 4.375 12.335 4.735 ;
      RECT 12.305 4.365 12.32 4.73 ;
      RECT 12.285 4.355 12.305 4.705 ;
      RECT 12.275 4.347 12.285 4.682 ;
      RECT 12.245 4.33 12.275 4.672 ;
      RECT 12.24 4.307 12.245 4.663 ;
      RECT 12.235 4.294 12.24 4.661 ;
      RECT 12.22 4.27 12.235 4.655 ;
      RECT 12.215 4.246 12.22 4.649 ;
      RECT 12.205 4.235 12.215 4.644 ;
      RECT 12.2 4.225 12.205 4.64 ;
      RECT 12.195 4.217 12.2 4.637 ;
      RECT 12.185 4.212 12.195 4.633 ;
      RECT 12.18 4.207 12.185 4.629 ;
      RECT 12.095 4.205 12.18 4.604 ;
      RECT 12.065 4.205 12.095 4.57 ;
      RECT 12.05 4.205 12.065 4.553 ;
      RECT 11.995 4.205 12.05 4.498 ;
      RECT 11.99 4.21 11.995 4.447 ;
      RECT 11.98 4.215 11.99 4.437 ;
      RECT 11.975 4.225 11.98 4.423 ;
      RECT 11.925 4.965 12.185 5.225 ;
      RECT 11.845 4.98 12.185 5.201 ;
      RECT 11.825 4.98 12.185 5.196 ;
      RECT 11.801 4.98 12.185 5.194 ;
      RECT 11.715 4.98 12.185 5.189 ;
      RECT 11.565 4.92 11.825 5.185 ;
      RECT 11.52 4.98 12.185 5.18 ;
      RECT 11.515 4.987 12.185 5.175 ;
      RECT 11.53 4.975 11.845 5.185 ;
      RECT 11.42 3.41 11.68 3.67 ;
      RECT 11.42 3.467 11.685 3.663 ;
      RECT 11.42 3.497 11.69 3.595 ;
      RECT 11.48 3.928 11.595 3.93 ;
      RECT 11.566 3.925 11.595 3.93 ;
      RECT 10.59 4.929 10.615 5.169 ;
      RECT 10.575 4.932 10.665 5.163 ;
      RECT 10.57 4.937 10.751 5.158 ;
      RECT 10.565 4.945 10.815 5.156 ;
      RECT 10.565 4.945 10.825 5.155 ;
      RECT 10.56 4.952 10.835 5.148 ;
      RECT 10.56 4.952 10.921 5.137 ;
      RECT 10.555 4.987 10.921 5.133 ;
      RECT 10.555 4.987 10.93 5.122 ;
      RECT 10.835 4.86 11.095 5.12 ;
      RECT 10.545 5.037 11.095 5.118 ;
      RECT 10.815 4.905 10.835 5.153 ;
      RECT 10.751 4.908 10.815 5.157 ;
      RECT 10.665 4.913 10.751 5.162 ;
      RECT 10.595 4.924 11.095 5.12 ;
      RECT 10.615 4.918 10.665 5.167 ;
      RECT 10.74 3.395 10.75 3.657 ;
      RECT 10.73 3.452 10.74 3.66 ;
      RECT 10.705 3.457 10.73 3.666 ;
      RECT 10.68 3.461 10.705 3.678 ;
      RECT 10.67 3.464 10.68 3.688 ;
      RECT 10.665 3.465 10.67 3.693 ;
      RECT 10.66 3.466 10.665 3.698 ;
      RECT 10.655 3.467 10.66 3.7 ;
      RECT 10.63 3.47 10.655 3.703 ;
      RECT 10.6 3.476 10.63 3.706 ;
      RECT 10.535 3.487 10.6 3.709 ;
      RECT 10.49 3.495 10.535 3.713 ;
      RECT 10.475 3.495 10.49 3.721 ;
      RECT 10.47 3.496 10.475 3.728 ;
      RECT 10.465 3.498 10.47 3.731 ;
      RECT 10.46 3.502 10.465 3.734 ;
      RECT 10.45 3.51 10.46 3.738 ;
      RECT 10.445 3.523 10.45 3.743 ;
      RECT 10.44 3.531 10.445 3.745 ;
      RECT 10.435 3.537 10.44 3.745 ;
      RECT 10.43 3.541 10.435 3.748 ;
      RECT 10.425 3.543 10.43 3.751 ;
      RECT 10.42 3.546 10.425 3.754 ;
      RECT 10.41 3.551 10.42 3.758 ;
      RECT 10.405 3.557 10.41 3.763 ;
      RECT 10.395 3.563 10.405 3.767 ;
      RECT 10.38 3.57 10.395 3.773 ;
      RECT 10.351 3.584 10.38 3.783 ;
      RECT 10.265 3.619 10.351 3.815 ;
      RECT 10.245 3.652 10.265 3.844 ;
      RECT 10.225 3.665 10.245 3.855 ;
      RECT 10.205 3.677 10.225 3.866 ;
      RECT 10.155 3.699 10.205 3.886 ;
      RECT 10.14 3.717 10.155 3.903 ;
      RECT 10.135 3.723 10.14 3.906 ;
      RECT 10.13 3.727 10.135 3.909 ;
      RECT 10.125 3.731 10.13 3.913 ;
      RECT 10.12 3.733 10.125 3.916 ;
      RECT 10.11 3.74 10.12 3.919 ;
      RECT 10.105 3.745 10.11 3.923 ;
      RECT 10.1 3.747 10.105 3.926 ;
      RECT 10.095 3.751 10.1 3.929 ;
      RECT 10.09 3.753 10.095 3.933 ;
      RECT 10.075 3.758 10.09 3.938 ;
      RECT 10.07 3.763 10.075 3.941 ;
      RECT 10.065 3.771 10.07 3.944 ;
      RECT 10.06 3.773 10.065 3.947 ;
      RECT 10.055 3.775 10.06 3.95 ;
      RECT 10.045 3.777 10.055 3.956 ;
      RECT 10.01 3.791 10.045 3.968 ;
      RECT 10 3.806 10.01 3.978 ;
      RECT 9.925 3.835 10 4.002 ;
      RECT 9.92 3.86 9.925 4.025 ;
      RECT 9.905 3.864 9.92 4.031 ;
      RECT 9.895 3.872 9.905 4.036 ;
      RECT 9.865 3.885 9.895 4.04 ;
      RECT 9.855 3.9 9.865 4.045 ;
      RECT 9.845 3.905 9.855 4.048 ;
      RECT 9.84 3.907 9.845 4.05 ;
      RECT 9.825 3.91 9.84 4.053 ;
      RECT 9.82 3.912 9.825 4.056 ;
      RECT 9.8 3.917 9.82 4.06 ;
      RECT 9.77 3.922 9.8 4.068 ;
      RECT 9.745 3.929 9.77 4.076 ;
      RECT 9.74 3.934 9.745 4.081 ;
      RECT 9.71 3.937 9.74 4.085 ;
      RECT 9.67 3.94 9.71 4.095 ;
      RECT 9.635 3.937 9.67 4.107 ;
      RECT 9.625 3.933 9.635 4.114 ;
      RECT 9.6 3.929 9.625 4.12 ;
      RECT 9.595 3.925 9.6 4.125 ;
      RECT 9.555 3.922 9.595 4.125 ;
      RECT 9.54 3.907 9.555 4.126 ;
      RECT 9.517 3.895 9.54 4.126 ;
      RECT 9.431 3.895 9.517 4.127 ;
      RECT 9.345 3.895 9.431 4.129 ;
      RECT 9.325 3.895 9.345 4.126 ;
      RECT 9.32 3.9 9.325 4.121 ;
      RECT 9.315 3.905 9.32 4.119 ;
      RECT 9.305 3.915 9.315 4.117 ;
      RECT 9.3 3.921 9.305 4.11 ;
      RECT 9.295 3.923 9.3 4.095 ;
      RECT 9.29 3.927 9.295 4.085 ;
      RECT 10.75 3.395 11 3.655 ;
      RECT 8.475 4.93 8.735 5.19 ;
      RECT 10.77 4.42 10.775 4.63 ;
      RECT 10.775 4.425 10.785 4.625 ;
      RECT 10.725 4.42 10.77 4.645 ;
      RECT 10.715 4.42 10.725 4.665 ;
      RECT 10.696 4.42 10.715 4.67 ;
      RECT 10.61 4.42 10.696 4.667 ;
      RECT 10.58 4.422 10.61 4.665 ;
      RECT 10.525 4.432 10.58 4.663 ;
      RECT 10.46 4.446 10.525 4.661 ;
      RECT 10.455 4.454 10.46 4.66 ;
      RECT 10.44 4.457 10.455 4.658 ;
      RECT 10.375 4.467 10.44 4.654 ;
      RECT 10.327 4.481 10.375 4.655 ;
      RECT 10.241 4.498 10.327 4.669 ;
      RECT 10.155 4.519 10.241 4.686 ;
      RECT 10.135 4.532 10.155 4.696 ;
      RECT 10.09 4.54 10.135 4.703 ;
      RECT 10.055 4.548 10.09 4.711 ;
      RECT 10.021 4.556 10.055 4.719 ;
      RECT 9.935 4.57 10.021 4.731 ;
      RECT 9.9 4.587 9.935 4.743 ;
      RECT 9.891 4.596 9.9 4.747 ;
      RECT 9.805 4.614 9.891 4.764 ;
      RECT 9.746 4.641 9.805 4.791 ;
      RECT 9.66 4.668 9.746 4.819 ;
      RECT 9.64 4.69 9.66 4.839 ;
      RECT 9.58 4.705 9.64 4.855 ;
      RECT 9.57 4.717 9.58 4.868 ;
      RECT 9.565 4.722 9.57 4.871 ;
      RECT 9.555 4.725 9.565 4.874 ;
      RECT 9.55 4.727 9.555 4.877 ;
      RECT 9.52 4.735 9.55 4.884 ;
      RECT 9.505 4.742 9.52 4.892 ;
      RECT 9.495 4.747 9.505 4.896 ;
      RECT 9.49 4.75 9.495 4.899 ;
      RECT 9.48 4.752 9.49 4.902 ;
      RECT 9.445 4.762 9.48 4.911 ;
      RECT 9.37 4.785 9.445 4.933 ;
      RECT 9.35 4.803 9.37 4.951 ;
      RECT 9.32 4.81 9.35 4.961 ;
      RECT 9.3 4.818 9.32 4.971 ;
      RECT 9.29 4.824 9.3 4.978 ;
      RECT 9.271 4.829 9.29 4.984 ;
      RECT 9.185 4.849 9.271 5.004 ;
      RECT 9.17 4.869 9.185 5.023 ;
      RECT 9.125 4.881 9.17 5.034 ;
      RECT 9.06 4.902 9.125 5.057 ;
      RECT 9.02 4.922 9.06 5.078 ;
      RECT 9.01 4.932 9.02 5.088 ;
      RECT 8.96 4.944 9.01 5.099 ;
      RECT 8.94 4.96 8.96 5.111 ;
      RECT 8.91 4.97 8.94 5.117 ;
      RECT 8.9 4.975 8.91 5.119 ;
      RECT 8.831 4.976 8.9 5.125 ;
      RECT 8.745 4.978 8.831 5.135 ;
      RECT 8.735 4.979 8.745 5.14 ;
      RECT 10.005 5.005 10.195 5.215 ;
      RECT 9.995 5.01 10.205 5.208 ;
      RECT 9.98 5.01 10.205 5.173 ;
      RECT 9.9 4.895 10.16 5.155 ;
      RECT 8.815 4.425 9 4.72 ;
      RECT 8.805 4.425 9 4.718 ;
      RECT 8.79 4.425 9.005 4.713 ;
      RECT 8.79 4.425 9.01 4.71 ;
      RECT 8.785 4.425 9.01 4.708 ;
      RECT 8.78 4.68 9.01 4.698 ;
      RECT 8.785 4.425 9.045 4.685 ;
      RECT 8.745 3.46 9.005 3.72 ;
      RECT 8.555 3.385 8.641 3.718 ;
      RECT 8.53 3.389 8.685 3.714 ;
      RECT 8.641 3.381 8.685 3.714 ;
      RECT 8.641 3.382 8.69 3.713 ;
      RECT 8.555 3.387 8.705 3.712 ;
      RECT 8.53 3.395 8.745 3.711 ;
      RECT 8.525 3.39 8.705 3.706 ;
      RECT 8.515 3.405 8.745 3.613 ;
      RECT 8.515 3.457 8.945 3.613 ;
      RECT 8.515 3.45 8.925 3.613 ;
      RECT 8.515 3.437 8.895 3.613 ;
      RECT 8.515 3.425 8.835 3.613 ;
      RECT 8.515 3.41 8.81 3.613 ;
      RECT 7.715 4.04 7.85 4.335 ;
      RECT 7.975 4.063 7.98 4.25 ;
      RECT 8.695 3.96 8.84 4.195 ;
      RECT 8.855 3.96 8.86 4.185 ;
      RECT 8.89 3.971 8.895 4.165 ;
      RECT 8.885 3.963 8.89 4.17 ;
      RECT 8.865 3.96 8.885 4.175 ;
      RECT 8.86 3.96 8.865 4.183 ;
      RECT 8.85 3.96 8.855 4.188 ;
      RECT 8.84 3.96 8.85 4.193 ;
      RECT 8.67 3.962 8.695 4.195 ;
      RECT 8.62 3.969 8.67 4.195 ;
      RECT 8.615 3.974 8.62 4.195 ;
      RECT 8.576 3.979 8.615 4.196 ;
      RECT 8.49 3.991 8.576 4.197 ;
      RECT 8.481 4.001 8.49 4.197 ;
      RECT 8.395 4.01 8.481 4.199 ;
      RECT 8.371 4.02 8.395 4.201 ;
      RECT 8.285 4.031 8.371 4.202 ;
      RECT 8.255 4.042 8.285 4.204 ;
      RECT 8.225 4.047 8.255 4.206 ;
      RECT 8.2 4.053 8.225 4.209 ;
      RECT 8.185 4.058 8.2 4.21 ;
      RECT 8.14 4.064 8.185 4.21 ;
      RECT 8.135 4.069 8.14 4.211 ;
      RECT 8.115 4.069 8.135 4.213 ;
      RECT 8.095 4.067 8.115 4.218 ;
      RECT 8.06 4.066 8.095 4.225 ;
      RECT 8.03 4.065 8.06 4.235 ;
      RECT 7.98 4.064 8.03 4.245 ;
      RECT 7.89 4.061 7.975 4.335 ;
      RECT 7.865 4.055 7.89 4.335 ;
      RECT 7.85 4.045 7.865 4.335 ;
      RECT 7.665 4.04 7.715 4.255 ;
      RECT 7.655 4.045 7.665 4.245 ;
      RECT 7.895 4.52 8.155 4.78 ;
      RECT 7.895 4.52 8.185 4.673 ;
      RECT 7.895 4.52 8.22 4.658 ;
      RECT 8.15 4.44 8.34 4.65 ;
      RECT 8.14 4.445 8.35 4.643 ;
      RECT 8.105 4.515 8.35 4.643 ;
      RECT 8.135 4.457 8.155 4.78 ;
      RECT 8.12 4.505 8.35 4.643 ;
      RECT 8.125 4.477 8.155 4.78 ;
      RECT 7.205 3.545 7.275 4.65 ;
      RECT 7.94 3.65 8.2 3.91 ;
      RECT 7.52 3.696 7.535 3.905 ;
      RECT 7.856 3.709 7.94 3.86 ;
      RECT 7.77 3.706 7.856 3.86 ;
      RECT 7.731 3.704 7.77 3.86 ;
      RECT 7.645 3.702 7.731 3.86 ;
      RECT 7.585 3.7 7.645 3.871 ;
      RECT 7.55 3.698 7.585 3.889 ;
      RECT 7.535 3.696 7.55 3.9 ;
      RECT 7.505 3.696 7.52 3.913 ;
      RECT 7.495 3.696 7.505 3.918 ;
      RECT 7.47 3.695 7.495 3.923 ;
      RECT 7.455 3.69 7.47 3.929 ;
      RECT 7.45 3.683 7.455 3.934 ;
      RECT 7.425 3.674 7.45 3.94 ;
      RECT 7.38 3.653 7.425 3.953 ;
      RECT 7.37 3.637 7.38 3.963 ;
      RECT 7.355 3.63 7.37 3.973 ;
      RECT 7.345 3.623 7.355 3.99 ;
      RECT 7.34 3.62 7.345 4.02 ;
      RECT 7.335 3.618 7.34 4.05 ;
      RECT 7.33 3.616 7.335 4.087 ;
      RECT 7.315 3.612 7.33 4.154 ;
      RECT 7.315 4.445 7.325 4.645 ;
      RECT 7.31 3.608 7.315 4.28 ;
      RECT 7.31 4.432 7.315 4.65 ;
      RECT 7.305 3.606 7.31 4.365 ;
      RECT 7.305 4.422 7.31 4.65 ;
      RECT 7.29 3.577 7.305 4.65 ;
      RECT 7.275 3.55 7.29 4.65 ;
      RECT 7.2 3.545 7.205 3.9 ;
      RECT 7.2 3.955 7.205 4.65 ;
      RECT 7.185 3.545 7.2 3.878 ;
      RECT 7.195 3.977 7.2 4.65 ;
      RECT 7.185 4.017 7.195 4.65 ;
      RECT 7.15 3.545 7.185 3.82 ;
      RECT 7.18 4.052 7.185 4.65 ;
      RECT 7.165 4.107 7.18 4.65 ;
      RECT 7.16 4.172 7.165 4.65 ;
      RECT 7.145 4.22 7.16 4.65 ;
      RECT 7.12 3.545 7.15 3.775 ;
      RECT 7.14 4.275 7.145 4.65 ;
      RECT 7.125 4.335 7.14 4.65 ;
      RECT 7.12 4.383 7.125 4.648 ;
      RECT 7.115 3.545 7.12 3.768 ;
      RECT 7.115 4.415 7.12 4.643 ;
      RECT 7.09 3.545 7.115 3.76 ;
      RECT 7.08 3.55 7.09 3.75 ;
      RECT 7.295 4.825 7.315 5.065 ;
      RECT 6.525 4.755 6.53 4.965 ;
      RECT 7.805 4.828 7.815 5.023 ;
      RECT 7.8 4.818 7.805 5.026 ;
      RECT 7.72 4.815 7.8 5.049 ;
      RECT 7.716 4.815 7.72 5.071 ;
      RECT 7.63 4.815 7.716 5.081 ;
      RECT 7.615 4.815 7.63 5.089 ;
      RECT 7.586 4.816 7.615 5.087 ;
      RECT 7.5 4.821 7.586 5.083 ;
      RECT 7.487 4.825 7.5 5.079 ;
      RECT 7.401 4.825 7.487 5.075 ;
      RECT 7.315 4.825 7.401 5.069 ;
      RECT 7.231 4.825 7.295 5.063 ;
      RECT 7.145 4.825 7.231 5.058 ;
      RECT 7.125 4.825 7.145 5.054 ;
      RECT 7.065 4.82 7.125 5.051 ;
      RECT 7.037 4.814 7.065 5.048 ;
      RECT 6.951 4.809 7.037 5.044 ;
      RECT 6.865 4.803 6.951 5.038 ;
      RECT 6.79 4.785 6.865 5.033 ;
      RECT 6.755 4.762 6.79 5.029 ;
      RECT 6.745 4.752 6.755 5.028 ;
      RECT 6.69 4.75 6.745 5.027 ;
      RECT 6.615 4.75 6.69 5.023 ;
      RECT 6.605 4.75 6.615 5.018 ;
      RECT 6.59 4.75 6.605 5.01 ;
      RECT 6.54 4.752 6.59 4.988 ;
      RECT 6.53 4.755 6.54 4.968 ;
      RECT 6.52 4.76 6.525 4.963 ;
      RECT 6.515 4.765 6.52 4.958 ;
      RECT 6.64 3.93 6.9 4.19 ;
      RECT 6.64 3.945 6.92 4.155 ;
      RECT 6.64 3.95 6.93 4.15 ;
      RECT 4.625 3.41 4.885 3.67 ;
      RECT 4.615 3.44 4.885 3.65 ;
      RECT 6.535 3.355 6.795 3.615 ;
      RECT 6.53 3.43 6.535 3.616 ;
      RECT 6.505 3.435 6.53 3.618 ;
      RECT 6.49 3.442 6.505 3.621 ;
      RECT 6.43 3.46 6.49 3.626 ;
      RECT 6.4 3.48 6.43 3.633 ;
      RECT 6.375 3.488 6.4 3.638 ;
      RECT 6.35 3.496 6.375 3.64 ;
      RECT 6.332 3.5 6.35 3.639 ;
      RECT 6.246 3.498 6.332 3.639 ;
      RECT 6.16 3.496 6.246 3.639 ;
      RECT 6.074 3.494 6.16 3.638 ;
      RECT 5.988 3.492 6.074 3.638 ;
      RECT 5.902 3.49 5.988 3.638 ;
      RECT 5.816 3.488 5.902 3.638 ;
      RECT 5.73 3.486 5.816 3.637 ;
      RECT 5.712 3.485 5.73 3.637 ;
      RECT 5.626 3.484 5.712 3.637 ;
      RECT 5.54 3.482 5.626 3.637 ;
      RECT 5.454 3.481 5.54 3.636 ;
      RECT 5.368 3.48 5.454 3.636 ;
      RECT 5.282 3.478 5.368 3.636 ;
      RECT 5.196 3.477 5.282 3.636 ;
      RECT 5.11 3.475 5.196 3.635 ;
      RECT 5.086 3.473 5.11 3.635 ;
      RECT 5 3.466 5.086 3.635 ;
      RECT 4.971 3.458 5 3.635 ;
      RECT 4.885 3.45 4.971 3.635 ;
      RECT 4.605 3.447 4.615 3.645 ;
      RECT 6.11 4.41 6.115 4.76 ;
      RECT 5.88 4.5 6.02 4.76 ;
      RECT 6.355 4.185 6.4 4.395 ;
      RECT 6.41 4.196 6.42 4.39 ;
      RECT 6.4 4.188 6.41 4.395 ;
      RECT 6.335 4.185 6.355 4.4 ;
      RECT 6.305 4.185 6.335 4.423 ;
      RECT 6.295 4.185 6.305 4.448 ;
      RECT 6.29 4.185 6.295 4.458 ;
      RECT 6.235 4.185 6.29 4.498 ;
      RECT 6.23 4.185 6.235 4.538 ;
      RECT 6.225 4.187 6.23 4.543 ;
      RECT 6.21 4.197 6.225 4.554 ;
      RECT 6.165 4.255 6.21 4.59 ;
      RECT 6.155 4.31 6.165 4.624 ;
      RECT 6.14 4.337 6.155 4.64 ;
      RECT 6.13 4.364 6.14 4.76 ;
      RECT 6.115 4.387 6.13 4.76 ;
      RECT 6.105 4.427 6.11 4.76 ;
      RECT 6.1 4.437 6.105 4.76 ;
      RECT 6.095 4.452 6.1 4.76 ;
      RECT 6.085 4.457 6.095 4.76 ;
      RECT 6.02 4.48 6.085 4.76 ;
      RECT 5.52 3.975 5.71 4.185 ;
      RECT 4.095 3.9 4.355 4.16 ;
      RECT 4.445 3.895 4.54 4.105 ;
      RECT 4.42 3.91 4.43 4.105 ;
      RECT 5.71 3.982 5.72 4.18 ;
      RECT 5.51 3.982 5.52 4.18 ;
      RECT 5.495 3.997 5.51 4.17 ;
      RECT 5.49 4.005 5.495 4.163 ;
      RECT 5.48 4.008 5.49 4.16 ;
      RECT 5.445 4.007 5.48 4.158 ;
      RECT 5.416 4.003 5.445 4.155 ;
      RECT 5.33 3.998 5.416 4.152 ;
      RECT 5.27 3.992 5.33 4.148 ;
      RECT 5.241 3.988 5.27 4.145 ;
      RECT 5.155 3.98 5.241 4.142 ;
      RECT 5.146 3.974 5.155 4.14 ;
      RECT 5.06 3.969 5.146 4.138 ;
      RECT 5.037 3.964 5.06 4.135 ;
      RECT 4.951 3.958 5.037 4.132 ;
      RECT 4.865 3.949 4.951 4.127 ;
      RECT 4.855 3.944 4.865 4.125 ;
      RECT 4.836 3.943 4.855 4.124 ;
      RECT 4.75 3.938 4.836 4.12 ;
      RECT 4.73 3.933 4.75 4.116 ;
      RECT 4.67 3.928 4.73 4.113 ;
      RECT 4.645 3.918 4.67 4.111 ;
      RECT 4.64 3.911 4.645 4.11 ;
      RECT 4.63 3.902 4.64 4.109 ;
      RECT 4.626 3.895 4.63 4.109 ;
      RECT 4.54 3.895 4.626 4.107 ;
      RECT 4.43 3.902 4.445 4.105 ;
      RECT 4.415 3.912 4.42 4.105 ;
      RECT 4.395 3.915 4.415 4.102 ;
      RECT 4.365 3.915 4.395 4.098 ;
      RECT 4.355 3.915 4.365 4.098 ;
      RECT 5.27 4.41 5.53 4.67 ;
      RECT 5.2 4.42 5.53 4.63 ;
      RECT 5.19 4.427 5.53 4.625 ;
      RECT 4.61 4.415 4.87 4.675 ;
      RECT 4.61 4.455 4.975 4.665 ;
      RECT 4.61 4.457 4.98 4.664 ;
      RECT 4.61 4.465 4.985 4.661 ;
      RECT 3.535 3.54 3.635 5.065 ;
      RECT 3.725 4.68 3.775 4.94 ;
      RECT 3.72 3.553 3.725 3.74 ;
      RECT 3.715 4.661 3.725 4.94 ;
      RECT 3.715 3.55 3.72 3.748 ;
      RECT 3.7 3.544 3.715 3.755 ;
      RECT 3.71 4.649 3.715 5.023 ;
      RECT 3.7 4.637 3.71 5.06 ;
      RECT 3.69 3.54 3.7 3.762 ;
      RECT 3.69 4.622 3.7 5.065 ;
      RECT 3.685 3.54 3.69 3.77 ;
      RECT 3.665 4.592 3.69 5.065 ;
      RECT 3.645 3.54 3.685 3.818 ;
      RECT 3.655 4.552 3.665 5.065 ;
      RECT 3.645 4.507 3.655 5.065 ;
      RECT 3.64 3.54 3.645 3.888 ;
      RECT 3.64 4.465 3.645 5.065 ;
      RECT 3.635 3.54 3.64 4.365 ;
      RECT 3.635 4.447 3.64 5.065 ;
      RECT 3.525 3.543 3.535 5.065 ;
      RECT 3.51 3.55 3.525 5.061 ;
      RECT 3.505 3.56 3.51 5.056 ;
      RECT 3.5 3.76 3.505 4.948 ;
      RECT 3.495 3.845 3.5 4.5 ;
      RECT 1.725 10.2 2.015 10.43 ;
      RECT 1.785 9.46 1.955 10.43 ;
      RECT 1.695 9.46 2.045 9.75 ;
      RECT 1.32 8.72 1.67 9.01 ;
      RECT 1.18 8.75 1.67 8.92 ;
      RECT 87.225 2.435 87.6 2.805 ;
      RECT 81.205 3.52 81.465 3.78 ;
      RECT 69.3 2.435 69.675 2.805 ;
      RECT 63.28 3.52 63.54 3.78 ;
      RECT 51.375 2.435 51.75 2.805 ;
      RECT 45.355 3.52 45.615 3.78 ;
      RECT 33.45 2.435 33.825 2.805 ;
      RECT 27.43 3.52 27.69 3.78 ;
      RECT 9.505 3.52 9.765 3.78 ;
    LAYER mcon ;
      RECT 92.055 8.755 92.225 8.925 ;
      RECT 92.055 10.235 92.225 10.405 ;
      RECT 91.705 1.395 91.875 1.565 ;
      RECT 91.685 4.055 91.855 4.225 ;
      RECT 91.685 8.385 91.855 8.555 ;
      RECT 91.065 2.205 91.235 2.375 ;
      RECT 91.065 3.685 91.235 3.855 ;
      RECT 91.065 8.755 91.235 8.925 ;
      RECT 91.065 10.235 91.235 10.405 ;
      RECT 90.715 1.395 90.885 1.565 ;
      RECT 90.695 4.055 90.865 4.225 ;
      RECT 90.695 8.385 90.865 8.555 ;
      RECT 90.015 1.4 90.185 1.57 ;
      RECT 89.705 3.32 89.875 3.49 ;
      RECT 89.705 9.12 89.875 9.29 ;
      RECT 89.335 1.4 89.505 1.57 ;
      RECT 89.275 2.21 89.445 2.38 ;
      RECT 89.275 2.95 89.445 3.12 ;
      RECT 89.275 9.49 89.445 9.66 ;
      RECT 89.275 10.23 89.445 10.4 ;
      RECT 88.9 3.69 89.07 3.86 ;
      RECT 88.9 8.75 89.07 8.92 ;
      RECT 88.655 1.4 88.825 1.57 ;
      RECT 87.975 1.4 88.145 1.57 ;
      RECT 86.695 2.86 86.865 3.03 ;
      RECT 86.235 2.86 86.405 3.03 ;
      RECT 85.84 4.2 86.01 4.37 ;
      RECT 85.775 2.86 85.945 3.03 ;
      RECT 85.63 3.54 85.8 3.71 ;
      RECT 85.315 2.86 85.485 3.03 ;
      RECT 85.315 4.45 85.485 4.62 ;
      RECT 84.945 9.12 85.115 9.29 ;
      RECT 84.93 4.045 85.1 4.215 ;
      RECT 84.855 2.86 85.025 3.03 ;
      RECT 84.715 4.61 84.885 4.78 ;
      RECT 84.695 5.01 84.865 5.18 ;
      RECT 84.52 3.565 84.69 3.735 ;
      RECT 84.515 9.49 84.685 9.66 ;
      RECT 84.515 10.23 84.685 10.4 ;
      RECT 84.395 2.86 84.565 3.03 ;
      RECT 84.025 4.545 84.195 4.715 ;
      RECT 83.935 2.86 84.105 3.03 ;
      RECT 83.7 4.23 83.87 4.4 ;
      RECT 83.635 5.01 83.805 5.18 ;
      RECT 83.475 2.86 83.645 3.03 ;
      RECT 83.235 4.995 83.405 5.165 ;
      RECT 83.195 3.48 83.365 3.65 ;
      RECT 83.015 2.86 83.185 3.03 ;
      RECT 82.555 2.86 82.725 3.03 ;
      RECT 82.295 3.98 82.465 4.15 ;
      RECT 82.295 4.44 82.465 4.61 ;
      RECT 82.295 4.955 82.465 5.125 ;
      RECT 82.18 3.515 82.35 3.685 ;
      RECT 82.095 2.86 82.265 3.03 ;
      RECT 81.715 5.025 81.885 5.195 ;
      RECT 81.635 2.86 81.805 3.03 ;
      RECT 81.235 3.555 81.405 3.725 ;
      RECT 81.175 2.86 81.345 3.03 ;
      RECT 81.02 3.93 81.19 4.1 ;
      RECT 80.715 2.86 80.885 3.03 ;
      RECT 80.52 4.53 80.69 4.7 ;
      RECT 80.405 3.98 80.575 4.15 ;
      RECT 80.255 2.86 80.425 3.03 ;
      RECT 80.235 3.43 80.405 3.6 ;
      RECT 79.86 4.46 80.03 4.63 ;
      RECT 79.795 2.86 79.965 3.03 ;
      RECT 79.375 4.06 79.545 4.23 ;
      RECT 79.335 2.86 79.505 3.03 ;
      RECT 79.325 4.835 79.495 5.005 ;
      RECT 78.875 2.86 79.045 3.03 ;
      RECT 78.835 4.46 79.005 4.63 ;
      RECT 78.8 3.565 78.97 3.735 ;
      RECT 78.44 3.965 78.61 4.135 ;
      RECT 78.415 2.86 78.585 3.03 ;
      RECT 78.235 4.775 78.405 4.945 ;
      RECT 77.955 2.86 78.125 3.03 ;
      RECT 77.93 4.205 78.1 4.375 ;
      RECT 77.495 2.86 77.665 3.03 ;
      RECT 77.23 3.995 77.4 4.165 ;
      RECT 77.035 2.86 77.205 3.03 ;
      RECT 76.91 4.44 77.08 4.61 ;
      RECT 76.575 2.86 76.745 3.03 ;
      RECT 76.495 4.475 76.665 4.645 ;
      RECT 76.325 3.46 76.495 3.63 ;
      RECT 76.15 3.915 76.32 4.085 ;
      RECT 76.115 2.86 76.285 3.03 ;
      RECT 75.655 2.86 75.825 3.03 ;
      RECT 75.23 3.565 75.4 3.735 ;
      RECT 75.225 4.88 75.395 5.05 ;
      RECT 75.195 2.86 75.365 3.03 ;
      RECT 74.13 8.755 74.3 8.925 ;
      RECT 74.13 10.235 74.3 10.405 ;
      RECT 73.78 1.395 73.95 1.565 ;
      RECT 73.76 4.055 73.93 4.225 ;
      RECT 73.76 8.385 73.93 8.555 ;
      RECT 73.14 2.205 73.31 2.375 ;
      RECT 73.14 3.685 73.31 3.855 ;
      RECT 73.14 8.755 73.31 8.925 ;
      RECT 73.14 10.235 73.31 10.405 ;
      RECT 72.79 1.395 72.96 1.565 ;
      RECT 72.77 4.055 72.94 4.225 ;
      RECT 72.77 8.385 72.94 8.555 ;
      RECT 72.09 1.4 72.26 1.57 ;
      RECT 71.78 3.32 71.95 3.49 ;
      RECT 71.78 9.12 71.95 9.29 ;
      RECT 71.41 1.4 71.58 1.57 ;
      RECT 71.35 2.21 71.52 2.38 ;
      RECT 71.35 2.95 71.52 3.12 ;
      RECT 71.35 9.49 71.52 9.66 ;
      RECT 71.35 10.23 71.52 10.4 ;
      RECT 70.975 3.69 71.145 3.86 ;
      RECT 70.975 8.75 71.145 8.92 ;
      RECT 70.73 1.4 70.9 1.57 ;
      RECT 70.05 1.4 70.22 1.57 ;
      RECT 68.77 2.86 68.94 3.03 ;
      RECT 68.31 2.86 68.48 3.03 ;
      RECT 67.915 4.2 68.085 4.37 ;
      RECT 67.85 2.86 68.02 3.03 ;
      RECT 67.705 3.54 67.875 3.71 ;
      RECT 67.39 2.86 67.56 3.03 ;
      RECT 67.39 4.45 67.56 4.62 ;
      RECT 67.02 9.12 67.19 9.29 ;
      RECT 67.005 4.045 67.175 4.215 ;
      RECT 66.93 2.86 67.1 3.03 ;
      RECT 66.79 4.61 66.96 4.78 ;
      RECT 66.77 5.01 66.94 5.18 ;
      RECT 66.595 3.565 66.765 3.735 ;
      RECT 66.59 9.49 66.76 9.66 ;
      RECT 66.59 10.23 66.76 10.4 ;
      RECT 66.47 2.86 66.64 3.03 ;
      RECT 66.1 4.545 66.27 4.715 ;
      RECT 66.01 2.86 66.18 3.03 ;
      RECT 65.775 4.23 65.945 4.4 ;
      RECT 65.71 5.01 65.88 5.18 ;
      RECT 65.55 2.86 65.72 3.03 ;
      RECT 65.31 4.995 65.48 5.165 ;
      RECT 65.27 3.48 65.44 3.65 ;
      RECT 65.09 2.86 65.26 3.03 ;
      RECT 64.63 2.86 64.8 3.03 ;
      RECT 64.37 3.98 64.54 4.15 ;
      RECT 64.37 4.44 64.54 4.61 ;
      RECT 64.37 4.955 64.54 5.125 ;
      RECT 64.255 3.515 64.425 3.685 ;
      RECT 64.17 2.86 64.34 3.03 ;
      RECT 63.79 5.025 63.96 5.195 ;
      RECT 63.71 2.86 63.88 3.03 ;
      RECT 63.31 3.555 63.48 3.725 ;
      RECT 63.25 2.86 63.42 3.03 ;
      RECT 63.095 3.93 63.265 4.1 ;
      RECT 62.79 2.86 62.96 3.03 ;
      RECT 62.595 4.53 62.765 4.7 ;
      RECT 62.48 3.98 62.65 4.15 ;
      RECT 62.33 2.86 62.5 3.03 ;
      RECT 62.31 3.43 62.48 3.6 ;
      RECT 61.935 4.46 62.105 4.63 ;
      RECT 61.87 2.86 62.04 3.03 ;
      RECT 61.45 4.06 61.62 4.23 ;
      RECT 61.41 2.86 61.58 3.03 ;
      RECT 61.4 4.835 61.57 5.005 ;
      RECT 60.95 2.86 61.12 3.03 ;
      RECT 60.91 4.46 61.08 4.63 ;
      RECT 60.875 3.565 61.045 3.735 ;
      RECT 60.515 3.965 60.685 4.135 ;
      RECT 60.49 2.86 60.66 3.03 ;
      RECT 60.31 4.775 60.48 4.945 ;
      RECT 60.03 2.86 60.2 3.03 ;
      RECT 60.005 4.205 60.175 4.375 ;
      RECT 59.57 2.86 59.74 3.03 ;
      RECT 59.305 3.995 59.475 4.165 ;
      RECT 59.11 2.86 59.28 3.03 ;
      RECT 58.985 4.44 59.155 4.61 ;
      RECT 58.65 2.86 58.82 3.03 ;
      RECT 58.57 4.475 58.74 4.645 ;
      RECT 58.4 3.46 58.57 3.63 ;
      RECT 58.225 3.915 58.395 4.085 ;
      RECT 58.19 2.86 58.36 3.03 ;
      RECT 57.73 2.86 57.9 3.03 ;
      RECT 57.305 3.565 57.475 3.735 ;
      RECT 57.3 4.88 57.47 5.05 ;
      RECT 57.27 2.86 57.44 3.03 ;
      RECT 56.205 8.755 56.375 8.925 ;
      RECT 56.205 10.235 56.375 10.405 ;
      RECT 55.855 1.395 56.025 1.565 ;
      RECT 55.835 4.055 56.005 4.225 ;
      RECT 55.835 8.385 56.005 8.555 ;
      RECT 55.215 2.205 55.385 2.375 ;
      RECT 55.215 3.685 55.385 3.855 ;
      RECT 55.215 8.755 55.385 8.925 ;
      RECT 55.215 10.235 55.385 10.405 ;
      RECT 54.865 1.395 55.035 1.565 ;
      RECT 54.845 4.055 55.015 4.225 ;
      RECT 54.845 8.385 55.015 8.555 ;
      RECT 54.165 1.4 54.335 1.57 ;
      RECT 53.855 3.32 54.025 3.49 ;
      RECT 53.855 9.12 54.025 9.29 ;
      RECT 53.485 1.4 53.655 1.57 ;
      RECT 53.425 2.21 53.595 2.38 ;
      RECT 53.425 2.95 53.595 3.12 ;
      RECT 53.425 9.49 53.595 9.66 ;
      RECT 53.425 10.23 53.595 10.4 ;
      RECT 53.05 3.69 53.22 3.86 ;
      RECT 53.05 8.75 53.22 8.92 ;
      RECT 52.805 1.4 52.975 1.57 ;
      RECT 52.125 1.4 52.295 1.57 ;
      RECT 50.845 2.86 51.015 3.03 ;
      RECT 50.385 2.86 50.555 3.03 ;
      RECT 49.99 4.2 50.16 4.37 ;
      RECT 49.925 2.86 50.095 3.03 ;
      RECT 49.78 3.54 49.95 3.71 ;
      RECT 49.465 2.86 49.635 3.03 ;
      RECT 49.465 4.45 49.635 4.62 ;
      RECT 49.095 9.12 49.265 9.29 ;
      RECT 49.08 4.045 49.25 4.215 ;
      RECT 49.005 2.86 49.175 3.03 ;
      RECT 48.865 4.61 49.035 4.78 ;
      RECT 48.845 5.01 49.015 5.18 ;
      RECT 48.67 3.565 48.84 3.735 ;
      RECT 48.665 9.49 48.835 9.66 ;
      RECT 48.665 10.23 48.835 10.4 ;
      RECT 48.545 2.86 48.715 3.03 ;
      RECT 48.175 4.545 48.345 4.715 ;
      RECT 48.085 2.86 48.255 3.03 ;
      RECT 47.85 4.23 48.02 4.4 ;
      RECT 47.785 5.01 47.955 5.18 ;
      RECT 47.625 2.86 47.795 3.03 ;
      RECT 47.385 4.995 47.555 5.165 ;
      RECT 47.345 3.48 47.515 3.65 ;
      RECT 47.165 2.86 47.335 3.03 ;
      RECT 46.705 2.86 46.875 3.03 ;
      RECT 46.445 3.98 46.615 4.15 ;
      RECT 46.445 4.44 46.615 4.61 ;
      RECT 46.445 4.955 46.615 5.125 ;
      RECT 46.33 3.515 46.5 3.685 ;
      RECT 46.245 2.86 46.415 3.03 ;
      RECT 45.865 5.025 46.035 5.195 ;
      RECT 45.785 2.86 45.955 3.03 ;
      RECT 45.385 3.555 45.555 3.725 ;
      RECT 45.325 2.86 45.495 3.03 ;
      RECT 45.17 3.93 45.34 4.1 ;
      RECT 44.865 2.86 45.035 3.03 ;
      RECT 44.67 4.53 44.84 4.7 ;
      RECT 44.555 3.98 44.725 4.15 ;
      RECT 44.405 2.86 44.575 3.03 ;
      RECT 44.385 3.43 44.555 3.6 ;
      RECT 44.01 4.46 44.18 4.63 ;
      RECT 43.945 2.86 44.115 3.03 ;
      RECT 43.525 4.06 43.695 4.23 ;
      RECT 43.485 2.86 43.655 3.03 ;
      RECT 43.475 4.835 43.645 5.005 ;
      RECT 43.025 2.86 43.195 3.03 ;
      RECT 42.985 4.46 43.155 4.63 ;
      RECT 42.95 3.565 43.12 3.735 ;
      RECT 42.59 3.965 42.76 4.135 ;
      RECT 42.565 2.86 42.735 3.03 ;
      RECT 42.385 4.775 42.555 4.945 ;
      RECT 42.105 2.86 42.275 3.03 ;
      RECT 42.08 4.205 42.25 4.375 ;
      RECT 41.645 2.86 41.815 3.03 ;
      RECT 41.38 3.995 41.55 4.165 ;
      RECT 41.185 2.86 41.355 3.03 ;
      RECT 41.06 4.44 41.23 4.61 ;
      RECT 40.725 2.86 40.895 3.03 ;
      RECT 40.645 4.475 40.815 4.645 ;
      RECT 40.475 3.46 40.645 3.63 ;
      RECT 40.3 3.915 40.47 4.085 ;
      RECT 40.265 2.86 40.435 3.03 ;
      RECT 39.805 2.86 39.975 3.03 ;
      RECT 39.38 3.565 39.55 3.735 ;
      RECT 39.375 4.88 39.545 5.05 ;
      RECT 39.345 2.86 39.515 3.03 ;
      RECT 38.28 8.755 38.45 8.925 ;
      RECT 38.28 10.235 38.45 10.405 ;
      RECT 37.93 1.395 38.1 1.565 ;
      RECT 37.91 4.055 38.08 4.225 ;
      RECT 37.91 8.385 38.08 8.555 ;
      RECT 37.29 2.205 37.46 2.375 ;
      RECT 37.29 3.685 37.46 3.855 ;
      RECT 37.29 8.755 37.46 8.925 ;
      RECT 37.29 10.235 37.46 10.405 ;
      RECT 36.94 1.395 37.11 1.565 ;
      RECT 36.92 4.055 37.09 4.225 ;
      RECT 36.92 8.385 37.09 8.555 ;
      RECT 36.24 1.4 36.41 1.57 ;
      RECT 35.93 3.32 36.1 3.49 ;
      RECT 35.93 9.12 36.1 9.29 ;
      RECT 35.56 1.4 35.73 1.57 ;
      RECT 35.5 2.21 35.67 2.38 ;
      RECT 35.5 2.95 35.67 3.12 ;
      RECT 35.5 9.49 35.67 9.66 ;
      RECT 35.5 10.23 35.67 10.4 ;
      RECT 35.125 3.69 35.295 3.86 ;
      RECT 35.125 8.75 35.295 8.92 ;
      RECT 34.88 1.4 35.05 1.57 ;
      RECT 34.2 1.4 34.37 1.57 ;
      RECT 32.92 2.86 33.09 3.03 ;
      RECT 32.46 2.86 32.63 3.03 ;
      RECT 32.065 4.2 32.235 4.37 ;
      RECT 32 2.86 32.17 3.03 ;
      RECT 31.855 3.54 32.025 3.71 ;
      RECT 31.54 2.86 31.71 3.03 ;
      RECT 31.54 4.45 31.71 4.62 ;
      RECT 31.17 9.12 31.34 9.29 ;
      RECT 31.155 4.045 31.325 4.215 ;
      RECT 31.08 2.86 31.25 3.03 ;
      RECT 30.94 4.61 31.11 4.78 ;
      RECT 30.92 5.01 31.09 5.18 ;
      RECT 30.745 3.565 30.915 3.735 ;
      RECT 30.74 9.49 30.91 9.66 ;
      RECT 30.74 10.23 30.91 10.4 ;
      RECT 30.62 2.86 30.79 3.03 ;
      RECT 30.25 4.545 30.42 4.715 ;
      RECT 30.16 2.86 30.33 3.03 ;
      RECT 29.925 4.23 30.095 4.4 ;
      RECT 29.86 5.01 30.03 5.18 ;
      RECT 29.7 2.86 29.87 3.03 ;
      RECT 29.46 4.995 29.63 5.165 ;
      RECT 29.42 3.48 29.59 3.65 ;
      RECT 29.24 2.86 29.41 3.03 ;
      RECT 28.78 2.86 28.95 3.03 ;
      RECT 28.52 3.98 28.69 4.15 ;
      RECT 28.52 4.44 28.69 4.61 ;
      RECT 28.52 4.955 28.69 5.125 ;
      RECT 28.405 3.515 28.575 3.685 ;
      RECT 28.32 2.86 28.49 3.03 ;
      RECT 27.94 5.025 28.11 5.195 ;
      RECT 27.86 2.86 28.03 3.03 ;
      RECT 27.46 3.555 27.63 3.725 ;
      RECT 27.4 2.86 27.57 3.03 ;
      RECT 27.245 3.93 27.415 4.1 ;
      RECT 26.94 2.86 27.11 3.03 ;
      RECT 26.745 4.53 26.915 4.7 ;
      RECT 26.63 3.98 26.8 4.15 ;
      RECT 26.48 2.86 26.65 3.03 ;
      RECT 26.46 3.43 26.63 3.6 ;
      RECT 26.085 4.46 26.255 4.63 ;
      RECT 26.02 2.86 26.19 3.03 ;
      RECT 25.6 4.06 25.77 4.23 ;
      RECT 25.56 2.86 25.73 3.03 ;
      RECT 25.55 4.835 25.72 5.005 ;
      RECT 25.1 2.86 25.27 3.03 ;
      RECT 25.06 4.46 25.23 4.63 ;
      RECT 25.025 3.565 25.195 3.735 ;
      RECT 24.665 3.965 24.835 4.135 ;
      RECT 24.64 2.86 24.81 3.03 ;
      RECT 24.46 4.775 24.63 4.945 ;
      RECT 24.18 2.86 24.35 3.03 ;
      RECT 24.155 4.205 24.325 4.375 ;
      RECT 23.72 2.86 23.89 3.03 ;
      RECT 23.455 3.995 23.625 4.165 ;
      RECT 23.26 2.86 23.43 3.03 ;
      RECT 23.135 4.44 23.305 4.61 ;
      RECT 22.8 2.86 22.97 3.03 ;
      RECT 22.72 4.475 22.89 4.645 ;
      RECT 22.55 3.46 22.72 3.63 ;
      RECT 22.375 3.915 22.545 4.085 ;
      RECT 22.34 2.86 22.51 3.03 ;
      RECT 21.88 2.86 22.05 3.03 ;
      RECT 21.455 3.565 21.625 3.735 ;
      RECT 21.45 4.88 21.62 5.05 ;
      RECT 21.42 2.86 21.59 3.03 ;
      RECT 20.355 8.755 20.525 8.925 ;
      RECT 20.355 10.235 20.525 10.405 ;
      RECT 20.005 1.395 20.175 1.565 ;
      RECT 19.985 4.055 20.155 4.225 ;
      RECT 19.985 8.385 20.155 8.555 ;
      RECT 19.365 2.205 19.535 2.375 ;
      RECT 19.365 3.685 19.535 3.855 ;
      RECT 19.365 8.755 19.535 8.925 ;
      RECT 19.365 10.235 19.535 10.405 ;
      RECT 19.015 1.395 19.185 1.565 ;
      RECT 18.995 4.055 19.165 4.225 ;
      RECT 18.995 8.385 19.165 8.555 ;
      RECT 18.315 1.4 18.485 1.57 ;
      RECT 18.005 3.32 18.175 3.49 ;
      RECT 18.005 9.12 18.175 9.29 ;
      RECT 17.635 1.4 17.805 1.57 ;
      RECT 17.575 2.21 17.745 2.38 ;
      RECT 17.575 2.95 17.745 3.12 ;
      RECT 17.575 9.49 17.745 9.66 ;
      RECT 17.575 10.23 17.745 10.4 ;
      RECT 17.2 3.69 17.37 3.86 ;
      RECT 17.2 8.75 17.37 8.92 ;
      RECT 16.955 1.4 17.125 1.57 ;
      RECT 16.275 1.4 16.445 1.57 ;
      RECT 14.995 2.86 15.165 3.03 ;
      RECT 14.535 2.86 14.705 3.03 ;
      RECT 14.14 4.2 14.31 4.37 ;
      RECT 14.075 2.86 14.245 3.03 ;
      RECT 13.93 3.54 14.1 3.71 ;
      RECT 13.615 2.86 13.785 3.03 ;
      RECT 13.615 4.45 13.785 4.62 ;
      RECT 13.245 9.12 13.415 9.29 ;
      RECT 13.23 4.045 13.4 4.215 ;
      RECT 13.155 2.86 13.325 3.03 ;
      RECT 13.015 4.61 13.185 4.78 ;
      RECT 12.995 5.01 13.165 5.18 ;
      RECT 12.82 3.565 12.99 3.735 ;
      RECT 12.815 9.49 12.985 9.66 ;
      RECT 12.815 10.23 12.985 10.4 ;
      RECT 12.695 2.86 12.865 3.03 ;
      RECT 12.325 4.545 12.495 4.715 ;
      RECT 12.235 2.86 12.405 3.03 ;
      RECT 12 4.23 12.17 4.4 ;
      RECT 11.935 5.01 12.105 5.18 ;
      RECT 11.775 2.86 11.945 3.03 ;
      RECT 11.535 4.995 11.705 5.165 ;
      RECT 11.495 3.48 11.665 3.65 ;
      RECT 11.315 2.86 11.485 3.03 ;
      RECT 10.855 2.86 11.025 3.03 ;
      RECT 10.595 3.98 10.765 4.15 ;
      RECT 10.595 4.44 10.765 4.61 ;
      RECT 10.595 4.955 10.765 5.125 ;
      RECT 10.48 3.515 10.65 3.685 ;
      RECT 10.395 2.86 10.565 3.03 ;
      RECT 10.015 5.025 10.185 5.195 ;
      RECT 9.935 2.86 10.105 3.03 ;
      RECT 9.535 3.555 9.705 3.725 ;
      RECT 9.475 2.86 9.645 3.03 ;
      RECT 9.32 3.93 9.49 4.1 ;
      RECT 9.015 2.86 9.185 3.03 ;
      RECT 8.82 4.53 8.99 4.7 ;
      RECT 8.705 3.98 8.875 4.15 ;
      RECT 8.555 2.86 8.725 3.03 ;
      RECT 8.535 3.43 8.705 3.6 ;
      RECT 8.16 4.46 8.33 4.63 ;
      RECT 8.095 2.86 8.265 3.03 ;
      RECT 7.675 4.06 7.845 4.23 ;
      RECT 7.635 2.86 7.805 3.03 ;
      RECT 7.625 4.835 7.795 5.005 ;
      RECT 7.175 2.86 7.345 3.03 ;
      RECT 7.135 4.46 7.305 4.63 ;
      RECT 7.1 3.565 7.27 3.735 ;
      RECT 6.74 3.965 6.91 4.135 ;
      RECT 6.715 2.86 6.885 3.03 ;
      RECT 6.535 4.775 6.705 4.945 ;
      RECT 6.255 2.86 6.425 3.03 ;
      RECT 6.23 4.205 6.4 4.375 ;
      RECT 5.795 2.86 5.965 3.03 ;
      RECT 5.53 3.995 5.7 4.165 ;
      RECT 5.335 2.86 5.505 3.03 ;
      RECT 5.21 4.44 5.38 4.61 ;
      RECT 4.875 2.86 5.045 3.03 ;
      RECT 4.795 4.475 4.965 4.645 ;
      RECT 4.625 3.46 4.795 3.63 ;
      RECT 4.45 3.915 4.62 4.085 ;
      RECT 4.415 2.86 4.585 3.03 ;
      RECT 3.955 2.86 4.125 3.03 ;
      RECT 3.53 3.565 3.7 3.735 ;
      RECT 3.525 4.88 3.695 5.05 ;
      RECT 3.495 2.86 3.665 3.03 ;
      RECT 1.785 9.49 1.955 9.66 ;
      RECT 1.785 10.23 1.955 10.4 ;
      RECT 1.41 8.75 1.58 8.92 ;
    LAYER li1 ;
      RECT 86.1 0 86.27 3.53 ;
      RECT 85.14 0 85.31 3.53 ;
      RECT 84.18 0 84.35 3.53 ;
      RECT 83.66 0 83.83 3.53 ;
      RECT 82.7 0 82.87 3.53 ;
      RECT 81.7 0 81.87 3.53 ;
      RECT 80.74 0 80.91 3.53 ;
      RECT 79.26 0 79.43 3.53 ;
      RECT 77.34 0 77.51 3.53 ;
      RECT 75.86 0 76.03 3.53 ;
      RECT 68.175 0 68.345 3.53 ;
      RECT 67.215 0 67.385 3.53 ;
      RECT 66.255 0 66.425 3.53 ;
      RECT 65.735 0 65.905 3.53 ;
      RECT 64.775 0 64.945 3.53 ;
      RECT 63.775 0 63.945 3.53 ;
      RECT 62.815 0 62.985 3.53 ;
      RECT 61.335 0 61.505 3.53 ;
      RECT 59.415 0 59.585 3.53 ;
      RECT 57.935 0 58.105 3.53 ;
      RECT 50.25 0 50.42 3.53 ;
      RECT 49.29 0 49.46 3.53 ;
      RECT 48.33 0 48.5 3.53 ;
      RECT 47.81 0 47.98 3.53 ;
      RECT 46.85 0 47.02 3.53 ;
      RECT 45.85 0 46.02 3.53 ;
      RECT 44.89 0 45.06 3.53 ;
      RECT 43.41 0 43.58 3.53 ;
      RECT 41.49 0 41.66 3.53 ;
      RECT 40.01 0 40.18 3.53 ;
      RECT 32.325 0 32.495 3.53 ;
      RECT 31.365 0 31.535 3.53 ;
      RECT 30.405 0 30.575 3.53 ;
      RECT 29.885 0 30.055 3.53 ;
      RECT 28.925 0 29.095 3.53 ;
      RECT 27.925 0 28.095 3.53 ;
      RECT 26.965 0 27.135 3.53 ;
      RECT 25.485 0 25.655 3.53 ;
      RECT 23.565 0 23.735 3.53 ;
      RECT 22.085 0 22.255 3.53 ;
      RECT 14.4 0 14.57 3.53 ;
      RECT 13.44 0 13.61 3.53 ;
      RECT 12.48 0 12.65 3.53 ;
      RECT 11.96 0 12.13 3.53 ;
      RECT 11 0 11.17 3.53 ;
      RECT 10 0 10.17 3.53 ;
      RECT 9.04 0 9.21 3.53 ;
      RECT 7.56 0 7.73 3.53 ;
      RECT 5.64 0 5.81 3.53 ;
      RECT 4.16 0 4.33 3.53 ;
      RECT 75.05 0 87.01 3.03 ;
      RECT 57.125 0 69.085 3.03 ;
      RECT 39.2 0 51.16 3.03 ;
      RECT 21.275 0 33.235 3.03 ;
      RECT 3.35 0 15.31 3.03 ;
      RECT 75.045 0 87.01 2.975 ;
      RECT 57.12 0 69.085 2.975 ;
      RECT 39.195 0 51.16 2.975 ;
      RECT 21.27 0 33.235 2.975 ;
      RECT 3.345 0 15.31 2.975 ;
      RECT 3.345 2.435 16.275 2.74 ;
      RECT 87.895 0 88.065 2.23 ;
      RECT 69.97 0 70.14 2.23 ;
      RECT 52.045 0 52.215 2.23 ;
      RECT 34.12 0 34.29 2.23 ;
      RECT 16.195 0 16.365 2.23 ;
      RECT 91.625 0 91.795 2.225 ;
      RECT 90.635 0 90.805 2.225 ;
      RECT 73.7 0 73.87 2.225 ;
      RECT 72.71 0 72.88 2.225 ;
      RECT 55.775 0 55.945 2.225 ;
      RECT 54.785 0 54.955 2.225 ;
      RECT 37.85 0 38.02 2.225 ;
      RECT 36.86 0 37.03 2.225 ;
      RECT 19.925 0 20.095 2.225 ;
      RECT 18.935 0 19.105 2.225 ;
      RECT 0.02 0 92.6 1.6 ;
      RECT 91.685 3.035 91.855 4.225 ;
      RECT 91.685 3.035 92.155 3.205 ;
      RECT 91.685 9.405 92.155 9.575 ;
      RECT 91.685 8.385 91.855 9.575 ;
      RECT 90.695 3.035 90.865 4.225 ;
      RECT 90.695 3.035 91.165 3.205 ;
      RECT 90.695 9.405 91.165 9.575 ;
      RECT 90.695 8.385 90.865 9.575 ;
      RECT 88.845 3.93 89.015 5.16 ;
      RECT 88.9 2.15 89.07 4.1 ;
      RECT 88.845 1.87 89.015 2.32 ;
      RECT 88.845 10.29 89.015 10.74 ;
      RECT 88.9 8.51 89.07 10.46 ;
      RECT 88.845 7.45 89.015 8.68 ;
      RECT 88.325 1.87 88.495 5.16 ;
      RECT 88.325 3.37 88.73 3.7 ;
      RECT 88.325 2.53 88.73 2.86 ;
      RECT 88.325 7.45 88.495 10.74 ;
      RECT 88.325 9.75 88.73 10.08 ;
      RECT 88.325 8.91 88.73 9.24 ;
      RECT 86.425 4.687 86.44 4.738 ;
      RECT 86.42 4.667 86.425 4.785 ;
      RECT 86.405 4.657 86.42 4.853 ;
      RECT 86.38 4.637 86.405 4.908 ;
      RECT 86.34 4.622 86.38 4.928 ;
      RECT 86.295 4.616 86.34 4.956 ;
      RECT 86.225 4.606 86.295 4.973 ;
      RECT 86.205 4.598 86.225 4.973 ;
      RECT 86.145 4.592 86.205 4.965 ;
      RECT 86.086 4.583 86.145 4.953 ;
      RECT 86 4.572 86.086 4.936 ;
      RECT 85.978 4.563 86 4.924 ;
      RECT 85.892 4.556 85.978 4.911 ;
      RECT 85.806 4.543 85.892 4.892 ;
      RECT 85.72 4.531 85.806 4.872 ;
      RECT 85.69 4.52 85.72 4.859 ;
      RECT 85.64 4.506 85.69 4.851 ;
      RECT 85.62 4.495 85.64 4.843 ;
      RECT 85.571 4.484 85.62 4.835 ;
      RECT 85.485 4.463 85.571 4.82 ;
      RECT 85.44 4.45 85.485 4.805 ;
      RECT 85.395 4.45 85.44 4.785 ;
      RECT 85.34 4.45 85.395 4.72 ;
      RECT 85.315 4.45 85.34 4.643 ;
      RECT 85.84 4.187 86.01 4.37 ;
      RECT 85.84 4.187 86.025 4.328 ;
      RECT 85.84 4.187 86.03 4.27 ;
      RECT 85.9 3.955 86.035 4.246 ;
      RECT 85.9 3.959 86.04 4.229 ;
      RECT 85.845 4.122 86.04 4.229 ;
      RECT 85.87 3.967 86.01 4.37 ;
      RECT 85.87 3.971 86.05 4.17 ;
      RECT 85.855 4.057 86.05 4.17 ;
      RECT 85.865 3.987 86.01 4.37 ;
      RECT 85.865 3.99 86.06 4.083 ;
      RECT 85.86 4.007 86.06 4.083 ;
      RECT 85.63 3.227 85.8 3.71 ;
      RECT 85.625 3.222 85.775 3.7 ;
      RECT 85.625 3.229 85.805 3.694 ;
      RECT 85.615 3.223 85.775 3.673 ;
      RECT 85.615 3.239 85.82 3.632 ;
      RECT 85.585 3.224 85.775 3.595 ;
      RECT 85.585 3.254 85.83 3.535 ;
      RECT 85.58 3.226 85.775 3.533 ;
      RECT 85.56 3.235 85.805 3.49 ;
      RECT 85.535 3.251 85.82 3.402 ;
      RECT 85.535 3.27 85.845 3.393 ;
      RECT 85.53 3.307 85.845 3.345 ;
      RECT 85.535 3.287 85.85 3.313 ;
      RECT 85.63 3.221 85.74 3.71 ;
      RECT 85.716 3.22 85.74 3.71 ;
      RECT 84.95 4.005 84.955 4.216 ;
      RECT 85.55 4.005 85.555 4.19 ;
      RECT 85.615 4.045 85.62 4.158 ;
      RECT 85.61 4.037 85.615 4.164 ;
      RECT 85.605 4.027 85.61 4.172 ;
      RECT 85.6 4.017 85.605 4.181 ;
      RECT 85.595 4.007 85.6 4.185 ;
      RECT 85.555 4.005 85.595 4.188 ;
      RECT 85.527 4.004 85.55 4.192 ;
      RECT 85.441 4.001 85.527 4.199 ;
      RECT 85.355 3.997 85.441 4.21 ;
      RECT 85.335 3.995 85.355 4.216 ;
      RECT 85.317 3.994 85.335 4.219 ;
      RECT 85.231 3.992 85.317 4.226 ;
      RECT 85.145 3.987 85.231 4.239 ;
      RECT 85.126 3.984 85.145 4.244 ;
      RECT 85.04 3.982 85.126 4.235 ;
      RECT 85.03 3.982 85.04 4.228 ;
      RECT 84.955 3.995 85.03 4.222 ;
      RECT 84.94 4.006 84.95 4.216 ;
      RECT 84.93 4.008 84.94 4.215 ;
      RECT 84.92 4.012 84.93 4.211 ;
      RECT 84.915 4.015 84.92 4.205 ;
      RECT 84.905 4.017 84.915 4.199 ;
      RECT 84.9 4.02 84.905 4.193 ;
      RECT 84.88 4.606 84.885 4.81 ;
      RECT 84.865 4.593 84.88 4.903 ;
      RECT 84.85 4.574 84.865 5.18 ;
      RECT 84.815 4.54 84.85 5.18 ;
      RECT 84.811 4.51 84.815 5.18 ;
      RECT 84.725 4.392 84.811 5.18 ;
      RECT 84.715 4.267 84.725 5.18 ;
      RECT 84.7 4.235 84.715 5.18 ;
      RECT 84.695 4.21 84.7 5.18 ;
      RECT 84.69 4.2 84.695 5.136 ;
      RECT 84.675 4.172 84.69 5.041 ;
      RECT 84.66 4.138 84.675 4.94 ;
      RECT 84.655 4.116 84.66 4.893 ;
      RECT 84.65 4.105 84.655 4.863 ;
      RECT 84.645 4.095 84.65 4.829 ;
      RECT 84.635 4.082 84.645 4.797 ;
      RECT 84.61 4.058 84.635 4.723 ;
      RECT 84.605 4.038 84.61 4.648 ;
      RECT 84.6 4.032 84.605 4.623 ;
      RECT 84.595 4.027 84.6 4.588 ;
      RECT 84.59 4.022 84.595 4.563 ;
      RECT 84.585 4.02 84.59 4.543 ;
      RECT 84.58 4.02 84.585 4.528 ;
      RECT 84.575 4.02 84.58 4.488 ;
      RECT 84.565 4.02 84.575 4.46 ;
      RECT 84.555 4.02 84.565 4.405 ;
      RECT 84.54 4.02 84.555 4.343 ;
      RECT 84.535 4.019 84.54 4.288 ;
      RECT 84.52 4.018 84.535 4.268 ;
      RECT 84.46 4.016 84.52 4.242 ;
      RECT 84.425 4.017 84.46 4.222 ;
      RECT 84.42 4.019 84.425 4.212 ;
      RECT 84.41 4.038 84.42 4.202 ;
      RECT 84.405 4.065 84.41 4.133 ;
      RECT 84.52 3.49 84.69 3.735 ;
      RECT 84.555 3.261 84.69 3.735 ;
      RECT 84.555 3.263 84.7 3.73 ;
      RECT 84.555 3.265 84.725 3.718 ;
      RECT 84.555 3.268 84.75 3.7 ;
      RECT 84.555 3.273 84.8 3.673 ;
      RECT 84.555 3.278 84.82 3.638 ;
      RECT 84.535 3.28 84.83 3.613 ;
      RECT 84.525 3.375 84.83 3.613 ;
      RECT 84.555 3.26 84.665 3.735 ;
      RECT 84.565 3.257 84.66 3.735 ;
      RECT 84.085 4.522 84.275 4.88 ;
      RECT 84.085 4.534 84.31 4.879 ;
      RECT 84.085 4.562 84.33 4.877 ;
      RECT 84.085 4.587 84.335 4.876 ;
      RECT 84.085 4.645 84.35 4.875 ;
      RECT 84.07 4.518 84.23 4.86 ;
      RECT 84.05 4.527 84.275 4.813 ;
      RECT 84.025 4.538 84.31 4.75 ;
      RECT 84.025 4.622 84.345 4.75 ;
      RECT 84.025 4.597 84.34 4.75 ;
      RECT 84.085 4.513 84.23 4.88 ;
      RECT 84.171 4.512 84.23 4.88 ;
      RECT 84.171 4.511 84.215 4.88 ;
      RECT 83.565 7.45 83.735 10.74 ;
      RECT 83.565 9.75 83.97 10.08 ;
      RECT 83.565 8.91 83.97 9.24 ;
      RECT 83.87 4.027 83.875 4.405 ;
      RECT 83.865 3.995 83.87 4.405 ;
      RECT 83.86 3.967 83.865 4.405 ;
      RECT 83.855 3.947 83.86 4.405 ;
      RECT 83.8 3.93 83.855 4.405 ;
      RECT 83.76 3.915 83.8 4.405 ;
      RECT 83.705 3.902 83.76 4.405 ;
      RECT 83.67 3.893 83.705 4.405 ;
      RECT 83.666 3.891 83.67 4.404 ;
      RECT 83.58 3.887 83.666 4.387 ;
      RECT 83.495 3.879 83.58 4.35 ;
      RECT 83.485 3.875 83.495 4.323 ;
      RECT 83.475 3.875 83.485 4.305 ;
      RECT 83.465 3.877 83.475 4.288 ;
      RECT 83.46 3.882 83.465 4.274 ;
      RECT 83.455 3.886 83.46 4.261 ;
      RECT 83.445 3.891 83.455 4.245 ;
      RECT 83.43 3.905 83.445 4.22 ;
      RECT 83.425 3.911 83.43 4.2 ;
      RECT 83.42 3.913 83.425 4.193 ;
      RECT 83.415 3.917 83.42 4.068 ;
      RECT 83.595 4.717 83.84 5.18 ;
      RECT 83.515 4.69 83.835 5.176 ;
      RECT 83.445 4.725 83.84 5.169 ;
      RECT 83.235 4.98 83.84 5.165 ;
      RECT 83.415 4.748 83.84 5.165 ;
      RECT 83.255 4.94 83.84 5.165 ;
      RECT 83.405 4.76 83.84 5.165 ;
      RECT 83.29 4.877 83.84 5.165 ;
      RECT 83.345 4.802 83.84 5.165 ;
      RECT 83.595 4.667 83.835 5.18 ;
      RECT 83.625 4.66 83.835 5.18 ;
      RECT 83.615 4.662 83.835 5.18 ;
      RECT 83.625 4.657 83.755 5.18 ;
      RECT 83.18 3.22 83.266 3.659 ;
      RECT 83.175 3.22 83.266 3.657 ;
      RECT 83.175 3.22 83.335 3.656 ;
      RECT 83.175 3.22 83.365 3.653 ;
      RECT 83.16 3.227 83.365 3.644 ;
      RECT 83.16 3.227 83.37 3.64 ;
      RECT 83.155 3.237 83.37 3.633 ;
      RECT 83.15 3.242 83.37 3.608 ;
      RECT 83.15 3.242 83.385 3.59 ;
      RECT 83.175 3.22 83.405 3.505 ;
      RECT 83.145 3.247 83.405 3.503 ;
      RECT 83.155 3.24 83.41 3.441 ;
      RECT 83.145 3.362 83.415 3.424 ;
      RECT 83.13 3.257 83.41 3.375 ;
      RECT 83.125 3.267 83.41 3.275 ;
      RECT 83.205 4.038 83.21 4.115 ;
      RECT 83.195 4.032 83.205 4.305 ;
      RECT 83.185 4.024 83.195 4.326 ;
      RECT 83.175 4.015 83.185 4.348 ;
      RECT 83.17 4.01 83.175 4.365 ;
      RECT 83.13 4.01 83.17 4.405 ;
      RECT 83.11 4.01 83.13 4.46 ;
      RECT 83.105 4.01 83.11 4.488 ;
      RECT 83.095 4.01 83.105 4.503 ;
      RECT 83.06 4.01 83.095 4.545 ;
      RECT 83.055 4.01 83.06 4.588 ;
      RECT 83.045 4.01 83.055 4.603 ;
      RECT 83.03 4.01 83.045 4.623 ;
      RECT 83.015 4.01 83.03 4.65 ;
      RECT 83.01 4.011 83.015 4.668 ;
      RECT 82.99 4.012 83.01 4.675 ;
      RECT 82.935 4.013 82.99 4.695 ;
      RECT 82.925 4.014 82.935 4.709 ;
      RECT 82.92 4.017 82.925 4.708 ;
      RECT 82.88 4.09 82.92 4.706 ;
      RECT 82.865 4.17 82.88 4.704 ;
      RECT 82.84 4.225 82.865 4.702 ;
      RECT 82.825 4.29 82.84 4.701 ;
      RECT 82.78 4.322 82.825 4.698 ;
      RECT 82.695 4.345 82.78 4.693 ;
      RECT 82.67 4.365 82.695 4.688 ;
      RECT 82.6 4.37 82.67 4.684 ;
      RECT 82.58 4.372 82.6 4.681 ;
      RECT 82.495 4.383 82.58 4.675 ;
      RECT 82.49 4.394 82.495 4.67 ;
      RECT 82.48 4.396 82.49 4.67 ;
      RECT 82.445 4.4 82.48 4.668 ;
      RECT 82.395 4.41 82.445 4.655 ;
      RECT 82.375 4.418 82.395 4.64 ;
      RECT 82.295 4.43 82.375 4.623 ;
      RECT 82.46 3.98 82.63 4.19 ;
      RECT 82.576 3.976 82.63 4.19 ;
      RECT 82.381 3.98 82.63 4.181 ;
      RECT 82.381 3.98 82.635 4.17 ;
      RECT 82.295 3.98 82.635 4.161 ;
      RECT 82.295 3.988 82.645 4.105 ;
      RECT 82.295 4 82.65 4.018 ;
      RECT 82.295 4.007 82.655 4.01 ;
      RECT 82.49 3.978 82.63 4.19 ;
      RECT 82.245 4.923 82.49 5.255 ;
      RECT 82.24 4.915 82.245 5.252 ;
      RECT 82.21 4.935 82.49 5.233 ;
      RECT 82.19 4.967 82.49 5.206 ;
      RECT 82.24 4.92 82.417 5.252 ;
      RECT 82.24 4.917 82.331 5.252 ;
      RECT 82.18 3.265 82.35 3.685 ;
      RECT 82.175 3.265 82.35 3.683 ;
      RECT 82.175 3.265 82.375 3.673 ;
      RECT 82.175 3.265 82.395 3.648 ;
      RECT 82.17 3.265 82.395 3.643 ;
      RECT 82.17 3.265 82.405 3.633 ;
      RECT 82.17 3.265 82.41 3.628 ;
      RECT 82.17 3.27 82.415 3.623 ;
      RECT 82.17 3.302 82.43 3.613 ;
      RECT 82.17 3.372 82.455 3.596 ;
      RECT 82.15 3.372 82.455 3.588 ;
      RECT 82.15 3.432 82.465 3.565 ;
      RECT 82.15 3.472 82.475 3.51 ;
      RECT 82.135 3.265 82.41 3.49 ;
      RECT 82.125 3.28 82.415 3.388 ;
      RECT 81.715 4.67 81.885 5.195 ;
      RECT 81.71 4.67 81.885 5.188 ;
      RECT 81.7 4.67 81.89 5.153 ;
      RECT 81.695 4.68 81.89 5.125 ;
      RECT 81.69 4.7 81.89 5.108 ;
      RECT 81.7 4.675 81.895 5.098 ;
      RECT 81.685 4.72 81.895 5.09 ;
      RECT 81.68 4.74 81.895 5.075 ;
      RECT 81.675 4.77 81.895 5.065 ;
      RECT 81.665 4.815 81.895 5.04 ;
      RECT 81.695 4.685 81.9 5.023 ;
      RECT 81.66 4.867 81.9 5.018 ;
      RECT 81.695 4.695 81.905 4.988 ;
      RECT 81.655 4.9 81.905 4.985 ;
      RECT 81.65 4.925 81.905 4.965 ;
      RECT 81.69 4.712 81.915 4.905 ;
      RECT 81.685 4.734 81.925 4.798 ;
      RECT 81.635 3.981 81.65 4.25 ;
      RECT 81.59 3.965 81.635 4.295 ;
      RECT 81.585 3.953 81.59 4.345 ;
      RECT 81.575 3.949 81.585 4.378 ;
      RECT 81.57 3.946 81.575 4.406 ;
      RECT 81.555 3.948 81.57 4.448 ;
      RECT 81.55 3.952 81.555 4.488 ;
      RECT 81.53 3.957 81.55 4.54 ;
      RECT 81.526 3.962 81.53 4.597 ;
      RECT 81.44 3.981 81.526 4.634 ;
      RECT 81.43 4.002 81.44 4.67 ;
      RECT 81.425 4.01 81.43 4.671 ;
      RECT 81.42 4.052 81.425 4.672 ;
      RECT 81.405 4.14 81.42 4.673 ;
      RECT 81.395 4.29 81.405 4.675 ;
      RECT 81.39 4.335 81.395 4.677 ;
      RECT 81.355 4.377 81.39 4.68 ;
      RECT 81.35 4.395 81.355 4.683 ;
      RECT 81.273 4.401 81.35 4.689 ;
      RECT 81.187 4.415 81.273 4.702 ;
      RECT 81.101 4.429 81.187 4.716 ;
      RECT 81.015 4.443 81.101 4.729 ;
      RECT 80.955 4.455 81.015 4.741 ;
      RECT 80.93 4.462 80.955 4.748 ;
      RECT 80.916 4.465 80.93 4.753 ;
      RECT 80.83 4.473 80.916 4.769 ;
      RECT 80.825 4.48 80.83 4.784 ;
      RECT 80.801 4.48 80.825 4.791 ;
      RECT 80.715 4.483 80.801 4.819 ;
      RECT 80.63 4.487 80.715 4.863 ;
      RECT 80.565 4.491 80.63 4.9 ;
      RECT 80.54 4.494 80.565 4.916 ;
      RECT 80.465 4.507 80.54 4.92 ;
      RECT 80.44 4.525 80.465 4.924 ;
      RECT 80.43 4.532 80.44 4.926 ;
      RECT 80.415 4.535 80.43 4.927 ;
      RECT 80.355 4.547 80.415 4.931 ;
      RECT 80.345 4.561 80.355 4.935 ;
      RECT 80.29 4.571 80.345 4.923 ;
      RECT 80.265 4.592 80.29 4.906 ;
      RECT 80.245 4.612 80.265 4.897 ;
      RECT 80.24 4.625 80.245 4.892 ;
      RECT 80.225 4.637 80.24 4.888 ;
      RECT 81.46 3.292 81.465 3.315 ;
      RECT 81.455 3.283 81.46 3.355 ;
      RECT 81.45 3.281 81.455 3.398 ;
      RECT 81.445 3.272 81.45 3.433 ;
      RECT 81.44 3.262 81.445 3.505 ;
      RECT 81.435 3.252 81.44 3.57 ;
      RECT 81.43 3.249 81.435 3.61 ;
      RECT 81.405 3.243 81.43 3.7 ;
      RECT 81.37 3.231 81.405 3.725 ;
      RECT 81.36 3.222 81.37 3.725 ;
      RECT 81.225 3.22 81.235 3.708 ;
      RECT 81.215 3.22 81.225 3.675 ;
      RECT 81.21 3.22 81.215 3.65 ;
      RECT 81.205 3.22 81.21 3.638 ;
      RECT 81.2 3.22 81.205 3.62 ;
      RECT 81.19 3.22 81.2 3.585 ;
      RECT 81.185 3.222 81.19 3.563 ;
      RECT 81.18 3.228 81.185 3.548 ;
      RECT 81.175 3.234 81.18 3.533 ;
      RECT 81.16 3.246 81.175 3.506 ;
      RECT 81.155 3.257 81.16 3.474 ;
      RECT 81.15 3.267 81.155 3.458 ;
      RECT 81.14 3.275 81.15 3.427 ;
      RECT 81.135 3.285 81.14 3.401 ;
      RECT 81.13 3.342 81.135 3.384 ;
      RECT 81.235 3.22 81.36 3.725 ;
      RECT 80.95 3.907 81.21 4.205 ;
      RECT 80.945 3.914 81.21 4.203 ;
      RECT 80.95 3.909 81.225 4.198 ;
      RECT 80.94 3.922 81.225 4.195 ;
      RECT 80.94 3.927 81.23 4.188 ;
      RECT 80.935 3.935 81.23 4.185 ;
      RECT 80.935 3.952 81.235 3.983 ;
      RECT 80.95 3.904 81.181 4.205 ;
      RECT 81.005 3.903 81.181 4.205 ;
      RECT 81.005 3.9 81.095 4.205 ;
      RECT 81.005 3.897 81.091 4.205 ;
      RECT 80.695 4.17 80.7 4.183 ;
      RECT 80.69 4.137 80.695 4.188 ;
      RECT 80.685 4.092 80.69 4.195 ;
      RECT 80.68 4.047 80.685 4.203 ;
      RECT 80.675 4.015 80.68 4.211 ;
      RECT 80.67 3.975 80.675 4.212 ;
      RECT 80.655 3.955 80.67 4.214 ;
      RECT 80.58 3.937 80.655 4.226 ;
      RECT 80.57 3.93 80.58 4.237 ;
      RECT 80.565 3.93 80.57 4.239 ;
      RECT 80.535 3.936 80.565 4.243 ;
      RECT 80.495 3.949 80.535 4.243 ;
      RECT 80.47 3.96 80.495 4.229 ;
      RECT 80.455 3.966 80.47 4.212 ;
      RECT 80.445 3.968 80.455 4.203 ;
      RECT 80.44 3.969 80.445 4.198 ;
      RECT 80.435 3.97 80.44 4.193 ;
      RECT 80.43 3.971 80.435 4.19 ;
      RECT 80.405 3.976 80.43 4.18 ;
      RECT 80.395 3.992 80.405 4.167 ;
      RECT 80.39 4.012 80.395 4.162 ;
      RECT 80.4 3.405 80.405 3.601 ;
      RECT 80.385 3.369 80.4 3.603 ;
      RECT 80.375 3.351 80.385 3.608 ;
      RECT 80.365 3.337 80.375 3.612 ;
      RECT 80.32 3.321 80.365 3.622 ;
      RECT 80.315 3.311 80.32 3.631 ;
      RECT 80.27 3.3 80.315 3.637 ;
      RECT 80.265 3.288 80.27 3.644 ;
      RECT 80.25 3.283 80.265 3.648 ;
      RECT 80.235 3.275 80.25 3.653 ;
      RECT 80.225 3.268 80.235 3.658 ;
      RECT 80.215 3.265 80.225 3.663 ;
      RECT 80.205 3.265 80.215 3.664 ;
      RECT 80.2 3.262 80.205 3.663 ;
      RECT 80.165 3.257 80.19 3.662 ;
      RECT 80.141 3.253 80.165 3.661 ;
      RECT 80.055 3.244 80.141 3.658 ;
      RECT 80.04 3.236 80.055 3.655 ;
      RECT 80.018 3.235 80.04 3.654 ;
      RECT 79.932 3.235 80.018 3.652 ;
      RECT 79.846 3.235 79.932 3.65 ;
      RECT 79.76 3.235 79.846 3.647 ;
      RECT 79.75 3.235 79.76 3.638 ;
      RECT 79.72 3.235 79.75 3.598 ;
      RECT 79.71 3.245 79.72 3.553 ;
      RECT 79.705 3.285 79.71 3.538 ;
      RECT 79.7 3.3 79.705 3.525 ;
      RECT 79.67 3.38 79.7 3.487 ;
      RECT 80.19 3.26 80.2 3.663 ;
      RECT 80.015 4.025 80.03 4.63 ;
      RECT 80.02 4.02 80.03 4.63 ;
      RECT 80.185 4.02 80.19 4.203 ;
      RECT 80.175 4.02 80.185 4.233 ;
      RECT 80.16 4.02 80.175 4.293 ;
      RECT 80.155 4.02 80.16 4.338 ;
      RECT 80.15 4.02 80.155 4.368 ;
      RECT 80.145 4.02 80.15 4.388 ;
      RECT 80.135 4.02 80.145 4.423 ;
      RECT 80.12 4.02 80.135 4.455 ;
      RECT 80.075 4.02 80.12 4.483 ;
      RECT 80.07 4.02 80.075 4.513 ;
      RECT 80.065 4.02 80.07 4.525 ;
      RECT 80.06 4.02 80.065 4.533 ;
      RECT 80.05 4.02 80.06 4.548 ;
      RECT 80.045 4.02 80.05 4.57 ;
      RECT 80.035 4.02 80.045 4.593 ;
      RECT 80.03 4.02 80.035 4.613 ;
      RECT 79.995 4.035 80.015 4.63 ;
      RECT 79.97 4.052 79.995 4.63 ;
      RECT 79.965 4.062 79.97 4.63 ;
      RECT 79.935 4.077 79.965 4.63 ;
      RECT 79.86 4.119 79.935 4.63 ;
      RECT 79.855 4.15 79.86 4.613 ;
      RECT 79.85 4.154 79.855 4.595 ;
      RECT 79.845 4.158 79.85 4.558 ;
      RECT 79.84 4.342 79.845 4.525 ;
      RECT 79.325 4.531 79.411 5.096 ;
      RECT 79.28 4.533 79.445 5.09 ;
      RECT 79.411 4.53 79.445 5.09 ;
      RECT 79.325 4.532 79.53 5.084 ;
      RECT 79.28 4.542 79.54 5.08 ;
      RECT 79.255 4.534 79.53 5.076 ;
      RECT 79.25 4.537 79.53 5.071 ;
      RECT 79.225 4.552 79.54 5.065 ;
      RECT 79.225 4.577 79.58 5.06 ;
      RECT 79.185 4.585 79.58 5.035 ;
      RECT 79.185 4.612 79.595 5.033 ;
      RECT 79.185 4.642 79.605 5.02 ;
      RECT 79.18 4.787 79.605 5.008 ;
      RECT 79.185 4.716 79.625 5.005 ;
      RECT 79.185 4.773 79.63 4.813 ;
      RECT 79.375 4.052 79.545 4.23 ;
      RECT 79.325 3.991 79.375 4.215 ;
      RECT 79.06 3.971 79.325 4.2 ;
      RECT 79.02 4.035 79.495 4.2 ;
      RECT 79.02 4.025 79.45 4.2 ;
      RECT 79.02 4.022 79.44 4.2 ;
      RECT 79.02 4.01 79.43 4.2 ;
      RECT 79.02 3.995 79.375 4.2 ;
      RECT 79.06 3.967 79.261 4.2 ;
      RECT 79.07 3.945 79.261 4.2 ;
      RECT 79.095 3.93 79.175 4.2 ;
      RECT 78.85 4.46 78.97 4.905 ;
      RECT 78.835 4.46 78.97 4.904 ;
      RECT 78.79 4.482 78.97 4.899 ;
      RECT 78.75 4.531 78.97 4.893 ;
      RECT 78.75 4.531 78.975 4.868 ;
      RECT 78.75 4.531 78.995 4.758 ;
      RECT 78.745 4.561 78.995 4.755 ;
      RECT 78.835 4.46 79.005 4.65 ;
      RECT 78.495 3.245 78.5 3.69 ;
      RECT 78.305 3.245 78.325 3.655 ;
      RECT 78.275 3.245 78.28 3.63 ;
      RECT 78.955 3.552 78.97 3.74 ;
      RECT 78.95 3.537 78.955 3.746 ;
      RECT 78.93 3.51 78.95 3.749 ;
      RECT 78.88 3.477 78.93 3.758 ;
      RECT 78.85 3.457 78.88 3.762 ;
      RECT 78.831 3.445 78.85 3.758 ;
      RECT 78.745 3.417 78.831 3.748 ;
      RECT 78.735 3.392 78.745 3.738 ;
      RECT 78.665 3.36 78.735 3.73 ;
      RECT 78.64 3.32 78.665 3.722 ;
      RECT 78.62 3.302 78.64 3.716 ;
      RECT 78.61 3.292 78.62 3.713 ;
      RECT 78.6 3.285 78.61 3.711 ;
      RECT 78.58 3.272 78.6 3.708 ;
      RECT 78.57 3.262 78.58 3.705 ;
      RECT 78.56 3.255 78.57 3.703 ;
      RECT 78.51 3.247 78.56 3.697 ;
      RECT 78.5 3.245 78.51 3.691 ;
      RECT 78.47 3.245 78.495 3.688 ;
      RECT 78.441 3.245 78.47 3.683 ;
      RECT 78.355 3.245 78.441 3.673 ;
      RECT 78.325 3.245 78.355 3.66 ;
      RECT 78.28 3.245 78.305 3.643 ;
      RECT 78.265 3.245 78.275 3.625 ;
      RECT 78.245 3.252 78.265 3.61 ;
      RECT 78.24 3.267 78.245 3.598 ;
      RECT 78.235 3.272 78.24 3.538 ;
      RECT 78.23 3.277 78.235 3.38 ;
      RECT 78.225 3.28 78.23 3.298 ;
      RECT 78.49 3.965 78.576 4.286 ;
      RECT 78.49 3.965 78.61 4.279 ;
      RECT 78.44 3.965 78.61 4.275 ;
      RECT 78.44 3.967 78.696 4.273 ;
      RECT 78.44 3.969 78.72 4.267 ;
      RECT 78.44 3.976 78.73 4.266 ;
      RECT 78.44 3.985 78.735 4.263 ;
      RECT 78.44 3.991 78.74 4.258 ;
      RECT 78.44 4.035 78.745 4.255 ;
      RECT 78.44 4.127 78.75 4.252 ;
      RECT 77.965 4.57 78 4.89 ;
      RECT 78.55 4.755 78.555 4.937 ;
      RECT 78.505 4.637 78.55 4.956 ;
      RECT 78.49 4.614 78.505 4.979 ;
      RECT 78.48 4.604 78.49 4.989 ;
      RECT 78.46 4.599 78.48 5.002 ;
      RECT 78.435 4.597 78.46 5.023 ;
      RECT 78.416 4.596 78.435 5.035 ;
      RECT 78.33 4.593 78.416 5.035 ;
      RECT 78.26 4.588 78.33 5.023 ;
      RECT 78.185 4.584 78.26 4.998 ;
      RECT 78.12 4.58 78.185 4.965 ;
      RECT 78.05 4.577 78.12 4.925 ;
      RECT 78.02 4.573 78.05 4.9 ;
      RECT 78 4.571 78.02 4.893 ;
      RECT 77.916 4.569 77.965 4.891 ;
      RECT 77.83 4.566 77.916 4.892 ;
      RECT 77.755 4.565 77.83 4.894 ;
      RECT 77.67 4.565 77.755 4.92 ;
      RECT 77.593 4.566 77.67 4.945 ;
      RECT 77.507 4.567 77.593 4.945 ;
      RECT 77.421 4.567 77.507 4.945 ;
      RECT 77.335 4.568 77.421 4.945 ;
      RECT 77.315 4.569 77.335 4.937 ;
      RECT 77.3 4.575 77.315 4.922 ;
      RECT 77.265 4.595 77.3 4.902 ;
      RECT 77.255 4.615 77.265 4.884 ;
      RECT 78.225 3.92 78.23 4.19 ;
      RECT 78.22 3.911 78.225 4.195 ;
      RECT 78.21 3.901 78.22 4.207 ;
      RECT 78.205 3.89 78.21 4.218 ;
      RECT 78.185 3.884 78.205 4.236 ;
      RECT 78.14 3.881 78.185 4.285 ;
      RECT 78.125 3.88 78.14 4.33 ;
      RECT 78.12 3.88 78.125 4.343 ;
      RECT 78.11 3.88 78.12 4.355 ;
      RECT 78.105 3.881 78.11 4.37 ;
      RECT 78.085 3.889 78.105 4.375 ;
      RECT 78.055 3.905 78.085 4.375 ;
      RECT 78.045 3.917 78.05 4.375 ;
      RECT 78.01 3.932 78.045 4.375 ;
      RECT 77.98 3.952 78.01 4.375 ;
      RECT 77.97 3.977 77.98 4.375 ;
      RECT 77.965 4.005 77.97 4.375 ;
      RECT 77.96 4.035 77.965 4.375 ;
      RECT 77.955 4.052 77.96 4.375 ;
      RECT 77.945 4.08 77.955 4.375 ;
      RECT 77.935 4.115 77.945 4.375 ;
      RECT 77.93 4.15 77.935 4.375 ;
      RECT 78.05 3.915 78.055 4.375 ;
      RECT 77.565 4.017 77.75 4.19 ;
      RECT 77.525 3.935 77.71 4.188 ;
      RECT 77.486 3.94 77.71 4.184 ;
      RECT 77.4 3.949 77.71 4.179 ;
      RECT 77.316 3.965 77.715 4.174 ;
      RECT 77.23 3.985 77.74 4.168 ;
      RECT 77.23 4.005 77.745 4.168 ;
      RECT 77.316 3.975 77.74 4.174 ;
      RECT 77.4 3.95 77.715 4.179 ;
      RECT 77.565 3.932 77.71 4.19 ;
      RECT 77.565 3.927 77.665 4.19 ;
      RECT 77.651 3.921 77.665 4.19 ;
      RECT 77.04 3.245 77.045 3.644 ;
      RECT 76.785 3.245 76.82 3.642 ;
      RECT 76.38 3.28 76.385 3.636 ;
      RECT 77.125 3.283 77.13 3.538 ;
      RECT 77.12 3.281 77.125 3.544 ;
      RECT 77.115 3.28 77.12 3.551 ;
      RECT 77.09 3.273 77.115 3.575 ;
      RECT 77.085 3.266 77.09 3.599 ;
      RECT 77.08 3.262 77.085 3.608 ;
      RECT 77.07 3.257 77.08 3.621 ;
      RECT 77.065 3.254 77.07 3.63 ;
      RECT 77.06 3.252 77.065 3.635 ;
      RECT 77.045 3.248 77.06 3.645 ;
      RECT 77.03 3.242 77.04 3.644 ;
      RECT 76.992 3.24 77.03 3.644 ;
      RECT 76.906 3.242 76.992 3.644 ;
      RECT 76.82 3.244 76.906 3.643 ;
      RECT 76.749 3.245 76.785 3.642 ;
      RECT 76.663 3.247 76.749 3.642 ;
      RECT 76.577 3.249 76.663 3.641 ;
      RECT 76.491 3.251 76.577 3.641 ;
      RECT 76.405 3.254 76.491 3.64 ;
      RECT 76.395 3.26 76.405 3.639 ;
      RECT 76.385 3.272 76.395 3.637 ;
      RECT 76.325 3.307 76.38 3.633 ;
      RECT 76.32 3.337 76.325 3.395 ;
      RECT 77.065 4.417 77.08 4.61 ;
      RECT 77.06 4.385 77.065 4.61 ;
      RECT 77.05 4.36 77.06 4.61 ;
      RECT 77.045 4.332 77.05 4.61 ;
      RECT 77.015 4.255 77.045 4.61 ;
      RECT 76.99 4.137 77.015 4.61 ;
      RECT 76.985 4.075 76.99 4.61 ;
      RECT 76.975 4.062 76.985 4.61 ;
      RECT 76.955 4.052 76.975 4.61 ;
      RECT 76.94 4.035 76.955 4.61 ;
      RECT 76.91 4.023 76.94 4.61 ;
      RECT 76.905 4.022 76.91 4.555 ;
      RECT 76.9 4.022 76.905 4.513 ;
      RECT 76.885 4.021 76.9 4.465 ;
      RECT 76.87 4.021 76.885 4.403 ;
      RECT 76.85 4.021 76.87 4.363 ;
      RECT 76.845 4.021 76.85 4.348 ;
      RECT 76.82 4.02 76.845 4.343 ;
      RECT 76.75 4.019 76.82 4.33 ;
      RECT 76.735 4.018 76.75 4.315 ;
      RECT 76.705 4.017 76.735 4.298 ;
      RECT 76.7 4.017 76.705 4.283 ;
      RECT 76.65 4.016 76.7 4.263 ;
      RECT 76.585 4.015 76.65 4.218 ;
      RECT 76.58 4.015 76.585 4.19 ;
      RECT 76.665 4.552 76.67 4.809 ;
      RECT 76.645 4.471 76.665 4.826 ;
      RECT 76.625 4.465 76.645 4.855 ;
      RECT 76.565 4.452 76.625 4.875 ;
      RECT 76.52 4.436 76.565 4.876 ;
      RECT 76.436 4.424 76.52 4.864 ;
      RECT 76.35 4.411 76.436 4.848 ;
      RECT 76.34 4.404 76.35 4.84 ;
      RECT 76.295 4.401 76.34 4.78 ;
      RECT 76.275 4.397 76.295 4.695 ;
      RECT 76.26 4.395 76.275 4.648 ;
      RECT 76.23 4.392 76.26 4.618 ;
      RECT 76.195 4.388 76.23 4.595 ;
      RECT 76.152 4.383 76.195 4.583 ;
      RECT 76.066 4.374 76.152 4.592 ;
      RECT 75.98 4.363 76.066 4.604 ;
      RECT 75.915 4.354 75.98 4.613 ;
      RECT 75.895 4.345 75.915 4.618 ;
      RECT 75.89 4.338 75.895 4.62 ;
      RECT 75.85 4.323 75.89 4.617 ;
      RECT 75.83 4.302 75.85 4.612 ;
      RECT 75.815 4.29 75.83 4.605 ;
      RECT 75.81 4.282 75.815 4.598 ;
      RECT 75.795 4.262 75.81 4.591 ;
      RECT 75.79 4.125 75.795 4.585 ;
      RECT 75.71 4.014 75.79 4.557 ;
      RECT 75.701 4.007 75.71 4.523 ;
      RECT 75.615 4.001 75.701 4.448 ;
      RECT 75.59 3.992 75.615 4.36 ;
      RECT 75.56 3.987 75.59 4.335 ;
      RECT 75.495 3.996 75.56 4.32 ;
      RECT 75.475 4.012 75.495 4.295 ;
      RECT 75.465 4.018 75.475 4.243 ;
      RECT 75.445 4.04 75.465 4.125 ;
      RECT 76.1 4.005 76.27 4.19 ;
      RECT 76.1 4.005 76.305 4.188 ;
      RECT 76.15 3.915 76.32 4.179 ;
      RECT 76.1 4.072 76.325 4.172 ;
      RECT 76.115 3.95 76.32 4.179 ;
      RECT 75.315 4.683 75.38 5.126 ;
      RECT 75.255 4.708 75.38 5.124 ;
      RECT 75.255 4.708 75.435 5.118 ;
      RECT 75.24 4.733 75.435 5.117 ;
      RECT 75.38 4.67 75.455 5.114 ;
      RECT 75.315 4.695 75.535 5.108 ;
      RECT 75.24 4.734 75.58 5.102 ;
      RECT 75.225 4.761 75.58 5.093 ;
      RECT 75.24 4.754 75.6 5.085 ;
      RECT 75.225 4.763 75.605 5.068 ;
      RECT 75.22 4.78 75.605 4.895 ;
      RECT 75.225 3.502 75.26 3.74 ;
      RECT 75.225 3.502 75.29 3.739 ;
      RECT 75.225 3.502 75.405 3.735 ;
      RECT 75.225 3.502 75.46 3.713 ;
      RECT 75.235 3.445 75.515 3.613 ;
      RECT 75.34 3.285 75.37 3.736 ;
      RECT 75.37 3.28 75.55 3.493 ;
      RECT 75.24 3.421 75.55 3.493 ;
      RECT 75.29 3.317 75.34 3.737 ;
      RECT 75.26 3.373 75.55 3.493 ;
      RECT 73.76 3.035 73.93 4.225 ;
      RECT 73.76 3.035 74.23 3.205 ;
      RECT 73.76 9.405 74.23 9.575 ;
      RECT 73.76 8.385 73.93 9.575 ;
      RECT 72.77 3.035 72.94 4.225 ;
      RECT 72.77 3.035 73.24 3.205 ;
      RECT 72.77 9.405 73.24 9.575 ;
      RECT 72.77 8.385 72.94 9.575 ;
      RECT 70.92 3.93 71.09 5.16 ;
      RECT 70.975 2.15 71.145 4.1 ;
      RECT 70.92 1.87 71.09 2.32 ;
      RECT 70.92 10.29 71.09 10.74 ;
      RECT 70.975 8.51 71.145 10.46 ;
      RECT 70.92 7.45 71.09 8.68 ;
      RECT 70.4 1.87 70.57 5.16 ;
      RECT 70.4 3.37 70.805 3.7 ;
      RECT 70.4 2.53 70.805 2.86 ;
      RECT 70.4 7.45 70.57 10.74 ;
      RECT 70.4 9.75 70.805 10.08 ;
      RECT 70.4 8.91 70.805 9.24 ;
      RECT 68.5 4.687 68.515 4.738 ;
      RECT 68.495 4.667 68.5 4.785 ;
      RECT 68.48 4.657 68.495 4.853 ;
      RECT 68.455 4.637 68.48 4.908 ;
      RECT 68.415 4.622 68.455 4.928 ;
      RECT 68.37 4.616 68.415 4.956 ;
      RECT 68.3 4.606 68.37 4.973 ;
      RECT 68.28 4.598 68.3 4.973 ;
      RECT 68.22 4.592 68.28 4.965 ;
      RECT 68.161 4.583 68.22 4.953 ;
      RECT 68.075 4.572 68.161 4.936 ;
      RECT 68.053 4.563 68.075 4.924 ;
      RECT 67.967 4.556 68.053 4.911 ;
      RECT 67.881 4.543 67.967 4.892 ;
      RECT 67.795 4.531 67.881 4.872 ;
      RECT 67.765 4.52 67.795 4.859 ;
      RECT 67.715 4.506 67.765 4.851 ;
      RECT 67.695 4.495 67.715 4.843 ;
      RECT 67.646 4.484 67.695 4.835 ;
      RECT 67.56 4.463 67.646 4.82 ;
      RECT 67.515 4.45 67.56 4.805 ;
      RECT 67.47 4.45 67.515 4.785 ;
      RECT 67.415 4.45 67.47 4.72 ;
      RECT 67.39 4.45 67.415 4.643 ;
      RECT 67.915 4.187 68.085 4.37 ;
      RECT 67.915 4.187 68.1 4.328 ;
      RECT 67.915 4.187 68.105 4.27 ;
      RECT 67.975 3.955 68.11 4.246 ;
      RECT 67.975 3.959 68.115 4.229 ;
      RECT 67.92 4.122 68.115 4.229 ;
      RECT 67.945 3.967 68.085 4.37 ;
      RECT 67.945 3.971 68.125 4.17 ;
      RECT 67.93 4.057 68.125 4.17 ;
      RECT 67.94 3.987 68.085 4.37 ;
      RECT 67.94 3.99 68.135 4.083 ;
      RECT 67.935 4.007 68.135 4.083 ;
      RECT 67.705 3.227 67.875 3.71 ;
      RECT 67.7 3.222 67.85 3.7 ;
      RECT 67.7 3.229 67.88 3.694 ;
      RECT 67.69 3.223 67.85 3.673 ;
      RECT 67.69 3.239 67.895 3.632 ;
      RECT 67.66 3.224 67.85 3.595 ;
      RECT 67.66 3.254 67.905 3.535 ;
      RECT 67.655 3.226 67.85 3.533 ;
      RECT 67.635 3.235 67.88 3.49 ;
      RECT 67.61 3.251 67.895 3.402 ;
      RECT 67.61 3.27 67.92 3.393 ;
      RECT 67.605 3.307 67.92 3.345 ;
      RECT 67.61 3.287 67.925 3.313 ;
      RECT 67.705 3.221 67.815 3.71 ;
      RECT 67.791 3.22 67.815 3.71 ;
      RECT 67.025 4.005 67.03 4.216 ;
      RECT 67.625 4.005 67.63 4.19 ;
      RECT 67.69 4.045 67.695 4.158 ;
      RECT 67.685 4.037 67.69 4.164 ;
      RECT 67.68 4.027 67.685 4.172 ;
      RECT 67.675 4.017 67.68 4.181 ;
      RECT 67.67 4.007 67.675 4.185 ;
      RECT 67.63 4.005 67.67 4.188 ;
      RECT 67.602 4.004 67.625 4.192 ;
      RECT 67.516 4.001 67.602 4.199 ;
      RECT 67.43 3.997 67.516 4.21 ;
      RECT 67.41 3.995 67.43 4.216 ;
      RECT 67.392 3.994 67.41 4.219 ;
      RECT 67.306 3.992 67.392 4.226 ;
      RECT 67.22 3.987 67.306 4.239 ;
      RECT 67.201 3.984 67.22 4.244 ;
      RECT 67.115 3.982 67.201 4.235 ;
      RECT 67.105 3.982 67.115 4.228 ;
      RECT 67.03 3.995 67.105 4.222 ;
      RECT 67.015 4.006 67.025 4.216 ;
      RECT 67.005 4.008 67.015 4.215 ;
      RECT 66.995 4.012 67.005 4.211 ;
      RECT 66.99 4.015 66.995 4.205 ;
      RECT 66.98 4.017 66.99 4.199 ;
      RECT 66.975 4.02 66.98 4.193 ;
      RECT 66.955 4.606 66.96 4.81 ;
      RECT 66.94 4.593 66.955 4.903 ;
      RECT 66.925 4.574 66.94 5.18 ;
      RECT 66.89 4.54 66.925 5.18 ;
      RECT 66.886 4.51 66.89 5.18 ;
      RECT 66.8 4.392 66.886 5.18 ;
      RECT 66.79 4.267 66.8 5.18 ;
      RECT 66.775 4.235 66.79 5.18 ;
      RECT 66.77 4.21 66.775 5.18 ;
      RECT 66.765 4.2 66.77 5.136 ;
      RECT 66.75 4.172 66.765 5.041 ;
      RECT 66.735 4.138 66.75 4.94 ;
      RECT 66.73 4.116 66.735 4.893 ;
      RECT 66.725 4.105 66.73 4.863 ;
      RECT 66.72 4.095 66.725 4.829 ;
      RECT 66.71 4.082 66.72 4.797 ;
      RECT 66.685 4.058 66.71 4.723 ;
      RECT 66.68 4.038 66.685 4.648 ;
      RECT 66.675 4.032 66.68 4.623 ;
      RECT 66.67 4.027 66.675 4.588 ;
      RECT 66.665 4.022 66.67 4.563 ;
      RECT 66.66 4.02 66.665 4.543 ;
      RECT 66.655 4.02 66.66 4.528 ;
      RECT 66.65 4.02 66.655 4.488 ;
      RECT 66.64 4.02 66.65 4.46 ;
      RECT 66.63 4.02 66.64 4.405 ;
      RECT 66.615 4.02 66.63 4.343 ;
      RECT 66.61 4.019 66.615 4.288 ;
      RECT 66.595 4.018 66.61 4.268 ;
      RECT 66.535 4.016 66.595 4.242 ;
      RECT 66.5 4.017 66.535 4.222 ;
      RECT 66.495 4.019 66.5 4.212 ;
      RECT 66.485 4.038 66.495 4.202 ;
      RECT 66.48 4.065 66.485 4.133 ;
      RECT 66.595 3.49 66.765 3.735 ;
      RECT 66.63 3.261 66.765 3.735 ;
      RECT 66.63 3.263 66.775 3.73 ;
      RECT 66.63 3.265 66.8 3.718 ;
      RECT 66.63 3.268 66.825 3.7 ;
      RECT 66.63 3.273 66.875 3.673 ;
      RECT 66.63 3.278 66.895 3.638 ;
      RECT 66.61 3.28 66.905 3.613 ;
      RECT 66.6 3.375 66.905 3.613 ;
      RECT 66.63 3.26 66.74 3.735 ;
      RECT 66.64 3.257 66.735 3.735 ;
      RECT 66.16 4.522 66.35 4.88 ;
      RECT 66.16 4.534 66.385 4.879 ;
      RECT 66.16 4.562 66.405 4.877 ;
      RECT 66.16 4.587 66.41 4.876 ;
      RECT 66.16 4.645 66.425 4.875 ;
      RECT 66.145 4.518 66.305 4.86 ;
      RECT 66.125 4.527 66.35 4.813 ;
      RECT 66.1 4.538 66.385 4.75 ;
      RECT 66.1 4.622 66.42 4.75 ;
      RECT 66.1 4.597 66.415 4.75 ;
      RECT 66.16 4.513 66.305 4.88 ;
      RECT 66.246 4.512 66.305 4.88 ;
      RECT 66.246 4.511 66.29 4.88 ;
      RECT 65.64 7.45 65.81 10.74 ;
      RECT 65.64 9.75 66.045 10.08 ;
      RECT 65.64 8.91 66.045 9.24 ;
      RECT 65.945 4.027 65.95 4.405 ;
      RECT 65.94 3.995 65.945 4.405 ;
      RECT 65.935 3.967 65.94 4.405 ;
      RECT 65.93 3.947 65.935 4.405 ;
      RECT 65.875 3.93 65.93 4.405 ;
      RECT 65.835 3.915 65.875 4.405 ;
      RECT 65.78 3.902 65.835 4.405 ;
      RECT 65.745 3.893 65.78 4.405 ;
      RECT 65.741 3.891 65.745 4.404 ;
      RECT 65.655 3.887 65.741 4.387 ;
      RECT 65.57 3.879 65.655 4.35 ;
      RECT 65.56 3.875 65.57 4.323 ;
      RECT 65.55 3.875 65.56 4.305 ;
      RECT 65.54 3.877 65.55 4.288 ;
      RECT 65.535 3.882 65.54 4.274 ;
      RECT 65.53 3.886 65.535 4.261 ;
      RECT 65.52 3.891 65.53 4.245 ;
      RECT 65.505 3.905 65.52 4.22 ;
      RECT 65.5 3.911 65.505 4.2 ;
      RECT 65.495 3.913 65.5 4.193 ;
      RECT 65.49 3.917 65.495 4.068 ;
      RECT 65.67 4.717 65.915 5.18 ;
      RECT 65.59 4.69 65.91 5.176 ;
      RECT 65.52 4.725 65.915 5.169 ;
      RECT 65.31 4.98 65.915 5.165 ;
      RECT 65.49 4.748 65.915 5.165 ;
      RECT 65.33 4.94 65.915 5.165 ;
      RECT 65.48 4.76 65.915 5.165 ;
      RECT 65.365 4.877 65.915 5.165 ;
      RECT 65.42 4.802 65.915 5.165 ;
      RECT 65.67 4.667 65.91 5.18 ;
      RECT 65.7 4.66 65.91 5.18 ;
      RECT 65.69 4.662 65.91 5.18 ;
      RECT 65.7 4.657 65.83 5.18 ;
      RECT 65.255 3.22 65.341 3.659 ;
      RECT 65.25 3.22 65.341 3.657 ;
      RECT 65.25 3.22 65.41 3.656 ;
      RECT 65.25 3.22 65.44 3.653 ;
      RECT 65.235 3.227 65.44 3.644 ;
      RECT 65.235 3.227 65.445 3.64 ;
      RECT 65.23 3.237 65.445 3.633 ;
      RECT 65.225 3.242 65.445 3.608 ;
      RECT 65.225 3.242 65.46 3.59 ;
      RECT 65.25 3.22 65.48 3.505 ;
      RECT 65.22 3.247 65.48 3.503 ;
      RECT 65.23 3.24 65.485 3.441 ;
      RECT 65.22 3.362 65.49 3.424 ;
      RECT 65.205 3.257 65.485 3.375 ;
      RECT 65.2 3.267 65.485 3.275 ;
      RECT 65.28 4.038 65.285 4.115 ;
      RECT 65.27 4.032 65.28 4.305 ;
      RECT 65.26 4.024 65.27 4.326 ;
      RECT 65.25 4.015 65.26 4.348 ;
      RECT 65.245 4.01 65.25 4.365 ;
      RECT 65.205 4.01 65.245 4.405 ;
      RECT 65.185 4.01 65.205 4.46 ;
      RECT 65.18 4.01 65.185 4.488 ;
      RECT 65.17 4.01 65.18 4.503 ;
      RECT 65.135 4.01 65.17 4.545 ;
      RECT 65.13 4.01 65.135 4.588 ;
      RECT 65.12 4.01 65.13 4.603 ;
      RECT 65.105 4.01 65.12 4.623 ;
      RECT 65.09 4.01 65.105 4.65 ;
      RECT 65.085 4.011 65.09 4.668 ;
      RECT 65.065 4.012 65.085 4.675 ;
      RECT 65.01 4.013 65.065 4.695 ;
      RECT 65 4.014 65.01 4.709 ;
      RECT 64.995 4.017 65 4.708 ;
      RECT 64.955 4.09 64.995 4.706 ;
      RECT 64.94 4.17 64.955 4.704 ;
      RECT 64.915 4.225 64.94 4.702 ;
      RECT 64.9 4.29 64.915 4.701 ;
      RECT 64.855 4.322 64.9 4.698 ;
      RECT 64.77 4.345 64.855 4.693 ;
      RECT 64.745 4.365 64.77 4.688 ;
      RECT 64.675 4.37 64.745 4.684 ;
      RECT 64.655 4.372 64.675 4.681 ;
      RECT 64.57 4.383 64.655 4.675 ;
      RECT 64.565 4.394 64.57 4.67 ;
      RECT 64.555 4.396 64.565 4.67 ;
      RECT 64.52 4.4 64.555 4.668 ;
      RECT 64.47 4.41 64.52 4.655 ;
      RECT 64.45 4.418 64.47 4.64 ;
      RECT 64.37 4.43 64.45 4.623 ;
      RECT 64.535 3.98 64.705 4.19 ;
      RECT 64.651 3.976 64.705 4.19 ;
      RECT 64.456 3.98 64.705 4.181 ;
      RECT 64.456 3.98 64.71 4.17 ;
      RECT 64.37 3.98 64.71 4.161 ;
      RECT 64.37 3.988 64.72 4.105 ;
      RECT 64.37 4 64.725 4.018 ;
      RECT 64.37 4.007 64.73 4.01 ;
      RECT 64.565 3.978 64.705 4.19 ;
      RECT 64.32 4.923 64.565 5.255 ;
      RECT 64.315 4.915 64.32 5.252 ;
      RECT 64.285 4.935 64.565 5.233 ;
      RECT 64.265 4.967 64.565 5.206 ;
      RECT 64.315 4.92 64.492 5.252 ;
      RECT 64.315 4.917 64.406 5.252 ;
      RECT 64.255 3.265 64.425 3.685 ;
      RECT 64.25 3.265 64.425 3.683 ;
      RECT 64.25 3.265 64.45 3.673 ;
      RECT 64.25 3.265 64.47 3.648 ;
      RECT 64.245 3.265 64.47 3.643 ;
      RECT 64.245 3.265 64.48 3.633 ;
      RECT 64.245 3.265 64.485 3.628 ;
      RECT 64.245 3.27 64.49 3.623 ;
      RECT 64.245 3.302 64.505 3.613 ;
      RECT 64.245 3.372 64.53 3.596 ;
      RECT 64.225 3.372 64.53 3.588 ;
      RECT 64.225 3.432 64.54 3.565 ;
      RECT 64.225 3.472 64.55 3.51 ;
      RECT 64.21 3.265 64.485 3.49 ;
      RECT 64.2 3.28 64.49 3.388 ;
      RECT 63.79 4.67 63.96 5.195 ;
      RECT 63.785 4.67 63.96 5.188 ;
      RECT 63.775 4.67 63.965 5.153 ;
      RECT 63.77 4.68 63.965 5.125 ;
      RECT 63.765 4.7 63.965 5.108 ;
      RECT 63.775 4.675 63.97 5.098 ;
      RECT 63.76 4.72 63.97 5.09 ;
      RECT 63.755 4.74 63.97 5.075 ;
      RECT 63.75 4.77 63.97 5.065 ;
      RECT 63.74 4.815 63.97 5.04 ;
      RECT 63.77 4.685 63.975 5.023 ;
      RECT 63.735 4.867 63.975 5.018 ;
      RECT 63.77 4.695 63.98 4.988 ;
      RECT 63.73 4.9 63.98 4.985 ;
      RECT 63.725 4.925 63.98 4.965 ;
      RECT 63.765 4.712 63.99 4.905 ;
      RECT 63.76 4.734 64 4.798 ;
      RECT 63.71 3.981 63.725 4.25 ;
      RECT 63.665 3.965 63.71 4.295 ;
      RECT 63.66 3.953 63.665 4.345 ;
      RECT 63.65 3.949 63.66 4.378 ;
      RECT 63.645 3.946 63.65 4.406 ;
      RECT 63.63 3.948 63.645 4.448 ;
      RECT 63.625 3.952 63.63 4.488 ;
      RECT 63.605 3.957 63.625 4.54 ;
      RECT 63.601 3.962 63.605 4.597 ;
      RECT 63.515 3.981 63.601 4.634 ;
      RECT 63.505 4.002 63.515 4.67 ;
      RECT 63.5 4.01 63.505 4.671 ;
      RECT 63.495 4.052 63.5 4.672 ;
      RECT 63.48 4.14 63.495 4.673 ;
      RECT 63.47 4.29 63.48 4.675 ;
      RECT 63.465 4.335 63.47 4.677 ;
      RECT 63.43 4.377 63.465 4.68 ;
      RECT 63.425 4.395 63.43 4.683 ;
      RECT 63.348 4.401 63.425 4.689 ;
      RECT 63.262 4.415 63.348 4.702 ;
      RECT 63.176 4.429 63.262 4.716 ;
      RECT 63.09 4.443 63.176 4.729 ;
      RECT 63.03 4.455 63.09 4.741 ;
      RECT 63.005 4.462 63.03 4.748 ;
      RECT 62.991 4.465 63.005 4.753 ;
      RECT 62.905 4.473 62.991 4.769 ;
      RECT 62.9 4.48 62.905 4.784 ;
      RECT 62.876 4.48 62.9 4.791 ;
      RECT 62.79 4.483 62.876 4.819 ;
      RECT 62.705 4.487 62.79 4.863 ;
      RECT 62.64 4.491 62.705 4.9 ;
      RECT 62.615 4.494 62.64 4.916 ;
      RECT 62.54 4.507 62.615 4.92 ;
      RECT 62.515 4.525 62.54 4.924 ;
      RECT 62.505 4.532 62.515 4.926 ;
      RECT 62.49 4.535 62.505 4.927 ;
      RECT 62.43 4.547 62.49 4.931 ;
      RECT 62.42 4.561 62.43 4.935 ;
      RECT 62.365 4.571 62.42 4.923 ;
      RECT 62.34 4.592 62.365 4.906 ;
      RECT 62.32 4.612 62.34 4.897 ;
      RECT 62.315 4.625 62.32 4.892 ;
      RECT 62.3 4.637 62.315 4.888 ;
      RECT 63.535 3.292 63.54 3.315 ;
      RECT 63.53 3.283 63.535 3.355 ;
      RECT 63.525 3.281 63.53 3.398 ;
      RECT 63.52 3.272 63.525 3.433 ;
      RECT 63.515 3.262 63.52 3.505 ;
      RECT 63.51 3.252 63.515 3.57 ;
      RECT 63.505 3.249 63.51 3.61 ;
      RECT 63.48 3.243 63.505 3.7 ;
      RECT 63.445 3.231 63.48 3.725 ;
      RECT 63.435 3.222 63.445 3.725 ;
      RECT 63.3 3.22 63.31 3.708 ;
      RECT 63.29 3.22 63.3 3.675 ;
      RECT 63.285 3.22 63.29 3.65 ;
      RECT 63.28 3.22 63.285 3.638 ;
      RECT 63.275 3.22 63.28 3.62 ;
      RECT 63.265 3.22 63.275 3.585 ;
      RECT 63.26 3.222 63.265 3.563 ;
      RECT 63.255 3.228 63.26 3.548 ;
      RECT 63.25 3.234 63.255 3.533 ;
      RECT 63.235 3.246 63.25 3.506 ;
      RECT 63.23 3.257 63.235 3.474 ;
      RECT 63.225 3.267 63.23 3.458 ;
      RECT 63.215 3.275 63.225 3.427 ;
      RECT 63.21 3.285 63.215 3.401 ;
      RECT 63.205 3.342 63.21 3.384 ;
      RECT 63.31 3.22 63.435 3.725 ;
      RECT 63.025 3.907 63.285 4.205 ;
      RECT 63.02 3.914 63.285 4.203 ;
      RECT 63.025 3.909 63.3 4.198 ;
      RECT 63.015 3.922 63.3 4.195 ;
      RECT 63.015 3.927 63.305 4.188 ;
      RECT 63.01 3.935 63.305 4.185 ;
      RECT 63.01 3.952 63.31 3.983 ;
      RECT 63.025 3.904 63.256 4.205 ;
      RECT 63.08 3.903 63.256 4.205 ;
      RECT 63.08 3.9 63.17 4.205 ;
      RECT 63.08 3.897 63.166 4.205 ;
      RECT 62.77 4.17 62.775 4.183 ;
      RECT 62.765 4.137 62.77 4.188 ;
      RECT 62.76 4.092 62.765 4.195 ;
      RECT 62.755 4.047 62.76 4.203 ;
      RECT 62.75 4.015 62.755 4.211 ;
      RECT 62.745 3.975 62.75 4.212 ;
      RECT 62.73 3.955 62.745 4.214 ;
      RECT 62.655 3.937 62.73 4.226 ;
      RECT 62.645 3.93 62.655 4.237 ;
      RECT 62.64 3.93 62.645 4.239 ;
      RECT 62.61 3.936 62.64 4.243 ;
      RECT 62.57 3.949 62.61 4.243 ;
      RECT 62.545 3.96 62.57 4.229 ;
      RECT 62.53 3.966 62.545 4.212 ;
      RECT 62.52 3.968 62.53 4.203 ;
      RECT 62.515 3.969 62.52 4.198 ;
      RECT 62.51 3.97 62.515 4.193 ;
      RECT 62.505 3.971 62.51 4.19 ;
      RECT 62.48 3.976 62.505 4.18 ;
      RECT 62.47 3.992 62.48 4.167 ;
      RECT 62.465 4.012 62.47 4.162 ;
      RECT 62.475 3.405 62.48 3.601 ;
      RECT 62.46 3.369 62.475 3.603 ;
      RECT 62.45 3.351 62.46 3.608 ;
      RECT 62.44 3.337 62.45 3.612 ;
      RECT 62.395 3.321 62.44 3.622 ;
      RECT 62.39 3.311 62.395 3.631 ;
      RECT 62.345 3.3 62.39 3.637 ;
      RECT 62.34 3.288 62.345 3.644 ;
      RECT 62.325 3.283 62.34 3.648 ;
      RECT 62.31 3.275 62.325 3.653 ;
      RECT 62.3 3.268 62.31 3.658 ;
      RECT 62.29 3.265 62.3 3.663 ;
      RECT 62.28 3.265 62.29 3.664 ;
      RECT 62.275 3.262 62.28 3.663 ;
      RECT 62.24 3.257 62.265 3.662 ;
      RECT 62.216 3.253 62.24 3.661 ;
      RECT 62.13 3.244 62.216 3.658 ;
      RECT 62.115 3.236 62.13 3.655 ;
      RECT 62.093 3.235 62.115 3.654 ;
      RECT 62.007 3.235 62.093 3.652 ;
      RECT 61.921 3.235 62.007 3.65 ;
      RECT 61.835 3.235 61.921 3.647 ;
      RECT 61.825 3.235 61.835 3.638 ;
      RECT 61.795 3.235 61.825 3.598 ;
      RECT 61.785 3.245 61.795 3.553 ;
      RECT 61.78 3.285 61.785 3.538 ;
      RECT 61.775 3.3 61.78 3.525 ;
      RECT 61.745 3.38 61.775 3.487 ;
      RECT 62.265 3.26 62.275 3.663 ;
      RECT 62.09 4.025 62.105 4.63 ;
      RECT 62.095 4.02 62.105 4.63 ;
      RECT 62.26 4.02 62.265 4.203 ;
      RECT 62.25 4.02 62.26 4.233 ;
      RECT 62.235 4.02 62.25 4.293 ;
      RECT 62.23 4.02 62.235 4.338 ;
      RECT 62.225 4.02 62.23 4.368 ;
      RECT 62.22 4.02 62.225 4.388 ;
      RECT 62.21 4.02 62.22 4.423 ;
      RECT 62.195 4.02 62.21 4.455 ;
      RECT 62.15 4.02 62.195 4.483 ;
      RECT 62.145 4.02 62.15 4.513 ;
      RECT 62.14 4.02 62.145 4.525 ;
      RECT 62.135 4.02 62.14 4.533 ;
      RECT 62.125 4.02 62.135 4.548 ;
      RECT 62.12 4.02 62.125 4.57 ;
      RECT 62.11 4.02 62.12 4.593 ;
      RECT 62.105 4.02 62.11 4.613 ;
      RECT 62.07 4.035 62.09 4.63 ;
      RECT 62.045 4.052 62.07 4.63 ;
      RECT 62.04 4.062 62.045 4.63 ;
      RECT 62.01 4.077 62.04 4.63 ;
      RECT 61.935 4.119 62.01 4.63 ;
      RECT 61.93 4.15 61.935 4.613 ;
      RECT 61.925 4.154 61.93 4.595 ;
      RECT 61.92 4.158 61.925 4.558 ;
      RECT 61.915 4.342 61.92 4.525 ;
      RECT 61.4 4.531 61.486 5.096 ;
      RECT 61.355 4.533 61.52 5.09 ;
      RECT 61.486 4.53 61.52 5.09 ;
      RECT 61.4 4.532 61.605 5.084 ;
      RECT 61.355 4.542 61.615 5.08 ;
      RECT 61.33 4.534 61.605 5.076 ;
      RECT 61.325 4.537 61.605 5.071 ;
      RECT 61.3 4.552 61.615 5.065 ;
      RECT 61.3 4.577 61.655 5.06 ;
      RECT 61.26 4.585 61.655 5.035 ;
      RECT 61.26 4.612 61.67 5.033 ;
      RECT 61.26 4.642 61.68 5.02 ;
      RECT 61.255 4.787 61.68 5.008 ;
      RECT 61.26 4.716 61.7 5.005 ;
      RECT 61.26 4.773 61.705 4.813 ;
      RECT 61.45 4.052 61.62 4.23 ;
      RECT 61.4 3.991 61.45 4.215 ;
      RECT 61.135 3.971 61.4 4.2 ;
      RECT 61.095 4.035 61.57 4.2 ;
      RECT 61.095 4.025 61.525 4.2 ;
      RECT 61.095 4.022 61.515 4.2 ;
      RECT 61.095 4.01 61.505 4.2 ;
      RECT 61.095 3.995 61.45 4.2 ;
      RECT 61.135 3.967 61.336 4.2 ;
      RECT 61.145 3.945 61.336 4.2 ;
      RECT 61.17 3.93 61.25 4.2 ;
      RECT 60.925 4.46 61.045 4.905 ;
      RECT 60.91 4.46 61.045 4.904 ;
      RECT 60.865 4.482 61.045 4.899 ;
      RECT 60.825 4.531 61.045 4.893 ;
      RECT 60.825 4.531 61.05 4.868 ;
      RECT 60.825 4.531 61.07 4.758 ;
      RECT 60.82 4.561 61.07 4.755 ;
      RECT 60.91 4.46 61.08 4.65 ;
      RECT 60.57 3.245 60.575 3.69 ;
      RECT 60.38 3.245 60.4 3.655 ;
      RECT 60.35 3.245 60.355 3.63 ;
      RECT 61.03 3.552 61.045 3.74 ;
      RECT 61.025 3.537 61.03 3.746 ;
      RECT 61.005 3.51 61.025 3.749 ;
      RECT 60.955 3.477 61.005 3.758 ;
      RECT 60.925 3.457 60.955 3.762 ;
      RECT 60.906 3.445 60.925 3.758 ;
      RECT 60.82 3.417 60.906 3.748 ;
      RECT 60.81 3.392 60.82 3.738 ;
      RECT 60.74 3.36 60.81 3.73 ;
      RECT 60.715 3.32 60.74 3.722 ;
      RECT 60.695 3.302 60.715 3.716 ;
      RECT 60.685 3.292 60.695 3.713 ;
      RECT 60.675 3.285 60.685 3.711 ;
      RECT 60.655 3.272 60.675 3.708 ;
      RECT 60.645 3.262 60.655 3.705 ;
      RECT 60.635 3.255 60.645 3.703 ;
      RECT 60.585 3.247 60.635 3.697 ;
      RECT 60.575 3.245 60.585 3.691 ;
      RECT 60.545 3.245 60.57 3.688 ;
      RECT 60.516 3.245 60.545 3.683 ;
      RECT 60.43 3.245 60.516 3.673 ;
      RECT 60.4 3.245 60.43 3.66 ;
      RECT 60.355 3.245 60.38 3.643 ;
      RECT 60.34 3.245 60.35 3.625 ;
      RECT 60.32 3.252 60.34 3.61 ;
      RECT 60.315 3.267 60.32 3.598 ;
      RECT 60.31 3.272 60.315 3.538 ;
      RECT 60.305 3.277 60.31 3.38 ;
      RECT 60.3 3.28 60.305 3.298 ;
      RECT 60.565 3.965 60.651 4.286 ;
      RECT 60.565 3.965 60.685 4.279 ;
      RECT 60.515 3.965 60.685 4.275 ;
      RECT 60.515 3.967 60.771 4.273 ;
      RECT 60.515 3.969 60.795 4.267 ;
      RECT 60.515 3.976 60.805 4.266 ;
      RECT 60.515 3.985 60.81 4.263 ;
      RECT 60.515 3.991 60.815 4.258 ;
      RECT 60.515 4.035 60.82 4.255 ;
      RECT 60.515 4.127 60.825 4.252 ;
      RECT 60.04 4.57 60.075 4.89 ;
      RECT 60.625 4.755 60.63 4.937 ;
      RECT 60.58 4.637 60.625 4.956 ;
      RECT 60.565 4.614 60.58 4.979 ;
      RECT 60.555 4.604 60.565 4.989 ;
      RECT 60.535 4.599 60.555 5.002 ;
      RECT 60.51 4.597 60.535 5.023 ;
      RECT 60.491 4.596 60.51 5.035 ;
      RECT 60.405 4.593 60.491 5.035 ;
      RECT 60.335 4.588 60.405 5.023 ;
      RECT 60.26 4.584 60.335 4.998 ;
      RECT 60.195 4.58 60.26 4.965 ;
      RECT 60.125 4.577 60.195 4.925 ;
      RECT 60.095 4.573 60.125 4.9 ;
      RECT 60.075 4.571 60.095 4.893 ;
      RECT 59.991 4.569 60.04 4.891 ;
      RECT 59.905 4.566 59.991 4.892 ;
      RECT 59.83 4.565 59.905 4.894 ;
      RECT 59.745 4.565 59.83 4.92 ;
      RECT 59.668 4.566 59.745 4.945 ;
      RECT 59.582 4.567 59.668 4.945 ;
      RECT 59.496 4.567 59.582 4.945 ;
      RECT 59.41 4.568 59.496 4.945 ;
      RECT 59.39 4.569 59.41 4.937 ;
      RECT 59.375 4.575 59.39 4.922 ;
      RECT 59.34 4.595 59.375 4.902 ;
      RECT 59.33 4.615 59.34 4.884 ;
      RECT 60.3 3.92 60.305 4.19 ;
      RECT 60.295 3.911 60.3 4.195 ;
      RECT 60.285 3.901 60.295 4.207 ;
      RECT 60.28 3.89 60.285 4.218 ;
      RECT 60.26 3.884 60.28 4.236 ;
      RECT 60.215 3.881 60.26 4.285 ;
      RECT 60.2 3.88 60.215 4.33 ;
      RECT 60.195 3.88 60.2 4.343 ;
      RECT 60.185 3.88 60.195 4.355 ;
      RECT 60.18 3.881 60.185 4.37 ;
      RECT 60.16 3.889 60.18 4.375 ;
      RECT 60.13 3.905 60.16 4.375 ;
      RECT 60.12 3.917 60.125 4.375 ;
      RECT 60.085 3.932 60.12 4.375 ;
      RECT 60.055 3.952 60.085 4.375 ;
      RECT 60.045 3.977 60.055 4.375 ;
      RECT 60.04 4.005 60.045 4.375 ;
      RECT 60.035 4.035 60.04 4.375 ;
      RECT 60.03 4.052 60.035 4.375 ;
      RECT 60.02 4.08 60.03 4.375 ;
      RECT 60.01 4.115 60.02 4.375 ;
      RECT 60.005 4.15 60.01 4.375 ;
      RECT 60.125 3.915 60.13 4.375 ;
      RECT 59.64 4.017 59.825 4.19 ;
      RECT 59.6 3.935 59.785 4.188 ;
      RECT 59.561 3.94 59.785 4.184 ;
      RECT 59.475 3.949 59.785 4.179 ;
      RECT 59.391 3.965 59.79 4.174 ;
      RECT 59.305 3.985 59.815 4.168 ;
      RECT 59.305 4.005 59.82 4.168 ;
      RECT 59.391 3.975 59.815 4.174 ;
      RECT 59.475 3.95 59.79 4.179 ;
      RECT 59.64 3.932 59.785 4.19 ;
      RECT 59.64 3.927 59.74 4.19 ;
      RECT 59.726 3.921 59.74 4.19 ;
      RECT 59.115 3.245 59.12 3.644 ;
      RECT 58.86 3.245 58.895 3.642 ;
      RECT 58.455 3.28 58.46 3.636 ;
      RECT 59.2 3.283 59.205 3.538 ;
      RECT 59.195 3.281 59.2 3.544 ;
      RECT 59.19 3.28 59.195 3.551 ;
      RECT 59.165 3.273 59.19 3.575 ;
      RECT 59.16 3.266 59.165 3.599 ;
      RECT 59.155 3.262 59.16 3.608 ;
      RECT 59.145 3.257 59.155 3.621 ;
      RECT 59.14 3.254 59.145 3.63 ;
      RECT 59.135 3.252 59.14 3.635 ;
      RECT 59.12 3.248 59.135 3.645 ;
      RECT 59.105 3.242 59.115 3.644 ;
      RECT 59.067 3.24 59.105 3.644 ;
      RECT 58.981 3.242 59.067 3.644 ;
      RECT 58.895 3.244 58.981 3.643 ;
      RECT 58.824 3.245 58.86 3.642 ;
      RECT 58.738 3.247 58.824 3.642 ;
      RECT 58.652 3.249 58.738 3.641 ;
      RECT 58.566 3.251 58.652 3.641 ;
      RECT 58.48 3.254 58.566 3.64 ;
      RECT 58.47 3.26 58.48 3.639 ;
      RECT 58.46 3.272 58.47 3.637 ;
      RECT 58.4 3.307 58.455 3.633 ;
      RECT 58.395 3.337 58.4 3.395 ;
      RECT 59.14 4.417 59.155 4.61 ;
      RECT 59.135 4.385 59.14 4.61 ;
      RECT 59.125 4.36 59.135 4.61 ;
      RECT 59.12 4.332 59.125 4.61 ;
      RECT 59.09 4.255 59.12 4.61 ;
      RECT 59.065 4.137 59.09 4.61 ;
      RECT 59.06 4.075 59.065 4.61 ;
      RECT 59.05 4.062 59.06 4.61 ;
      RECT 59.03 4.052 59.05 4.61 ;
      RECT 59.015 4.035 59.03 4.61 ;
      RECT 58.985 4.023 59.015 4.61 ;
      RECT 58.98 4.022 58.985 4.555 ;
      RECT 58.975 4.022 58.98 4.513 ;
      RECT 58.96 4.021 58.975 4.465 ;
      RECT 58.945 4.021 58.96 4.403 ;
      RECT 58.925 4.021 58.945 4.363 ;
      RECT 58.92 4.021 58.925 4.348 ;
      RECT 58.895 4.02 58.92 4.343 ;
      RECT 58.825 4.019 58.895 4.33 ;
      RECT 58.81 4.018 58.825 4.315 ;
      RECT 58.78 4.017 58.81 4.298 ;
      RECT 58.775 4.017 58.78 4.283 ;
      RECT 58.725 4.016 58.775 4.263 ;
      RECT 58.66 4.015 58.725 4.218 ;
      RECT 58.655 4.015 58.66 4.19 ;
      RECT 58.74 4.552 58.745 4.809 ;
      RECT 58.72 4.471 58.74 4.826 ;
      RECT 58.7 4.465 58.72 4.855 ;
      RECT 58.64 4.452 58.7 4.875 ;
      RECT 58.595 4.436 58.64 4.876 ;
      RECT 58.511 4.424 58.595 4.864 ;
      RECT 58.425 4.411 58.511 4.848 ;
      RECT 58.415 4.404 58.425 4.84 ;
      RECT 58.37 4.401 58.415 4.78 ;
      RECT 58.35 4.397 58.37 4.695 ;
      RECT 58.335 4.395 58.35 4.648 ;
      RECT 58.305 4.392 58.335 4.618 ;
      RECT 58.27 4.388 58.305 4.595 ;
      RECT 58.227 4.383 58.27 4.583 ;
      RECT 58.141 4.374 58.227 4.592 ;
      RECT 58.055 4.363 58.141 4.604 ;
      RECT 57.99 4.354 58.055 4.613 ;
      RECT 57.97 4.345 57.99 4.618 ;
      RECT 57.965 4.338 57.97 4.62 ;
      RECT 57.925 4.323 57.965 4.617 ;
      RECT 57.905 4.302 57.925 4.612 ;
      RECT 57.89 4.29 57.905 4.605 ;
      RECT 57.885 4.282 57.89 4.598 ;
      RECT 57.87 4.262 57.885 4.591 ;
      RECT 57.865 4.125 57.87 4.585 ;
      RECT 57.785 4.014 57.865 4.557 ;
      RECT 57.776 4.007 57.785 4.523 ;
      RECT 57.69 4.001 57.776 4.448 ;
      RECT 57.665 3.992 57.69 4.36 ;
      RECT 57.635 3.987 57.665 4.335 ;
      RECT 57.57 3.996 57.635 4.32 ;
      RECT 57.55 4.012 57.57 4.295 ;
      RECT 57.54 4.018 57.55 4.243 ;
      RECT 57.52 4.04 57.54 4.125 ;
      RECT 58.175 4.005 58.345 4.19 ;
      RECT 58.175 4.005 58.38 4.188 ;
      RECT 58.225 3.915 58.395 4.179 ;
      RECT 58.175 4.072 58.4 4.172 ;
      RECT 58.19 3.95 58.395 4.179 ;
      RECT 57.39 4.683 57.455 5.126 ;
      RECT 57.33 4.708 57.455 5.124 ;
      RECT 57.33 4.708 57.51 5.118 ;
      RECT 57.315 4.733 57.51 5.117 ;
      RECT 57.455 4.67 57.53 5.114 ;
      RECT 57.39 4.695 57.61 5.108 ;
      RECT 57.315 4.734 57.655 5.102 ;
      RECT 57.3 4.761 57.655 5.093 ;
      RECT 57.315 4.754 57.675 5.085 ;
      RECT 57.3 4.763 57.68 5.068 ;
      RECT 57.295 4.78 57.68 4.895 ;
      RECT 57.3 3.502 57.335 3.74 ;
      RECT 57.3 3.502 57.365 3.739 ;
      RECT 57.3 3.502 57.48 3.735 ;
      RECT 57.3 3.502 57.535 3.713 ;
      RECT 57.31 3.445 57.59 3.613 ;
      RECT 57.415 3.285 57.445 3.736 ;
      RECT 57.445 3.28 57.625 3.493 ;
      RECT 57.315 3.421 57.625 3.493 ;
      RECT 57.365 3.317 57.415 3.737 ;
      RECT 57.335 3.373 57.625 3.493 ;
      RECT 55.835 3.035 56.005 4.225 ;
      RECT 55.835 3.035 56.305 3.205 ;
      RECT 55.835 9.405 56.305 9.575 ;
      RECT 55.835 8.385 56.005 9.575 ;
      RECT 54.845 3.035 55.015 4.225 ;
      RECT 54.845 3.035 55.315 3.205 ;
      RECT 54.845 9.405 55.315 9.575 ;
      RECT 54.845 8.385 55.015 9.575 ;
      RECT 52.995 3.93 53.165 5.16 ;
      RECT 53.05 2.15 53.22 4.1 ;
      RECT 52.995 1.87 53.165 2.32 ;
      RECT 52.995 10.29 53.165 10.74 ;
      RECT 53.05 8.51 53.22 10.46 ;
      RECT 52.995 7.45 53.165 8.68 ;
      RECT 52.475 1.87 52.645 5.16 ;
      RECT 52.475 3.37 52.88 3.7 ;
      RECT 52.475 2.53 52.88 2.86 ;
      RECT 52.475 7.45 52.645 10.74 ;
      RECT 52.475 9.75 52.88 10.08 ;
      RECT 52.475 8.91 52.88 9.24 ;
      RECT 50.575 4.687 50.59 4.738 ;
      RECT 50.57 4.667 50.575 4.785 ;
      RECT 50.555 4.657 50.57 4.853 ;
      RECT 50.53 4.637 50.555 4.908 ;
      RECT 50.49 4.622 50.53 4.928 ;
      RECT 50.445 4.616 50.49 4.956 ;
      RECT 50.375 4.606 50.445 4.973 ;
      RECT 50.355 4.598 50.375 4.973 ;
      RECT 50.295 4.592 50.355 4.965 ;
      RECT 50.236 4.583 50.295 4.953 ;
      RECT 50.15 4.572 50.236 4.936 ;
      RECT 50.128 4.563 50.15 4.924 ;
      RECT 50.042 4.556 50.128 4.911 ;
      RECT 49.956 4.543 50.042 4.892 ;
      RECT 49.87 4.531 49.956 4.872 ;
      RECT 49.84 4.52 49.87 4.859 ;
      RECT 49.79 4.506 49.84 4.851 ;
      RECT 49.77 4.495 49.79 4.843 ;
      RECT 49.721 4.484 49.77 4.835 ;
      RECT 49.635 4.463 49.721 4.82 ;
      RECT 49.59 4.45 49.635 4.805 ;
      RECT 49.545 4.45 49.59 4.785 ;
      RECT 49.49 4.45 49.545 4.72 ;
      RECT 49.465 4.45 49.49 4.643 ;
      RECT 49.99 4.187 50.16 4.37 ;
      RECT 49.99 4.187 50.175 4.328 ;
      RECT 49.99 4.187 50.18 4.27 ;
      RECT 50.05 3.955 50.185 4.246 ;
      RECT 50.05 3.959 50.19 4.229 ;
      RECT 49.995 4.122 50.19 4.229 ;
      RECT 50.02 3.967 50.16 4.37 ;
      RECT 50.02 3.971 50.2 4.17 ;
      RECT 50.005 4.057 50.2 4.17 ;
      RECT 50.015 3.987 50.16 4.37 ;
      RECT 50.015 3.99 50.21 4.083 ;
      RECT 50.01 4.007 50.21 4.083 ;
      RECT 49.78 3.227 49.95 3.71 ;
      RECT 49.775 3.222 49.925 3.7 ;
      RECT 49.775 3.229 49.955 3.694 ;
      RECT 49.765 3.223 49.925 3.673 ;
      RECT 49.765 3.239 49.97 3.632 ;
      RECT 49.735 3.224 49.925 3.595 ;
      RECT 49.735 3.254 49.98 3.535 ;
      RECT 49.73 3.226 49.925 3.533 ;
      RECT 49.71 3.235 49.955 3.49 ;
      RECT 49.685 3.251 49.97 3.402 ;
      RECT 49.685 3.27 49.995 3.393 ;
      RECT 49.68 3.307 49.995 3.345 ;
      RECT 49.685 3.287 50 3.313 ;
      RECT 49.78 3.221 49.89 3.71 ;
      RECT 49.866 3.22 49.89 3.71 ;
      RECT 49.1 4.005 49.105 4.216 ;
      RECT 49.7 4.005 49.705 4.19 ;
      RECT 49.765 4.045 49.77 4.158 ;
      RECT 49.76 4.037 49.765 4.164 ;
      RECT 49.755 4.027 49.76 4.172 ;
      RECT 49.75 4.017 49.755 4.181 ;
      RECT 49.745 4.007 49.75 4.185 ;
      RECT 49.705 4.005 49.745 4.188 ;
      RECT 49.677 4.004 49.7 4.192 ;
      RECT 49.591 4.001 49.677 4.199 ;
      RECT 49.505 3.997 49.591 4.21 ;
      RECT 49.485 3.995 49.505 4.216 ;
      RECT 49.467 3.994 49.485 4.219 ;
      RECT 49.381 3.992 49.467 4.226 ;
      RECT 49.295 3.987 49.381 4.239 ;
      RECT 49.276 3.984 49.295 4.244 ;
      RECT 49.19 3.982 49.276 4.235 ;
      RECT 49.18 3.982 49.19 4.228 ;
      RECT 49.105 3.995 49.18 4.222 ;
      RECT 49.09 4.006 49.1 4.216 ;
      RECT 49.08 4.008 49.09 4.215 ;
      RECT 49.07 4.012 49.08 4.211 ;
      RECT 49.065 4.015 49.07 4.205 ;
      RECT 49.055 4.017 49.065 4.199 ;
      RECT 49.05 4.02 49.055 4.193 ;
      RECT 49.03 4.606 49.035 4.81 ;
      RECT 49.015 4.593 49.03 4.903 ;
      RECT 49 4.574 49.015 5.18 ;
      RECT 48.965 4.54 49 5.18 ;
      RECT 48.961 4.51 48.965 5.18 ;
      RECT 48.875 4.392 48.961 5.18 ;
      RECT 48.865 4.267 48.875 5.18 ;
      RECT 48.85 4.235 48.865 5.18 ;
      RECT 48.845 4.21 48.85 5.18 ;
      RECT 48.84 4.2 48.845 5.136 ;
      RECT 48.825 4.172 48.84 5.041 ;
      RECT 48.81 4.138 48.825 4.94 ;
      RECT 48.805 4.116 48.81 4.893 ;
      RECT 48.8 4.105 48.805 4.863 ;
      RECT 48.795 4.095 48.8 4.829 ;
      RECT 48.785 4.082 48.795 4.797 ;
      RECT 48.76 4.058 48.785 4.723 ;
      RECT 48.755 4.038 48.76 4.648 ;
      RECT 48.75 4.032 48.755 4.623 ;
      RECT 48.745 4.027 48.75 4.588 ;
      RECT 48.74 4.022 48.745 4.563 ;
      RECT 48.735 4.02 48.74 4.543 ;
      RECT 48.73 4.02 48.735 4.528 ;
      RECT 48.725 4.02 48.73 4.488 ;
      RECT 48.715 4.02 48.725 4.46 ;
      RECT 48.705 4.02 48.715 4.405 ;
      RECT 48.69 4.02 48.705 4.343 ;
      RECT 48.685 4.019 48.69 4.288 ;
      RECT 48.67 4.018 48.685 4.268 ;
      RECT 48.61 4.016 48.67 4.242 ;
      RECT 48.575 4.017 48.61 4.222 ;
      RECT 48.57 4.019 48.575 4.212 ;
      RECT 48.56 4.038 48.57 4.202 ;
      RECT 48.555 4.065 48.56 4.133 ;
      RECT 48.67 3.49 48.84 3.735 ;
      RECT 48.705 3.261 48.84 3.735 ;
      RECT 48.705 3.263 48.85 3.73 ;
      RECT 48.705 3.265 48.875 3.718 ;
      RECT 48.705 3.268 48.9 3.7 ;
      RECT 48.705 3.273 48.95 3.673 ;
      RECT 48.705 3.278 48.97 3.638 ;
      RECT 48.685 3.28 48.98 3.613 ;
      RECT 48.675 3.375 48.98 3.613 ;
      RECT 48.705 3.26 48.815 3.735 ;
      RECT 48.715 3.257 48.81 3.735 ;
      RECT 48.235 4.522 48.425 4.88 ;
      RECT 48.235 4.534 48.46 4.879 ;
      RECT 48.235 4.562 48.48 4.877 ;
      RECT 48.235 4.587 48.485 4.876 ;
      RECT 48.235 4.645 48.5 4.875 ;
      RECT 48.22 4.518 48.38 4.86 ;
      RECT 48.2 4.527 48.425 4.813 ;
      RECT 48.175 4.538 48.46 4.75 ;
      RECT 48.175 4.622 48.495 4.75 ;
      RECT 48.175 4.597 48.49 4.75 ;
      RECT 48.235 4.513 48.38 4.88 ;
      RECT 48.321 4.512 48.38 4.88 ;
      RECT 48.321 4.511 48.365 4.88 ;
      RECT 47.715 7.45 47.885 10.74 ;
      RECT 47.715 9.75 48.12 10.08 ;
      RECT 47.715 8.91 48.12 9.24 ;
      RECT 48.02 4.027 48.025 4.405 ;
      RECT 48.015 3.995 48.02 4.405 ;
      RECT 48.01 3.967 48.015 4.405 ;
      RECT 48.005 3.947 48.01 4.405 ;
      RECT 47.95 3.93 48.005 4.405 ;
      RECT 47.91 3.915 47.95 4.405 ;
      RECT 47.855 3.902 47.91 4.405 ;
      RECT 47.82 3.893 47.855 4.405 ;
      RECT 47.816 3.891 47.82 4.404 ;
      RECT 47.73 3.887 47.816 4.387 ;
      RECT 47.645 3.879 47.73 4.35 ;
      RECT 47.635 3.875 47.645 4.323 ;
      RECT 47.625 3.875 47.635 4.305 ;
      RECT 47.615 3.877 47.625 4.288 ;
      RECT 47.61 3.882 47.615 4.274 ;
      RECT 47.605 3.886 47.61 4.261 ;
      RECT 47.595 3.891 47.605 4.245 ;
      RECT 47.58 3.905 47.595 4.22 ;
      RECT 47.575 3.911 47.58 4.2 ;
      RECT 47.57 3.913 47.575 4.193 ;
      RECT 47.565 3.917 47.57 4.068 ;
      RECT 47.745 4.717 47.99 5.18 ;
      RECT 47.665 4.69 47.985 5.176 ;
      RECT 47.595 4.725 47.99 5.169 ;
      RECT 47.385 4.98 47.99 5.165 ;
      RECT 47.565 4.748 47.99 5.165 ;
      RECT 47.405 4.94 47.99 5.165 ;
      RECT 47.555 4.76 47.99 5.165 ;
      RECT 47.44 4.877 47.99 5.165 ;
      RECT 47.495 4.802 47.99 5.165 ;
      RECT 47.745 4.667 47.985 5.18 ;
      RECT 47.775 4.66 47.985 5.18 ;
      RECT 47.765 4.662 47.985 5.18 ;
      RECT 47.775 4.657 47.905 5.18 ;
      RECT 47.33 3.22 47.416 3.659 ;
      RECT 47.325 3.22 47.416 3.657 ;
      RECT 47.325 3.22 47.485 3.656 ;
      RECT 47.325 3.22 47.515 3.653 ;
      RECT 47.31 3.227 47.515 3.644 ;
      RECT 47.31 3.227 47.52 3.64 ;
      RECT 47.305 3.237 47.52 3.633 ;
      RECT 47.3 3.242 47.52 3.608 ;
      RECT 47.3 3.242 47.535 3.59 ;
      RECT 47.325 3.22 47.555 3.505 ;
      RECT 47.295 3.247 47.555 3.503 ;
      RECT 47.305 3.24 47.56 3.441 ;
      RECT 47.295 3.362 47.565 3.424 ;
      RECT 47.28 3.257 47.56 3.375 ;
      RECT 47.275 3.267 47.56 3.275 ;
      RECT 47.355 4.038 47.36 4.115 ;
      RECT 47.345 4.032 47.355 4.305 ;
      RECT 47.335 4.024 47.345 4.326 ;
      RECT 47.325 4.015 47.335 4.348 ;
      RECT 47.32 4.01 47.325 4.365 ;
      RECT 47.28 4.01 47.32 4.405 ;
      RECT 47.26 4.01 47.28 4.46 ;
      RECT 47.255 4.01 47.26 4.488 ;
      RECT 47.245 4.01 47.255 4.503 ;
      RECT 47.21 4.01 47.245 4.545 ;
      RECT 47.205 4.01 47.21 4.588 ;
      RECT 47.195 4.01 47.205 4.603 ;
      RECT 47.18 4.01 47.195 4.623 ;
      RECT 47.165 4.01 47.18 4.65 ;
      RECT 47.16 4.011 47.165 4.668 ;
      RECT 47.14 4.012 47.16 4.675 ;
      RECT 47.085 4.013 47.14 4.695 ;
      RECT 47.075 4.014 47.085 4.709 ;
      RECT 47.07 4.017 47.075 4.708 ;
      RECT 47.03 4.09 47.07 4.706 ;
      RECT 47.015 4.17 47.03 4.704 ;
      RECT 46.99 4.225 47.015 4.702 ;
      RECT 46.975 4.29 46.99 4.701 ;
      RECT 46.93 4.322 46.975 4.698 ;
      RECT 46.845 4.345 46.93 4.693 ;
      RECT 46.82 4.365 46.845 4.688 ;
      RECT 46.75 4.37 46.82 4.684 ;
      RECT 46.73 4.372 46.75 4.681 ;
      RECT 46.645 4.383 46.73 4.675 ;
      RECT 46.64 4.394 46.645 4.67 ;
      RECT 46.63 4.396 46.64 4.67 ;
      RECT 46.595 4.4 46.63 4.668 ;
      RECT 46.545 4.41 46.595 4.655 ;
      RECT 46.525 4.418 46.545 4.64 ;
      RECT 46.445 4.43 46.525 4.623 ;
      RECT 46.61 3.98 46.78 4.19 ;
      RECT 46.726 3.976 46.78 4.19 ;
      RECT 46.531 3.98 46.78 4.181 ;
      RECT 46.531 3.98 46.785 4.17 ;
      RECT 46.445 3.98 46.785 4.161 ;
      RECT 46.445 3.988 46.795 4.105 ;
      RECT 46.445 4 46.8 4.018 ;
      RECT 46.445 4.007 46.805 4.01 ;
      RECT 46.64 3.978 46.78 4.19 ;
      RECT 46.395 4.923 46.64 5.255 ;
      RECT 46.39 4.915 46.395 5.252 ;
      RECT 46.36 4.935 46.64 5.233 ;
      RECT 46.34 4.967 46.64 5.206 ;
      RECT 46.39 4.92 46.567 5.252 ;
      RECT 46.39 4.917 46.481 5.252 ;
      RECT 46.33 3.265 46.5 3.685 ;
      RECT 46.325 3.265 46.5 3.683 ;
      RECT 46.325 3.265 46.525 3.673 ;
      RECT 46.325 3.265 46.545 3.648 ;
      RECT 46.32 3.265 46.545 3.643 ;
      RECT 46.32 3.265 46.555 3.633 ;
      RECT 46.32 3.265 46.56 3.628 ;
      RECT 46.32 3.27 46.565 3.623 ;
      RECT 46.32 3.302 46.58 3.613 ;
      RECT 46.32 3.372 46.605 3.596 ;
      RECT 46.3 3.372 46.605 3.588 ;
      RECT 46.3 3.432 46.615 3.565 ;
      RECT 46.3 3.472 46.625 3.51 ;
      RECT 46.285 3.265 46.56 3.49 ;
      RECT 46.275 3.28 46.565 3.388 ;
      RECT 45.865 4.67 46.035 5.195 ;
      RECT 45.86 4.67 46.035 5.188 ;
      RECT 45.85 4.67 46.04 5.153 ;
      RECT 45.845 4.68 46.04 5.125 ;
      RECT 45.84 4.7 46.04 5.108 ;
      RECT 45.85 4.675 46.045 5.098 ;
      RECT 45.835 4.72 46.045 5.09 ;
      RECT 45.83 4.74 46.045 5.075 ;
      RECT 45.825 4.77 46.045 5.065 ;
      RECT 45.815 4.815 46.045 5.04 ;
      RECT 45.845 4.685 46.05 5.023 ;
      RECT 45.81 4.867 46.05 5.018 ;
      RECT 45.845 4.695 46.055 4.988 ;
      RECT 45.805 4.9 46.055 4.985 ;
      RECT 45.8 4.925 46.055 4.965 ;
      RECT 45.84 4.712 46.065 4.905 ;
      RECT 45.835 4.734 46.075 4.798 ;
      RECT 45.785 3.981 45.8 4.25 ;
      RECT 45.74 3.965 45.785 4.295 ;
      RECT 45.735 3.953 45.74 4.345 ;
      RECT 45.725 3.949 45.735 4.378 ;
      RECT 45.72 3.946 45.725 4.406 ;
      RECT 45.705 3.948 45.72 4.448 ;
      RECT 45.7 3.952 45.705 4.488 ;
      RECT 45.68 3.957 45.7 4.54 ;
      RECT 45.676 3.962 45.68 4.597 ;
      RECT 45.59 3.981 45.676 4.634 ;
      RECT 45.58 4.002 45.59 4.67 ;
      RECT 45.575 4.01 45.58 4.671 ;
      RECT 45.57 4.052 45.575 4.672 ;
      RECT 45.555 4.14 45.57 4.673 ;
      RECT 45.545 4.29 45.555 4.675 ;
      RECT 45.54 4.335 45.545 4.677 ;
      RECT 45.505 4.377 45.54 4.68 ;
      RECT 45.5 4.395 45.505 4.683 ;
      RECT 45.423 4.401 45.5 4.689 ;
      RECT 45.337 4.415 45.423 4.702 ;
      RECT 45.251 4.429 45.337 4.716 ;
      RECT 45.165 4.443 45.251 4.729 ;
      RECT 45.105 4.455 45.165 4.741 ;
      RECT 45.08 4.462 45.105 4.748 ;
      RECT 45.066 4.465 45.08 4.753 ;
      RECT 44.98 4.473 45.066 4.769 ;
      RECT 44.975 4.48 44.98 4.784 ;
      RECT 44.951 4.48 44.975 4.791 ;
      RECT 44.865 4.483 44.951 4.819 ;
      RECT 44.78 4.487 44.865 4.863 ;
      RECT 44.715 4.491 44.78 4.9 ;
      RECT 44.69 4.494 44.715 4.916 ;
      RECT 44.615 4.507 44.69 4.92 ;
      RECT 44.59 4.525 44.615 4.924 ;
      RECT 44.58 4.532 44.59 4.926 ;
      RECT 44.565 4.535 44.58 4.927 ;
      RECT 44.505 4.547 44.565 4.931 ;
      RECT 44.495 4.561 44.505 4.935 ;
      RECT 44.44 4.571 44.495 4.923 ;
      RECT 44.415 4.592 44.44 4.906 ;
      RECT 44.395 4.612 44.415 4.897 ;
      RECT 44.39 4.625 44.395 4.892 ;
      RECT 44.375 4.637 44.39 4.888 ;
      RECT 45.61 3.292 45.615 3.315 ;
      RECT 45.605 3.283 45.61 3.355 ;
      RECT 45.6 3.281 45.605 3.398 ;
      RECT 45.595 3.272 45.6 3.433 ;
      RECT 45.59 3.262 45.595 3.505 ;
      RECT 45.585 3.252 45.59 3.57 ;
      RECT 45.58 3.249 45.585 3.61 ;
      RECT 45.555 3.243 45.58 3.7 ;
      RECT 45.52 3.231 45.555 3.725 ;
      RECT 45.51 3.222 45.52 3.725 ;
      RECT 45.375 3.22 45.385 3.708 ;
      RECT 45.365 3.22 45.375 3.675 ;
      RECT 45.36 3.22 45.365 3.65 ;
      RECT 45.355 3.22 45.36 3.638 ;
      RECT 45.35 3.22 45.355 3.62 ;
      RECT 45.34 3.22 45.35 3.585 ;
      RECT 45.335 3.222 45.34 3.563 ;
      RECT 45.33 3.228 45.335 3.548 ;
      RECT 45.325 3.234 45.33 3.533 ;
      RECT 45.31 3.246 45.325 3.506 ;
      RECT 45.305 3.257 45.31 3.474 ;
      RECT 45.3 3.267 45.305 3.458 ;
      RECT 45.29 3.275 45.3 3.427 ;
      RECT 45.285 3.285 45.29 3.401 ;
      RECT 45.28 3.342 45.285 3.384 ;
      RECT 45.385 3.22 45.51 3.725 ;
      RECT 45.1 3.907 45.36 4.205 ;
      RECT 45.095 3.914 45.36 4.203 ;
      RECT 45.1 3.909 45.375 4.198 ;
      RECT 45.09 3.922 45.375 4.195 ;
      RECT 45.09 3.927 45.38 4.188 ;
      RECT 45.085 3.935 45.38 4.185 ;
      RECT 45.085 3.952 45.385 3.983 ;
      RECT 45.1 3.904 45.331 4.205 ;
      RECT 45.155 3.903 45.331 4.205 ;
      RECT 45.155 3.9 45.245 4.205 ;
      RECT 45.155 3.897 45.241 4.205 ;
      RECT 44.845 4.17 44.85 4.183 ;
      RECT 44.84 4.137 44.845 4.188 ;
      RECT 44.835 4.092 44.84 4.195 ;
      RECT 44.83 4.047 44.835 4.203 ;
      RECT 44.825 4.015 44.83 4.211 ;
      RECT 44.82 3.975 44.825 4.212 ;
      RECT 44.805 3.955 44.82 4.214 ;
      RECT 44.73 3.937 44.805 4.226 ;
      RECT 44.72 3.93 44.73 4.237 ;
      RECT 44.715 3.93 44.72 4.239 ;
      RECT 44.685 3.936 44.715 4.243 ;
      RECT 44.645 3.949 44.685 4.243 ;
      RECT 44.62 3.96 44.645 4.229 ;
      RECT 44.605 3.966 44.62 4.212 ;
      RECT 44.595 3.968 44.605 4.203 ;
      RECT 44.59 3.969 44.595 4.198 ;
      RECT 44.585 3.97 44.59 4.193 ;
      RECT 44.58 3.971 44.585 4.19 ;
      RECT 44.555 3.976 44.58 4.18 ;
      RECT 44.545 3.992 44.555 4.167 ;
      RECT 44.54 4.012 44.545 4.162 ;
      RECT 44.55 3.405 44.555 3.601 ;
      RECT 44.535 3.369 44.55 3.603 ;
      RECT 44.525 3.351 44.535 3.608 ;
      RECT 44.515 3.337 44.525 3.612 ;
      RECT 44.47 3.321 44.515 3.622 ;
      RECT 44.465 3.311 44.47 3.631 ;
      RECT 44.42 3.3 44.465 3.637 ;
      RECT 44.415 3.288 44.42 3.644 ;
      RECT 44.4 3.283 44.415 3.648 ;
      RECT 44.385 3.275 44.4 3.653 ;
      RECT 44.375 3.268 44.385 3.658 ;
      RECT 44.365 3.265 44.375 3.663 ;
      RECT 44.355 3.265 44.365 3.664 ;
      RECT 44.35 3.262 44.355 3.663 ;
      RECT 44.315 3.257 44.34 3.662 ;
      RECT 44.291 3.253 44.315 3.661 ;
      RECT 44.205 3.244 44.291 3.658 ;
      RECT 44.19 3.236 44.205 3.655 ;
      RECT 44.168 3.235 44.19 3.654 ;
      RECT 44.082 3.235 44.168 3.652 ;
      RECT 43.996 3.235 44.082 3.65 ;
      RECT 43.91 3.235 43.996 3.647 ;
      RECT 43.9 3.235 43.91 3.638 ;
      RECT 43.87 3.235 43.9 3.598 ;
      RECT 43.86 3.245 43.87 3.553 ;
      RECT 43.855 3.285 43.86 3.538 ;
      RECT 43.85 3.3 43.855 3.525 ;
      RECT 43.82 3.38 43.85 3.487 ;
      RECT 44.34 3.26 44.35 3.663 ;
      RECT 44.165 4.025 44.18 4.63 ;
      RECT 44.17 4.02 44.18 4.63 ;
      RECT 44.335 4.02 44.34 4.203 ;
      RECT 44.325 4.02 44.335 4.233 ;
      RECT 44.31 4.02 44.325 4.293 ;
      RECT 44.305 4.02 44.31 4.338 ;
      RECT 44.3 4.02 44.305 4.368 ;
      RECT 44.295 4.02 44.3 4.388 ;
      RECT 44.285 4.02 44.295 4.423 ;
      RECT 44.27 4.02 44.285 4.455 ;
      RECT 44.225 4.02 44.27 4.483 ;
      RECT 44.22 4.02 44.225 4.513 ;
      RECT 44.215 4.02 44.22 4.525 ;
      RECT 44.21 4.02 44.215 4.533 ;
      RECT 44.2 4.02 44.21 4.548 ;
      RECT 44.195 4.02 44.2 4.57 ;
      RECT 44.185 4.02 44.195 4.593 ;
      RECT 44.18 4.02 44.185 4.613 ;
      RECT 44.145 4.035 44.165 4.63 ;
      RECT 44.12 4.052 44.145 4.63 ;
      RECT 44.115 4.062 44.12 4.63 ;
      RECT 44.085 4.077 44.115 4.63 ;
      RECT 44.01 4.119 44.085 4.63 ;
      RECT 44.005 4.15 44.01 4.613 ;
      RECT 44 4.154 44.005 4.595 ;
      RECT 43.995 4.158 44 4.558 ;
      RECT 43.99 4.342 43.995 4.525 ;
      RECT 43.475 4.531 43.561 5.096 ;
      RECT 43.43 4.533 43.595 5.09 ;
      RECT 43.561 4.53 43.595 5.09 ;
      RECT 43.475 4.532 43.68 5.084 ;
      RECT 43.43 4.542 43.69 5.08 ;
      RECT 43.405 4.534 43.68 5.076 ;
      RECT 43.4 4.537 43.68 5.071 ;
      RECT 43.375 4.552 43.69 5.065 ;
      RECT 43.375 4.577 43.73 5.06 ;
      RECT 43.335 4.585 43.73 5.035 ;
      RECT 43.335 4.612 43.745 5.033 ;
      RECT 43.335 4.642 43.755 5.02 ;
      RECT 43.33 4.787 43.755 5.008 ;
      RECT 43.335 4.716 43.775 5.005 ;
      RECT 43.335 4.773 43.78 4.813 ;
      RECT 43.525 4.052 43.695 4.23 ;
      RECT 43.475 3.991 43.525 4.215 ;
      RECT 43.21 3.971 43.475 4.2 ;
      RECT 43.17 4.035 43.645 4.2 ;
      RECT 43.17 4.025 43.6 4.2 ;
      RECT 43.17 4.022 43.59 4.2 ;
      RECT 43.17 4.01 43.58 4.2 ;
      RECT 43.17 3.995 43.525 4.2 ;
      RECT 43.21 3.967 43.411 4.2 ;
      RECT 43.22 3.945 43.411 4.2 ;
      RECT 43.245 3.93 43.325 4.2 ;
      RECT 43 4.46 43.12 4.905 ;
      RECT 42.985 4.46 43.12 4.904 ;
      RECT 42.94 4.482 43.12 4.899 ;
      RECT 42.9 4.531 43.12 4.893 ;
      RECT 42.9 4.531 43.125 4.868 ;
      RECT 42.9 4.531 43.145 4.758 ;
      RECT 42.895 4.561 43.145 4.755 ;
      RECT 42.985 4.46 43.155 4.65 ;
      RECT 42.645 3.245 42.65 3.69 ;
      RECT 42.455 3.245 42.475 3.655 ;
      RECT 42.425 3.245 42.43 3.63 ;
      RECT 43.105 3.552 43.12 3.74 ;
      RECT 43.1 3.537 43.105 3.746 ;
      RECT 43.08 3.51 43.1 3.749 ;
      RECT 43.03 3.477 43.08 3.758 ;
      RECT 43 3.457 43.03 3.762 ;
      RECT 42.981 3.445 43 3.758 ;
      RECT 42.895 3.417 42.981 3.748 ;
      RECT 42.885 3.392 42.895 3.738 ;
      RECT 42.815 3.36 42.885 3.73 ;
      RECT 42.79 3.32 42.815 3.722 ;
      RECT 42.77 3.302 42.79 3.716 ;
      RECT 42.76 3.292 42.77 3.713 ;
      RECT 42.75 3.285 42.76 3.711 ;
      RECT 42.73 3.272 42.75 3.708 ;
      RECT 42.72 3.262 42.73 3.705 ;
      RECT 42.71 3.255 42.72 3.703 ;
      RECT 42.66 3.247 42.71 3.697 ;
      RECT 42.65 3.245 42.66 3.691 ;
      RECT 42.62 3.245 42.645 3.688 ;
      RECT 42.591 3.245 42.62 3.683 ;
      RECT 42.505 3.245 42.591 3.673 ;
      RECT 42.475 3.245 42.505 3.66 ;
      RECT 42.43 3.245 42.455 3.643 ;
      RECT 42.415 3.245 42.425 3.625 ;
      RECT 42.395 3.252 42.415 3.61 ;
      RECT 42.39 3.267 42.395 3.598 ;
      RECT 42.385 3.272 42.39 3.538 ;
      RECT 42.38 3.277 42.385 3.38 ;
      RECT 42.375 3.28 42.38 3.298 ;
      RECT 42.64 3.965 42.726 4.286 ;
      RECT 42.64 3.965 42.76 4.279 ;
      RECT 42.59 3.965 42.76 4.275 ;
      RECT 42.59 3.967 42.846 4.273 ;
      RECT 42.59 3.969 42.87 4.267 ;
      RECT 42.59 3.976 42.88 4.266 ;
      RECT 42.59 3.985 42.885 4.263 ;
      RECT 42.59 3.991 42.89 4.258 ;
      RECT 42.59 4.035 42.895 4.255 ;
      RECT 42.59 4.127 42.9 4.252 ;
      RECT 42.115 4.57 42.15 4.89 ;
      RECT 42.7 4.755 42.705 4.937 ;
      RECT 42.655 4.637 42.7 4.956 ;
      RECT 42.64 4.614 42.655 4.979 ;
      RECT 42.63 4.604 42.64 4.989 ;
      RECT 42.61 4.599 42.63 5.002 ;
      RECT 42.585 4.597 42.61 5.023 ;
      RECT 42.566 4.596 42.585 5.035 ;
      RECT 42.48 4.593 42.566 5.035 ;
      RECT 42.41 4.588 42.48 5.023 ;
      RECT 42.335 4.584 42.41 4.998 ;
      RECT 42.27 4.58 42.335 4.965 ;
      RECT 42.2 4.577 42.27 4.925 ;
      RECT 42.17 4.573 42.2 4.9 ;
      RECT 42.15 4.571 42.17 4.893 ;
      RECT 42.066 4.569 42.115 4.891 ;
      RECT 41.98 4.566 42.066 4.892 ;
      RECT 41.905 4.565 41.98 4.894 ;
      RECT 41.82 4.565 41.905 4.92 ;
      RECT 41.743 4.566 41.82 4.945 ;
      RECT 41.657 4.567 41.743 4.945 ;
      RECT 41.571 4.567 41.657 4.945 ;
      RECT 41.485 4.568 41.571 4.945 ;
      RECT 41.465 4.569 41.485 4.937 ;
      RECT 41.45 4.575 41.465 4.922 ;
      RECT 41.415 4.595 41.45 4.902 ;
      RECT 41.405 4.615 41.415 4.884 ;
      RECT 42.375 3.92 42.38 4.19 ;
      RECT 42.37 3.911 42.375 4.195 ;
      RECT 42.36 3.901 42.37 4.207 ;
      RECT 42.355 3.89 42.36 4.218 ;
      RECT 42.335 3.884 42.355 4.236 ;
      RECT 42.29 3.881 42.335 4.285 ;
      RECT 42.275 3.88 42.29 4.33 ;
      RECT 42.27 3.88 42.275 4.343 ;
      RECT 42.26 3.88 42.27 4.355 ;
      RECT 42.255 3.881 42.26 4.37 ;
      RECT 42.235 3.889 42.255 4.375 ;
      RECT 42.205 3.905 42.235 4.375 ;
      RECT 42.195 3.917 42.2 4.375 ;
      RECT 42.16 3.932 42.195 4.375 ;
      RECT 42.13 3.952 42.16 4.375 ;
      RECT 42.12 3.977 42.13 4.375 ;
      RECT 42.115 4.005 42.12 4.375 ;
      RECT 42.11 4.035 42.115 4.375 ;
      RECT 42.105 4.052 42.11 4.375 ;
      RECT 42.095 4.08 42.105 4.375 ;
      RECT 42.085 4.115 42.095 4.375 ;
      RECT 42.08 4.15 42.085 4.375 ;
      RECT 42.2 3.915 42.205 4.375 ;
      RECT 41.715 4.017 41.9 4.19 ;
      RECT 41.675 3.935 41.86 4.188 ;
      RECT 41.636 3.94 41.86 4.184 ;
      RECT 41.55 3.949 41.86 4.179 ;
      RECT 41.466 3.965 41.865 4.174 ;
      RECT 41.38 3.985 41.89 4.168 ;
      RECT 41.38 4.005 41.895 4.168 ;
      RECT 41.466 3.975 41.89 4.174 ;
      RECT 41.55 3.95 41.865 4.179 ;
      RECT 41.715 3.932 41.86 4.19 ;
      RECT 41.715 3.927 41.815 4.19 ;
      RECT 41.801 3.921 41.815 4.19 ;
      RECT 41.19 3.245 41.195 3.644 ;
      RECT 40.935 3.245 40.97 3.642 ;
      RECT 40.53 3.28 40.535 3.636 ;
      RECT 41.275 3.283 41.28 3.538 ;
      RECT 41.27 3.281 41.275 3.544 ;
      RECT 41.265 3.28 41.27 3.551 ;
      RECT 41.24 3.273 41.265 3.575 ;
      RECT 41.235 3.266 41.24 3.599 ;
      RECT 41.23 3.262 41.235 3.608 ;
      RECT 41.22 3.257 41.23 3.621 ;
      RECT 41.215 3.254 41.22 3.63 ;
      RECT 41.21 3.252 41.215 3.635 ;
      RECT 41.195 3.248 41.21 3.645 ;
      RECT 41.18 3.242 41.19 3.644 ;
      RECT 41.142 3.24 41.18 3.644 ;
      RECT 41.056 3.242 41.142 3.644 ;
      RECT 40.97 3.244 41.056 3.643 ;
      RECT 40.899 3.245 40.935 3.642 ;
      RECT 40.813 3.247 40.899 3.642 ;
      RECT 40.727 3.249 40.813 3.641 ;
      RECT 40.641 3.251 40.727 3.641 ;
      RECT 40.555 3.254 40.641 3.64 ;
      RECT 40.545 3.26 40.555 3.639 ;
      RECT 40.535 3.272 40.545 3.637 ;
      RECT 40.475 3.307 40.53 3.633 ;
      RECT 40.47 3.337 40.475 3.395 ;
      RECT 41.215 4.417 41.23 4.61 ;
      RECT 41.21 4.385 41.215 4.61 ;
      RECT 41.2 4.36 41.21 4.61 ;
      RECT 41.195 4.332 41.2 4.61 ;
      RECT 41.165 4.255 41.195 4.61 ;
      RECT 41.14 4.137 41.165 4.61 ;
      RECT 41.135 4.075 41.14 4.61 ;
      RECT 41.125 4.062 41.135 4.61 ;
      RECT 41.105 4.052 41.125 4.61 ;
      RECT 41.09 4.035 41.105 4.61 ;
      RECT 41.06 4.023 41.09 4.61 ;
      RECT 41.055 4.022 41.06 4.555 ;
      RECT 41.05 4.022 41.055 4.513 ;
      RECT 41.035 4.021 41.05 4.465 ;
      RECT 41.02 4.021 41.035 4.403 ;
      RECT 41 4.021 41.02 4.363 ;
      RECT 40.995 4.021 41 4.348 ;
      RECT 40.97 4.02 40.995 4.343 ;
      RECT 40.9 4.019 40.97 4.33 ;
      RECT 40.885 4.018 40.9 4.315 ;
      RECT 40.855 4.017 40.885 4.298 ;
      RECT 40.85 4.017 40.855 4.283 ;
      RECT 40.8 4.016 40.85 4.263 ;
      RECT 40.735 4.015 40.8 4.218 ;
      RECT 40.73 4.015 40.735 4.19 ;
      RECT 40.815 4.552 40.82 4.809 ;
      RECT 40.795 4.471 40.815 4.826 ;
      RECT 40.775 4.465 40.795 4.855 ;
      RECT 40.715 4.452 40.775 4.875 ;
      RECT 40.67 4.436 40.715 4.876 ;
      RECT 40.586 4.424 40.67 4.864 ;
      RECT 40.5 4.411 40.586 4.848 ;
      RECT 40.49 4.404 40.5 4.84 ;
      RECT 40.445 4.401 40.49 4.78 ;
      RECT 40.425 4.397 40.445 4.695 ;
      RECT 40.41 4.395 40.425 4.648 ;
      RECT 40.38 4.392 40.41 4.618 ;
      RECT 40.345 4.388 40.38 4.595 ;
      RECT 40.302 4.383 40.345 4.583 ;
      RECT 40.216 4.374 40.302 4.592 ;
      RECT 40.13 4.363 40.216 4.604 ;
      RECT 40.065 4.354 40.13 4.613 ;
      RECT 40.045 4.345 40.065 4.618 ;
      RECT 40.04 4.338 40.045 4.62 ;
      RECT 40 4.323 40.04 4.617 ;
      RECT 39.98 4.302 40 4.612 ;
      RECT 39.965 4.29 39.98 4.605 ;
      RECT 39.96 4.282 39.965 4.598 ;
      RECT 39.945 4.262 39.96 4.591 ;
      RECT 39.94 4.125 39.945 4.585 ;
      RECT 39.86 4.014 39.94 4.557 ;
      RECT 39.851 4.007 39.86 4.523 ;
      RECT 39.765 4.001 39.851 4.448 ;
      RECT 39.74 3.992 39.765 4.36 ;
      RECT 39.71 3.987 39.74 4.335 ;
      RECT 39.645 3.996 39.71 4.32 ;
      RECT 39.625 4.012 39.645 4.295 ;
      RECT 39.615 4.018 39.625 4.243 ;
      RECT 39.595 4.04 39.615 4.125 ;
      RECT 40.25 4.005 40.42 4.19 ;
      RECT 40.25 4.005 40.455 4.188 ;
      RECT 40.3 3.915 40.47 4.179 ;
      RECT 40.25 4.072 40.475 4.172 ;
      RECT 40.265 3.95 40.47 4.179 ;
      RECT 39.465 4.683 39.53 5.126 ;
      RECT 39.405 4.708 39.53 5.124 ;
      RECT 39.405 4.708 39.585 5.118 ;
      RECT 39.39 4.733 39.585 5.117 ;
      RECT 39.53 4.67 39.605 5.114 ;
      RECT 39.465 4.695 39.685 5.108 ;
      RECT 39.39 4.734 39.73 5.102 ;
      RECT 39.375 4.761 39.73 5.093 ;
      RECT 39.39 4.754 39.75 5.085 ;
      RECT 39.375 4.763 39.755 5.068 ;
      RECT 39.37 4.78 39.755 4.895 ;
      RECT 39.375 3.502 39.41 3.74 ;
      RECT 39.375 3.502 39.44 3.739 ;
      RECT 39.375 3.502 39.555 3.735 ;
      RECT 39.375 3.502 39.61 3.713 ;
      RECT 39.385 3.445 39.665 3.613 ;
      RECT 39.49 3.285 39.52 3.736 ;
      RECT 39.52 3.28 39.7 3.493 ;
      RECT 39.39 3.421 39.7 3.493 ;
      RECT 39.44 3.317 39.49 3.737 ;
      RECT 39.41 3.373 39.7 3.493 ;
      RECT 37.91 3.035 38.08 4.225 ;
      RECT 37.91 3.035 38.38 3.205 ;
      RECT 37.91 9.405 38.38 9.575 ;
      RECT 37.91 8.385 38.08 9.575 ;
      RECT 36.92 3.035 37.09 4.225 ;
      RECT 36.92 3.035 37.39 3.205 ;
      RECT 36.92 9.405 37.39 9.575 ;
      RECT 36.92 8.385 37.09 9.575 ;
      RECT 35.07 3.93 35.24 5.16 ;
      RECT 35.125 2.15 35.295 4.1 ;
      RECT 35.07 1.87 35.24 2.32 ;
      RECT 35.07 10.29 35.24 10.74 ;
      RECT 35.125 8.51 35.295 10.46 ;
      RECT 35.07 7.45 35.24 8.68 ;
      RECT 34.55 1.87 34.72 5.16 ;
      RECT 34.55 3.37 34.955 3.7 ;
      RECT 34.55 2.53 34.955 2.86 ;
      RECT 34.55 7.45 34.72 10.74 ;
      RECT 34.55 9.75 34.955 10.08 ;
      RECT 34.55 8.91 34.955 9.24 ;
      RECT 32.65 4.687 32.665 4.738 ;
      RECT 32.645 4.667 32.65 4.785 ;
      RECT 32.63 4.657 32.645 4.853 ;
      RECT 32.605 4.637 32.63 4.908 ;
      RECT 32.565 4.622 32.605 4.928 ;
      RECT 32.52 4.616 32.565 4.956 ;
      RECT 32.45 4.606 32.52 4.973 ;
      RECT 32.43 4.598 32.45 4.973 ;
      RECT 32.37 4.592 32.43 4.965 ;
      RECT 32.311 4.583 32.37 4.953 ;
      RECT 32.225 4.572 32.311 4.936 ;
      RECT 32.203 4.563 32.225 4.924 ;
      RECT 32.117 4.556 32.203 4.911 ;
      RECT 32.031 4.543 32.117 4.892 ;
      RECT 31.945 4.531 32.031 4.872 ;
      RECT 31.915 4.52 31.945 4.859 ;
      RECT 31.865 4.506 31.915 4.851 ;
      RECT 31.845 4.495 31.865 4.843 ;
      RECT 31.796 4.484 31.845 4.835 ;
      RECT 31.71 4.463 31.796 4.82 ;
      RECT 31.665 4.45 31.71 4.805 ;
      RECT 31.62 4.45 31.665 4.785 ;
      RECT 31.565 4.45 31.62 4.72 ;
      RECT 31.54 4.45 31.565 4.643 ;
      RECT 32.065 4.187 32.235 4.37 ;
      RECT 32.065 4.187 32.25 4.328 ;
      RECT 32.065 4.187 32.255 4.27 ;
      RECT 32.125 3.955 32.26 4.246 ;
      RECT 32.125 3.959 32.265 4.229 ;
      RECT 32.07 4.122 32.265 4.229 ;
      RECT 32.095 3.967 32.235 4.37 ;
      RECT 32.095 3.971 32.275 4.17 ;
      RECT 32.08 4.057 32.275 4.17 ;
      RECT 32.09 3.987 32.235 4.37 ;
      RECT 32.09 3.99 32.285 4.083 ;
      RECT 32.085 4.007 32.285 4.083 ;
      RECT 31.855 3.227 32.025 3.71 ;
      RECT 31.85 3.222 32 3.7 ;
      RECT 31.85 3.229 32.03 3.694 ;
      RECT 31.84 3.223 32 3.673 ;
      RECT 31.84 3.239 32.045 3.632 ;
      RECT 31.81 3.224 32 3.595 ;
      RECT 31.81 3.254 32.055 3.535 ;
      RECT 31.805 3.226 32 3.533 ;
      RECT 31.785 3.235 32.03 3.49 ;
      RECT 31.76 3.251 32.045 3.402 ;
      RECT 31.76 3.27 32.07 3.393 ;
      RECT 31.755 3.307 32.07 3.345 ;
      RECT 31.76 3.287 32.075 3.313 ;
      RECT 31.855 3.221 31.965 3.71 ;
      RECT 31.941 3.22 31.965 3.71 ;
      RECT 31.175 4.005 31.18 4.216 ;
      RECT 31.775 4.005 31.78 4.19 ;
      RECT 31.84 4.045 31.845 4.158 ;
      RECT 31.835 4.037 31.84 4.164 ;
      RECT 31.83 4.027 31.835 4.172 ;
      RECT 31.825 4.017 31.83 4.181 ;
      RECT 31.82 4.007 31.825 4.185 ;
      RECT 31.78 4.005 31.82 4.188 ;
      RECT 31.752 4.004 31.775 4.192 ;
      RECT 31.666 4.001 31.752 4.199 ;
      RECT 31.58 3.997 31.666 4.21 ;
      RECT 31.56 3.995 31.58 4.216 ;
      RECT 31.542 3.994 31.56 4.219 ;
      RECT 31.456 3.992 31.542 4.226 ;
      RECT 31.37 3.987 31.456 4.239 ;
      RECT 31.351 3.984 31.37 4.244 ;
      RECT 31.265 3.982 31.351 4.235 ;
      RECT 31.255 3.982 31.265 4.228 ;
      RECT 31.18 3.995 31.255 4.222 ;
      RECT 31.165 4.006 31.175 4.216 ;
      RECT 31.155 4.008 31.165 4.215 ;
      RECT 31.145 4.012 31.155 4.211 ;
      RECT 31.14 4.015 31.145 4.205 ;
      RECT 31.13 4.017 31.14 4.199 ;
      RECT 31.125 4.02 31.13 4.193 ;
      RECT 31.105 4.606 31.11 4.81 ;
      RECT 31.09 4.593 31.105 4.903 ;
      RECT 31.075 4.574 31.09 5.18 ;
      RECT 31.04 4.54 31.075 5.18 ;
      RECT 31.036 4.51 31.04 5.18 ;
      RECT 30.95 4.392 31.036 5.18 ;
      RECT 30.94 4.267 30.95 5.18 ;
      RECT 30.925 4.235 30.94 5.18 ;
      RECT 30.92 4.21 30.925 5.18 ;
      RECT 30.915 4.2 30.92 5.136 ;
      RECT 30.9 4.172 30.915 5.041 ;
      RECT 30.885 4.138 30.9 4.94 ;
      RECT 30.88 4.116 30.885 4.893 ;
      RECT 30.875 4.105 30.88 4.863 ;
      RECT 30.87 4.095 30.875 4.829 ;
      RECT 30.86 4.082 30.87 4.797 ;
      RECT 30.835 4.058 30.86 4.723 ;
      RECT 30.83 4.038 30.835 4.648 ;
      RECT 30.825 4.032 30.83 4.623 ;
      RECT 30.82 4.027 30.825 4.588 ;
      RECT 30.815 4.022 30.82 4.563 ;
      RECT 30.81 4.02 30.815 4.543 ;
      RECT 30.805 4.02 30.81 4.528 ;
      RECT 30.8 4.02 30.805 4.488 ;
      RECT 30.79 4.02 30.8 4.46 ;
      RECT 30.78 4.02 30.79 4.405 ;
      RECT 30.765 4.02 30.78 4.343 ;
      RECT 30.76 4.019 30.765 4.288 ;
      RECT 30.745 4.018 30.76 4.268 ;
      RECT 30.685 4.016 30.745 4.242 ;
      RECT 30.65 4.017 30.685 4.222 ;
      RECT 30.645 4.019 30.65 4.212 ;
      RECT 30.635 4.038 30.645 4.202 ;
      RECT 30.63 4.065 30.635 4.133 ;
      RECT 30.745 3.49 30.915 3.735 ;
      RECT 30.78 3.261 30.915 3.735 ;
      RECT 30.78 3.263 30.925 3.73 ;
      RECT 30.78 3.265 30.95 3.718 ;
      RECT 30.78 3.268 30.975 3.7 ;
      RECT 30.78 3.273 31.025 3.673 ;
      RECT 30.78 3.278 31.045 3.638 ;
      RECT 30.76 3.28 31.055 3.613 ;
      RECT 30.75 3.375 31.055 3.613 ;
      RECT 30.78 3.26 30.89 3.735 ;
      RECT 30.79 3.257 30.885 3.735 ;
      RECT 30.31 4.522 30.5 4.88 ;
      RECT 30.31 4.534 30.535 4.879 ;
      RECT 30.31 4.562 30.555 4.877 ;
      RECT 30.31 4.587 30.56 4.876 ;
      RECT 30.31 4.645 30.575 4.875 ;
      RECT 30.295 4.518 30.455 4.86 ;
      RECT 30.275 4.527 30.5 4.813 ;
      RECT 30.25 4.538 30.535 4.75 ;
      RECT 30.25 4.622 30.57 4.75 ;
      RECT 30.25 4.597 30.565 4.75 ;
      RECT 30.31 4.513 30.455 4.88 ;
      RECT 30.396 4.512 30.455 4.88 ;
      RECT 30.396 4.511 30.44 4.88 ;
      RECT 29.79 7.45 29.96 10.74 ;
      RECT 29.79 9.75 30.195 10.08 ;
      RECT 29.79 8.91 30.195 9.24 ;
      RECT 30.095 4.027 30.1 4.405 ;
      RECT 30.09 3.995 30.095 4.405 ;
      RECT 30.085 3.967 30.09 4.405 ;
      RECT 30.08 3.947 30.085 4.405 ;
      RECT 30.025 3.93 30.08 4.405 ;
      RECT 29.985 3.915 30.025 4.405 ;
      RECT 29.93 3.902 29.985 4.405 ;
      RECT 29.895 3.893 29.93 4.405 ;
      RECT 29.891 3.891 29.895 4.404 ;
      RECT 29.805 3.887 29.891 4.387 ;
      RECT 29.72 3.879 29.805 4.35 ;
      RECT 29.71 3.875 29.72 4.323 ;
      RECT 29.7 3.875 29.71 4.305 ;
      RECT 29.69 3.877 29.7 4.288 ;
      RECT 29.685 3.882 29.69 4.274 ;
      RECT 29.68 3.886 29.685 4.261 ;
      RECT 29.67 3.891 29.68 4.245 ;
      RECT 29.655 3.905 29.67 4.22 ;
      RECT 29.65 3.911 29.655 4.2 ;
      RECT 29.645 3.913 29.65 4.193 ;
      RECT 29.64 3.917 29.645 4.068 ;
      RECT 29.82 4.717 30.065 5.18 ;
      RECT 29.74 4.69 30.06 5.176 ;
      RECT 29.67 4.725 30.065 5.169 ;
      RECT 29.46 4.98 30.065 5.165 ;
      RECT 29.64 4.748 30.065 5.165 ;
      RECT 29.48 4.94 30.065 5.165 ;
      RECT 29.63 4.76 30.065 5.165 ;
      RECT 29.515 4.877 30.065 5.165 ;
      RECT 29.57 4.802 30.065 5.165 ;
      RECT 29.82 4.667 30.06 5.18 ;
      RECT 29.85 4.66 30.06 5.18 ;
      RECT 29.84 4.662 30.06 5.18 ;
      RECT 29.85 4.657 29.98 5.18 ;
      RECT 29.405 3.22 29.491 3.659 ;
      RECT 29.4 3.22 29.491 3.657 ;
      RECT 29.4 3.22 29.56 3.656 ;
      RECT 29.4 3.22 29.59 3.653 ;
      RECT 29.385 3.227 29.59 3.644 ;
      RECT 29.385 3.227 29.595 3.64 ;
      RECT 29.38 3.237 29.595 3.633 ;
      RECT 29.375 3.242 29.595 3.608 ;
      RECT 29.375 3.242 29.61 3.59 ;
      RECT 29.4 3.22 29.63 3.505 ;
      RECT 29.37 3.247 29.63 3.503 ;
      RECT 29.38 3.24 29.635 3.441 ;
      RECT 29.37 3.362 29.64 3.424 ;
      RECT 29.355 3.257 29.635 3.375 ;
      RECT 29.35 3.267 29.635 3.275 ;
      RECT 29.43 4.038 29.435 4.115 ;
      RECT 29.42 4.032 29.43 4.305 ;
      RECT 29.41 4.024 29.42 4.326 ;
      RECT 29.4 4.015 29.41 4.348 ;
      RECT 29.395 4.01 29.4 4.365 ;
      RECT 29.355 4.01 29.395 4.405 ;
      RECT 29.335 4.01 29.355 4.46 ;
      RECT 29.33 4.01 29.335 4.488 ;
      RECT 29.32 4.01 29.33 4.503 ;
      RECT 29.285 4.01 29.32 4.545 ;
      RECT 29.28 4.01 29.285 4.588 ;
      RECT 29.27 4.01 29.28 4.603 ;
      RECT 29.255 4.01 29.27 4.623 ;
      RECT 29.24 4.01 29.255 4.65 ;
      RECT 29.235 4.011 29.24 4.668 ;
      RECT 29.215 4.012 29.235 4.675 ;
      RECT 29.16 4.013 29.215 4.695 ;
      RECT 29.15 4.014 29.16 4.709 ;
      RECT 29.145 4.017 29.15 4.708 ;
      RECT 29.105 4.09 29.145 4.706 ;
      RECT 29.09 4.17 29.105 4.704 ;
      RECT 29.065 4.225 29.09 4.702 ;
      RECT 29.05 4.29 29.065 4.701 ;
      RECT 29.005 4.322 29.05 4.698 ;
      RECT 28.92 4.345 29.005 4.693 ;
      RECT 28.895 4.365 28.92 4.688 ;
      RECT 28.825 4.37 28.895 4.684 ;
      RECT 28.805 4.372 28.825 4.681 ;
      RECT 28.72 4.383 28.805 4.675 ;
      RECT 28.715 4.394 28.72 4.67 ;
      RECT 28.705 4.396 28.715 4.67 ;
      RECT 28.67 4.4 28.705 4.668 ;
      RECT 28.62 4.41 28.67 4.655 ;
      RECT 28.6 4.418 28.62 4.64 ;
      RECT 28.52 4.43 28.6 4.623 ;
      RECT 28.685 3.98 28.855 4.19 ;
      RECT 28.801 3.976 28.855 4.19 ;
      RECT 28.606 3.98 28.855 4.181 ;
      RECT 28.606 3.98 28.86 4.17 ;
      RECT 28.52 3.98 28.86 4.161 ;
      RECT 28.52 3.988 28.87 4.105 ;
      RECT 28.52 4 28.875 4.018 ;
      RECT 28.52 4.007 28.88 4.01 ;
      RECT 28.715 3.978 28.855 4.19 ;
      RECT 28.47 4.923 28.715 5.255 ;
      RECT 28.465 4.915 28.47 5.252 ;
      RECT 28.435 4.935 28.715 5.233 ;
      RECT 28.415 4.967 28.715 5.206 ;
      RECT 28.465 4.92 28.642 5.252 ;
      RECT 28.465 4.917 28.556 5.252 ;
      RECT 28.405 3.265 28.575 3.685 ;
      RECT 28.4 3.265 28.575 3.683 ;
      RECT 28.4 3.265 28.6 3.673 ;
      RECT 28.4 3.265 28.62 3.648 ;
      RECT 28.395 3.265 28.62 3.643 ;
      RECT 28.395 3.265 28.63 3.633 ;
      RECT 28.395 3.265 28.635 3.628 ;
      RECT 28.395 3.27 28.64 3.623 ;
      RECT 28.395 3.302 28.655 3.613 ;
      RECT 28.395 3.372 28.68 3.596 ;
      RECT 28.375 3.372 28.68 3.588 ;
      RECT 28.375 3.432 28.69 3.565 ;
      RECT 28.375 3.472 28.7 3.51 ;
      RECT 28.36 3.265 28.635 3.49 ;
      RECT 28.35 3.28 28.64 3.388 ;
      RECT 27.94 4.67 28.11 5.195 ;
      RECT 27.935 4.67 28.11 5.188 ;
      RECT 27.925 4.67 28.115 5.153 ;
      RECT 27.92 4.68 28.115 5.125 ;
      RECT 27.915 4.7 28.115 5.108 ;
      RECT 27.925 4.675 28.12 5.098 ;
      RECT 27.91 4.72 28.12 5.09 ;
      RECT 27.905 4.74 28.12 5.075 ;
      RECT 27.9 4.77 28.12 5.065 ;
      RECT 27.89 4.815 28.12 5.04 ;
      RECT 27.92 4.685 28.125 5.023 ;
      RECT 27.885 4.867 28.125 5.018 ;
      RECT 27.92 4.695 28.13 4.988 ;
      RECT 27.88 4.9 28.13 4.985 ;
      RECT 27.875 4.925 28.13 4.965 ;
      RECT 27.915 4.712 28.14 4.905 ;
      RECT 27.91 4.734 28.15 4.798 ;
      RECT 27.86 3.981 27.875 4.25 ;
      RECT 27.815 3.965 27.86 4.295 ;
      RECT 27.81 3.953 27.815 4.345 ;
      RECT 27.8 3.949 27.81 4.378 ;
      RECT 27.795 3.946 27.8 4.406 ;
      RECT 27.78 3.948 27.795 4.448 ;
      RECT 27.775 3.952 27.78 4.488 ;
      RECT 27.755 3.957 27.775 4.54 ;
      RECT 27.751 3.962 27.755 4.597 ;
      RECT 27.665 3.981 27.751 4.634 ;
      RECT 27.655 4.002 27.665 4.67 ;
      RECT 27.65 4.01 27.655 4.671 ;
      RECT 27.645 4.052 27.65 4.672 ;
      RECT 27.63 4.14 27.645 4.673 ;
      RECT 27.62 4.29 27.63 4.675 ;
      RECT 27.615 4.335 27.62 4.677 ;
      RECT 27.58 4.377 27.615 4.68 ;
      RECT 27.575 4.395 27.58 4.683 ;
      RECT 27.498 4.401 27.575 4.689 ;
      RECT 27.412 4.415 27.498 4.702 ;
      RECT 27.326 4.429 27.412 4.716 ;
      RECT 27.24 4.443 27.326 4.729 ;
      RECT 27.18 4.455 27.24 4.741 ;
      RECT 27.155 4.462 27.18 4.748 ;
      RECT 27.141 4.465 27.155 4.753 ;
      RECT 27.055 4.473 27.141 4.769 ;
      RECT 27.05 4.48 27.055 4.784 ;
      RECT 27.026 4.48 27.05 4.791 ;
      RECT 26.94 4.483 27.026 4.819 ;
      RECT 26.855 4.487 26.94 4.863 ;
      RECT 26.79 4.491 26.855 4.9 ;
      RECT 26.765 4.494 26.79 4.916 ;
      RECT 26.69 4.507 26.765 4.92 ;
      RECT 26.665 4.525 26.69 4.924 ;
      RECT 26.655 4.532 26.665 4.926 ;
      RECT 26.64 4.535 26.655 4.927 ;
      RECT 26.58 4.547 26.64 4.931 ;
      RECT 26.57 4.561 26.58 4.935 ;
      RECT 26.515 4.571 26.57 4.923 ;
      RECT 26.49 4.592 26.515 4.906 ;
      RECT 26.47 4.612 26.49 4.897 ;
      RECT 26.465 4.625 26.47 4.892 ;
      RECT 26.45 4.637 26.465 4.888 ;
      RECT 27.685 3.292 27.69 3.315 ;
      RECT 27.68 3.283 27.685 3.355 ;
      RECT 27.675 3.281 27.68 3.398 ;
      RECT 27.67 3.272 27.675 3.433 ;
      RECT 27.665 3.262 27.67 3.505 ;
      RECT 27.66 3.252 27.665 3.57 ;
      RECT 27.655 3.249 27.66 3.61 ;
      RECT 27.63 3.243 27.655 3.7 ;
      RECT 27.595 3.231 27.63 3.725 ;
      RECT 27.585 3.222 27.595 3.725 ;
      RECT 27.45 3.22 27.46 3.708 ;
      RECT 27.44 3.22 27.45 3.675 ;
      RECT 27.435 3.22 27.44 3.65 ;
      RECT 27.43 3.22 27.435 3.638 ;
      RECT 27.425 3.22 27.43 3.62 ;
      RECT 27.415 3.22 27.425 3.585 ;
      RECT 27.41 3.222 27.415 3.563 ;
      RECT 27.405 3.228 27.41 3.548 ;
      RECT 27.4 3.234 27.405 3.533 ;
      RECT 27.385 3.246 27.4 3.506 ;
      RECT 27.38 3.257 27.385 3.474 ;
      RECT 27.375 3.267 27.38 3.458 ;
      RECT 27.365 3.275 27.375 3.427 ;
      RECT 27.36 3.285 27.365 3.401 ;
      RECT 27.355 3.342 27.36 3.384 ;
      RECT 27.46 3.22 27.585 3.725 ;
      RECT 27.175 3.907 27.435 4.205 ;
      RECT 27.17 3.914 27.435 4.203 ;
      RECT 27.175 3.909 27.45 4.198 ;
      RECT 27.165 3.922 27.45 4.195 ;
      RECT 27.165 3.927 27.455 4.188 ;
      RECT 27.16 3.935 27.455 4.185 ;
      RECT 27.16 3.952 27.46 3.983 ;
      RECT 27.175 3.904 27.406 4.205 ;
      RECT 27.23 3.903 27.406 4.205 ;
      RECT 27.23 3.9 27.32 4.205 ;
      RECT 27.23 3.897 27.316 4.205 ;
      RECT 26.92 4.17 26.925 4.183 ;
      RECT 26.915 4.137 26.92 4.188 ;
      RECT 26.91 4.092 26.915 4.195 ;
      RECT 26.905 4.047 26.91 4.203 ;
      RECT 26.9 4.015 26.905 4.211 ;
      RECT 26.895 3.975 26.9 4.212 ;
      RECT 26.88 3.955 26.895 4.214 ;
      RECT 26.805 3.937 26.88 4.226 ;
      RECT 26.795 3.93 26.805 4.237 ;
      RECT 26.79 3.93 26.795 4.239 ;
      RECT 26.76 3.936 26.79 4.243 ;
      RECT 26.72 3.949 26.76 4.243 ;
      RECT 26.695 3.96 26.72 4.229 ;
      RECT 26.68 3.966 26.695 4.212 ;
      RECT 26.67 3.968 26.68 4.203 ;
      RECT 26.665 3.969 26.67 4.198 ;
      RECT 26.66 3.97 26.665 4.193 ;
      RECT 26.655 3.971 26.66 4.19 ;
      RECT 26.63 3.976 26.655 4.18 ;
      RECT 26.62 3.992 26.63 4.167 ;
      RECT 26.615 4.012 26.62 4.162 ;
      RECT 26.625 3.405 26.63 3.601 ;
      RECT 26.61 3.369 26.625 3.603 ;
      RECT 26.6 3.351 26.61 3.608 ;
      RECT 26.59 3.337 26.6 3.612 ;
      RECT 26.545 3.321 26.59 3.622 ;
      RECT 26.54 3.311 26.545 3.631 ;
      RECT 26.495 3.3 26.54 3.637 ;
      RECT 26.49 3.288 26.495 3.644 ;
      RECT 26.475 3.283 26.49 3.648 ;
      RECT 26.46 3.275 26.475 3.653 ;
      RECT 26.45 3.268 26.46 3.658 ;
      RECT 26.44 3.265 26.45 3.663 ;
      RECT 26.43 3.265 26.44 3.664 ;
      RECT 26.425 3.262 26.43 3.663 ;
      RECT 26.39 3.257 26.415 3.662 ;
      RECT 26.366 3.253 26.39 3.661 ;
      RECT 26.28 3.244 26.366 3.658 ;
      RECT 26.265 3.236 26.28 3.655 ;
      RECT 26.243 3.235 26.265 3.654 ;
      RECT 26.157 3.235 26.243 3.652 ;
      RECT 26.071 3.235 26.157 3.65 ;
      RECT 25.985 3.235 26.071 3.647 ;
      RECT 25.975 3.235 25.985 3.638 ;
      RECT 25.945 3.235 25.975 3.598 ;
      RECT 25.935 3.245 25.945 3.553 ;
      RECT 25.93 3.285 25.935 3.538 ;
      RECT 25.925 3.3 25.93 3.525 ;
      RECT 25.895 3.38 25.925 3.487 ;
      RECT 26.415 3.26 26.425 3.663 ;
      RECT 26.24 4.025 26.255 4.63 ;
      RECT 26.245 4.02 26.255 4.63 ;
      RECT 26.41 4.02 26.415 4.203 ;
      RECT 26.4 4.02 26.41 4.233 ;
      RECT 26.385 4.02 26.4 4.293 ;
      RECT 26.38 4.02 26.385 4.338 ;
      RECT 26.375 4.02 26.38 4.368 ;
      RECT 26.37 4.02 26.375 4.388 ;
      RECT 26.36 4.02 26.37 4.423 ;
      RECT 26.345 4.02 26.36 4.455 ;
      RECT 26.3 4.02 26.345 4.483 ;
      RECT 26.295 4.02 26.3 4.513 ;
      RECT 26.29 4.02 26.295 4.525 ;
      RECT 26.285 4.02 26.29 4.533 ;
      RECT 26.275 4.02 26.285 4.548 ;
      RECT 26.27 4.02 26.275 4.57 ;
      RECT 26.26 4.02 26.27 4.593 ;
      RECT 26.255 4.02 26.26 4.613 ;
      RECT 26.22 4.035 26.24 4.63 ;
      RECT 26.195 4.052 26.22 4.63 ;
      RECT 26.19 4.062 26.195 4.63 ;
      RECT 26.16 4.077 26.19 4.63 ;
      RECT 26.085 4.119 26.16 4.63 ;
      RECT 26.08 4.15 26.085 4.613 ;
      RECT 26.075 4.154 26.08 4.595 ;
      RECT 26.07 4.158 26.075 4.558 ;
      RECT 26.065 4.342 26.07 4.525 ;
      RECT 25.55 4.531 25.636 5.096 ;
      RECT 25.505 4.533 25.67 5.09 ;
      RECT 25.636 4.53 25.67 5.09 ;
      RECT 25.55 4.532 25.755 5.084 ;
      RECT 25.505 4.542 25.765 5.08 ;
      RECT 25.48 4.534 25.755 5.076 ;
      RECT 25.475 4.537 25.755 5.071 ;
      RECT 25.45 4.552 25.765 5.065 ;
      RECT 25.45 4.577 25.805 5.06 ;
      RECT 25.41 4.585 25.805 5.035 ;
      RECT 25.41 4.612 25.82 5.033 ;
      RECT 25.41 4.642 25.83 5.02 ;
      RECT 25.405 4.787 25.83 5.008 ;
      RECT 25.41 4.716 25.85 5.005 ;
      RECT 25.41 4.773 25.855 4.813 ;
      RECT 25.6 4.052 25.77 4.23 ;
      RECT 25.55 3.991 25.6 4.215 ;
      RECT 25.285 3.971 25.55 4.2 ;
      RECT 25.245 4.035 25.72 4.2 ;
      RECT 25.245 4.025 25.675 4.2 ;
      RECT 25.245 4.022 25.665 4.2 ;
      RECT 25.245 4.01 25.655 4.2 ;
      RECT 25.245 3.995 25.6 4.2 ;
      RECT 25.285 3.967 25.486 4.2 ;
      RECT 25.295 3.945 25.486 4.2 ;
      RECT 25.32 3.93 25.4 4.2 ;
      RECT 25.075 4.46 25.195 4.905 ;
      RECT 25.06 4.46 25.195 4.904 ;
      RECT 25.015 4.482 25.195 4.899 ;
      RECT 24.975 4.531 25.195 4.893 ;
      RECT 24.975 4.531 25.2 4.868 ;
      RECT 24.975 4.531 25.22 4.758 ;
      RECT 24.97 4.561 25.22 4.755 ;
      RECT 25.06 4.46 25.23 4.65 ;
      RECT 24.72 3.245 24.725 3.69 ;
      RECT 24.53 3.245 24.55 3.655 ;
      RECT 24.5 3.245 24.505 3.63 ;
      RECT 25.18 3.552 25.195 3.74 ;
      RECT 25.175 3.537 25.18 3.746 ;
      RECT 25.155 3.51 25.175 3.749 ;
      RECT 25.105 3.477 25.155 3.758 ;
      RECT 25.075 3.457 25.105 3.762 ;
      RECT 25.056 3.445 25.075 3.758 ;
      RECT 24.97 3.417 25.056 3.748 ;
      RECT 24.96 3.392 24.97 3.738 ;
      RECT 24.89 3.36 24.96 3.73 ;
      RECT 24.865 3.32 24.89 3.722 ;
      RECT 24.845 3.302 24.865 3.716 ;
      RECT 24.835 3.292 24.845 3.713 ;
      RECT 24.825 3.285 24.835 3.711 ;
      RECT 24.805 3.272 24.825 3.708 ;
      RECT 24.795 3.262 24.805 3.705 ;
      RECT 24.785 3.255 24.795 3.703 ;
      RECT 24.735 3.247 24.785 3.697 ;
      RECT 24.725 3.245 24.735 3.691 ;
      RECT 24.695 3.245 24.72 3.688 ;
      RECT 24.666 3.245 24.695 3.683 ;
      RECT 24.58 3.245 24.666 3.673 ;
      RECT 24.55 3.245 24.58 3.66 ;
      RECT 24.505 3.245 24.53 3.643 ;
      RECT 24.49 3.245 24.5 3.625 ;
      RECT 24.47 3.252 24.49 3.61 ;
      RECT 24.465 3.267 24.47 3.598 ;
      RECT 24.46 3.272 24.465 3.538 ;
      RECT 24.455 3.277 24.46 3.38 ;
      RECT 24.45 3.28 24.455 3.298 ;
      RECT 24.715 3.965 24.801 4.286 ;
      RECT 24.715 3.965 24.835 4.279 ;
      RECT 24.665 3.965 24.835 4.275 ;
      RECT 24.665 3.967 24.921 4.273 ;
      RECT 24.665 3.969 24.945 4.267 ;
      RECT 24.665 3.976 24.955 4.266 ;
      RECT 24.665 3.985 24.96 4.263 ;
      RECT 24.665 3.991 24.965 4.258 ;
      RECT 24.665 4.035 24.97 4.255 ;
      RECT 24.665 4.127 24.975 4.252 ;
      RECT 24.19 4.57 24.225 4.89 ;
      RECT 24.775 4.755 24.78 4.937 ;
      RECT 24.73 4.637 24.775 4.956 ;
      RECT 24.715 4.614 24.73 4.979 ;
      RECT 24.705 4.604 24.715 4.989 ;
      RECT 24.685 4.599 24.705 5.002 ;
      RECT 24.66 4.597 24.685 5.023 ;
      RECT 24.641 4.596 24.66 5.035 ;
      RECT 24.555 4.593 24.641 5.035 ;
      RECT 24.485 4.588 24.555 5.023 ;
      RECT 24.41 4.584 24.485 4.998 ;
      RECT 24.345 4.58 24.41 4.965 ;
      RECT 24.275 4.577 24.345 4.925 ;
      RECT 24.245 4.573 24.275 4.9 ;
      RECT 24.225 4.571 24.245 4.893 ;
      RECT 24.141 4.569 24.19 4.891 ;
      RECT 24.055 4.566 24.141 4.892 ;
      RECT 23.98 4.565 24.055 4.894 ;
      RECT 23.895 4.565 23.98 4.92 ;
      RECT 23.818 4.566 23.895 4.945 ;
      RECT 23.732 4.567 23.818 4.945 ;
      RECT 23.646 4.567 23.732 4.945 ;
      RECT 23.56 4.568 23.646 4.945 ;
      RECT 23.54 4.569 23.56 4.937 ;
      RECT 23.525 4.575 23.54 4.922 ;
      RECT 23.49 4.595 23.525 4.902 ;
      RECT 23.48 4.615 23.49 4.884 ;
      RECT 24.45 3.92 24.455 4.19 ;
      RECT 24.445 3.911 24.45 4.195 ;
      RECT 24.435 3.901 24.445 4.207 ;
      RECT 24.43 3.89 24.435 4.218 ;
      RECT 24.41 3.884 24.43 4.236 ;
      RECT 24.365 3.881 24.41 4.285 ;
      RECT 24.35 3.88 24.365 4.33 ;
      RECT 24.345 3.88 24.35 4.343 ;
      RECT 24.335 3.88 24.345 4.355 ;
      RECT 24.33 3.881 24.335 4.37 ;
      RECT 24.31 3.889 24.33 4.375 ;
      RECT 24.28 3.905 24.31 4.375 ;
      RECT 24.27 3.917 24.275 4.375 ;
      RECT 24.235 3.932 24.27 4.375 ;
      RECT 24.205 3.952 24.235 4.375 ;
      RECT 24.195 3.977 24.205 4.375 ;
      RECT 24.19 4.005 24.195 4.375 ;
      RECT 24.185 4.035 24.19 4.375 ;
      RECT 24.18 4.052 24.185 4.375 ;
      RECT 24.17 4.08 24.18 4.375 ;
      RECT 24.16 4.115 24.17 4.375 ;
      RECT 24.155 4.15 24.16 4.375 ;
      RECT 24.275 3.915 24.28 4.375 ;
      RECT 23.79 4.017 23.975 4.19 ;
      RECT 23.75 3.935 23.935 4.188 ;
      RECT 23.711 3.94 23.935 4.184 ;
      RECT 23.625 3.949 23.935 4.179 ;
      RECT 23.541 3.965 23.94 4.174 ;
      RECT 23.455 3.985 23.965 4.168 ;
      RECT 23.455 4.005 23.97 4.168 ;
      RECT 23.541 3.975 23.965 4.174 ;
      RECT 23.625 3.95 23.94 4.179 ;
      RECT 23.79 3.932 23.935 4.19 ;
      RECT 23.79 3.927 23.89 4.19 ;
      RECT 23.876 3.921 23.89 4.19 ;
      RECT 23.265 3.245 23.27 3.644 ;
      RECT 23.01 3.245 23.045 3.642 ;
      RECT 22.605 3.28 22.61 3.636 ;
      RECT 23.35 3.283 23.355 3.538 ;
      RECT 23.345 3.281 23.35 3.544 ;
      RECT 23.34 3.28 23.345 3.551 ;
      RECT 23.315 3.273 23.34 3.575 ;
      RECT 23.31 3.266 23.315 3.599 ;
      RECT 23.305 3.262 23.31 3.608 ;
      RECT 23.295 3.257 23.305 3.621 ;
      RECT 23.29 3.254 23.295 3.63 ;
      RECT 23.285 3.252 23.29 3.635 ;
      RECT 23.27 3.248 23.285 3.645 ;
      RECT 23.255 3.242 23.265 3.644 ;
      RECT 23.217 3.24 23.255 3.644 ;
      RECT 23.131 3.242 23.217 3.644 ;
      RECT 23.045 3.244 23.131 3.643 ;
      RECT 22.974 3.245 23.01 3.642 ;
      RECT 22.888 3.247 22.974 3.642 ;
      RECT 22.802 3.249 22.888 3.641 ;
      RECT 22.716 3.251 22.802 3.641 ;
      RECT 22.63 3.254 22.716 3.64 ;
      RECT 22.62 3.26 22.63 3.639 ;
      RECT 22.61 3.272 22.62 3.637 ;
      RECT 22.55 3.307 22.605 3.633 ;
      RECT 22.545 3.337 22.55 3.395 ;
      RECT 23.29 4.417 23.305 4.61 ;
      RECT 23.285 4.385 23.29 4.61 ;
      RECT 23.275 4.36 23.285 4.61 ;
      RECT 23.27 4.332 23.275 4.61 ;
      RECT 23.24 4.255 23.27 4.61 ;
      RECT 23.215 4.137 23.24 4.61 ;
      RECT 23.21 4.075 23.215 4.61 ;
      RECT 23.2 4.062 23.21 4.61 ;
      RECT 23.18 4.052 23.2 4.61 ;
      RECT 23.165 4.035 23.18 4.61 ;
      RECT 23.135 4.023 23.165 4.61 ;
      RECT 23.13 4.022 23.135 4.555 ;
      RECT 23.125 4.022 23.13 4.513 ;
      RECT 23.11 4.021 23.125 4.465 ;
      RECT 23.095 4.021 23.11 4.403 ;
      RECT 23.075 4.021 23.095 4.363 ;
      RECT 23.07 4.021 23.075 4.348 ;
      RECT 23.045 4.02 23.07 4.343 ;
      RECT 22.975 4.019 23.045 4.33 ;
      RECT 22.96 4.018 22.975 4.315 ;
      RECT 22.93 4.017 22.96 4.298 ;
      RECT 22.925 4.017 22.93 4.283 ;
      RECT 22.875 4.016 22.925 4.263 ;
      RECT 22.81 4.015 22.875 4.218 ;
      RECT 22.805 4.015 22.81 4.19 ;
      RECT 22.89 4.552 22.895 4.809 ;
      RECT 22.87 4.471 22.89 4.826 ;
      RECT 22.85 4.465 22.87 4.855 ;
      RECT 22.79 4.452 22.85 4.875 ;
      RECT 22.745 4.436 22.79 4.876 ;
      RECT 22.661 4.424 22.745 4.864 ;
      RECT 22.575 4.411 22.661 4.848 ;
      RECT 22.565 4.404 22.575 4.84 ;
      RECT 22.52 4.401 22.565 4.78 ;
      RECT 22.5 4.397 22.52 4.695 ;
      RECT 22.485 4.395 22.5 4.648 ;
      RECT 22.455 4.392 22.485 4.618 ;
      RECT 22.42 4.388 22.455 4.595 ;
      RECT 22.377 4.383 22.42 4.583 ;
      RECT 22.291 4.374 22.377 4.592 ;
      RECT 22.205 4.363 22.291 4.604 ;
      RECT 22.14 4.354 22.205 4.613 ;
      RECT 22.12 4.345 22.14 4.618 ;
      RECT 22.115 4.338 22.12 4.62 ;
      RECT 22.075 4.323 22.115 4.617 ;
      RECT 22.055 4.302 22.075 4.612 ;
      RECT 22.04 4.29 22.055 4.605 ;
      RECT 22.035 4.282 22.04 4.598 ;
      RECT 22.02 4.262 22.035 4.591 ;
      RECT 22.015 4.125 22.02 4.585 ;
      RECT 21.935 4.014 22.015 4.557 ;
      RECT 21.926 4.007 21.935 4.523 ;
      RECT 21.84 4.001 21.926 4.448 ;
      RECT 21.815 3.992 21.84 4.36 ;
      RECT 21.785 3.987 21.815 4.335 ;
      RECT 21.72 3.996 21.785 4.32 ;
      RECT 21.7 4.012 21.72 4.295 ;
      RECT 21.69 4.018 21.7 4.243 ;
      RECT 21.67 4.04 21.69 4.125 ;
      RECT 22.325 4.005 22.495 4.19 ;
      RECT 22.325 4.005 22.53 4.188 ;
      RECT 22.375 3.915 22.545 4.179 ;
      RECT 22.325 4.072 22.55 4.172 ;
      RECT 22.34 3.95 22.545 4.179 ;
      RECT 21.54 4.683 21.605 5.126 ;
      RECT 21.48 4.708 21.605 5.124 ;
      RECT 21.48 4.708 21.66 5.118 ;
      RECT 21.465 4.733 21.66 5.117 ;
      RECT 21.605 4.67 21.68 5.114 ;
      RECT 21.54 4.695 21.76 5.108 ;
      RECT 21.465 4.734 21.805 5.102 ;
      RECT 21.45 4.761 21.805 5.093 ;
      RECT 21.465 4.754 21.825 5.085 ;
      RECT 21.45 4.763 21.83 5.068 ;
      RECT 21.445 4.78 21.83 4.895 ;
      RECT 21.45 3.502 21.485 3.74 ;
      RECT 21.45 3.502 21.515 3.739 ;
      RECT 21.45 3.502 21.63 3.735 ;
      RECT 21.45 3.502 21.685 3.713 ;
      RECT 21.46 3.445 21.74 3.613 ;
      RECT 21.565 3.285 21.595 3.736 ;
      RECT 21.595 3.28 21.775 3.493 ;
      RECT 21.465 3.421 21.775 3.493 ;
      RECT 21.515 3.317 21.565 3.737 ;
      RECT 21.485 3.373 21.775 3.493 ;
      RECT 19.985 3.035 20.155 4.225 ;
      RECT 19.985 3.035 20.455 3.205 ;
      RECT 19.985 9.405 20.455 9.575 ;
      RECT 19.985 8.385 20.155 9.575 ;
      RECT 18.995 3.035 19.165 4.225 ;
      RECT 18.995 3.035 19.465 3.205 ;
      RECT 18.995 9.405 19.465 9.575 ;
      RECT 18.995 8.385 19.165 9.575 ;
      RECT 17.145 3.93 17.315 5.16 ;
      RECT 17.2 2.15 17.37 4.1 ;
      RECT 17.145 1.87 17.315 2.32 ;
      RECT 17.145 10.29 17.315 10.74 ;
      RECT 17.2 8.51 17.37 10.46 ;
      RECT 17.145 7.45 17.315 8.68 ;
      RECT 16.625 1.87 16.795 5.16 ;
      RECT 16.625 3.37 17.03 3.7 ;
      RECT 16.625 2.53 17.03 2.86 ;
      RECT 16.625 7.45 16.795 10.74 ;
      RECT 16.625 9.75 17.03 10.08 ;
      RECT 16.625 8.91 17.03 9.24 ;
      RECT 14.725 4.687 14.74 4.738 ;
      RECT 14.72 4.667 14.725 4.785 ;
      RECT 14.705 4.657 14.72 4.853 ;
      RECT 14.68 4.637 14.705 4.908 ;
      RECT 14.64 4.622 14.68 4.928 ;
      RECT 14.595 4.616 14.64 4.956 ;
      RECT 14.525 4.606 14.595 4.973 ;
      RECT 14.505 4.598 14.525 4.973 ;
      RECT 14.445 4.592 14.505 4.965 ;
      RECT 14.386 4.583 14.445 4.953 ;
      RECT 14.3 4.572 14.386 4.936 ;
      RECT 14.278 4.563 14.3 4.924 ;
      RECT 14.192 4.556 14.278 4.911 ;
      RECT 14.106 4.543 14.192 4.892 ;
      RECT 14.02 4.531 14.106 4.872 ;
      RECT 13.99 4.52 14.02 4.859 ;
      RECT 13.94 4.506 13.99 4.851 ;
      RECT 13.92 4.495 13.94 4.843 ;
      RECT 13.871 4.484 13.92 4.835 ;
      RECT 13.785 4.463 13.871 4.82 ;
      RECT 13.74 4.45 13.785 4.805 ;
      RECT 13.695 4.45 13.74 4.785 ;
      RECT 13.64 4.45 13.695 4.72 ;
      RECT 13.615 4.45 13.64 4.643 ;
      RECT 14.14 4.187 14.31 4.37 ;
      RECT 14.14 4.187 14.325 4.328 ;
      RECT 14.14 4.187 14.33 4.27 ;
      RECT 14.2 3.955 14.335 4.246 ;
      RECT 14.2 3.959 14.34 4.229 ;
      RECT 14.145 4.122 14.34 4.229 ;
      RECT 14.17 3.967 14.31 4.37 ;
      RECT 14.17 3.971 14.35 4.17 ;
      RECT 14.155 4.057 14.35 4.17 ;
      RECT 14.165 3.987 14.31 4.37 ;
      RECT 14.165 3.99 14.36 4.083 ;
      RECT 14.16 4.007 14.36 4.083 ;
      RECT 13.93 3.227 14.1 3.71 ;
      RECT 13.925 3.222 14.075 3.7 ;
      RECT 13.925 3.229 14.105 3.694 ;
      RECT 13.915 3.223 14.075 3.673 ;
      RECT 13.915 3.239 14.12 3.632 ;
      RECT 13.885 3.224 14.075 3.595 ;
      RECT 13.885 3.254 14.13 3.535 ;
      RECT 13.88 3.226 14.075 3.533 ;
      RECT 13.86 3.235 14.105 3.49 ;
      RECT 13.835 3.251 14.12 3.402 ;
      RECT 13.835 3.27 14.145 3.393 ;
      RECT 13.83 3.307 14.145 3.345 ;
      RECT 13.835 3.287 14.15 3.313 ;
      RECT 13.93 3.221 14.04 3.71 ;
      RECT 14.016 3.22 14.04 3.71 ;
      RECT 13.25 4.005 13.255 4.216 ;
      RECT 13.85 4.005 13.855 4.19 ;
      RECT 13.915 4.045 13.92 4.158 ;
      RECT 13.91 4.037 13.915 4.164 ;
      RECT 13.905 4.027 13.91 4.172 ;
      RECT 13.9 4.017 13.905 4.181 ;
      RECT 13.895 4.007 13.9 4.185 ;
      RECT 13.855 4.005 13.895 4.188 ;
      RECT 13.827 4.004 13.85 4.192 ;
      RECT 13.741 4.001 13.827 4.199 ;
      RECT 13.655 3.997 13.741 4.21 ;
      RECT 13.635 3.995 13.655 4.216 ;
      RECT 13.617 3.994 13.635 4.219 ;
      RECT 13.531 3.992 13.617 4.226 ;
      RECT 13.445 3.987 13.531 4.239 ;
      RECT 13.426 3.984 13.445 4.244 ;
      RECT 13.34 3.982 13.426 4.235 ;
      RECT 13.33 3.982 13.34 4.228 ;
      RECT 13.255 3.995 13.33 4.222 ;
      RECT 13.24 4.006 13.25 4.216 ;
      RECT 13.23 4.008 13.24 4.215 ;
      RECT 13.22 4.012 13.23 4.211 ;
      RECT 13.215 4.015 13.22 4.205 ;
      RECT 13.205 4.017 13.215 4.199 ;
      RECT 13.2 4.02 13.205 4.193 ;
      RECT 13.18 4.606 13.185 4.81 ;
      RECT 13.165 4.593 13.18 4.903 ;
      RECT 13.15 4.574 13.165 5.18 ;
      RECT 13.115 4.54 13.15 5.18 ;
      RECT 13.111 4.51 13.115 5.18 ;
      RECT 13.025 4.392 13.111 5.18 ;
      RECT 13.015 4.267 13.025 5.18 ;
      RECT 13 4.235 13.015 5.18 ;
      RECT 12.995 4.21 13 5.18 ;
      RECT 12.99 4.2 12.995 5.136 ;
      RECT 12.975 4.172 12.99 5.041 ;
      RECT 12.96 4.138 12.975 4.94 ;
      RECT 12.955 4.116 12.96 4.893 ;
      RECT 12.95 4.105 12.955 4.863 ;
      RECT 12.945 4.095 12.95 4.829 ;
      RECT 12.935 4.082 12.945 4.797 ;
      RECT 12.91 4.058 12.935 4.723 ;
      RECT 12.905 4.038 12.91 4.648 ;
      RECT 12.9 4.032 12.905 4.623 ;
      RECT 12.895 4.027 12.9 4.588 ;
      RECT 12.89 4.022 12.895 4.563 ;
      RECT 12.885 4.02 12.89 4.543 ;
      RECT 12.88 4.02 12.885 4.528 ;
      RECT 12.875 4.02 12.88 4.488 ;
      RECT 12.865 4.02 12.875 4.46 ;
      RECT 12.855 4.02 12.865 4.405 ;
      RECT 12.84 4.02 12.855 4.343 ;
      RECT 12.835 4.019 12.84 4.288 ;
      RECT 12.82 4.018 12.835 4.268 ;
      RECT 12.76 4.016 12.82 4.242 ;
      RECT 12.725 4.017 12.76 4.222 ;
      RECT 12.72 4.019 12.725 4.212 ;
      RECT 12.71 4.038 12.72 4.202 ;
      RECT 12.705 4.065 12.71 4.133 ;
      RECT 12.82 3.49 12.99 3.735 ;
      RECT 12.855 3.261 12.99 3.735 ;
      RECT 12.855 3.263 13 3.73 ;
      RECT 12.855 3.265 13.025 3.718 ;
      RECT 12.855 3.268 13.05 3.7 ;
      RECT 12.855 3.273 13.1 3.673 ;
      RECT 12.855 3.278 13.12 3.638 ;
      RECT 12.835 3.28 13.13 3.613 ;
      RECT 12.825 3.375 13.13 3.613 ;
      RECT 12.855 3.26 12.965 3.735 ;
      RECT 12.865 3.257 12.96 3.735 ;
      RECT 12.385 4.522 12.575 4.88 ;
      RECT 12.385 4.534 12.61 4.879 ;
      RECT 12.385 4.562 12.63 4.877 ;
      RECT 12.385 4.587 12.635 4.876 ;
      RECT 12.385 4.645 12.65 4.875 ;
      RECT 12.37 4.518 12.53 4.86 ;
      RECT 12.35 4.527 12.575 4.813 ;
      RECT 12.325 4.538 12.61 4.75 ;
      RECT 12.325 4.622 12.645 4.75 ;
      RECT 12.325 4.597 12.64 4.75 ;
      RECT 12.385 4.513 12.53 4.88 ;
      RECT 12.471 4.512 12.53 4.88 ;
      RECT 12.471 4.511 12.515 4.88 ;
      RECT 11.865 7.45 12.035 10.74 ;
      RECT 11.865 9.75 12.27 10.08 ;
      RECT 11.865 8.91 12.27 9.24 ;
      RECT 12.17 4.027 12.175 4.405 ;
      RECT 12.165 3.995 12.17 4.405 ;
      RECT 12.16 3.967 12.165 4.405 ;
      RECT 12.155 3.947 12.16 4.405 ;
      RECT 12.1 3.93 12.155 4.405 ;
      RECT 12.06 3.915 12.1 4.405 ;
      RECT 12.005 3.902 12.06 4.405 ;
      RECT 11.97 3.893 12.005 4.405 ;
      RECT 11.966 3.891 11.97 4.404 ;
      RECT 11.88 3.887 11.966 4.387 ;
      RECT 11.795 3.879 11.88 4.35 ;
      RECT 11.785 3.875 11.795 4.323 ;
      RECT 11.775 3.875 11.785 4.305 ;
      RECT 11.765 3.877 11.775 4.288 ;
      RECT 11.76 3.882 11.765 4.274 ;
      RECT 11.755 3.886 11.76 4.261 ;
      RECT 11.745 3.891 11.755 4.245 ;
      RECT 11.73 3.905 11.745 4.22 ;
      RECT 11.725 3.911 11.73 4.2 ;
      RECT 11.72 3.913 11.725 4.193 ;
      RECT 11.715 3.917 11.72 4.068 ;
      RECT 11.895 4.717 12.14 5.18 ;
      RECT 11.815 4.69 12.135 5.176 ;
      RECT 11.745 4.725 12.14 5.169 ;
      RECT 11.535 4.98 12.14 5.165 ;
      RECT 11.715 4.748 12.14 5.165 ;
      RECT 11.555 4.94 12.14 5.165 ;
      RECT 11.705 4.76 12.14 5.165 ;
      RECT 11.59 4.877 12.14 5.165 ;
      RECT 11.645 4.802 12.14 5.165 ;
      RECT 11.895 4.667 12.135 5.18 ;
      RECT 11.925 4.66 12.135 5.18 ;
      RECT 11.915 4.662 12.135 5.18 ;
      RECT 11.925 4.657 12.055 5.18 ;
      RECT 11.48 3.22 11.566 3.659 ;
      RECT 11.475 3.22 11.566 3.657 ;
      RECT 11.475 3.22 11.635 3.656 ;
      RECT 11.475 3.22 11.665 3.653 ;
      RECT 11.46 3.227 11.665 3.644 ;
      RECT 11.46 3.227 11.67 3.64 ;
      RECT 11.455 3.237 11.67 3.633 ;
      RECT 11.45 3.242 11.67 3.608 ;
      RECT 11.45 3.242 11.685 3.59 ;
      RECT 11.475 3.22 11.705 3.505 ;
      RECT 11.445 3.247 11.705 3.503 ;
      RECT 11.455 3.24 11.71 3.441 ;
      RECT 11.445 3.362 11.715 3.424 ;
      RECT 11.43 3.257 11.71 3.375 ;
      RECT 11.425 3.267 11.71 3.275 ;
      RECT 11.505 4.038 11.51 4.115 ;
      RECT 11.495 4.032 11.505 4.305 ;
      RECT 11.485 4.024 11.495 4.326 ;
      RECT 11.475 4.015 11.485 4.348 ;
      RECT 11.47 4.01 11.475 4.365 ;
      RECT 11.43 4.01 11.47 4.405 ;
      RECT 11.41 4.01 11.43 4.46 ;
      RECT 11.405 4.01 11.41 4.488 ;
      RECT 11.395 4.01 11.405 4.503 ;
      RECT 11.36 4.01 11.395 4.545 ;
      RECT 11.355 4.01 11.36 4.588 ;
      RECT 11.345 4.01 11.355 4.603 ;
      RECT 11.33 4.01 11.345 4.623 ;
      RECT 11.315 4.01 11.33 4.65 ;
      RECT 11.31 4.011 11.315 4.668 ;
      RECT 11.29 4.012 11.31 4.675 ;
      RECT 11.235 4.013 11.29 4.695 ;
      RECT 11.225 4.014 11.235 4.709 ;
      RECT 11.22 4.017 11.225 4.708 ;
      RECT 11.18 4.09 11.22 4.706 ;
      RECT 11.165 4.17 11.18 4.704 ;
      RECT 11.14 4.225 11.165 4.702 ;
      RECT 11.125 4.29 11.14 4.701 ;
      RECT 11.08 4.322 11.125 4.698 ;
      RECT 10.995 4.345 11.08 4.693 ;
      RECT 10.97 4.365 10.995 4.688 ;
      RECT 10.9 4.37 10.97 4.684 ;
      RECT 10.88 4.372 10.9 4.681 ;
      RECT 10.795 4.383 10.88 4.675 ;
      RECT 10.79 4.394 10.795 4.67 ;
      RECT 10.78 4.396 10.79 4.67 ;
      RECT 10.745 4.4 10.78 4.668 ;
      RECT 10.695 4.41 10.745 4.655 ;
      RECT 10.675 4.418 10.695 4.64 ;
      RECT 10.595 4.43 10.675 4.623 ;
      RECT 10.76 3.98 10.93 4.19 ;
      RECT 10.876 3.976 10.93 4.19 ;
      RECT 10.681 3.98 10.93 4.181 ;
      RECT 10.681 3.98 10.935 4.17 ;
      RECT 10.595 3.98 10.935 4.161 ;
      RECT 10.595 3.988 10.945 4.105 ;
      RECT 10.595 4 10.95 4.018 ;
      RECT 10.595 4.007 10.955 4.01 ;
      RECT 10.79 3.978 10.93 4.19 ;
      RECT 10.545 4.923 10.79 5.255 ;
      RECT 10.54 4.915 10.545 5.252 ;
      RECT 10.51 4.935 10.79 5.233 ;
      RECT 10.49 4.967 10.79 5.206 ;
      RECT 10.54 4.92 10.717 5.252 ;
      RECT 10.54 4.917 10.631 5.252 ;
      RECT 10.48 3.265 10.65 3.685 ;
      RECT 10.475 3.265 10.65 3.683 ;
      RECT 10.475 3.265 10.675 3.673 ;
      RECT 10.475 3.265 10.695 3.648 ;
      RECT 10.47 3.265 10.695 3.643 ;
      RECT 10.47 3.265 10.705 3.633 ;
      RECT 10.47 3.265 10.71 3.628 ;
      RECT 10.47 3.27 10.715 3.623 ;
      RECT 10.47 3.302 10.73 3.613 ;
      RECT 10.47 3.372 10.755 3.596 ;
      RECT 10.45 3.372 10.755 3.588 ;
      RECT 10.45 3.432 10.765 3.565 ;
      RECT 10.45 3.472 10.775 3.51 ;
      RECT 10.435 3.265 10.71 3.49 ;
      RECT 10.425 3.28 10.715 3.388 ;
      RECT 10.015 4.67 10.185 5.195 ;
      RECT 10.01 4.67 10.185 5.188 ;
      RECT 10 4.67 10.19 5.153 ;
      RECT 9.995 4.68 10.19 5.125 ;
      RECT 9.99 4.7 10.19 5.108 ;
      RECT 10 4.675 10.195 5.098 ;
      RECT 9.985 4.72 10.195 5.09 ;
      RECT 9.98 4.74 10.195 5.075 ;
      RECT 9.975 4.77 10.195 5.065 ;
      RECT 9.965 4.815 10.195 5.04 ;
      RECT 9.995 4.685 10.2 5.023 ;
      RECT 9.96 4.867 10.2 5.018 ;
      RECT 9.995 4.695 10.205 4.988 ;
      RECT 9.955 4.9 10.205 4.985 ;
      RECT 9.95 4.925 10.205 4.965 ;
      RECT 9.99 4.712 10.215 4.905 ;
      RECT 9.985 4.734 10.225 4.798 ;
      RECT 9.935 3.981 9.95 4.25 ;
      RECT 9.89 3.965 9.935 4.295 ;
      RECT 9.885 3.953 9.89 4.345 ;
      RECT 9.875 3.949 9.885 4.378 ;
      RECT 9.87 3.946 9.875 4.406 ;
      RECT 9.855 3.948 9.87 4.448 ;
      RECT 9.85 3.952 9.855 4.488 ;
      RECT 9.83 3.957 9.85 4.54 ;
      RECT 9.826 3.962 9.83 4.597 ;
      RECT 9.74 3.981 9.826 4.634 ;
      RECT 9.73 4.002 9.74 4.67 ;
      RECT 9.725 4.01 9.73 4.671 ;
      RECT 9.72 4.052 9.725 4.672 ;
      RECT 9.705 4.14 9.72 4.673 ;
      RECT 9.695 4.29 9.705 4.675 ;
      RECT 9.69 4.335 9.695 4.677 ;
      RECT 9.655 4.377 9.69 4.68 ;
      RECT 9.65 4.395 9.655 4.683 ;
      RECT 9.573 4.401 9.65 4.689 ;
      RECT 9.487 4.415 9.573 4.702 ;
      RECT 9.401 4.429 9.487 4.716 ;
      RECT 9.315 4.443 9.401 4.729 ;
      RECT 9.255 4.455 9.315 4.741 ;
      RECT 9.23 4.462 9.255 4.748 ;
      RECT 9.216 4.465 9.23 4.753 ;
      RECT 9.13 4.473 9.216 4.769 ;
      RECT 9.125 4.48 9.13 4.784 ;
      RECT 9.101 4.48 9.125 4.791 ;
      RECT 9.015 4.483 9.101 4.819 ;
      RECT 8.93 4.487 9.015 4.863 ;
      RECT 8.865 4.491 8.93 4.9 ;
      RECT 8.84 4.494 8.865 4.916 ;
      RECT 8.765 4.507 8.84 4.92 ;
      RECT 8.74 4.525 8.765 4.924 ;
      RECT 8.73 4.532 8.74 4.926 ;
      RECT 8.715 4.535 8.73 4.927 ;
      RECT 8.655 4.547 8.715 4.931 ;
      RECT 8.645 4.561 8.655 4.935 ;
      RECT 8.59 4.571 8.645 4.923 ;
      RECT 8.565 4.592 8.59 4.906 ;
      RECT 8.545 4.612 8.565 4.897 ;
      RECT 8.54 4.625 8.545 4.892 ;
      RECT 8.525 4.637 8.54 4.888 ;
      RECT 9.76 3.292 9.765 3.315 ;
      RECT 9.755 3.283 9.76 3.355 ;
      RECT 9.75 3.281 9.755 3.398 ;
      RECT 9.745 3.272 9.75 3.433 ;
      RECT 9.74 3.262 9.745 3.505 ;
      RECT 9.735 3.252 9.74 3.57 ;
      RECT 9.73 3.249 9.735 3.61 ;
      RECT 9.705 3.243 9.73 3.7 ;
      RECT 9.67 3.231 9.705 3.725 ;
      RECT 9.66 3.222 9.67 3.725 ;
      RECT 9.525 3.22 9.535 3.708 ;
      RECT 9.515 3.22 9.525 3.675 ;
      RECT 9.51 3.22 9.515 3.65 ;
      RECT 9.505 3.22 9.51 3.638 ;
      RECT 9.5 3.22 9.505 3.62 ;
      RECT 9.49 3.22 9.5 3.585 ;
      RECT 9.485 3.222 9.49 3.563 ;
      RECT 9.48 3.228 9.485 3.548 ;
      RECT 9.475 3.234 9.48 3.533 ;
      RECT 9.46 3.246 9.475 3.506 ;
      RECT 9.455 3.257 9.46 3.474 ;
      RECT 9.45 3.267 9.455 3.458 ;
      RECT 9.44 3.275 9.45 3.427 ;
      RECT 9.435 3.285 9.44 3.401 ;
      RECT 9.43 3.342 9.435 3.384 ;
      RECT 9.535 3.22 9.66 3.725 ;
      RECT 9.25 3.907 9.51 4.205 ;
      RECT 9.245 3.914 9.51 4.203 ;
      RECT 9.25 3.909 9.525 4.198 ;
      RECT 9.24 3.922 9.525 4.195 ;
      RECT 9.24 3.927 9.53 4.188 ;
      RECT 9.235 3.935 9.53 4.185 ;
      RECT 9.235 3.952 9.535 3.983 ;
      RECT 9.25 3.904 9.481 4.205 ;
      RECT 9.305 3.903 9.481 4.205 ;
      RECT 9.305 3.9 9.395 4.205 ;
      RECT 9.305 3.897 9.391 4.205 ;
      RECT 8.995 4.17 9 4.183 ;
      RECT 8.99 4.137 8.995 4.188 ;
      RECT 8.985 4.092 8.99 4.195 ;
      RECT 8.98 4.047 8.985 4.203 ;
      RECT 8.975 4.015 8.98 4.211 ;
      RECT 8.97 3.975 8.975 4.212 ;
      RECT 8.955 3.955 8.97 4.214 ;
      RECT 8.88 3.937 8.955 4.226 ;
      RECT 8.87 3.93 8.88 4.237 ;
      RECT 8.865 3.93 8.87 4.239 ;
      RECT 8.835 3.936 8.865 4.243 ;
      RECT 8.795 3.949 8.835 4.243 ;
      RECT 8.77 3.96 8.795 4.229 ;
      RECT 8.755 3.966 8.77 4.212 ;
      RECT 8.745 3.968 8.755 4.203 ;
      RECT 8.74 3.969 8.745 4.198 ;
      RECT 8.735 3.97 8.74 4.193 ;
      RECT 8.73 3.971 8.735 4.19 ;
      RECT 8.705 3.976 8.73 4.18 ;
      RECT 8.695 3.992 8.705 4.167 ;
      RECT 8.69 4.012 8.695 4.162 ;
      RECT 8.7 3.405 8.705 3.601 ;
      RECT 8.685 3.369 8.7 3.603 ;
      RECT 8.675 3.351 8.685 3.608 ;
      RECT 8.665 3.337 8.675 3.612 ;
      RECT 8.62 3.321 8.665 3.622 ;
      RECT 8.615 3.311 8.62 3.631 ;
      RECT 8.57 3.3 8.615 3.637 ;
      RECT 8.565 3.288 8.57 3.644 ;
      RECT 8.55 3.283 8.565 3.648 ;
      RECT 8.535 3.275 8.55 3.653 ;
      RECT 8.525 3.268 8.535 3.658 ;
      RECT 8.515 3.265 8.525 3.663 ;
      RECT 8.505 3.265 8.515 3.664 ;
      RECT 8.5 3.262 8.505 3.663 ;
      RECT 8.465 3.257 8.49 3.662 ;
      RECT 8.441 3.253 8.465 3.661 ;
      RECT 8.355 3.244 8.441 3.658 ;
      RECT 8.34 3.236 8.355 3.655 ;
      RECT 8.318 3.235 8.34 3.654 ;
      RECT 8.232 3.235 8.318 3.652 ;
      RECT 8.146 3.235 8.232 3.65 ;
      RECT 8.06 3.235 8.146 3.647 ;
      RECT 8.05 3.235 8.06 3.638 ;
      RECT 8.02 3.235 8.05 3.598 ;
      RECT 8.01 3.245 8.02 3.553 ;
      RECT 8.005 3.285 8.01 3.538 ;
      RECT 8 3.3 8.005 3.525 ;
      RECT 7.97 3.38 8 3.487 ;
      RECT 8.49 3.26 8.5 3.663 ;
      RECT 8.315 4.025 8.33 4.63 ;
      RECT 8.32 4.02 8.33 4.63 ;
      RECT 8.485 4.02 8.49 4.203 ;
      RECT 8.475 4.02 8.485 4.233 ;
      RECT 8.46 4.02 8.475 4.293 ;
      RECT 8.455 4.02 8.46 4.338 ;
      RECT 8.45 4.02 8.455 4.368 ;
      RECT 8.445 4.02 8.45 4.388 ;
      RECT 8.435 4.02 8.445 4.423 ;
      RECT 8.42 4.02 8.435 4.455 ;
      RECT 8.375 4.02 8.42 4.483 ;
      RECT 8.37 4.02 8.375 4.513 ;
      RECT 8.365 4.02 8.37 4.525 ;
      RECT 8.36 4.02 8.365 4.533 ;
      RECT 8.35 4.02 8.36 4.548 ;
      RECT 8.345 4.02 8.35 4.57 ;
      RECT 8.335 4.02 8.345 4.593 ;
      RECT 8.33 4.02 8.335 4.613 ;
      RECT 8.295 4.035 8.315 4.63 ;
      RECT 8.27 4.052 8.295 4.63 ;
      RECT 8.265 4.062 8.27 4.63 ;
      RECT 8.235 4.077 8.265 4.63 ;
      RECT 8.16 4.119 8.235 4.63 ;
      RECT 8.155 4.15 8.16 4.613 ;
      RECT 8.15 4.154 8.155 4.595 ;
      RECT 8.145 4.158 8.15 4.558 ;
      RECT 8.14 4.342 8.145 4.525 ;
      RECT 7.625 4.531 7.711 5.096 ;
      RECT 7.58 4.533 7.745 5.09 ;
      RECT 7.711 4.53 7.745 5.09 ;
      RECT 7.625 4.532 7.83 5.084 ;
      RECT 7.58 4.542 7.84 5.08 ;
      RECT 7.555 4.534 7.83 5.076 ;
      RECT 7.55 4.537 7.83 5.071 ;
      RECT 7.525 4.552 7.84 5.065 ;
      RECT 7.525 4.577 7.88 5.06 ;
      RECT 7.485 4.585 7.88 5.035 ;
      RECT 7.485 4.612 7.895 5.033 ;
      RECT 7.485 4.642 7.905 5.02 ;
      RECT 7.48 4.787 7.905 5.008 ;
      RECT 7.485 4.716 7.925 5.005 ;
      RECT 7.485 4.773 7.93 4.813 ;
      RECT 7.675 4.052 7.845 4.23 ;
      RECT 7.625 3.991 7.675 4.215 ;
      RECT 7.36 3.971 7.625 4.2 ;
      RECT 7.32 4.035 7.795 4.2 ;
      RECT 7.32 4.025 7.75 4.2 ;
      RECT 7.32 4.022 7.74 4.2 ;
      RECT 7.32 4.01 7.73 4.2 ;
      RECT 7.32 3.995 7.675 4.2 ;
      RECT 7.36 3.967 7.561 4.2 ;
      RECT 7.37 3.945 7.561 4.2 ;
      RECT 7.395 3.93 7.475 4.2 ;
      RECT 7.15 4.46 7.27 4.905 ;
      RECT 7.135 4.46 7.27 4.904 ;
      RECT 7.09 4.482 7.27 4.899 ;
      RECT 7.05 4.531 7.27 4.893 ;
      RECT 7.05 4.531 7.275 4.868 ;
      RECT 7.05 4.531 7.295 4.758 ;
      RECT 7.045 4.561 7.295 4.755 ;
      RECT 7.135 4.46 7.305 4.65 ;
      RECT 6.795 3.245 6.8 3.69 ;
      RECT 6.605 3.245 6.625 3.655 ;
      RECT 6.575 3.245 6.58 3.63 ;
      RECT 7.255 3.552 7.27 3.74 ;
      RECT 7.25 3.537 7.255 3.746 ;
      RECT 7.23 3.51 7.25 3.749 ;
      RECT 7.18 3.477 7.23 3.758 ;
      RECT 7.15 3.457 7.18 3.762 ;
      RECT 7.131 3.445 7.15 3.758 ;
      RECT 7.045 3.417 7.131 3.748 ;
      RECT 7.035 3.392 7.045 3.738 ;
      RECT 6.965 3.36 7.035 3.73 ;
      RECT 6.94 3.32 6.965 3.722 ;
      RECT 6.92 3.302 6.94 3.716 ;
      RECT 6.91 3.292 6.92 3.713 ;
      RECT 6.9 3.285 6.91 3.711 ;
      RECT 6.88 3.272 6.9 3.708 ;
      RECT 6.87 3.262 6.88 3.705 ;
      RECT 6.86 3.255 6.87 3.703 ;
      RECT 6.81 3.247 6.86 3.697 ;
      RECT 6.8 3.245 6.81 3.691 ;
      RECT 6.77 3.245 6.795 3.688 ;
      RECT 6.741 3.245 6.77 3.683 ;
      RECT 6.655 3.245 6.741 3.673 ;
      RECT 6.625 3.245 6.655 3.66 ;
      RECT 6.58 3.245 6.605 3.643 ;
      RECT 6.565 3.245 6.575 3.625 ;
      RECT 6.545 3.252 6.565 3.61 ;
      RECT 6.54 3.267 6.545 3.598 ;
      RECT 6.535 3.272 6.54 3.538 ;
      RECT 6.53 3.277 6.535 3.38 ;
      RECT 6.525 3.28 6.53 3.298 ;
      RECT 6.79 3.965 6.876 4.286 ;
      RECT 6.79 3.965 6.91 4.279 ;
      RECT 6.74 3.965 6.91 4.275 ;
      RECT 6.74 3.967 6.996 4.273 ;
      RECT 6.74 3.969 7.02 4.267 ;
      RECT 6.74 3.976 7.03 4.266 ;
      RECT 6.74 3.985 7.035 4.263 ;
      RECT 6.74 3.991 7.04 4.258 ;
      RECT 6.74 4.035 7.045 4.255 ;
      RECT 6.74 4.127 7.05 4.252 ;
      RECT 6.265 4.57 6.3 4.89 ;
      RECT 6.85 4.755 6.855 4.937 ;
      RECT 6.805 4.637 6.85 4.956 ;
      RECT 6.79 4.614 6.805 4.979 ;
      RECT 6.78 4.604 6.79 4.989 ;
      RECT 6.76 4.599 6.78 5.002 ;
      RECT 6.735 4.597 6.76 5.023 ;
      RECT 6.716 4.596 6.735 5.035 ;
      RECT 6.63 4.593 6.716 5.035 ;
      RECT 6.56 4.588 6.63 5.023 ;
      RECT 6.485 4.584 6.56 4.998 ;
      RECT 6.42 4.58 6.485 4.965 ;
      RECT 6.35 4.577 6.42 4.925 ;
      RECT 6.32 4.573 6.35 4.9 ;
      RECT 6.3 4.571 6.32 4.893 ;
      RECT 6.216 4.569 6.265 4.891 ;
      RECT 6.13 4.566 6.216 4.892 ;
      RECT 6.055 4.565 6.13 4.894 ;
      RECT 5.97 4.565 6.055 4.92 ;
      RECT 5.893 4.566 5.97 4.945 ;
      RECT 5.807 4.567 5.893 4.945 ;
      RECT 5.721 4.567 5.807 4.945 ;
      RECT 5.635 4.568 5.721 4.945 ;
      RECT 5.615 4.569 5.635 4.937 ;
      RECT 5.6 4.575 5.615 4.922 ;
      RECT 5.565 4.595 5.6 4.902 ;
      RECT 5.555 4.615 5.565 4.884 ;
      RECT 6.525 3.92 6.53 4.19 ;
      RECT 6.52 3.911 6.525 4.195 ;
      RECT 6.51 3.901 6.52 4.207 ;
      RECT 6.505 3.89 6.51 4.218 ;
      RECT 6.485 3.884 6.505 4.236 ;
      RECT 6.44 3.881 6.485 4.285 ;
      RECT 6.425 3.88 6.44 4.33 ;
      RECT 6.42 3.88 6.425 4.343 ;
      RECT 6.41 3.88 6.42 4.355 ;
      RECT 6.405 3.881 6.41 4.37 ;
      RECT 6.385 3.889 6.405 4.375 ;
      RECT 6.355 3.905 6.385 4.375 ;
      RECT 6.345 3.917 6.35 4.375 ;
      RECT 6.31 3.932 6.345 4.375 ;
      RECT 6.28 3.952 6.31 4.375 ;
      RECT 6.27 3.977 6.28 4.375 ;
      RECT 6.265 4.005 6.27 4.375 ;
      RECT 6.26 4.035 6.265 4.375 ;
      RECT 6.255 4.052 6.26 4.375 ;
      RECT 6.245 4.08 6.255 4.375 ;
      RECT 6.235 4.115 6.245 4.375 ;
      RECT 6.23 4.15 6.235 4.375 ;
      RECT 6.35 3.915 6.355 4.375 ;
      RECT 5.865 4.017 6.05 4.19 ;
      RECT 5.825 3.935 6.01 4.188 ;
      RECT 5.786 3.94 6.01 4.184 ;
      RECT 5.7 3.949 6.01 4.179 ;
      RECT 5.616 3.965 6.015 4.174 ;
      RECT 5.53 3.985 6.04 4.168 ;
      RECT 5.53 4.005 6.045 4.168 ;
      RECT 5.616 3.975 6.04 4.174 ;
      RECT 5.7 3.95 6.015 4.179 ;
      RECT 5.865 3.932 6.01 4.19 ;
      RECT 5.865 3.927 5.965 4.19 ;
      RECT 5.951 3.921 5.965 4.19 ;
      RECT 5.34 3.245 5.345 3.644 ;
      RECT 5.085 3.245 5.12 3.642 ;
      RECT 4.68 3.28 4.685 3.636 ;
      RECT 5.425 3.283 5.43 3.538 ;
      RECT 5.42 3.281 5.425 3.544 ;
      RECT 5.415 3.28 5.42 3.551 ;
      RECT 5.39 3.273 5.415 3.575 ;
      RECT 5.385 3.266 5.39 3.599 ;
      RECT 5.38 3.262 5.385 3.608 ;
      RECT 5.37 3.257 5.38 3.621 ;
      RECT 5.365 3.254 5.37 3.63 ;
      RECT 5.36 3.252 5.365 3.635 ;
      RECT 5.345 3.248 5.36 3.645 ;
      RECT 5.33 3.242 5.34 3.644 ;
      RECT 5.292 3.24 5.33 3.644 ;
      RECT 5.206 3.242 5.292 3.644 ;
      RECT 5.12 3.244 5.206 3.643 ;
      RECT 5.049 3.245 5.085 3.642 ;
      RECT 4.963 3.247 5.049 3.642 ;
      RECT 4.877 3.249 4.963 3.641 ;
      RECT 4.791 3.251 4.877 3.641 ;
      RECT 4.705 3.254 4.791 3.64 ;
      RECT 4.695 3.26 4.705 3.639 ;
      RECT 4.685 3.272 4.695 3.637 ;
      RECT 4.625 3.307 4.68 3.633 ;
      RECT 4.62 3.337 4.625 3.395 ;
      RECT 5.365 4.417 5.38 4.61 ;
      RECT 5.36 4.385 5.365 4.61 ;
      RECT 5.35 4.36 5.36 4.61 ;
      RECT 5.345 4.332 5.35 4.61 ;
      RECT 5.315 4.255 5.345 4.61 ;
      RECT 5.29 4.137 5.315 4.61 ;
      RECT 5.285 4.075 5.29 4.61 ;
      RECT 5.275 4.062 5.285 4.61 ;
      RECT 5.255 4.052 5.275 4.61 ;
      RECT 5.24 4.035 5.255 4.61 ;
      RECT 5.21 4.023 5.24 4.61 ;
      RECT 5.205 4.022 5.21 4.555 ;
      RECT 5.2 4.022 5.205 4.513 ;
      RECT 5.185 4.021 5.2 4.465 ;
      RECT 5.17 4.021 5.185 4.403 ;
      RECT 5.15 4.021 5.17 4.363 ;
      RECT 5.145 4.021 5.15 4.348 ;
      RECT 5.12 4.02 5.145 4.343 ;
      RECT 5.05 4.019 5.12 4.33 ;
      RECT 5.035 4.018 5.05 4.315 ;
      RECT 5.005 4.017 5.035 4.298 ;
      RECT 5 4.017 5.005 4.283 ;
      RECT 4.95 4.016 5 4.263 ;
      RECT 4.885 4.015 4.95 4.218 ;
      RECT 4.88 4.015 4.885 4.19 ;
      RECT 4.965 4.552 4.97 4.809 ;
      RECT 4.945 4.471 4.965 4.826 ;
      RECT 4.925 4.465 4.945 4.855 ;
      RECT 4.865 4.452 4.925 4.875 ;
      RECT 4.82 4.436 4.865 4.876 ;
      RECT 4.736 4.424 4.82 4.864 ;
      RECT 4.65 4.411 4.736 4.848 ;
      RECT 4.64 4.404 4.65 4.84 ;
      RECT 4.595 4.401 4.64 4.78 ;
      RECT 4.575 4.397 4.595 4.695 ;
      RECT 4.56 4.395 4.575 4.648 ;
      RECT 4.53 4.392 4.56 4.618 ;
      RECT 4.495 4.388 4.53 4.595 ;
      RECT 4.452 4.383 4.495 4.583 ;
      RECT 4.366 4.374 4.452 4.592 ;
      RECT 4.28 4.363 4.366 4.604 ;
      RECT 4.215 4.354 4.28 4.613 ;
      RECT 4.195 4.345 4.215 4.618 ;
      RECT 4.19 4.338 4.195 4.62 ;
      RECT 4.15 4.323 4.19 4.617 ;
      RECT 4.13 4.302 4.15 4.612 ;
      RECT 4.115 4.29 4.13 4.605 ;
      RECT 4.11 4.282 4.115 4.598 ;
      RECT 4.095 4.262 4.11 4.591 ;
      RECT 4.09 4.125 4.095 4.585 ;
      RECT 4.01 4.014 4.09 4.557 ;
      RECT 4.001 4.007 4.01 4.523 ;
      RECT 3.915 4.001 4.001 4.448 ;
      RECT 3.89 3.992 3.915 4.36 ;
      RECT 3.86 3.987 3.89 4.335 ;
      RECT 3.795 3.996 3.86 4.32 ;
      RECT 3.775 4.012 3.795 4.295 ;
      RECT 3.765 4.018 3.775 4.243 ;
      RECT 3.745 4.04 3.765 4.125 ;
      RECT 4.4 4.005 4.57 4.19 ;
      RECT 4.4 4.005 4.605 4.188 ;
      RECT 4.45 3.915 4.62 4.179 ;
      RECT 4.4 4.072 4.625 4.172 ;
      RECT 4.415 3.95 4.62 4.179 ;
      RECT 3.615 4.683 3.68 5.126 ;
      RECT 3.555 4.708 3.68 5.124 ;
      RECT 3.555 4.708 3.735 5.118 ;
      RECT 3.54 4.733 3.735 5.117 ;
      RECT 3.68 4.67 3.755 5.114 ;
      RECT 3.615 4.695 3.835 5.108 ;
      RECT 3.54 4.734 3.88 5.102 ;
      RECT 3.525 4.761 3.88 5.093 ;
      RECT 3.54 4.754 3.9 5.085 ;
      RECT 3.525 4.763 3.905 5.068 ;
      RECT 3.52 4.78 3.905 4.895 ;
      RECT 3.525 3.502 3.56 3.74 ;
      RECT 3.525 3.502 3.59 3.739 ;
      RECT 3.525 3.502 3.705 3.735 ;
      RECT 3.525 3.502 3.76 3.713 ;
      RECT 3.535 3.445 3.815 3.613 ;
      RECT 3.64 3.285 3.67 3.736 ;
      RECT 3.67 3.28 3.85 3.493 ;
      RECT 3.54 3.421 3.85 3.493 ;
      RECT 3.59 3.317 3.64 3.737 ;
      RECT 3.56 3.373 3.85 3.493 ;
      RECT 1.355 10.29 1.525 10.74 ;
      RECT 1.41 8.51 1.58 10.46 ;
      RECT 1.355 7.45 1.525 8.68 ;
      RECT 0.835 7.45 1.005 10.74 ;
      RECT 0.835 9.75 1.24 10.08 ;
      RECT 0.835 8.91 1.24 9.24 ;
      RECT 92.055 7.455 92.225 8.925 ;
      RECT 92.055 10.235 92.225 10.745 ;
      RECT 91.065 1.865 91.235 2.375 ;
      RECT 91.065 3.685 91.235 5.155 ;
      RECT 91.065 7.455 91.235 8.925 ;
      RECT 91.065 10.235 91.235 10.745 ;
      RECT 89.705 1.87 89.875 5.16 ;
      RECT 89.705 7.45 89.875 10.74 ;
      RECT 89.275 1.87 89.445 2.38 ;
      RECT 89.275 2.95 89.445 5.16 ;
      RECT 89.275 7.45 89.445 9.66 ;
      RECT 89.275 10.23 89.445 10.74 ;
      RECT 84.945 7.45 85.115 10.74 ;
      RECT 84.515 7.45 84.685 9.66 ;
      RECT 84.515 10.23 84.685 10.74 ;
      RECT 74.13 7.455 74.3 8.925 ;
      RECT 74.13 10.235 74.3 10.745 ;
      RECT 73.14 1.865 73.31 2.375 ;
      RECT 73.14 3.685 73.31 5.155 ;
      RECT 73.14 7.455 73.31 8.925 ;
      RECT 73.14 10.235 73.31 10.745 ;
      RECT 71.78 1.87 71.95 5.16 ;
      RECT 71.78 7.45 71.95 10.74 ;
      RECT 71.35 1.87 71.52 2.38 ;
      RECT 71.35 2.95 71.52 5.16 ;
      RECT 71.35 7.45 71.52 9.66 ;
      RECT 71.35 10.23 71.52 10.74 ;
      RECT 67.02 7.45 67.19 10.74 ;
      RECT 66.59 7.45 66.76 9.66 ;
      RECT 66.59 10.23 66.76 10.74 ;
      RECT 56.205 7.455 56.375 8.925 ;
      RECT 56.205 10.235 56.375 10.745 ;
      RECT 55.215 1.865 55.385 2.375 ;
      RECT 55.215 3.685 55.385 5.155 ;
      RECT 55.215 7.455 55.385 8.925 ;
      RECT 55.215 10.235 55.385 10.745 ;
      RECT 53.855 1.87 54.025 5.16 ;
      RECT 53.855 7.45 54.025 10.74 ;
      RECT 53.425 1.87 53.595 2.38 ;
      RECT 53.425 2.95 53.595 5.16 ;
      RECT 53.425 7.45 53.595 9.66 ;
      RECT 53.425 10.23 53.595 10.74 ;
      RECT 49.095 7.45 49.265 10.74 ;
      RECT 48.665 7.45 48.835 9.66 ;
      RECT 48.665 10.23 48.835 10.74 ;
      RECT 38.28 7.455 38.45 8.925 ;
      RECT 38.28 10.235 38.45 10.745 ;
      RECT 37.29 1.865 37.46 2.375 ;
      RECT 37.29 3.685 37.46 5.155 ;
      RECT 37.29 7.455 37.46 8.925 ;
      RECT 37.29 10.235 37.46 10.745 ;
      RECT 35.93 1.87 36.1 5.16 ;
      RECT 35.93 7.45 36.1 10.74 ;
      RECT 35.5 1.87 35.67 2.38 ;
      RECT 35.5 2.95 35.67 5.16 ;
      RECT 35.5 7.45 35.67 9.66 ;
      RECT 35.5 10.23 35.67 10.74 ;
      RECT 31.17 7.45 31.34 10.74 ;
      RECT 30.74 7.45 30.91 9.66 ;
      RECT 30.74 10.23 30.91 10.74 ;
      RECT 20.355 7.455 20.525 8.925 ;
      RECT 20.355 10.235 20.525 10.745 ;
      RECT 19.365 1.865 19.535 2.375 ;
      RECT 19.365 3.685 19.535 5.155 ;
      RECT 19.365 7.455 19.535 8.925 ;
      RECT 19.365 10.235 19.535 10.745 ;
      RECT 18.005 1.87 18.175 5.16 ;
      RECT 18.005 7.45 18.175 10.74 ;
      RECT 17.575 1.87 17.745 2.38 ;
      RECT 17.575 2.95 17.745 5.16 ;
      RECT 17.575 7.45 17.745 9.66 ;
      RECT 17.575 10.23 17.745 10.74 ;
      RECT 13.245 7.45 13.415 10.74 ;
      RECT 12.815 7.45 12.985 9.66 ;
      RECT 12.815 10.23 12.985 10.74 ;
      RECT 1.785 7.45 1.955 9.66 ;
      RECT 1.785 10.23 1.955 10.74 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  SIZE 85.77 BY 12.455 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 18.86 1.865 19.03 2.375 ;
        RECT 18.86 3.685 19.03 5.155 ;
      LAYER met1 ;
        RECT 18.8 3.655 19.09 3.885 ;
        RECT 18.8 2.175 19.09 2.405 ;
        RECT 18.86 2.175 19.03 3.885 ;
      LAYER mcon ;
        RECT 18.86 3.685 19.03 3.855 ;
        RECT 18.86 2.205 19.03 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 35.445 1.865 35.615 2.375 ;
        RECT 35.445 3.685 35.615 5.155 ;
      LAYER met1 ;
        RECT 35.385 3.655 35.675 3.885 ;
        RECT 35.385 2.175 35.675 2.405 ;
        RECT 35.445 2.175 35.615 3.885 ;
      LAYER mcon ;
        RECT 35.445 3.685 35.615 3.855 ;
        RECT 35.445 2.205 35.615 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 52.03 1.865 52.2 2.375 ;
        RECT 52.03 3.685 52.2 5.155 ;
      LAYER met1 ;
        RECT 51.97 3.655 52.26 3.885 ;
        RECT 51.97 2.175 52.26 2.405 ;
        RECT 52.03 2.175 52.2 3.885 ;
      LAYER mcon ;
        RECT 52.03 3.685 52.2 3.855 ;
        RECT 52.03 2.205 52.2 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 68.615 1.865 68.785 2.375 ;
        RECT 68.615 3.685 68.785 5.155 ;
      LAYER met1 ;
        RECT 68.555 3.655 68.845 3.885 ;
        RECT 68.555 2.175 68.845 2.405 ;
        RECT 68.615 2.175 68.785 3.885 ;
      LAYER mcon ;
        RECT 68.615 3.685 68.785 3.855 ;
        RECT 68.615 2.205 68.785 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 85.195 1.865 85.365 2.375 ;
        RECT 85.195 3.685 85.365 5.155 ;
      LAYER met1 ;
        RECT 85.135 3.655 85.425 3.885 ;
        RECT 85.135 2.175 85.425 2.405 ;
        RECT 85.195 2.175 85.365 3.885 ;
      LAYER mcon ;
        RECT 85.195 3.685 85.365 3.855 ;
        RECT 85.195 2.205 85.365 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 14.71 2.955 14.88 4.23 ;
        RECT 14.71 8.23 14.88 9.505 ;
        RECT 3.485 8.23 3.655 9.505 ;
      LAYER met2 ;
        RECT 14.635 8.15 14.96 8.475 ;
        RECT 14.63 4.93 14.955 5.255 ;
        RECT 5.79 9.315 14.875 9.485 ;
        RECT 14.7 4.93 14.875 9.485 ;
        RECT 5.735 8.145 6.015 8.485 ;
        RECT 5.79 8.145 5.96 9.485 ;
      LAYER met1 ;
        RECT 14.65 4.06 15.11 4.23 ;
        RECT 14.63 4.93 14.955 5.255 ;
        RECT 14.65 4.03 14.94 4.26 ;
        RECT 14.705 4.03 14.885 5.255 ;
        RECT 14.635 8.23 15.11 8.4 ;
        RECT 14.635 8.15 14.96 8.475 ;
        RECT 5.705 8.175 6.045 8.455 ;
        RECT 3.425 8.23 6.045 8.4 ;
        RECT 3.425 8.2 3.715 8.43 ;
      LAYER via1 ;
        RECT 5.8 8.24 5.95 8.39 ;
        RECT 14.72 5.015 14.87 5.165 ;
        RECT 14.725 8.235 14.875 8.385 ;
      LAYER mcon ;
        RECT 3.485 8.23 3.655 8.4 ;
        RECT 14.71 8.23 14.88 8.4 ;
        RECT 14.71 4.06 14.88 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 31.295 2.955 31.465 4.23 ;
        RECT 31.295 8.23 31.465 9.505 ;
        RECT 20.07 8.23 20.24 9.505 ;
      LAYER met2 ;
        RECT 31.22 8.15 31.545 8.475 ;
        RECT 31.215 4.93 31.54 5.255 ;
        RECT 22.375 9.315 31.46 9.485 ;
        RECT 31.285 4.93 31.46 9.485 ;
        RECT 22.32 8.145 22.6 8.485 ;
        RECT 22.375 8.145 22.545 9.485 ;
      LAYER met1 ;
        RECT 31.235 4.06 31.695 4.23 ;
        RECT 31.215 4.93 31.54 5.255 ;
        RECT 31.235 4.03 31.525 4.26 ;
        RECT 31.29 4.03 31.47 5.255 ;
        RECT 31.22 8.23 31.695 8.4 ;
        RECT 31.22 8.15 31.545 8.475 ;
        RECT 22.29 8.175 22.63 8.455 ;
        RECT 20.01 8.23 22.63 8.4 ;
        RECT 20.01 8.2 20.3 8.43 ;
      LAYER via1 ;
        RECT 22.385 8.24 22.535 8.39 ;
        RECT 31.305 5.015 31.455 5.165 ;
        RECT 31.31 8.235 31.46 8.385 ;
      LAYER mcon ;
        RECT 20.07 8.23 20.24 8.4 ;
        RECT 31.295 8.23 31.465 8.4 ;
        RECT 31.295 4.06 31.465 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 47.88 2.955 48.05 4.23 ;
        RECT 47.88 8.23 48.05 9.505 ;
        RECT 36.655 8.23 36.825 9.505 ;
      LAYER met2 ;
        RECT 47.805 8.15 48.13 8.475 ;
        RECT 47.8 4.93 48.125 5.255 ;
        RECT 38.96 9.315 48.045 9.485 ;
        RECT 47.87 4.93 48.045 9.485 ;
        RECT 38.905 8.145 39.185 8.485 ;
        RECT 38.96 8.145 39.13 9.485 ;
      LAYER met1 ;
        RECT 47.82 4.06 48.28 4.23 ;
        RECT 47.8 4.93 48.125 5.255 ;
        RECT 47.82 4.03 48.11 4.26 ;
        RECT 47.875 4.03 48.055 5.255 ;
        RECT 47.805 8.23 48.28 8.4 ;
        RECT 47.805 8.15 48.13 8.475 ;
        RECT 38.875 8.175 39.215 8.455 ;
        RECT 36.595 8.23 39.215 8.4 ;
        RECT 36.595 8.2 36.885 8.43 ;
      LAYER via1 ;
        RECT 38.97 8.24 39.12 8.39 ;
        RECT 47.89 5.015 48.04 5.165 ;
        RECT 47.895 8.235 48.045 8.385 ;
      LAYER mcon ;
        RECT 36.655 8.23 36.825 8.4 ;
        RECT 47.88 8.23 48.05 8.4 ;
        RECT 47.88 4.06 48.05 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 64.465 2.955 64.635 4.23 ;
        RECT 64.465 8.23 64.635 9.505 ;
        RECT 53.24 8.23 53.41 9.505 ;
      LAYER met2 ;
        RECT 64.39 8.15 64.715 8.475 ;
        RECT 64.385 4.93 64.71 5.255 ;
        RECT 55.545 9.315 64.63 9.485 ;
        RECT 64.455 4.93 64.63 9.485 ;
        RECT 55.49 8.145 55.77 8.485 ;
        RECT 55.545 8.145 55.715 9.485 ;
      LAYER met1 ;
        RECT 64.405 4.06 64.865 4.23 ;
        RECT 64.385 4.93 64.71 5.255 ;
        RECT 64.405 4.03 64.695 4.26 ;
        RECT 64.46 4.03 64.64 5.255 ;
        RECT 64.39 8.23 64.865 8.4 ;
        RECT 64.39 8.15 64.715 8.475 ;
        RECT 55.46 8.175 55.8 8.455 ;
        RECT 53.18 8.23 55.8 8.4 ;
        RECT 53.18 8.2 53.47 8.43 ;
      LAYER via1 ;
        RECT 55.555 8.24 55.705 8.39 ;
        RECT 64.475 5.015 64.625 5.165 ;
        RECT 64.48 8.235 64.63 8.385 ;
      LAYER mcon ;
        RECT 53.24 8.23 53.41 8.4 ;
        RECT 64.465 8.23 64.635 8.4 ;
        RECT 64.465 4.06 64.635 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 81.045 2.955 81.215 4.23 ;
        RECT 81.045 8.23 81.215 9.505 ;
        RECT 69.82 8.23 69.99 9.505 ;
      LAYER met2 ;
        RECT 80.97 8.15 81.295 8.475 ;
        RECT 80.965 4.93 81.29 5.255 ;
        RECT 72.125 9.315 81.21 9.485 ;
        RECT 81.035 4.93 81.21 9.485 ;
        RECT 72.07 8.145 72.35 8.485 ;
        RECT 72.125 8.145 72.295 9.485 ;
      LAYER met1 ;
        RECT 80.985 4.06 81.445 4.23 ;
        RECT 80.965 4.93 81.29 5.255 ;
        RECT 80.985 4.03 81.275 4.26 ;
        RECT 81.04 4.03 81.22 5.255 ;
        RECT 80.97 8.23 81.445 8.4 ;
        RECT 80.97 8.15 81.295 8.475 ;
        RECT 72.04 8.175 72.38 8.455 ;
        RECT 69.76 8.23 72.38 8.4 ;
        RECT 69.76 8.2 70.05 8.43 ;
      LAYER via1 ;
        RECT 72.135 8.24 72.285 8.39 ;
        RECT 81.055 5.015 81.205 5.165 ;
        RECT 81.06 8.235 81.21 8.385 ;
      LAYER mcon ;
        RECT 69.82 8.23 69.99 8.4 ;
        RECT 81.045 8.23 81.215 8.4 ;
        RECT 81.045 4.06 81.215 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.255 8.225 0.425 9.5 ;
      LAYER met1 ;
        RECT 0.195 8.225 0.655 8.395 ;
        RECT 0.195 8.195 0.485 8.425 ;
      LAYER mcon ;
        RECT 0.255 8.225 0.425 8.395 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 79.8 5.43 85.74 7.03 ;
        RECT 83.605 5.425 85.585 7.035 ;
        RECT 84.765 4.695 84.935 7.765 ;
        RECT 83.775 4.695 83.945 7.765 ;
        RECT 81.035 4.7 81.205 7.76 ;
        RECT 79.67 5.43 85.74 5.965 ;
        RECT 79.34 4.495 79.67 5.805 ;
        RECT 0.015 5.635 85.74 5.805 ;
        RECT 77.6 5.095 77.86 5.805 ;
        RECT 77.04 5.635 77.41 6.185 ;
        RECT 76.6 4.715 76.93 4.955 ;
        RECT 76.6 4.715 76.79 5.085 ;
        RECT 76.17 4.985 76.78 5.805 ;
        RECT 76.22 4.985 76.49 6.585 ;
        RECT 75.3 5.095 75.52 5.805 ;
        RECT 75.06 5.635 75.34 6.475 ;
        RECT 74.29 4.765 74.62 4.955 ;
        RECT 73.87 5.135 74.49 5.805 ;
        RECT 74.29 4.765 74.49 5.805 ;
        RECT 74.06 5.135 74.39 6.525 ;
        RECT 72.95 5.125 73.21 5.805 ;
        RECT 63.22 5.43 72.975 7.03 ;
        RECT 69.155 5.425 73.21 5.805 ;
        RECT 69.81 5.425 69.98 7.76 ;
        RECT 67.025 5.425 69.005 7.035 ;
        RECT 68.185 4.695 68.355 7.765 ;
        RECT 67.195 4.695 67.365 7.765 ;
        RECT 64.455 4.7 64.625 7.76 ;
        RECT 63.09 5.43 72.975 5.965 ;
        RECT 62.76 4.495 63.09 5.805 ;
        RECT 61.02 5.095 61.28 5.805 ;
        RECT 60.46 5.635 60.83 6.185 ;
        RECT 60.02 4.715 60.35 4.955 ;
        RECT 60.02 4.715 60.21 5.085 ;
        RECT 59.59 4.985 60.2 5.805 ;
        RECT 59.64 4.985 59.91 6.585 ;
        RECT 58.72 5.095 58.94 5.805 ;
        RECT 58.48 5.635 58.76 6.475 ;
        RECT 57.71 4.765 58.04 4.955 ;
        RECT 57.29 5.135 57.91 5.805 ;
        RECT 57.71 4.765 57.91 5.805 ;
        RECT 57.48 5.135 57.81 6.525 ;
        RECT 56.37 5.125 56.63 5.805 ;
        RECT 46.635 5.43 56.39 7.03 ;
        RECT 52.575 5.425 56.63 5.805 ;
        RECT 53.23 5.425 53.4 7.76 ;
        RECT 50.44 5.425 52.42 7.035 ;
        RECT 51.6 4.695 51.77 7.765 ;
        RECT 50.61 4.695 50.78 7.765 ;
        RECT 47.87 4.7 48.04 7.76 ;
        RECT 46.505 5.43 56.39 5.965 ;
        RECT 46.175 4.495 46.505 5.805 ;
        RECT 44.435 5.095 44.695 5.805 ;
        RECT 43.875 5.635 44.245 6.185 ;
        RECT 43.435 4.715 43.765 4.955 ;
        RECT 43.435 4.715 43.625 5.085 ;
        RECT 43.005 4.985 43.615 5.805 ;
        RECT 43.055 4.985 43.325 6.585 ;
        RECT 42.135 5.095 42.355 5.805 ;
        RECT 41.895 5.635 42.175 6.475 ;
        RECT 41.125 4.765 41.455 4.955 ;
        RECT 40.705 5.135 41.325 5.805 ;
        RECT 41.125 4.765 41.325 5.805 ;
        RECT 40.895 5.135 41.225 6.525 ;
        RECT 39.785 5.125 40.045 5.805 ;
        RECT 30.05 5.43 39.805 7.03 ;
        RECT 35.99 5.425 40.045 5.805 ;
        RECT 36.645 5.425 36.815 7.76 ;
        RECT 33.855 5.425 35.835 7.035 ;
        RECT 35.015 4.695 35.185 7.765 ;
        RECT 34.025 4.695 34.195 7.765 ;
        RECT 31.285 4.7 31.455 7.76 ;
        RECT 29.92 5.43 39.805 5.965 ;
        RECT 29.59 4.495 29.92 5.805 ;
        RECT 27.85 5.095 28.11 5.805 ;
        RECT 27.29 5.635 27.66 6.185 ;
        RECT 26.85 4.715 27.18 4.955 ;
        RECT 26.85 4.715 27.04 5.085 ;
        RECT 26.42 4.985 27.03 5.805 ;
        RECT 26.47 4.985 26.74 6.585 ;
        RECT 25.55 5.095 25.77 5.805 ;
        RECT 25.31 5.635 25.59 6.475 ;
        RECT 24.54 4.765 24.87 4.955 ;
        RECT 24.12 5.135 24.74 5.805 ;
        RECT 24.54 4.765 24.74 5.805 ;
        RECT 24.31 5.135 24.64 6.525 ;
        RECT 23.2 5.125 23.46 5.805 ;
        RECT 13.465 5.43 23.22 7.03 ;
        RECT 19.405 5.425 23.46 5.805 ;
        RECT 20.06 5.425 20.23 7.76 ;
        RECT 17.27 5.425 19.25 7.035 ;
        RECT 18.43 4.695 18.6 7.765 ;
        RECT 17.44 4.695 17.61 7.765 ;
        RECT 14.7 4.7 14.87 7.76 ;
        RECT 13.335 5.43 23.22 5.965 ;
        RECT 13.005 4.495 13.335 5.805 ;
        RECT 11.265 5.095 11.525 5.805 ;
        RECT 10.705 5.635 11.075 6.185 ;
        RECT 10.265 4.715 10.595 4.955 ;
        RECT 10.265 4.715 10.455 5.085 ;
        RECT 9.835 4.985 10.445 5.805 ;
        RECT 9.885 4.985 10.155 6.585 ;
        RECT 8.965 5.095 9.185 5.805 ;
        RECT 8.725 5.635 9.005 6.475 ;
        RECT 7.955 4.765 8.285 4.955 ;
        RECT 7.535 5.135 8.155 5.805 ;
        RECT 7.955 4.765 8.155 5.805 ;
        RECT 7.725 5.135 8.055 6.525 ;
        RECT 6.615 5.125 6.875 5.805 ;
        RECT 0.015 5.425 6.635 7.025 ;
        RECT 3.3 5.425 6.05 7.03 ;
        RECT 3.475 5.425 3.645 7.76 ;
        RECT 2.055 5.425 2.225 10.585 ;
        RECT 0.245 5.425 0.415 7.755 ;
        RECT 0.015 5.415 0.22 7.025 ;
      LAYER met1 ;
        RECT 79.8 5.43 85.74 7.03 ;
        RECT 83.605 5.425 85.585 7.035 ;
        RECT 0.015 5.485 85.74 5.965 ;
        RECT 79.67 5.43 85.74 5.965 ;
        RECT 63.22 5.43 72.975 7.03 ;
        RECT 69.155 5.425 72.97 7.03 ;
        RECT 67.025 5.425 69.005 7.035 ;
        RECT 63.09 5.43 72.975 5.965 ;
        RECT 46.635 5.43 56.39 7.03 ;
        RECT 52.575 5.425 56.39 7.03 ;
        RECT 50.44 5.425 52.42 7.035 ;
        RECT 46.505 5.43 56.39 5.965 ;
        RECT 30.05 5.43 39.805 7.03 ;
        RECT 35.99 5.425 39.805 7.03 ;
        RECT 33.855 5.425 35.835 7.035 ;
        RECT 29.92 5.43 39.805 5.965 ;
        RECT 13.465 5.43 23.22 7.03 ;
        RECT 19.405 5.425 23.22 7.03 ;
        RECT 17.27 5.425 19.25 7.035 ;
        RECT 13.335 5.43 23.22 5.965 ;
        RECT 0.015 5.425 6.635 7.025 ;
        RECT 3.3 5.425 6.05 7.03 ;
        RECT 0.015 5.415 0.22 7.025 ;
        RECT 1.995 8.935 2.285 9.165 ;
        RECT 1.825 8.965 2.285 9.135 ;
      LAYER mcon ;
        RECT 2.055 8.965 2.225 9.135 ;
        RECT 2.365 6.825 2.535 6.995 ;
        RECT 5.595 6.83 5.765 7 ;
        RECT 6.675 5.635 6.845 5.805 ;
        RECT 7.135 5.635 7.305 5.805 ;
        RECT 7.595 5.635 7.765 5.805 ;
        RECT 8.055 5.635 8.225 5.805 ;
        RECT 8.515 5.635 8.685 5.805 ;
        RECT 8.975 5.635 9.145 5.805 ;
        RECT 9.435 5.635 9.605 5.805 ;
        RECT 9.895 5.635 10.065 5.805 ;
        RECT 10.355 5.635 10.525 5.805 ;
        RECT 10.815 5.635 10.985 5.805 ;
        RECT 11.275 5.635 11.445 5.805 ;
        RECT 11.735 5.635 11.905 5.805 ;
        RECT 12.195 5.635 12.365 5.805 ;
        RECT 12.655 5.635 12.825 5.805 ;
        RECT 13.115 5.635 13.285 5.805 ;
        RECT 16.82 6.83 16.99 7 ;
        RECT 16.82 5.46 16.99 5.63 ;
        RECT 17.52 6.835 17.69 7.005 ;
        RECT 17.52 5.455 17.69 5.625 ;
        RECT 18.51 6.835 18.68 7.005 ;
        RECT 18.51 5.455 18.68 5.625 ;
        RECT 22.18 6.83 22.35 7 ;
        RECT 23.26 5.635 23.43 5.805 ;
        RECT 23.72 5.635 23.89 5.805 ;
        RECT 24.18 5.635 24.35 5.805 ;
        RECT 24.64 5.635 24.81 5.805 ;
        RECT 25.1 5.635 25.27 5.805 ;
        RECT 25.56 5.635 25.73 5.805 ;
        RECT 26.02 5.635 26.19 5.805 ;
        RECT 26.48 5.635 26.65 5.805 ;
        RECT 26.94 5.635 27.11 5.805 ;
        RECT 27.4 5.635 27.57 5.805 ;
        RECT 27.86 5.635 28.03 5.805 ;
        RECT 28.32 5.635 28.49 5.805 ;
        RECT 28.78 5.635 28.95 5.805 ;
        RECT 29.24 5.635 29.41 5.805 ;
        RECT 29.7 5.635 29.87 5.805 ;
        RECT 33.405 6.83 33.575 7 ;
        RECT 33.405 5.46 33.575 5.63 ;
        RECT 34.105 6.835 34.275 7.005 ;
        RECT 34.105 5.455 34.275 5.625 ;
        RECT 35.095 6.835 35.265 7.005 ;
        RECT 35.095 5.455 35.265 5.625 ;
        RECT 38.765 6.83 38.935 7 ;
        RECT 39.845 5.635 40.015 5.805 ;
        RECT 40.305 5.635 40.475 5.805 ;
        RECT 40.765 5.635 40.935 5.805 ;
        RECT 41.225 5.635 41.395 5.805 ;
        RECT 41.685 5.635 41.855 5.805 ;
        RECT 42.145 5.635 42.315 5.805 ;
        RECT 42.605 5.635 42.775 5.805 ;
        RECT 43.065 5.635 43.235 5.805 ;
        RECT 43.525 5.635 43.695 5.805 ;
        RECT 43.985 5.635 44.155 5.805 ;
        RECT 44.445 5.635 44.615 5.805 ;
        RECT 44.905 5.635 45.075 5.805 ;
        RECT 45.365 5.635 45.535 5.805 ;
        RECT 45.825 5.635 45.995 5.805 ;
        RECT 46.285 5.635 46.455 5.805 ;
        RECT 49.99 6.83 50.16 7 ;
        RECT 49.99 5.46 50.16 5.63 ;
        RECT 50.69 6.835 50.86 7.005 ;
        RECT 50.69 5.455 50.86 5.625 ;
        RECT 51.68 6.835 51.85 7.005 ;
        RECT 51.68 5.455 51.85 5.625 ;
        RECT 55.35 6.83 55.52 7 ;
        RECT 56.43 5.635 56.6 5.805 ;
        RECT 56.89 5.635 57.06 5.805 ;
        RECT 57.35 5.635 57.52 5.805 ;
        RECT 57.81 5.635 57.98 5.805 ;
        RECT 58.27 5.635 58.44 5.805 ;
        RECT 58.73 5.635 58.9 5.805 ;
        RECT 59.19 5.635 59.36 5.805 ;
        RECT 59.65 5.635 59.82 5.805 ;
        RECT 60.11 5.635 60.28 5.805 ;
        RECT 60.57 5.635 60.74 5.805 ;
        RECT 61.03 5.635 61.2 5.805 ;
        RECT 61.49 5.635 61.66 5.805 ;
        RECT 61.95 5.635 62.12 5.805 ;
        RECT 62.41 5.635 62.58 5.805 ;
        RECT 62.87 5.635 63.04 5.805 ;
        RECT 66.575 6.83 66.745 7 ;
        RECT 66.575 5.46 66.745 5.63 ;
        RECT 67.275 6.835 67.445 7.005 ;
        RECT 67.275 5.455 67.445 5.625 ;
        RECT 68.265 6.835 68.435 7.005 ;
        RECT 68.265 5.455 68.435 5.625 ;
        RECT 71.93 6.83 72.1 7 ;
        RECT 73.01 5.635 73.18 5.805 ;
        RECT 73.47 5.635 73.64 5.805 ;
        RECT 73.93 5.635 74.1 5.805 ;
        RECT 74.39 5.635 74.56 5.805 ;
        RECT 74.85 5.635 75.02 5.805 ;
        RECT 75.31 5.635 75.48 5.805 ;
        RECT 75.77 5.635 75.94 5.805 ;
        RECT 76.23 5.635 76.4 5.805 ;
        RECT 76.69 5.635 76.86 5.805 ;
        RECT 77.15 5.635 77.32 5.805 ;
        RECT 77.61 5.635 77.78 5.805 ;
        RECT 78.07 5.635 78.24 5.805 ;
        RECT 78.53 5.635 78.7 5.805 ;
        RECT 78.99 5.635 79.16 5.805 ;
        RECT 79.45 5.635 79.62 5.805 ;
        RECT 83.155 6.83 83.325 7 ;
        RECT 83.155 5.46 83.325 5.63 ;
        RECT 83.855 6.835 84.025 7.005 ;
        RECT 83.855 5.455 84.025 5.625 ;
        RECT 84.845 6.835 85.015 7.005 ;
        RECT 84.845 5.455 85.015 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.07 10.855 85.77 11.165 ;
        RECT 0.07 10.855 85.74 12.455 ;
        RECT 84.765 10.235 84.935 12.455 ;
        RECT 83.775 10.235 83.945 12.455 ;
        RECT 81.035 10.23 81.205 12.455 ;
        RECT 72.87 8.36 79.785 9.605 ;
        RECT 72.865 9.465 79.775 12.455 ;
        RECT 72.87 8.355 79.77 12.455 ;
        RECT 78.3 7.845 78.75 12.455 ;
        RECT 76.21 7.955 76.54 12.455 ;
        RECT 74.14 7.895 74.39 12.455 ;
        RECT 69.81 10.23 69.98 12.455 ;
        RECT 68.185 10.235 68.355 12.455 ;
        RECT 67.195 10.235 67.365 12.455 ;
        RECT 64.455 10.23 64.625 12.455 ;
        RECT 56.29 8.36 63.205 9.605 ;
        RECT 56.285 9.465 63.195 12.455 ;
        RECT 56.29 8.355 63.19 12.455 ;
        RECT 61.72 7.845 62.17 12.455 ;
        RECT 59.63 7.955 59.96 12.455 ;
        RECT 57.56 7.895 57.81 12.455 ;
        RECT 53.23 10.23 53.4 12.455 ;
        RECT 51.6 10.235 51.77 12.455 ;
        RECT 50.61 10.235 50.78 12.455 ;
        RECT 47.87 10.23 48.04 12.455 ;
        RECT 39.705 8.36 46.62 9.605 ;
        RECT 39.7 9.465 46.61 12.455 ;
        RECT 39.705 8.355 46.605 12.455 ;
        RECT 45.135 7.845 45.585 12.455 ;
        RECT 43.045 7.955 43.375 12.455 ;
        RECT 40.975 7.895 41.225 12.455 ;
        RECT 36.645 10.23 36.815 12.455 ;
        RECT 35.015 10.235 35.185 12.455 ;
        RECT 34.025 10.235 34.195 12.455 ;
        RECT 31.285 10.23 31.455 12.455 ;
        RECT 23.12 8.36 30.035 9.605 ;
        RECT 23.115 9.465 30.025 12.455 ;
        RECT 23.12 8.355 30.02 12.455 ;
        RECT 28.55 7.845 29 12.455 ;
        RECT 26.46 7.955 26.79 12.455 ;
        RECT 24.39 7.895 24.64 12.455 ;
        RECT 20.06 10.23 20.23 12.455 ;
        RECT 18.43 10.235 18.6 12.455 ;
        RECT 17.44 10.235 17.61 12.455 ;
        RECT 14.7 10.23 14.87 12.455 ;
        RECT 6.535 8.36 13.45 9.605 ;
        RECT 6.53 9.465 13.44 12.455 ;
        RECT 6.535 8.355 13.435 12.455 ;
        RECT 11.965 7.845 12.415 12.455 ;
        RECT 9.875 7.955 10.205 12.455 ;
        RECT 7.805 7.895 8.055 12.455 ;
        RECT 3.475 10.23 3.645 12.455 ;
        RECT 0.245 10.225 0.415 12.455 ;
        RECT 0.015 0 85.74 1.6 ;
        RECT 84.765 0 84.935 2.225 ;
        RECT 83.775 0 83.945 2.225 ;
        RECT 81.035 0 81.205 2.23 ;
        RECT 79.765 0 79.96 3.09 ;
        RECT 72.87 0 79.96 3.085 ;
        RECT 79.4 0 79.67 3.895 ;
        RECT 78.49 0 78.73 3.895 ;
        RECT 77.62 0 77.87 3.625 ;
        RECT 75.24 0 75.57 3.545 ;
        RECT 72.95 0 73.21 3.905 ;
        RECT 72.615 0 79.96 2.95 ;
        RECT 68.185 0 68.355 2.225 ;
        RECT 67.195 0 67.365 2.225 ;
        RECT 64.455 0 64.625 2.23 ;
        RECT 63.185 0 63.38 3.09 ;
        RECT 56.29 0 63.38 3.085 ;
        RECT 62.82 0 63.09 3.895 ;
        RECT 61.91 0 62.15 3.895 ;
        RECT 61.04 0 61.29 3.625 ;
        RECT 58.66 0 58.99 3.545 ;
        RECT 56.37 0 56.63 3.905 ;
        RECT 56.035 0 63.38 2.95 ;
        RECT 51.6 0 51.77 2.225 ;
        RECT 50.61 0 50.78 2.225 ;
        RECT 47.87 0 48.04 2.23 ;
        RECT 46.6 0 46.795 3.09 ;
        RECT 39.705 0 46.795 3.085 ;
        RECT 46.235 0 46.505 3.895 ;
        RECT 45.325 0 45.565 3.895 ;
        RECT 44.455 0 44.705 3.625 ;
        RECT 42.075 0 42.405 3.545 ;
        RECT 39.785 0 40.045 3.905 ;
        RECT 39.45 0 46.795 2.95 ;
        RECT 35.015 0 35.185 2.225 ;
        RECT 34.025 0 34.195 2.225 ;
        RECT 31.285 0 31.455 2.23 ;
        RECT 30.015 0 30.21 3.09 ;
        RECT 23.12 0 30.21 3.085 ;
        RECT 29.65 0 29.92 3.895 ;
        RECT 28.74 0 28.98 3.895 ;
        RECT 27.87 0 28.12 3.625 ;
        RECT 25.49 0 25.82 3.545 ;
        RECT 23.2 0 23.46 3.905 ;
        RECT 22.865 0 30.21 2.95 ;
        RECT 18.43 0 18.6 2.225 ;
        RECT 17.44 0 17.61 2.225 ;
        RECT 14.7 0 14.87 2.23 ;
        RECT 13.43 0 13.625 3.09 ;
        RECT 6.535 0 13.625 3.085 ;
        RECT 13.065 0 13.335 3.895 ;
        RECT 12.155 0 12.395 3.895 ;
        RECT 11.285 0 11.535 3.625 ;
        RECT 8.905 0 9.235 3.545 ;
        RECT 6.615 0 6.875 3.905 ;
        RECT 6.28 0 13.625 2.95 ;
        RECT 70.815 8.36 70.985 10.31 ;
        RECT 70.76 10.14 70.93 10.59 ;
        RECT 70.76 7.3 70.93 8.53 ;
        RECT 54.235 8.36 54.405 10.31 ;
        RECT 54.18 10.14 54.35 10.59 ;
        RECT 54.18 7.3 54.35 8.53 ;
        RECT 37.65 8.36 37.82 10.31 ;
        RECT 37.595 10.14 37.765 10.59 ;
        RECT 37.595 7.3 37.765 8.53 ;
        RECT 21.065 8.36 21.235 10.31 ;
        RECT 21.01 10.14 21.18 10.59 ;
        RECT 21.01 7.3 21.18 8.53 ;
        RECT 4.48 8.36 4.65 10.31 ;
        RECT 4.425 10.14 4.595 10.59 ;
        RECT 4.425 7.3 4.595 8.53 ;
      LAYER met1 ;
        RECT 0.07 10.855 85.77 11.165 ;
        RECT 0.07 10.855 85.74 12.455 ;
        RECT 72.87 8.36 79.785 9.605 ;
        RECT 72.865 9.465 79.775 12.455 ;
        RECT 72.87 8.205 79.77 12.455 ;
        RECT 70.755 8.57 71.045 8.8 ;
        RECT 70.595 8.6 70.765 12.455 ;
        RECT 70.585 8.6 71.045 8.77 ;
        RECT 56.29 8.36 63.205 9.605 ;
        RECT 56.285 9.465 63.195 12.455 ;
        RECT 56.29 8.205 63.19 12.455 ;
        RECT 54.175 8.57 54.465 8.8 ;
        RECT 54.015 8.6 54.185 12.455 ;
        RECT 54.005 8.6 54.465 8.77 ;
        RECT 39.705 8.36 46.62 9.605 ;
        RECT 39.7 9.465 46.61 12.455 ;
        RECT 39.705 8.205 46.605 12.455 ;
        RECT 37.59 8.57 37.88 8.8 ;
        RECT 37.43 8.6 37.6 12.455 ;
        RECT 37.42 8.6 37.88 8.77 ;
        RECT 23.12 8.36 30.035 9.605 ;
        RECT 23.115 9.465 30.025 12.455 ;
        RECT 23.12 8.205 30.02 12.455 ;
        RECT 21.005 8.57 21.295 8.8 ;
        RECT 20.845 8.6 21.015 12.455 ;
        RECT 20.835 8.6 21.295 8.77 ;
        RECT 6.535 8.36 13.45 9.605 ;
        RECT 6.53 9.465 13.44 12.455 ;
        RECT 6.535 8.205 13.435 12.455 ;
        RECT 4.42 8.57 4.71 8.8 ;
        RECT 4.26 8.6 4.43 12.455 ;
        RECT 4.25 8.6 4.71 8.77 ;
        RECT 0.015 0 85.74 1.6 ;
        RECT 72.87 0 79.96 3.09 ;
        RECT 72.87 0 79.77 3.245 ;
        RECT 72.615 0 79.96 2.95 ;
        RECT 56.29 0 63.38 3.09 ;
        RECT 56.29 0 63.19 3.245 ;
        RECT 56.035 0 63.38 2.95 ;
        RECT 39.705 0 46.795 3.09 ;
        RECT 39.705 0 46.605 3.245 ;
        RECT 39.45 0 46.795 2.95 ;
        RECT 23.12 0 30.21 3.09 ;
        RECT 23.12 0 30.02 3.245 ;
        RECT 22.865 0 30.21 2.95 ;
        RECT 6.535 0 13.625 3.09 ;
        RECT 6.535 0 13.435 3.245 ;
        RECT 6.28 0 13.625 2.95 ;
      LAYER mcon ;
        RECT 0.325 10.885 0.495 11.055 ;
        RECT 1.005 10.885 1.175 11.055 ;
        RECT 1.685 10.885 1.855 11.055 ;
        RECT 2.365 10.885 2.535 11.055 ;
        RECT 3.555 10.89 3.725 11.06 ;
        RECT 4.235 10.89 4.405 11.06 ;
        RECT 4.48 8.6 4.65 8.77 ;
        RECT 4.915 10.89 5.085 11.06 ;
        RECT 5.595 10.89 5.765 11.06 ;
        RECT 6.675 8.355 6.845 8.525 ;
        RECT 7.135 8.355 7.305 8.525 ;
        RECT 7.595 8.355 7.765 8.525 ;
        RECT 8.055 8.355 8.225 8.525 ;
        RECT 8.515 8.355 8.685 8.525 ;
        RECT 8.975 8.355 9.145 8.525 ;
        RECT 9.435 8.355 9.605 8.525 ;
        RECT 9.895 8.355 10.065 8.525 ;
        RECT 10.355 8.355 10.525 8.525 ;
        RECT 10.815 8.355 10.985 8.525 ;
        RECT 11.275 8.355 11.445 8.525 ;
        RECT 11.735 8.355 11.905 8.525 ;
        RECT 12.195 8.355 12.365 8.525 ;
        RECT 12.655 8.355 12.825 8.525 ;
        RECT 13.115 8.355 13.285 8.525 ;
        RECT 14.78 10.89 14.95 11.06 ;
        RECT 14.78 1.4 14.95 1.57 ;
        RECT 15.46 10.89 15.63 11.06 ;
        RECT 15.46 1.4 15.63 1.57 ;
        RECT 16.14 10.89 16.31 11.06 ;
        RECT 16.14 1.4 16.31 1.57 ;
        RECT 16.82 10.89 16.99 11.06 ;
        RECT 16.82 1.4 16.99 1.57 ;
        RECT 17.52 10.895 17.69 11.065 ;
        RECT 17.52 1.395 17.69 1.565 ;
        RECT 18.51 10.895 18.68 11.065 ;
        RECT 18.51 1.395 18.68 1.565 ;
        RECT 20.14 10.89 20.31 11.06 ;
        RECT 20.82 10.89 20.99 11.06 ;
        RECT 21.065 8.6 21.235 8.77 ;
        RECT 21.5 10.89 21.67 11.06 ;
        RECT 22.18 10.89 22.35 11.06 ;
        RECT 23.26 8.355 23.43 8.525 ;
        RECT 23.72 8.355 23.89 8.525 ;
        RECT 24.18 8.355 24.35 8.525 ;
        RECT 24.64 8.355 24.81 8.525 ;
        RECT 25.1 8.355 25.27 8.525 ;
        RECT 25.56 8.355 25.73 8.525 ;
        RECT 26.02 8.355 26.19 8.525 ;
        RECT 26.48 8.355 26.65 8.525 ;
        RECT 26.94 8.355 27.11 8.525 ;
        RECT 27.4 8.355 27.57 8.525 ;
        RECT 27.86 8.355 28.03 8.525 ;
        RECT 28.32 8.355 28.49 8.525 ;
        RECT 28.78 8.355 28.95 8.525 ;
        RECT 29.24 8.355 29.41 8.525 ;
        RECT 29.7 8.355 29.87 8.525 ;
        RECT 31.365 10.89 31.535 11.06 ;
        RECT 31.365 1.4 31.535 1.57 ;
        RECT 32.045 10.89 32.215 11.06 ;
        RECT 32.045 1.4 32.215 1.57 ;
        RECT 32.725 10.89 32.895 11.06 ;
        RECT 32.725 1.4 32.895 1.57 ;
        RECT 33.405 10.89 33.575 11.06 ;
        RECT 33.405 1.4 33.575 1.57 ;
        RECT 34.105 10.895 34.275 11.065 ;
        RECT 34.105 1.395 34.275 1.565 ;
        RECT 35.095 10.895 35.265 11.065 ;
        RECT 35.095 1.395 35.265 1.565 ;
        RECT 36.725 10.89 36.895 11.06 ;
        RECT 37.405 10.89 37.575 11.06 ;
        RECT 37.65 8.6 37.82 8.77 ;
        RECT 38.085 10.89 38.255 11.06 ;
        RECT 38.765 10.89 38.935 11.06 ;
        RECT 39.845 8.355 40.015 8.525 ;
        RECT 40.305 8.355 40.475 8.525 ;
        RECT 40.765 8.355 40.935 8.525 ;
        RECT 41.225 8.355 41.395 8.525 ;
        RECT 41.685 8.355 41.855 8.525 ;
        RECT 42.145 8.355 42.315 8.525 ;
        RECT 42.605 8.355 42.775 8.525 ;
        RECT 43.065 8.355 43.235 8.525 ;
        RECT 43.525 8.355 43.695 8.525 ;
        RECT 43.985 8.355 44.155 8.525 ;
        RECT 44.445 8.355 44.615 8.525 ;
        RECT 44.905 8.355 45.075 8.525 ;
        RECT 45.365 8.355 45.535 8.525 ;
        RECT 45.825 8.355 45.995 8.525 ;
        RECT 46.285 8.355 46.455 8.525 ;
        RECT 47.95 10.89 48.12 11.06 ;
        RECT 47.95 1.4 48.12 1.57 ;
        RECT 48.63 10.89 48.8 11.06 ;
        RECT 48.63 1.4 48.8 1.57 ;
        RECT 49.31 10.89 49.48 11.06 ;
        RECT 49.31 1.4 49.48 1.57 ;
        RECT 49.99 10.89 50.16 11.06 ;
        RECT 49.99 1.4 50.16 1.57 ;
        RECT 50.69 10.895 50.86 11.065 ;
        RECT 50.69 1.395 50.86 1.565 ;
        RECT 51.68 10.895 51.85 11.065 ;
        RECT 51.68 1.395 51.85 1.565 ;
        RECT 53.31 10.89 53.48 11.06 ;
        RECT 53.99 10.89 54.16 11.06 ;
        RECT 54.235 8.6 54.405 8.77 ;
        RECT 54.67 10.89 54.84 11.06 ;
        RECT 55.35 10.89 55.52 11.06 ;
        RECT 56.43 8.355 56.6 8.525 ;
        RECT 56.89 8.355 57.06 8.525 ;
        RECT 57.35 8.355 57.52 8.525 ;
        RECT 57.81 8.355 57.98 8.525 ;
        RECT 58.27 8.355 58.44 8.525 ;
        RECT 58.73 8.355 58.9 8.525 ;
        RECT 59.19 8.355 59.36 8.525 ;
        RECT 59.65 8.355 59.82 8.525 ;
        RECT 60.11 8.355 60.28 8.525 ;
        RECT 60.57 8.355 60.74 8.525 ;
        RECT 61.03 8.355 61.2 8.525 ;
        RECT 61.49 8.355 61.66 8.525 ;
        RECT 61.95 8.355 62.12 8.525 ;
        RECT 62.41 8.355 62.58 8.525 ;
        RECT 62.87 8.355 63.04 8.525 ;
        RECT 64.535 10.89 64.705 11.06 ;
        RECT 64.535 1.4 64.705 1.57 ;
        RECT 65.215 10.89 65.385 11.06 ;
        RECT 65.215 1.4 65.385 1.57 ;
        RECT 65.895 10.89 66.065 11.06 ;
        RECT 65.895 1.4 66.065 1.57 ;
        RECT 66.575 10.89 66.745 11.06 ;
        RECT 66.575 1.4 66.745 1.57 ;
        RECT 67.275 10.895 67.445 11.065 ;
        RECT 67.275 1.395 67.445 1.565 ;
        RECT 68.265 10.895 68.435 11.065 ;
        RECT 68.265 1.395 68.435 1.565 ;
        RECT 69.89 10.89 70.06 11.06 ;
        RECT 70.57 10.89 70.74 11.06 ;
        RECT 70.815 8.6 70.985 8.77 ;
        RECT 71.25 10.89 71.42 11.06 ;
        RECT 71.93 10.89 72.1 11.06 ;
        RECT 73.01 8.355 73.18 8.525 ;
        RECT 73.47 8.355 73.64 8.525 ;
        RECT 73.93 8.355 74.1 8.525 ;
        RECT 74.39 8.355 74.56 8.525 ;
        RECT 74.85 8.355 75.02 8.525 ;
        RECT 75.31 8.355 75.48 8.525 ;
        RECT 75.77 8.355 75.94 8.525 ;
        RECT 76.23 8.355 76.4 8.525 ;
        RECT 76.69 8.355 76.86 8.525 ;
        RECT 77.15 8.355 77.32 8.525 ;
        RECT 77.61 8.355 77.78 8.525 ;
        RECT 78.07 8.355 78.24 8.525 ;
        RECT 78.53 8.355 78.7 8.525 ;
        RECT 78.99 8.355 79.16 8.525 ;
        RECT 79.45 8.355 79.62 8.525 ;
        RECT 81.115 10.89 81.285 11.06 ;
        RECT 81.115 1.4 81.285 1.57 ;
        RECT 81.795 10.89 81.965 11.06 ;
        RECT 81.795 1.4 81.965 1.57 ;
        RECT 82.475 10.89 82.645 11.06 ;
        RECT 82.475 1.4 82.645 1.57 ;
        RECT 83.155 10.89 83.325 11.06 ;
        RECT 83.155 1.4 83.325 1.57 ;
        RECT 83.855 10.895 84.025 11.065 ;
        RECT 83.855 1.395 84.025 1.565 ;
        RECT 84.845 10.895 85.015 11.065 ;
        RECT 84.845 1.395 85.015 1.565 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 77.665 4.025 77.965 4.36 ;
      RECT 77.64 4.025 77.97 4.355 ;
      RECT 77.64 4.045 78.44 4.345 ;
      RECT 71.09 9.28 71.46 9.65 ;
      RECT 71.09 9.315 76.245 9.615 ;
      RECT 75.94 7.085 76.24 9.615 ;
      RECT 75.315 7.105 76.25 7.425 ;
      RECT 75.92 7.085 76.25 7.425 ;
      RECT 76.96 7.085 77.29 7.415 ;
      RECT 75.315 7.11 77.29 7.41 ;
      RECT 76.745 7.095 77.29 7.41 ;
      RECT 76.745 7.105 77.76 7.405 ;
      RECT 75.315 5.06 75.62 7.425 ;
      RECT 75.315 6.12 75.645 6.42 ;
      RECT 75.315 5.06 75.645 5.805 ;
      RECT 75.315 5.06 77.61 5.39 ;
      RECT 75.315 5.06 77.965 5.38 ;
      RECT 77.64 5.045 77.97 5.375 ;
      RECT 75.315 5.065 78.44 5.365 ;
      RECT 77.65 4.995 77.95 5.38 ;
      RECT 76.94 4.365 77.27 4.695 ;
      RECT 76.97 4.355 77.27 4.695 ;
      RECT 76.47 4.385 77.27 4.685 ;
      RECT 76.275 6.08 76.31 6.4 ;
      RECT 76.28 6.065 76.61 6.395 ;
      RECT 76.275 6.085 77.08 6.385 ;
      RECT 75.6 3.685 75.93 4.015 ;
      RECT 75.13 3.705 75.49 4.005 ;
      RECT 75.49 3.695 75.93 3.995 ;
      RECT 75.21 7.785 75.51 8.195 ;
      RECT 75.24 7.765 75.57 8.095 ;
      RECT 74.77 7.785 75.57 8.085 ;
      RECT 61.085 4.025 61.385 4.36 ;
      RECT 61.06 4.025 61.39 4.355 ;
      RECT 61.06 4.045 61.86 4.345 ;
      RECT 54.51 9.28 54.88 9.65 ;
      RECT 54.51 9.315 59.665 9.615 ;
      RECT 59.36 7.085 59.66 9.615 ;
      RECT 58.735 7.105 59.67 7.425 ;
      RECT 59.34 7.085 59.67 7.425 ;
      RECT 60.38 7.085 60.71 7.415 ;
      RECT 58.735 7.11 60.71 7.41 ;
      RECT 60.165 7.095 60.71 7.41 ;
      RECT 60.165 7.105 61.18 7.405 ;
      RECT 58.735 5.06 59.04 7.425 ;
      RECT 58.735 6.12 59.065 6.42 ;
      RECT 58.735 5.06 59.065 5.805 ;
      RECT 58.735 5.06 61.03 5.39 ;
      RECT 58.735 5.06 61.385 5.38 ;
      RECT 61.06 5.045 61.39 5.375 ;
      RECT 58.735 5.065 61.86 5.365 ;
      RECT 61.07 4.995 61.37 5.38 ;
      RECT 60.36 4.365 60.69 4.695 ;
      RECT 60.39 4.355 60.69 4.695 ;
      RECT 59.89 4.385 60.69 4.685 ;
      RECT 59.695 6.08 59.73 6.4 ;
      RECT 59.7 6.065 60.03 6.395 ;
      RECT 59.695 6.085 60.5 6.385 ;
      RECT 59.02 3.685 59.35 4.015 ;
      RECT 58.55 3.705 58.91 4.005 ;
      RECT 58.91 3.695 59.35 3.995 ;
      RECT 58.63 7.785 58.93 8.195 ;
      RECT 58.66 7.765 58.99 8.095 ;
      RECT 58.19 7.785 58.99 8.085 ;
      RECT 44.5 4.025 44.8 4.36 ;
      RECT 44.475 4.025 44.805 4.355 ;
      RECT 44.475 4.045 45.275 4.345 ;
      RECT 37.925 9.28 38.295 9.65 ;
      RECT 37.925 9.315 43.08 9.615 ;
      RECT 42.775 7.085 43.075 9.615 ;
      RECT 42.15 7.105 43.085 7.425 ;
      RECT 42.755 7.085 43.085 7.425 ;
      RECT 43.795 7.085 44.125 7.415 ;
      RECT 42.15 7.11 44.125 7.41 ;
      RECT 43.58 7.095 44.125 7.41 ;
      RECT 43.58 7.105 44.595 7.405 ;
      RECT 42.15 5.06 42.455 7.425 ;
      RECT 42.15 6.12 42.48 6.42 ;
      RECT 42.15 5.06 42.48 5.805 ;
      RECT 42.15 5.06 44.445 5.39 ;
      RECT 42.15 5.06 44.8 5.38 ;
      RECT 44.475 5.045 44.805 5.375 ;
      RECT 42.15 5.065 45.275 5.365 ;
      RECT 44.485 4.995 44.785 5.38 ;
      RECT 43.775 4.365 44.105 4.695 ;
      RECT 43.805 4.355 44.105 4.695 ;
      RECT 43.305 4.385 44.105 4.685 ;
      RECT 43.11 6.08 43.145 6.4 ;
      RECT 43.115 6.065 43.445 6.395 ;
      RECT 43.11 6.085 43.915 6.385 ;
      RECT 42.435 3.685 42.765 4.015 ;
      RECT 41.965 3.705 42.325 4.005 ;
      RECT 42.325 3.695 42.765 3.995 ;
      RECT 42.045 7.785 42.345 8.195 ;
      RECT 42.075 7.765 42.405 8.095 ;
      RECT 41.605 7.785 42.405 8.085 ;
      RECT 27.915 4.025 28.215 4.36 ;
      RECT 27.89 4.025 28.22 4.355 ;
      RECT 27.89 4.045 28.69 4.345 ;
      RECT 21.34 9.28 21.71 9.65 ;
      RECT 21.34 9.315 26.495 9.615 ;
      RECT 26.19 7.085 26.49 9.615 ;
      RECT 25.565 7.105 26.5 7.425 ;
      RECT 26.17 7.085 26.5 7.425 ;
      RECT 27.21 7.085 27.54 7.415 ;
      RECT 25.565 7.11 27.54 7.41 ;
      RECT 26.995 7.095 27.54 7.41 ;
      RECT 26.995 7.105 28.01 7.405 ;
      RECT 25.565 5.06 25.87 7.425 ;
      RECT 25.565 6.12 25.895 6.42 ;
      RECT 25.565 5.06 25.895 5.805 ;
      RECT 25.565 5.06 27.86 5.39 ;
      RECT 25.565 5.06 28.215 5.38 ;
      RECT 27.89 5.045 28.22 5.375 ;
      RECT 25.565 5.065 28.69 5.365 ;
      RECT 27.9 4.995 28.2 5.38 ;
      RECT 27.19 4.365 27.52 4.695 ;
      RECT 27.22 4.355 27.52 4.695 ;
      RECT 26.72 4.385 27.52 4.685 ;
      RECT 26.525 6.08 26.56 6.4 ;
      RECT 26.53 6.065 26.86 6.395 ;
      RECT 26.525 6.085 27.33 6.385 ;
      RECT 25.85 3.685 26.18 4.015 ;
      RECT 25.38 3.705 25.74 4.005 ;
      RECT 25.74 3.695 26.18 3.995 ;
      RECT 25.46 7.785 25.76 8.195 ;
      RECT 25.49 7.765 25.82 8.095 ;
      RECT 25.02 7.785 25.82 8.085 ;
      RECT 11.33 4.025 11.63 4.36 ;
      RECT 11.305 4.025 11.635 4.355 ;
      RECT 11.305 4.045 12.105 4.345 ;
      RECT 4.755 9.28 5.125 9.65 ;
      RECT 4.755 9.315 9.91 9.615 ;
      RECT 9.605 7.085 9.905 9.615 ;
      RECT 8.98 7.105 9.915 7.425 ;
      RECT 9.585 7.085 9.915 7.425 ;
      RECT 10.625 7.085 10.955 7.415 ;
      RECT 8.98 7.11 10.955 7.41 ;
      RECT 10.41 7.095 10.955 7.41 ;
      RECT 10.41 7.105 11.425 7.405 ;
      RECT 8.98 5.06 9.285 7.425 ;
      RECT 8.98 6.12 9.31 6.42 ;
      RECT 8.98 5.06 9.31 5.805 ;
      RECT 8.98 5.06 11.275 5.39 ;
      RECT 8.98 5.06 11.63 5.38 ;
      RECT 11.305 5.045 11.635 5.375 ;
      RECT 8.98 5.065 12.105 5.365 ;
      RECT 11.315 4.995 11.615 5.38 ;
      RECT 10.605 4.365 10.935 4.695 ;
      RECT 10.635 4.355 10.935 4.695 ;
      RECT 10.135 4.385 10.935 4.685 ;
      RECT 9.94 6.08 9.975 6.4 ;
      RECT 9.945 6.065 10.275 6.395 ;
      RECT 9.94 6.085 10.745 6.385 ;
      RECT 9.265 3.685 9.595 4.015 ;
      RECT 8.795 3.705 9.155 4.005 ;
      RECT 9.155 3.695 9.595 3.995 ;
      RECT 8.875 7.785 9.175 8.195 ;
      RECT 8.905 7.765 9.235 8.095 ;
      RECT 8.435 7.785 9.235 8.085 ;
    LAYER via2 ;
      RECT 77.71 4.095 77.91 4.295 ;
      RECT 77.71 5.115 77.91 5.315 ;
      RECT 77.03 7.155 77.23 7.355 ;
      RECT 77.01 4.435 77.21 4.635 ;
      RECT 76.35 6.135 76.55 6.335 ;
      RECT 75.98 7.155 76.18 7.355 ;
      RECT 75.67 3.745 75.87 3.945 ;
      RECT 75.31 7.835 75.51 8.035 ;
      RECT 71.175 9.365 71.375 9.565 ;
      RECT 61.13 4.095 61.33 4.295 ;
      RECT 61.13 5.115 61.33 5.315 ;
      RECT 60.45 7.155 60.65 7.355 ;
      RECT 60.43 4.435 60.63 4.635 ;
      RECT 59.77 6.135 59.97 6.335 ;
      RECT 59.4 7.155 59.6 7.355 ;
      RECT 59.09 3.745 59.29 3.945 ;
      RECT 58.73 7.835 58.93 8.035 ;
      RECT 54.595 9.365 54.795 9.565 ;
      RECT 44.545 4.095 44.745 4.295 ;
      RECT 44.545 5.115 44.745 5.315 ;
      RECT 43.865 7.155 44.065 7.355 ;
      RECT 43.845 4.435 44.045 4.635 ;
      RECT 43.185 6.135 43.385 6.335 ;
      RECT 42.815 7.155 43.015 7.355 ;
      RECT 42.505 3.745 42.705 3.945 ;
      RECT 42.145 7.835 42.345 8.035 ;
      RECT 38.01 9.365 38.21 9.565 ;
      RECT 27.96 4.095 28.16 4.295 ;
      RECT 27.96 5.115 28.16 5.315 ;
      RECT 27.28 7.155 27.48 7.355 ;
      RECT 27.26 4.435 27.46 4.635 ;
      RECT 26.6 6.135 26.8 6.335 ;
      RECT 26.23 7.155 26.43 7.355 ;
      RECT 25.92 3.745 26.12 3.945 ;
      RECT 25.56 7.835 25.76 8.035 ;
      RECT 21.425 9.365 21.625 9.565 ;
      RECT 11.375 4.095 11.575 4.295 ;
      RECT 11.375 5.115 11.575 5.315 ;
      RECT 10.695 7.155 10.895 7.355 ;
      RECT 10.675 4.435 10.875 4.635 ;
      RECT 10.015 6.135 10.215 6.335 ;
      RECT 9.645 7.155 9.845 7.355 ;
      RECT 9.335 3.745 9.535 3.945 ;
      RECT 8.975 7.835 9.175 8.035 ;
      RECT 4.84 9.365 5.04 9.565 ;
    LAYER met2 ;
      RECT 2.78 10.12 85.37 10.29 ;
      RECT 85.2 9.585 85.37 10.29 ;
      RECT 1.245 10.115 2.78 10.285 ;
      RECT 1.245 8.535 1.415 10.285 ;
      RECT 85.165 9.585 85.49 9.91 ;
      RECT 1.19 8.535 1.47 8.875 ;
      RECT 82.01 8.565 82.33 8.89 ;
      RECT 82.04 7.98 82.21 8.89 ;
      RECT 82.04 7.98 82.215 8.33 ;
      RECT 82.04 7.98 83.015 8.155 ;
      RECT 82.84 3.26 83.015 8.155 ;
      RECT 82.785 3.26 83.135 3.61 ;
      RECT 71.675 9.72 81.855 9.89 ;
      RECT 81.695 3.69 81.855 9.89 ;
      RECT 71.675 8.885 71.845 9.89 ;
      RECT 82.81 8.94 83.135 9.265 ;
      RECT 68.62 8.94 68.945 9.265 ;
      RECT 71.62 8.885 71.9 9.225 ;
      RECT 81.695 9.03 83.135 9.2 ;
      RECT 68.62 8.97 71.9 9.14 ;
      RECT 82.01 3.66 82.33 3.98 ;
      RECT 81.695 3.69 82.33 3.86 ;
      RECT 79.755 4.48 80.08 4.805 ;
      RECT 79.755 4.51 80.585 4.695 ;
      RECT 80.415 3.29 80.585 4.695 ;
      RECT 80.34 3.29 80.665 3.615 ;
      RECT 79.37 6.075 79.63 6.395 ;
      RECT 79.43 4.035 79.57 6.395 ;
      RECT 79.37 4.035 79.63 4.355 ;
      RECT 78.35 7.095 78.61 7.415 ;
      RECT 77.73 7.185 78.61 7.325 ;
      RECT 77.73 5.025 77.87 7.325 ;
      RECT 77.67 5.025 77.95 5.395 ;
      RECT 76.99 7.065 77.27 7.435 ;
      RECT 77.05 5.145 77.19 7.435 ;
      RECT 77.05 5.145 77.53 5.285 ;
      RECT 77.39 3.355 77.53 5.285 ;
      RECT 77.33 3.355 77.59 3.675 ;
      RECT 76.31 6.045 76.59 6.415 ;
      RECT 76.37 3.695 76.51 6.415 ;
      RECT 76.31 3.695 76.57 4.015 ;
      RECT 75.94 7.065 76.22 7.435 ;
      RECT 75.94 7.095 76.23 7.415 ;
      RECT 65.43 8.565 65.75 8.89 ;
      RECT 65.46 7.98 65.63 8.89 ;
      RECT 65.46 7.98 65.635 8.33 ;
      RECT 65.46 7.98 66.435 8.155 ;
      RECT 66.26 3.26 66.435 8.155 ;
      RECT 66.205 3.26 66.555 3.61 ;
      RECT 55.095 9.72 65.275 9.89 ;
      RECT 65.115 3.69 65.275 9.89 ;
      RECT 55.095 8.885 55.265 9.89 ;
      RECT 66.23 8.94 66.555 9.265 ;
      RECT 52.035 8.94 52.36 9.265 ;
      RECT 55.04 8.885 55.32 9.225 ;
      RECT 65.115 9.03 66.555 9.2 ;
      RECT 52.035 8.97 55.32 9.14 ;
      RECT 65.43 3.66 65.75 3.98 ;
      RECT 65.115 3.69 65.75 3.86 ;
      RECT 63.175 4.48 63.5 4.805 ;
      RECT 63.175 4.51 64.005 4.695 ;
      RECT 63.835 3.29 64.005 4.695 ;
      RECT 63.76 3.29 64.085 3.615 ;
      RECT 62.79 6.075 63.05 6.395 ;
      RECT 62.85 4.035 62.99 6.395 ;
      RECT 62.79 4.035 63.05 4.355 ;
      RECT 61.77 7.095 62.03 7.415 ;
      RECT 61.15 7.185 62.03 7.325 ;
      RECT 61.15 5.025 61.29 7.325 ;
      RECT 61.09 5.025 61.37 5.395 ;
      RECT 60.41 7.065 60.69 7.435 ;
      RECT 60.47 5.145 60.61 7.435 ;
      RECT 60.47 5.145 60.95 5.285 ;
      RECT 60.81 3.355 60.95 5.285 ;
      RECT 60.75 3.355 61.01 3.675 ;
      RECT 59.73 6.045 60.01 6.415 ;
      RECT 59.79 3.695 59.93 6.415 ;
      RECT 59.73 3.695 59.99 4.015 ;
      RECT 59.36 7.065 59.64 7.435 ;
      RECT 59.36 7.095 59.65 7.415 ;
      RECT 48.845 8.565 49.165 8.89 ;
      RECT 48.875 7.98 49.045 8.89 ;
      RECT 48.875 7.98 49.05 8.33 ;
      RECT 48.875 7.98 49.85 8.155 ;
      RECT 49.675 3.26 49.85 8.155 ;
      RECT 49.62 3.26 49.97 3.61 ;
      RECT 38.51 9.72 48.69 9.89 ;
      RECT 48.53 3.69 48.69 9.89 ;
      RECT 38.51 8.885 38.68 9.89 ;
      RECT 49.645 8.94 49.97 9.265 ;
      RECT 35.45 8.94 35.775 9.265 ;
      RECT 38.455 8.885 38.735 9.225 ;
      RECT 48.53 9.03 49.97 9.2 ;
      RECT 35.45 8.97 38.735 9.14 ;
      RECT 48.845 3.66 49.165 3.98 ;
      RECT 48.53 3.69 49.165 3.86 ;
      RECT 46.59 4.48 46.915 4.805 ;
      RECT 46.59 4.51 47.42 4.695 ;
      RECT 47.25 3.29 47.42 4.695 ;
      RECT 47.175 3.29 47.5 3.615 ;
      RECT 46.205 6.075 46.465 6.395 ;
      RECT 46.265 4.035 46.405 6.395 ;
      RECT 46.205 4.035 46.465 4.355 ;
      RECT 45.185 7.095 45.445 7.415 ;
      RECT 44.565 7.185 45.445 7.325 ;
      RECT 44.565 5.025 44.705 7.325 ;
      RECT 44.505 5.025 44.785 5.395 ;
      RECT 43.825 7.065 44.105 7.435 ;
      RECT 43.885 5.145 44.025 7.435 ;
      RECT 43.885 5.145 44.365 5.285 ;
      RECT 44.225 3.355 44.365 5.285 ;
      RECT 44.165 3.355 44.425 3.675 ;
      RECT 43.145 6.045 43.425 6.415 ;
      RECT 43.205 3.695 43.345 6.415 ;
      RECT 43.145 3.695 43.405 4.015 ;
      RECT 42.775 7.065 43.055 7.435 ;
      RECT 42.775 7.095 43.065 7.415 ;
      RECT 32.26 8.565 32.58 8.89 ;
      RECT 32.29 7.98 32.46 8.89 ;
      RECT 32.29 7.98 32.465 8.33 ;
      RECT 32.29 7.98 33.265 8.155 ;
      RECT 33.09 3.26 33.265 8.155 ;
      RECT 33.035 3.26 33.385 3.61 ;
      RECT 21.925 9.72 32.105 9.89 ;
      RECT 31.945 3.69 32.105 9.89 ;
      RECT 21.925 8.885 22.095 9.89 ;
      RECT 33.06 8.94 33.385 9.265 ;
      RECT 18.865 8.94 19.19 9.265 ;
      RECT 21.87 8.885 22.15 9.225 ;
      RECT 31.945 9.03 33.385 9.2 ;
      RECT 18.865 8.97 22.15 9.14 ;
      RECT 32.26 3.66 32.58 3.98 ;
      RECT 31.945 3.69 32.58 3.86 ;
      RECT 30.005 4.48 30.33 4.805 ;
      RECT 30.005 4.51 30.835 4.695 ;
      RECT 30.665 3.29 30.835 4.695 ;
      RECT 30.59 3.29 30.915 3.615 ;
      RECT 29.62 6.075 29.88 6.395 ;
      RECT 29.68 4.035 29.82 6.395 ;
      RECT 29.62 4.035 29.88 4.355 ;
      RECT 28.6 7.095 28.86 7.415 ;
      RECT 27.98 7.185 28.86 7.325 ;
      RECT 27.98 5.025 28.12 7.325 ;
      RECT 27.92 5.025 28.2 5.395 ;
      RECT 27.24 7.065 27.52 7.435 ;
      RECT 27.3 5.145 27.44 7.435 ;
      RECT 27.3 5.145 27.78 5.285 ;
      RECT 27.64 3.355 27.78 5.285 ;
      RECT 27.58 3.355 27.84 3.675 ;
      RECT 26.56 6.045 26.84 6.415 ;
      RECT 26.62 3.695 26.76 6.415 ;
      RECT 26.56 3.695 26.82 4.015 ;
      RECT 26.19 7.065 26.47 7.435 ;
      RECT 26.19 7.095 26.48 7.415 ;
      RECT 15.675 8.565 15.995 8.89 ;
      RECT 15.705 7.98 15.875 8.89 ;
      RECT 15.705 7.98 15.88 8.33 ;
      RECT 15.705 7.98 16.68 8.155 ;
      RECT 16.505 3.26 16.68 8.155 ;
      RECT 16.45 3.26 16.8 3.61 ;
      RECT 5.34 9.72 15.52 9.89 ;
      RECT 15.36 3.69 15.52 9.89 ;
      RECT 5.34 8.885 5.51 9.89 ;
      RECT 1.565 9.275 1.845 9.615 ;
      RECT 1.565 9.34 2.73 9.51 ;
      RECT 2.56 8.97 2.73 9.51 ;
      RECT 16.475 8.94 16.8 9.265 ;
      RECT 5.285 8.885 5.565 9.225 ;
      RECT 15.36 9.03 16.8 9.2 ;
      RECT 2.56 8.97 2.88 9.145 ;
      RECT 2.56 8.97 5.565 9.14 ;
      RECT 15.675 3.66 15.995 3.98 ;
      RECT 15.36 3.69 15.995 3.86 ;
      RECT 13.42 4.48 13.745 4.805 ;
      RECT 13.42 4.51 14.25 4.695 ;
      RECT 14.08 3.29 14.25 4.695 ;
      RECT 14.005 3.29 14.33 3.615 ;
      RECT 13.035 6.075 13.295 6.395 ;
      RECT 13.095 4.035 13.235 6.395 ;
      RECT 13.035 4.035 13.295 4.355 ;
      RECT 12.015 7.095 12.275 7.415 ;
      RECT 11.395 7.185 12.275 7.325 ;
      RECT 11.395 5.025 11.535 7.325 ;
      RECT 11.335 5.025 11.615 5.395 ;
      RECT 10.655 7.065 10.935 7.435 ;
      RECT 10.715 5.145 10.855 7.435 ;
      RECT 10.715 5.145 11.195 5.285 ;
      RECT 11.055 3.355 11.195 5.285 ;
      RECT 10.995 3.355 11.255 3.675 ;
      RECT 9.975 6.045 10.255 6.415 ;
      RECT 10.035 3.695 10.175 6.415 ;
      RECT 9.975 3.695 10.235 4.015 ;
      RECT 9.605 7.065 9.885 7.435 ;
      RECT 9.605 7.095 9.895 7.415 ;
      RECT 77.67 4.005 77.95 4.375 ;
      RECT 76.97 4.345 77.25 4.715 ;
      RECT 75.63 3.665 75.91 4.035 ;
      RECT 75.27 7.745 75.55 8.115 ;
      RECT 71.09 9.28 71.465 9.65 ;
      RECT 61.09 4.005 61.37 4.375 ;
      RECT 60.39 4.345 60.67 4.715 ;
      RECT 59.05 3.665 59.33 4.035 ;
      RECT 58.69 7.745 58.97 8.115 ;
      RECT 54.51 9.28 54.88 9.65 ;
      RECT 44.505 4.005 44.785 4.375 ;
      RECT 43.805 4.345 44.085 4.715 ;
      RECT 42.465 3.665 42.745 4.035 ;
      RECT 42.105 7.745 42.385 8.115 ;
      RECT 37.925 9.28 38.295 9.65 ;
      RECT 27.92 4.005 28.2 4.375 ;
      RECT 27.22 4.345 27.5 4.715 ;
      RECT 25.88 3.665 26.16 4.035 ;
      RECT 25.52 7.745 25.8 8.115 ;
      RECT 21.34 9.28 21.71 9.65 ;
      RECT 11.335 4.005 11.615 4.375 ;
      RECT 10.635 4.345 10.915 4.715 ;
      RECT 9.295 3.665 9.575 4.035 ;
      RECT 8.935 7.745 9.215 8.115 ;
      RECT 4.755 9.28 5.125 9.65 ;
    LAYER via1 ;
      RECT 85.255 9.67 85.405 9.82 ;
      RECT 82.9 9.025 83.05 9.175 ;
      RECT 82.885 3.36 83.035 3.51 ;
      RECT 82.095 3.745 82.245 3.895 ;
      RECT 82.095 8.655 82.245 8.805 ;
      RECT 80.43 3.375 80.58 3.525 ;
      RECT 79.845 4.565 79.995 4.715 ;
      RECT 79.425 4.12 79.575 4.27 ;
      RECT 79.425 6.16 79.575 6.31 ;
      RECT 78.405 7.18 78.555 7.33 ;
      RECT 77.725 4.12 77.875 4.27 ;
      RECT 77.725 5.14 77.875 5.29 ;
      RECT 77.385 3.44 77.535 3.59 ;
      RECT 77.045 4.46 77.195 4.61 ;
      RECT 77.045 7.18 77.195 7.33 ;
      RECT 76.365 3.78 76.515 3.93 ;
      RECT 76.365 6.16 76.515 6.31 ;
      RECT 76.025 7.18 76.175 7.33 ;
      RECT 75.685 3.77 75.835 3.92 ;
      RECT 75.345 7.86 75.495 8.01 ;
      RECT 71.685 8.98 71.835 9.13 ;
      RECT 71.2 9.39 71.35 9.54 ;
      RECT 68.71 9.025 68.86 9.175 ;
      RECT 66.32 9.025 66.47 9.175 ;
      RECT 66.305 3.36 66.455 3.51 ;
      RECT 65.515 3.745 65.665 3.895 ;
      RECT 65.515 8.655 65.665 8.805 ;
      RECT 63.85 3.375 64 3.525 ;
      RECT 63.265 4.565 63.415 4.715 ;
      RECT 62.845 4.12 62.995 4.27 ;
      RECT 62.845 6.16 62.995 6.31 ;
      RECT 61.825 7.18 61.975 7.33 ;
      RECT 61.145 4.12 61.295 4.27 ;
      RECT 61.145 5.14 61.295 5.29 ;
      RECT 60.805 3.44 60.955 3.59 ;
      RECT 60.465 4.46 60.615 4.61 ;
      RECT 60.465 7.18 60.615 7.33 ;
      RECT 59.785 3.78 59.935 3.93 ;
      RECT 59.785 6.16 59.935 6.31 ;
      RECT 59.445 7.18 59.595 7.33 ;
      RECT 59.105 3.77 59.255 3.92 ;
      RECT 58.765 7.86 58.915 8.01 ;
      RECT 55.105 8.98 55.255 9.13 ;
      RECT 54.62 9.39 54.77 9.54 ;
      RECT 52.125 9.025 52.275 9.175 ;
      RECT 49.735 9.025 49.885 9.175 ;
      RECT 49.72 3.36 49.87 3.51 ;
      RECT 48.93 3.745 49.08 3.895 ;
      RECT 48.93 8.655 49.08 8.805 ;
      RECT 47.265 3.375 47.415 3.525 ;
      RECT 46.68 4.565 46.83 4.715 ;
      RECT 46.26 4.12 46.41 4.27 ;
      RECT 46.26 6.16 46.41 6.31 ;
      RECT 45.24 7.18 45.39 7.33 ;
      RECT 44.56 4.12 44.71 4.27 ;
      RECT 44.56 5.14 44.71 5.29 ;
      RECT 44.22 3.44 44.37 3.59 ;
      RECT 43.88 4.46 44.03 4.61 ;
      RECT 43.88 7.18 44.03 7.33 ;
      RECT 43.2 3.78 43.35 3.93 ;
      RECT 43.2 6.16 43.35 6.31 ;
      RECT 42.86 7.18 43.01 7.33 ;
      RECT 42.52 3.77 42.67 3.92 ;
      RECT 42.18 7.86 42.33 8.01 ;
      RECT 38.52 8.98 38.67 9.13 ;
      RECT 38.035 9.39 38.185 9.54 ;
      RECT 35.54 9.025 35.69 9.175 ;
      RECT 33.15 9.025 33.3 9.175 ;
      RECT 33.135 3.36 33.285 3.51 ;
      RECT 32.345 3.745 32.495 3.895 ;
      RECT 32.345 8.655 32.495 8.805 ;
      RECT 30.68 3.375 30.83 3.525 ;
      RECT 30.095 4.565 30.245 4.715 ;
      RECT 29.675 4.12 29.825 4.27 ;
      RECT 29.675 6.16 29.825 6.31 ;
      RECT 28.655 7.18 28.805 7.33 ;
      RECT 27.975 4.12 28.125 4.27 ;
      RECT 27.975 5.14 28.125 5.29 ;
      RECT 27.635 3.44 27.785 3.59 ;
      RECT 27.295 4.46 27.445 4.61 ;
      RECT 27.295 7.18 27.445 7.33 ;
      RECT 26.615 3.78 26.765 3.93 ;
      RECT 26.615 6.16 26.765 6.31 ;
      RECT 26.275 7.18 26.425 7.33 ;
      RECT 25.935 3.77 26.085 3.92 ;
      RECT 25.595 7.86 25.745 8.01 ;
      RECT 21.935 8.98 22.085 9.13 ;
      RECT 21.45 9.39 21.6 9.54 ;
      RECT 18.955 9.025 19.105 9.175 ;
      RECT 16.565 9.025 16.715 9.175 ;
      RECT 16.55 3.36 16.7 3.51 ;
      RECT 15.76 3.745 15.91 3.895 ;
      RECT 15.76 8.655 15.91 8.805 ;
      RECT 14.095 3.375 14.245 3.525 ;
      RECT 13.51 4.565 13.66 4.715 ;
      RECT 13.09 4.12 13.24 4.27 ;
      RECT 13.09 6.16 13.24 6.31 ;
      RECT 12.07 7.18 12.22 7.33 ;
      RECT 11.39 4.12 11.54 4.27 ;
      RECT 11.39 5.14 11.54 5.29 ;
      RECT 11.05 3.44 11.2 3.59 ;
      RECT 10.71 4.46 10.86 4.61 ;
      RECT 10.71 7.18 10.86 7.33 ;
      RECT 10.03 3.78 10.18 3.93 ;
      RECT 10.03 6.16 10.18 6.31 ;
      RECT 9.69 7.18 9.84 7.33 ;
      RECT 9.35 3.77 9.5 3.92 ;
      RECT 9.01 7.86 9.16 8.01 ;
      RECT 5.35 8.98 5.5 9.13 ;
      RECT 4.865 9.39 5.015 9.54 ;
      RECT 1.63 9.37 1.78 9.52 ;
      RECT 1.255 8.63 1.405 8.78 ;
    LAYER met1 ;
      RECT 85.135 10.055 85.425 10.285 ;
      RECT 85.195 8.575 85.365 10.285 ;
      RECT 85.165 9.585 85.49 9.91 ;
      RECT 85.135 8.575 85.425 8.805 ;
      RECT 84.73 3.69 84.835 4.26 ;
      RECT 84.73 4.025 85.055 4.255 ;
      RECT 84.73 4.055 85.225 4.225 ;
      RECT 84.73 3.69 84.92 4.255 ;
      RECT 84.145 3.655 84.435 3.885 ;
      RECT 84.145 3.69 84.92 3.86 ;
      RECT 84.205 2.175 84.375 3.885 ;
      RECT 84.145 2.175 84.435 2.405 ;
      RECT 84.145 10.055 84.435 10.285 ;
      RECT 84.205 8.575 84.375 10.285 ;
      RECT 84.145 8.575 84.435 8.805 ;
      RECT 84.145 8.61 85 8.77 ;
      RECT 84.83 8.205 85 8.77 ;
      RECT 84.145 8.605 84.54 8.77 ;
      RECT 84.765 8.205 85.055 8.435 ;
      RECT 84.765 8.235 85.225 8.405 ;
      RECT 83.775 4.025 84.065 4.255 ;
      RECT 83.775 4.055 84.235 4.225 ;
      RECT 83.84 2.95 84.005 4.255 ;
      RECT 82.355 2.92 82.645 3.15 ;
      RECT 82.355 2.95 84.005 3.12 ;
      RECT 82.415 2.18 82.585 3.15 ;
      RECT 82.355 2.18 82.645 2.41 ;
      RECT 82.355 10.05 82.645 10.28 ;
      RECT 82.415 9.31 82.585 10.28 ;
      RECT 82.415 9.405 84.005 9.575 ;
      RECT 83.835 8.205 84.005 9.575 ;
      RECT 82.355 9.31 82.645 9.54 ;
      RECT 83.775 8.205 84.065 8.435 ;
      RECT 83.775 8.235 84.235 8.405 ;
      RECT 80.34 3.29 80.665 3.615 ;
      RECT 82.785 3.26 83.135 3.61 ;
      RECT 80.34 3.32 83.135 3.49 ;
      RECT 82.81 8.94 83.135 9.265 ;
      RECT 82.785 8.94 83.135 9.17 ;
      RECT 82.615 8.97 83.135 9.14 ;
      RECT 82.01 3.66 82.33 3.98 ;
      RECT 81.98 3.66 82.33 3.89 ;
      RECT 81.695 3.69 82.33 3.86 ;
      RECT 82.01 8.565 82.33 8.89 ;
      RECT 81.98 8.57 82.33 8.8 ;
      RECT 81.81 8.6 82.33 8.77 ;
      RECT 79.755 4.48 80.08 4.805 ;
      RECT 76.96 4.405 77.28 4.665 ;
      RECT 78.93 4.415 79.22 4.645 ;
      RECT 79.655 4.48 80.08 4.62 ;
      RECT 76.96 4.465 79.795 4.605 ;
      RECT 79.34 4.065 79.66 4.325 ;
      RECT 79.06 4.125 79.66 4.265 ;
      RECT 78.32 7.125 78.64 7.385 ;
      RECT 78.32 7.185 78.91 7.325 ;
      RECT 77.64 4.065 77.96 4.325 ;
      RECT 72.9 4.075 73.19 4.305 ;
      RECT 72.9 4.125 77.96 4.265 ;
      RECT 77.73 3.785 77.87 4.325 ;
      RECT 77.73 3.785 78.21 3.925 ;
      RECT 78.07 3.395 78.21 3.925 ;
      RECT 77.99 3.395 78.28 3.625 ;
      RECT 77.64 5.085 77.96 5.345 ;
      RECT 76.97 5.095 77.26 5.325 ;
      RECT 74.76 5.095 75.05 5.325 ;
      RECT 74.76 5.145 77.96 5.285 ;
      RECT 75.94 7.125 76.26 7.385 ;
      RECT 77.65 7.135 77.94 7.365 ;
      RECT 75.27 7.135 75.56 7.365 ;
      RECT 75.27 7.185 76.26 7.325 ;
      RECT 77.73 6.845 77.87 7.365 ;
      RECT 76.03 6.845 76.17 7.385 ;
      RECT 76.03 6.845 77.87 6.985 ;
      RECT 74.93 3.735 75.22 3.965 ;
      RECT 75.01 3.445 75.15 3.965 ;
      RECT 77.3 3.385 77.62 3.645 ;
      RECT 77.2 3.395 77.62 3.625 ;
      RECT 75.01 3.445 77.62 3.585 ;
      RECT 76.28 3.725 76.6 3.985 ;
      RECT 76.28 3.785 76.87 3.925 ;
      RECT 75.26 7.805 75.58 8.065 ;
      RECT 74.33 7.805 76.68 7.945 ;
      RECT 76.54 7.135 76.68 7.945 ;
      RECT 74.33 7.135 74.47 7.945 ;
      RECT 76.46 7.135 76.75 7.365 ;
      RECT 74.25 7.135 74.54 7.365 ;
      RECT 76.28 6.105 76.6 6.365 ;
      RECT 73.57 6.115 73.86 6.345 ;
      RECT 73.57 6.165 76.6 6.305 ;
      RECT 75.6 3.685 75.93 4.015 ;
      RECT 75.6 3.735 76.06 3.965 ;
      RECT 75.6 3.785 76.08 3.925 ;
      RECT 75.48 3.785 75.49 3.925 ;
      RECT 75.49 3.775 76.06 3.915 ;
      RECT 71.59 8.915 71.93 9.195 ;
      RECT 71.56 8.94 71.93 9.17 ;
      RECT 71.39 8.97 71.93 9.14 ;
      RECT 71.13 10.05 71.42 10.28 ;
      RECT 71.19 9.28 71.36 10.28 ;
      RECT 71.09 9.28 71.46 9.65 ;
      RECT 68.555 10.055 68.845 10.285 ;
      RECT 68.615 8.575 68.785 10.285 ;
      RECT 68.615 8.94 68.945 9.265 ;
      RECT 68.555 8.575 68.845 8.805 ;
      RECT 68.15 3.69 68.255 4.26 ;
      RECT 68.15 4.025 68.475 4.255 ;
      RECT 68.15 4.055 68.645 4.225 ;
      RECT 68.15 3.69 68.34 4.255 ;
      RECT 67.565 3.655 67.855 3.885 ;
      RECT 67.565 3.69 68.34 3.86 ;
      RECT 67.625 2.175 67.795 3.885 ;
      RECT 67.565 2.175 67.855 2.405 ;
      RECT 67.565 10.055 67.855 10.285 ;
      RECT 67.625 8.575 67.795 10.285 ;
      RECT 67.565 8.575 67.855 8.805 ;
      RECT 67.565 8.61 68.42 8.77 ;
      RECT 68.25 8.205 68.42 8.77 ;
      RECT 67.565 8.605 67.96 8.77 ;
      RECT 68.185 8.205 68.475 8.435 ;
      RECT 68.185 8.235 68.645 8.405 ;
      RECT 67.195 4.025 67.485 4.255 ;
      RECT 67.195 4.055 67.655 4.225 ;
      RECT 67.26 2.95 67.425 4.255 ;
      RECT 65.775 2.92 66.065 3.15 ;
      RECT 65.775 2.95 67.425 3.12 ;
      RECT 65.835 2.18 66.005 3.15 ;
      RECT 65.775 2.18 66.065 2.41 ;
      RECT 65.775 10.05 66.065 10.28 ;
      RECT 65.835 9.31 66.005 10.28 ;
      RECT 65.835 9.405 67.425 9.575 ;
      RECT 67.255 8.205 67.425 9.575 ;
      RECT 65.775 9.31 66.065 9.54 ;
      RECT 67.195 8.205 67.485 8.435 ;
      RECT 67.195 8.235 67.655 8.405 ;
      RECT 63.76 3.29 64.085 3.615 ;
      RECT 66.205 3.26 66.555 3.61 ;
      RECT 63.76 3.32 66.555 3.49 ;
      RECT 66.23 8.94 66.555 9.265 ;
      RECT 66.205 8.94 66.555 9.17 ;
      RECT 66.035 8.97 66.555 9.14 ;
      RECT 65.43 3.66 65.75 3.98 ;
      RECT 65.4 3.66 65.75 3.89 ;
      RECT 65.115 3.69 65.75 3.86 ;
      RECT 65.43 8.565 65.75 8.89 ;
      RECT 65.4 8.57 65.75 8.8 ;
      RECT 65.23 8.6 65.75 8.77 ;
      RECT 63.175 4.48 63.5 4.805 ;
      RECT 60.38 4.405 60.7 4.665 ;
      RECT 62.35 4.415 62.64 4.645 ;
      RECT 63.075 4.48 63.5 4.62 ;
      RECT 60.38 4.465 63.215 4.605 ;
      RECT 62.76 4.065 63.08 4.325 ;
      RECT 62.48 4.125 63.08 4.265 ;
      RECT 61.74 7.125 62.06 7.385 ;
      RECT 61.74 7.185 62.33 7.325 ;
      RECT 61.06 4.065 61.38 4.325 ;
      RECT 56.32 4.075 56.61 4.305 ;
      RECT 56.32 4.125 61.38 4.265 ;
      RECT 61.15 3.785 61.29 4.325 ;
      RECT 61.15 3.785 61.63 3.925 ;
      RECT 61.49 3.395 61.63 3.925 ;
      RECT 61.41 3.395 61.7 3.625 ;
      RECT 61.06 5.085 61.38 5.345 ;
      RECT 60.39 5.095 60.68 5.325 ;
      RECT 58.18 5.095 58.47 5.325 ;
      RECT 58.18 5.145 61.38 5.285 ;
      RECT 59.36 7.125 59.68 7.385 ;
      RECT 61.07 7.135 61.36 7.365 ;
      RECT 58.69 7.135 58.98 7.365 ;
      RECT 58.69 7.185 59.68 7.325 ;
      RECT 61.15 6.845 61.29 7.365 ;
      RECT 59.45 6.845 59.59 7.385 ;
      RECT 59.45 6.845 61.29 6.985 ;
      RECT 58.35 3.735 58.64 3.965 ;
      RECT 58.43 3.445 58.57 3.965 ;
      RECT 60.72 3.385 61.04 3.645 ;
      RECT 60.62 3.395 61.04 3.625 ;
      RECT 58.43 3.445 61.04 3.585 ;
      RECT 59.7 3.725 60.02 3.985 ;
      RECT 59.7 3.785 60.29 3.925 ;
      RECT 58.68 7.805 59 8.065 ;
      RECT 57.75 7.805 60.1 7.945 ;
      RECT 59.96 7.135 60.1 7.945 ;
      RECT 57.75 7.135 57.89 7.945 ;
      RECT 59.88 7.135 60.17 7.365 ;
      RECT 57.67 7.135 57.96 7.365 ;
      RECT 59.7 6.105 60.02 6.365 ;
      RECT 56.99 6.115 57.28 6.345 ;
      RECT 56.99 6.165 60.02 6.305 ;
      RECT 59.02 3.685 59.35 4.015 ;
      RECT 59.02 3.735 59.48 3.965 ;
      RECT 59.02 3.785 59.5 3.925 ;
      RECT 58.9 3.785 58.91 3.925 ;
      RECT 58.91 3.775 59.48 3.915 ;
      RECT 55.01 8.915 55.35 9.195 ;
      RECT 54.98 8.94 55.35 9.17 ;
      RECT 54.81 8.97 55.35 9.14 ;
      RECT 54.55 10.05 54.84 10.28 ;
      RECT 54.61 9.28 54.78 10.28 ;
      RECT 54.51 9.28 54.88 9.65 ;
      RECT 51.97 10.055 52.26 10.285 ;
      RECT 52.03 8.575 52.2 10.285 ;
      RECT 52.03 8.94 52.36 9.265 ;
      RECT 51.97 8.575 52.26 8.805 ;
      RECT 51.565 3.69 51.67 4.26 ;
      RECT 51.565 4.025 51.89 4.255 ;
      RECT 51.565 4.055 52.06 4.225 ;
      RECT 51.565 3.69 51.755 4.255 ;
      RECT 50.98 3.655 51.27 3.885 ;
      RECT 50.98 3.69 51.755 3.86 ;
      RECT 51.04 2.175 51.21 3.885 ;
      RECT 50.98 2.175 51.27 2.405 ;
      RECT 50.98 10.055 51.27 10.285 ;
      RECT 51.04 8.575 51.21 10.285 ;
      RECT 50.98 8.575 51.27 8.805 ;
      RECT 50.98 8.61 51.835 8.77 ;
      RECT 51.665 8.205 51.835 8.77 ;
      RECT 50.98 8.605 51.375 8.77 ;
      RECT 51.6 8.205 51.89 8.435 ;
      RECT 51.6 8.235 52.06 8.405 ;
      RECT 50.61 4.025 50.9 4.255 ;
      RECT 50.61 4.055 51.07 4.225 ;
      RECT 50.675 2.95 50.84 4.255 ;
      RECT 49.19 2.92 49.48 3.15 ;
      RECT 49.19 2.95 50.84 3.12 ;
      RECT 49.25 2.18 49.42 3.15 ;
      RECT 49.19 2.18 49.48 2.41 ;
      RECT 49.19 10.05 49.48 10.28 ;
      RECT 49.25 9.31 49.42 10.28 ;
      RECT 49.25 9.405 50.84 9.575 ;
      RECT 50.67 8.205 50.84 9.575 ;
      RECT 49.19 9.31 49.48 9.54 ;
      RECT 50.61 8.205 50.9 8.435 ;
      RECT 50.61 8.235 51.07 8.405 ;
      RECT 47.175 3.29 47.5 3.615 ;
      RECT 49.62 3.26 49.97 3.61 ;
      RECT 47.175 3.32 49.97 3.49 ;
      RECT 49.645 8.94 49.97 9.265 ;
      RECT 49.62 8.94 49.97 9.17 ;
      RECT 49.45 8.97 49.97 9.14 ;
      RECT 48.845 3.66 49.165 3.98 ;
      RECT 48.815 3.66 49.165 3.89 ;
      RECT 48.53 3.69 49.165 3.86 ;
      RECT 48.845 8.565 49.165 8.89 ;
      RECT 48.815 8.57 49.165 8.8 ;
      RECT 48.645 8.6 49.165 8.77 ;
      RECT 46.59 4.48 46.915 4.805 ;
      RECT 43.795 4.405 44.115 4.665 ;
      RECT 45.765 4.415 46.055 4.645 ;
      RECT 46.49 4.48 46.915 4.62 ;
      RECT 43.795 4.465 46.63 4.605 ;
      RECT 46.175 4.065 46.495 4.325 ;
      RECT 45.895 4.125 46.495 4.265 ;
      RECT 45.155 7.125 45.475 7.385 ;
      RECT 45.155 7.185 45.745 7.325 ;
      RECT 44.475 4.065 44.795 4.325 ;
      RECT 39.735 4.075 40.025 4.305 ;
      RECT 39.735 4.125 44.795 4.265 ;
      RECT 44.565 3.785 44.705 4.325 ;
      RECT 44.565 3.785 45.045 3.925 ;
      RECT 44.905 3.395 45.045 3.925 ;
      RECT 44.825 3.395 45.115 3.625 ;
      RECT 44.475 5.085 44.795 5.345 ;
      RECT 43.805 5.095 44.095 5.325 ;
      RECT 41.595 5.095 41.885 5.325 ;
      RECT 41.595 5.145 44.795 5.285 ;
      RECT 42.775 7.125 43.095 7.385 ;
      RECT 44.485 7.135 44.775 7.365 ;
      RECT 42.105 7.135 42.395 7.365 ;
      RECT 42.105 7.185 43.095 7.325 ;
      RECT 44.565 6.845 44.705 7.365 ;
      RECT 42.865 6.845 43.005 7.385 ;
      RECT 42.865 6.845 44.705 6.985 ;
      RECT 41.765 3.735 42.055 3.965 ;
      RECT 41.845 3.445 41.985 3.965 ;
      RECT 44.135 3.385 44.455 3.645 ;
      RECT 44.035 3.395 44.455 3.625 ;
      RECT 41.845 3.445 44.455 3.585 ;
      RECT 43.115 3.725 43.435 3.985 ;
      RECT 43.115 3.785 43.705 3.925 ;
      RECT 42.095 7.805 42.415 8.065 ;
      RECT 41.165 7.805 43.515 7.945 ;
      RECT 43.375 7.135 43.515 7.945 ;
      RECT 41.165 7.135 41.305 7.945 ;
      RECT 43.295 7.135 43.585 7.365 ;
      RECT 41.085 7.135 41.375 7.365 ;
      RECT 43.115 6.105 43.435 6.365 ;
      RECT 40.405 6.115 40.695 6.345 ;
      RECT 40.405 6.165 43.435 6.305 ;
      RECT 42.435 3.685 42.765 4.015 ;
      RECT 42.435 3.735 42.895 3.965 ;
      RECT 42.435 3.785 42.915 3.925 ;
      RECT 42.315 3.785 42.325 3.925 ;
      RECT 42.325 3.775 42.895 3.915 ;
      RECT 38.425 8.915 38.765 9.195 ;
      RECT 38.395 8.94 38.765 9.17 ;
      RECT 38.225 8.97 38.765 9.14 ;
      RECT 37.965 10.05 38.255 10.28 ;
      RECT 38.025 9.28 38.195 10.28 ;
      RECT 37.925 9.28 38.295 9.65 ;
      RECT 35.385 10.055 35.675 10.285 ;
      RECT 35.445 8.575 35.615 10.285 ;
      RECT 35.445 8.94 35.775 9.265 ;
      RECT 35.385 8.575 35.675 8.805 ;
      RECT 34.98 3.69 35.085 4.26 ;
      RECT 34.98 4.025 35.305 4.255 ;
      RECT 34.98 4.055 35.475 4.225 ;
      RECT 34.98 3.69 35.17 4.255 ;
      RECT 34.395 3.655 34.685 3.885 ;
      RECT 34.395 3.69 35.17 3.86 ;
      RECT 34.455 2.175 34.625 3.885 ;
      RECT 34.395 2.175 34.685 2.405 ;
      RECT 34.395 10.055 34.685 10.285 ;
      RECT 34.455 8.575 34.625 10.285 ;
      RECT 34.395 8.575 34.685 8.805 ;
      RECT 34.395 8.61 35.25 8.77 ;
      RECT 35.08 8.205 35.25 8.77 ;
      RECT 34.395 8.605 34.79 8.77 ;
      RECT 35.015 8.205 35.305 8.435 ;
      RECT 35.015 8.235 35.475 8.405 ;
      RECT 34.025 4.025 34.315 4.255 ;
      RECT 34.025 4.055 34.485 4.225 ;
      RECT 34.09 2.95 34.255 4.255 ;
      RECT 32.605 2.92 32.895 3.15 ;
      RECT 32.605 2.95 34.255 3.12 ;
      RECT 32.665 2.18 32.835 3.15 ;
      RECT 32.605 2.18 32.895 2.41 ;
      RECT 32.605 10.05 32.895 10.28 ;
      RECT 32.665 9.31 32.835 10.28 ;
      RECT 32.665 9.405 34.255 9.575 ;
      RECT 34.085 8.205 34.255 9.575 ;
      RECT 32.605 9.31 32.895 9.54 ;
      RECT 34.025 8.205 34.315 8.435 ;
      RECT 34.025 8.235 34.485 8.405 ;
      RECT 30.59 3.29 30.915 3.615 ;
      RECT 33.035 3.26 33.385 3.61 ;
      RECT 30.59 3.32 33.385 3.49 ;
      RECT 33.06 8.94 33.385 9.265 ;
      RECT 33.035 8.94 33.385 9.17 ;
      RECT 32.865 8.97 33.385 9.14 ;
      RECT 32.26 3.66 32.58 3.98 ;
      RECT 32.23 3.66 32.58 3.89 ;
      RECT 31.945 3.69 32.58 3.86 ;
      RECT 32.26 8.565 32.58 8.89 ;
      RECT 32.23 8.57 32.58 8.8 ;
      RECT 32.06 8.6 32.58 8.77 ;
      RECT 30.005 4.48 30.33 4.805 ;
      RECT 27.21 4.405 27.53 4.665 ;
      RECT 29.18 4.415 29.47 4.645 ;
      RECT 29.905 4.48 30.33 4.62 ;
      RECT 27.21 4.465 30.045 4.605 ;
      RECT 29.59 4.065 29.91 4.325 ;
      RECT 29.31 4.125 29.91 4.265 ;
      RECT 28.57 7.125 28.89 7.385 ;
      RECT 28.57 7.185 29.16 7.325 ;
      RECT 27.89 4.065 28.21 4.325 ;
      RECT 23.15 4.075 23.44 4.305 ;
      RECT 23.15 4.125 28.21 4.265 ;
      RECT 27.98 3.785 28.12 4.325 ;
      RECT 27.98 3.785 28.46 3.925 ;
      RECT 28.32 3.395 28.46 3.925 ;
      RECT 28.24 3.395 28.53 3.625 ;
      RECT 27.89 5.085 28.21 5.345 ;
      RECT 27.22 5.095 27.51 5.325 ;
      RECT 25.01 5.095 25.3 5.325 ;
      RECT 25.01 5.145 28.21 5.285 ;
      RECT 26.19 7.125 26.51 7.385 ;
      RECT 27.9 7.135 28.19 7.365 ;
      RECT 25.52 7.135 25.81 7.365 ;
      RECT 25.52 7.185 26.51 7.325 ;
      RECT 27.98 6.845 28.12 7.365 ;
      RECT 26.28 6.845 26.42 7.385 ;
      RECT 26.28 6.845 28.12 6.985 ;
      RECT 25.18 3.735 25.47 3.965 ;
      RECT 25.26 3.445 25.4 3.965 ;
      RECT 27.55 3.385 27.87 3.645 ;
      RECT 27.45 3.395 27.87 3.625 ;
      RECT 25.26 3.445 27.87 3.585 ;
      RECT 26.53 3.725 26.85 3.985 ;
      RECT 26.53 3.785 27.12 3.925 ;
      RECT 25.51 7.805 25.83 8.065 ;
      RECT 24.58 7.805 26.93 7.945 ;
      RECT 26.79 7.135 26.93 7.945 ;
      RECT 24.58 7.135 24.72 7.945 ;
      RECT 26.71 7.135 27 7.365 ;
      RECT 24.5 7.135 24.79 7.365 ;
      RECT 26.53 6.105 26.85 6.365 ;
      RECT 23.82 6.115 24.11 6.345 ;
      RECT 23.82 6.165 26.85 6.305 ;
      RECT 25.85 3.685 26.18 4.015 ;
      RECT 25.85 3.735 26.31 3.965 ;
      RECT 25.85 3.785 26.33 3.925 ;
      RECT 25.73 3.785 25.74 3.925 ;
      RECT 25.74 3.775 26.31 3.915 ;
      RECT 21.84 8.915 22.18 9.195 ;
      RECT 21.81 8.94 22.18 9.17 ;
      RECT 21.64 8.97 22.18 9.14 ;
      RECT 21.38 10.05 21.67 10.28 ;
      RECT 21.44 9.28 21.61 10.28 ;
      RECT 21.34 9.28 21.71 9.65 ;
      RECT 18.8 10.055 19.09 10.285 ;
      RECT 18.86 8.575 19.03 10.285 ;
      RECT 18.86 8.94 19.19 9.265 ;
      RECT 18.8 8.575 19.09 8.805 ;
      RECT 18.395 3.69 18.5 4.26 ;
      RECT 18.395 4.025 18.72 4.255 ;
      RECT 18.395 4.055 18.89 4.225 ;
      RECT 18.395 3.69 18.585 4.255 ;
      RECT 17.81 3.655 18.1 3.885 ;
      RECT 17.81 3.69 18.585 3.86 ;
      RECT 17.87 2.175 18.04 3.885 ;
      RECT 17.81 2.175 18.1 2.405 ;
      RECT 17.81 10.055 18.1 10.285 ;
      RECT 17.87 8.575 18.04 10.285 ;
      RECT 17.81 8.575 18.1 8.805 ;
      RECT 17.81 8.61 18.665 8.77 ;
      RECT 18.495 8.205 18.665 8.77 ;
      RECT 17.81 8.605 18.205 8.77 ;
      RECT 18.43 8.205 18.72 8.435 ;
      RECT 18.43 8.235 18.89 8.405 ;
      RECT 17.44 4.025 17.73 4.255 ;
      RECT 17.44 4.055 17.9 4.225 ;
      RECT 17.505 2.95 17.67 4.255 ;
      RECT 16.02 2.92 16.31 3.15 ;
      RECT 16.02 2.95 17.67 3.12 ;
      RECT 16.08 2.18 16.25 3.15 ;
      RECT 16.02 2.18 16.31 2.41 ;
      RECT 16.02 10.05 16.31 10.28 ;
      RECT 16.08 9.31 16.25 10.28 ;
      RECT 16.08 9.405 17.67 9.575 ;
      RECT 17.5 8.205 17.67 9.575 ;
      RECT 16.02 9.31 16.31 9.54 ;
      RECT 17.44 8.205 17.73 8.435 ;
      RECT 17.44 8.235 17.9 8.405 ;
      RECT 14.005 3.29 14.33 3.615 ;
      RECT 16.45 3.26 16.8 3.61 ;
      RECT 14.005 3.32 16.8 3.49 ;
      RECT 16.475 8.94 16.8 9.265 ;
      RECT 16.45 8.94 16.8 9.17 ;
      RECT 16.28 8.97 16.8 9.14 ;
      RECT 15.675 3.66 15.995 3.98 ;
      RECT 15.645 3.66 15.995 3.89 ;
      RECT 15.36 3.69 15.995 3.86 ;
      RECT 15.675 8.565 15.995 8.89 ;
      RECT 15.645 8.57 15.995 8.8 ;
      RECT 15.475 8.6 15.995 8.77 ;
      RECT 13.42 4.48 13.745 4.805 ;
      RECT 10.625 4.405 10.945 4.665 ;
      RECT 12.595 4.415 12.885 4.645 ;
      RECT 13.32 4.48 13.745 4.62 ;
      RECT 10.625 4.465 13.46 4.605 ;
      RECT 13.005 4.065 13.325 4.325 ;
      RECT 12.725 4.125 13.325 4.265 ;
      RECT 11.985 7.125 12.305 7.385 ;
      RECT 11.985 7.185 12.575 7.325 ;
      RECT 11.305 4.065 11.625 4.325 ;
      RECT 6.565 4.075 6.855 4.305 ;
      RECT 6.565 4.125 11.625 4.265 ;
      RECT 11.395 3.785 11.535 4.325 ;
      RECT 11.395 3.785 11.875 3.925 ;
      RECT 11.735 3.395 11.875 3.925 ;
      RECT 11.655 3.395 11.945 3.625 ;
      RECT 11.305 5.085 11.625 5.345 ;
      RECT 10.635 5.095 10.925 5.325 ;
      RECT 8.425 5.095 8.715 5.325 ;
      RECT 8.425 5.145 11.625 5.285 ;
      RECT 9.605 7.125 9.925 7.385 ;
      RECT 11.315 7.135 11.605 7.365 ;
      RECT 8.935 7.135 9.225 7.365 ;
      RECT 8.935 7.185 9.925 7.325 ;
      RECT 11.395 6.845 11.535 7.365 ;
      RECT 9.695 6.845 9.835 7.385 ;
      RECT 9.695 6.845 11.535 6.985 ;
      RECT 8.595 3.735 8.885 3.965 ;
      RECT 8.675 3.445 8.815 3.965 ;
      RECT 10.965 3.385 11.285 3.645 ;
      RECT 10.865 3.395 11.285 3.625 ;
      RECT 8.675 3.445 11.285 3.585 ;
      RECT 9.945 3.725 10.265 3.985 ;
      RECT 9.945 3.785 10.535 3.925 ;
      RECT 8.925 7.805 9.245 8.065 ;
      RECT 7.995 7.805 10.345 7.945 ;
      RECT 10.205 7.135 10.345 7.945 ;
      RECT 7.995 7.135 8.135 7.945 ;
      RECT 10.125 7.135 10.415 7.365 ;
      RECT 7.915 7.135 8.205 7.365 ;
      RECT 9.945 6.105 10.265 6.365 ;
      RECT 7.235 6.115 7.525 6.345 ;
      RECT 7.235 6.165 10.265 6.305 ;
      RECT 9.265 3.685 9.595 4.015 ;
      RECT 9.265 3.735 9.725 3.965 ;
      RECT 9.265 3.785 9.745 3.925 ;
      RECT 9.145 3.785 9.155 3.925 ;
      RECT 9.155 3.775 9.725 3.915 ;
      RECT 5.255 8.915 5.595 9.195 ;
      RECT 5.225 8.94 5.595 9.17 ;
      RECT 5.055 8.97 5.595 9.14 ;
      RECT 4.795 10.05 5.085 10.28 ;
      RECT 4.855 9.28 5.025 10.28 ;
      RECT 4.755 9.28 5.125 9.65 ;
      RECT 1.565 10.045 1.855 10.275 ;
      RECT 1.625 9.305 1.795 10.275 ;
      RECT 1.535 9.305 1.875 9.585 ;
      RECT 1.16 8.565 1.5 8.845 ;
      RECT 1.02 8.595 1.5 8.765 ;
      RECT 79.01 6.105 79.66 6.365 ;
      RECT 76.96 7.125 77.28 7.385 ;
      RECT 62.43 6.105 63.08 6.365 ;
      RECT 60.38 7.125 60.7 7.385 ;
      RECT 45.845 6.105 46.495 6.365 ;
      RECT 43.795 7.125 44.115 7.385 ;
      RECT 29.26 6.105 29.91 6.365 ;
      RECT 27.21 7.125 27.53 7.385 ;
      RECT 12.675 6.105 13.325 6.365 ;
      RECT 10.625 7.125 10.945 7.385 ;
    LAYER mcon ;
      RECT 85.195 8.605 85.365 8.775 ;
      RECT 85.195 10.085 85.365 10.255 ;
      RECT 84.825 4.055 84.995 4.225 ;
      RECT 84.825 8.235 84.995 8.405 ;
      RECT 84.205 2.205 84.375 2.375 ;
      RECT 84.205 3.685 84.375 3.855 ;
      RECT 84.205 8.605 84.375 8.775 ;
      RECT 84.205 10.085 84.375 10.255 ;
      RECT 83.835 4.055 84.005 4.225 ;
      RECT 83.835 8.235 84.005 8.405 ;
      RECT 82.845 3.32 83.015 3.49 ;
      RECT 82.845 8.97 83.015 9.14 ;
      RECT 82.415 2.21 82.585 2.38 ;
      RECT 82.415 2.95 82.585 3.12 ;
      RECT 82.415 9.34 82.585 9.51 ;
      RECT 82.415 10.08 82.585 10.25 ;
      RECT 82.04 3.69 82.21 3.86 ;
      RECT 82.04 8.6 82.21 8.77 ;
      RECT 79.41 4.105 79.58 4.275 ;
      RECT 79.07 6.145 79.24 6.315 ;
      RECT 78.99 4.445 79.16 4.615 ;
      RECT 78.39 7.165 78.56 7.335 ;
      RECT 78.05 3.425 78.22 3.595 ;
      RECT 77.71 7.165 77.88 7.335 ;
      RECT 77.26 3.425 77.43 3.595 ;
      RECT 77.03 5.125 77.2 5.295 ;
      RECT 77.03 7.165 77.2 7.335 ;
      RECT 76.52 7.165 76.69 7.335 ;
      RECT 76.35 3.765 76.52 3.935 ;
      RECT 75.83 3.765 76 3.935 ;
      RECT 75.33 7.165 75.5 7.335 ;
      RECT 74.99 3.765 75.16 3.935 ;
      RECT 74.82 5.125 74.99 5.295 ;
      RECT 74.31 7.165 74.48 7.335 ;
      RECT 73.63 6.145 73.8 6.315 ;
      RECT 72.96 4.105 73.13 4.275 ;
      RECT 71.62 8.97 71.79 9.14 ;
      RECT 71.19 9.34 71.36 9.51 ;
      RECT 71.19 10.08 71.36 10.25 ;
      RECT 68.615 8.605 68.785 8.775 ;
      RECT 68.615 10.085 68.785 10.255 ;
      RECT 68.245 4.055 68.415 4.225 ;
      RECT 68.245 8.235 68.415 8.405 ;
      RECT 67.625 2.205 67.795 2.375 ;
      RECT 67.625 3.685 67.795 3.855 ;
      RECT 67.625 8.605 67.795 8.775 ;
      RECT 67.625 10.085 67.795 10.255 ;
      RECT 67.255 4.055 67.425 4.225 ;
      RECT 67.255 8.235 67.425 8.405 ;
      RECT 66.265 3.32 66.435 3.49 ;
      RECT 66.265 8.97 66.435 9.14 ;
      RECT 65.835 2.21 66.005 2.38 ;
      RECT 65.835 2.95 66.005 3.12 ;
      RECT 65.835 9.34 66.005 9.51 ;
      RECT 65.835 10.08 66.005 10.25 ;
      RECT 65.46 3.69 65.63 3.86 ;
      RECT 65.46 8.6 65.63 8.77 ;
      RECT 62.83 4.105 63 4.275 ;
      RECT 62.49 6.145 62.66 6.315 ;
      RECT 62.41 4.445 62.58 4.615 ;
      RECT 61.81 7.165 61.98 7.335 ;
      RECT 61.47 3.425 61.64 3.595 ;
      RECT 61.13 7.165 61.3 7.335 ;
      RECT 60.68 3.425 60.85 3.595 ;
      RECT 60.45 5.125 60.62 5.295 ;
      RECT 60.45 7.165 60.62 7.335 ;
      RECT 59.94 7.165 60.11 7.335 ;
      RECT 59.77 3.765 59.94 3.935 ;
      RECT 59.25 3.765 59.42 3.935 ;
      RECT 58.75 7.165 58.92 7.335 ;
      RECT 58.41 3.765 58.58 3.935 ;
      RECT 58.24 5.125 58.41 5.295 ;
      RECT 57.73 7.165 57.9 7.335 ;
      RECT 57.05 6.145 57.22 6.315 ;
      RECT 56.38 4.105 56.55 4.275 ;
      RECT 55.04 8.97 55.21 9.14 ;
      RECT 54.61 9.34 54.78 9.51 ;
      RECT 54.61 10.08 54.78 10.25 ;
      RECT 52.03 8.605 52.2 8.775 ;
      RECT 52.03 10.085 52.2 10.255 ;
      RECT 51.66 4.055 51.83 4.225 ;
      RECT 51.66 8.235 51.83 8.405 ;
      RECT 51.04 2.205 51.21 2.375 ;
      RECT 51.04 3.685 51.21 3.855 ;
      RECT 51.04 8.605 51.21 8.775 ;
      RECT 51.04 10.085 51.21 10.255 ;
      RECT 50.67 4.055 50.84 4.225 ;
      RECT 50.67 8.235 50.84 8.405 ;
      RECT 49.68 3.32 49.85 3.49 ;
      RECT 49.68 8.97 49.85 9.14 ;
      RECT 49.25 2.21 49.42 2.38 ;
      RECT 49.25 2.95 49.42 3.12 ;
      RECT 49.25 9.34 49.42 9.51 ;
      RECT 49.25 10.08 49.42 10.25 ;
      RECT 48.875 3.69 49.045 3.86 ;
      RECT 48.875 8.6 49.045 8.77 ;
      RECT 46.245 4.105 46.415 4.275 ;
      RECT 45.905 6.145 46.075 6.315 ;
      RECT 45.825 4.445 45.995 4.615 ;
      RECT 45.225 7.165 45.395 7.335 ;
      RECT 44.885 3.425 45.055 3.595 ;
      RECT 44.545 7.165 44.715 7.335 ;
      RECT 44.095 3.425 44.265 3.595 ;
      RECT 43.865 5.125 44.035 5.295 ;
      RECT 43.865 7.165 44.035 7.335 ;
      RECT 43.355 7.165 43.525 7.335 ;
      RECT 43.185 3.765 43.355 3.935 ;
      RECT 42.665 3.765 42.835 3.935 ;
      RECT 42.165 7.165 42.335 7.335 ;
      RECT 41.825 3.765 41.995 3.935 ;
      RECT 41.655 5.125 41.825 5.295 ;
      RECT 41.145 7.165 41.315 7.335 ;
      RECT 40.465 6.145 40.635 6.315 ;
      RECT 39.795 4.105 39.965 4.275 ;
      RECT 38.455 8.97 38.625 9.14 ;
      RECT 38.025 9.34 38.195 9.51 ;
      RECT 38.025 10.08 38.195 10.25 ;
      RECT 35.445 8.605 35.615 8.775 ;
      RECT 35.445 10.085 35.615 10.255 ;
      RECT 35.075 4.055 35.245 4.225 ;
      RECT 35.075 8.235 35.245 8.405 ;
      RECT 34.455 2.205 34.625 2.375 ;
      RECT 34.455 3.685 34.625 3.855 ;
      RECT 34.455 8.605 34.625 8.775 ;
      RECT 34.455 10.085 34.625 10.255 ;
      RECT 34.085 4.055 34.255 4.225 ;
      RECT 34.085 8.235 34.255 8.405 ;
      RECT 33.095 3.32 33.265 3.49 ;
      RECT 33.095 8.97 33.265 9.14 ;
      RECT 32.665 2.21 32.835 2.38 ;
      RECT 32.665 2.95 32.835 3.12 ;
      RECT 32.665 9.34 32.835 9.51 ;
      RECT 32.665 10.08 32.835 10.25 ;
      RECT 32.29 3.69 32.46 3.86 ;
      RECT 32.29 8.6 32.46 8.77 ;
      RECT 29.66 4.105 29.83 4.275 ;
      RECT 29.32 6.145 29.49 6.315 ;
      RECT 29.24 4.445 29.41 4.615 ;
      RECT 28.64 7.165 28.81 7.335 ;
      RECT 28.3 3.425 28.47 3.595 ;
      RECT 27.96 7.165 28.13 7.335 ;
      RECT 27.51 3.425 27.68 3.595 ;
      RECT 27.28 5.125 27.45 5.295 ;
      RECT 27.28 7.165 27.45 7.335 ;
      RECT 26.77 7.165 26.94 7.335 ;
      RECT 26.6 3.765 26.77 3.935 ;
      RECT 26.08 3.765 26.25 3.935 ;
      RECT 25.58 7.165 25.75 7.335 ;
      RECT 25.24 3.765 25.41 3.935 ;
      RECT 25.07 5.125 25.24 5.295 ;
      RECT 24.56 7.165 24.73 7.335 ;
      RECT 23.88 6.145 24.05 6.315 ;
      RECT 23.21 4.105 23.38 4.275 ;
      RECT 21.87 8.97 22.04 9.14 ;
      RECT 21.44 9.34 21.61 9.51 ;
      RECT 21.44 10.08 21.61 10.25 ;
      RECT 18.86 8.605 19.03 8.775 ;
      RECT 18.86 10.085 19.03 10.255 ;
      RECT 18.49 4.055 18.66 4.225 ;
      RECT 18.49 8.235 18.66 8.405 ;
      RECT 17.87 2.205 18.04 2.375 ;
      RECT 17.87 3.685 18.04 3.855 ;
      RECT 17.87 8.605 18.04 8.775 ;
      RECT 17.87 10.085 18.04 10.255 ;
      RECT 17.5 4.055 17.67 4.225 ;
      RECT 17.5 8.235 17.67 8.405 ;
      RECT 16.51 3.32 16.68 3.49 ;
      RECT 16.51 8.97 16.68 9.14 ;
      RECT 16.08 2.21 16.25 2.38 ;
      RECT 16.08 2.95 16.25 3.12 ;
      RECT 16.08 9.34 16.25 9.51 ;
      RECT 16.08 10.08 16.25 10.25 ;
      RECT 15.705 3.69 15.875 3.86 ;
      RECT 15.705 8.6 15.875 8.77 ;
      RECT 13.075 4.105 13.245 4.275 ;
      RECT 12.735 6.145 12.905 6.315 ;
      RECT 12.655 4.445 12.825 4.615 ;
      RECT 12.055 7.165 12.225 7.335 ;
      RECT 11.715 3.425 11.885 3.595 ;
      RECT 11.375 7.165 11.545 7.335 ;
      RECT 10.925 3.425 11.095 3.595 ;
      RECT 10.695 5.125 10.865 5.295 ;
      RECT 10.695 7.165 10.865 7.335 ;
      RECT 10.185 7.165 10.355 7.335 ;
      RECT 10.015 3.765 10.185 3.935 ;
      RECT 9.495 3.765 9.665 3.935 ;
      RECT 8.995 7.165 9.165 7.335 ;
      RECT 8.655 3.765 8.825 3.935 ;
      RECT 8.485 5.125 8.655 5.295 ;
      RECT 7.975 7.165 8.145 7.335 ;
      RECT 7.295 6.145 7.465 6.315 ;
      RECT 6.625 4.105 6.795 4.275 ;
      RECT 5.285 8.97 5.455 9.14 ;
      RECT 4.855 9.34 5.025 9.51 ;
      RECT 4.855 10.08 5.025 10.25 ;
      RECT 1.625 9.335 1.795 9.505 ;
      RECT 1.625 10.075 1.795 10.245 ;
      RECT 1.25 8.595 1.42 8.765 ;
    LAYER li1 ;
      RECT 84.825 3.035 84.995 4.225 ;
      RECT 84.825 3.035 85.295 3.205 ;
      RECT 84.825 9.255 85.295 9.425 ;
      RECT 84.825 8.235 84.995 9.425 ;
      RECT 83.835 3.035 84.005 4.225 ;
      RECT 83.835 3.035 84.305 3.205 ;
      RECT 83.835 9.255 84.305 9.425 ;
      RECT 83.835 8.235 84.005 9.425 ;
      RECT 81.985 3.93 82.155 5.16 ;
      RECT 82.04 2.15 82.21 4.1 ;
      RECT 81.985 1.87 82.155 2.32 ;
      RECT 81.985 10.14 82.155 10.59 ;
      RECT 82.04 8.36 82.21 10.31 ;
      RECT 81.985 7.3 82.155 8.53 ;
      RECT 81.465 1.87 81.635 5.16 ;
      RECT 81.465 3.37 81.87 3.7 ;
      RECT 81.465 2.53 81.87 2.86 ;
      RECT 81.465 7.3 81.635 10.59 ;
      RECT 81.465 9.6 81.87 9.93 ;
      RECT 81.465 8.76 81.87 9.09 ;
      RECT 76.72 7.935 78.03 8.185 ;
      RECT 76.72 7.615 76.9 8.185 ;
      RECT 76.17 7.615 76.9 7.785 ;
      RECT 76.17 6.775 76.34 7.785 ;
      RECT 77.01 6.815 78.75 6.995 ;
      RECT 78.42 5.975 78.75 6.995 ;
      RECT 76.17 6.775 77.23 6.945 ;
      RECT 78.42 6.145 79.24 6.315 ;
      RECT 77.58 5.975 77.91 6.185 ;
      RECT 77.58 5.975 78.75 6.145 ;
      RECT 78.48 4.495 78.81 5.455 ;
      RECT 78.48 4.495 79.16 4.665 ;
      RECT 78.99 3.255 79.16 4.665 ;
      RECT 78.9 3.255 79.23 3.895 ;
      RECT 78.03 4.765 78.3 5.465 ;
      RECT 78.13 3.255 78.3 5.465 ;
      RECT 78.47 4.075 78.82 4.325 ;
      RECT 78.13 4.105 78.82 4.275 ;
      RECT 78.04 3.255 78.3 3.735 ;
      RECT 77.37 6.405 78.25 6.645 ;
      RECT 78.02 6.315 78.25 6.645 ;
      RECT 76.72 6.405 78.25 6.605 ;
      RECT 77.64 6.355 78.25 6.645 ;
      RECT 76.72 6.275 76.89 6.605 ;
      RECT 77.61 7.165 77.86 7.765 ;
      RECT 77.61 7.165 78.08 7.365 ;
      RECT 77.1 4.385 77.86 4.885 ;
      RECT 76.17 4.195 76.43 4.815 ;
      RECT 77.09 4.325 77.1 4.635 ;
      RECT 77.07 4.315 77.09 4.605 ;
      RECT 77.73 3.995 77.96 4.595 ;
      RECT 77.05 4.265 77.07 4.575 ;
      RECT 77.03 4.385 77.96 4.565 ;
      RECT 77 4.385 77.96 4.555 ;
      RECT 76.93 4.385 77.96 4.545 ;
      RECT 76.91 4.385 77.96 4.515 ;
      RECT 76.89 3.295 77.06 4.485 ;
      RECT 76.86 4.385 77.96 4.455 ;
      RECT 76.83 4.385 77.96 4.425 ;
      RECT 76.8 4.375 77.16 4.395 ;
      RECT 76.8 4.365 77.15 4.395 ;
      RECT 76.17 4.195 77.06 4.365 ;
      RECT 76.17 4.355 77.13 4.365 ;
      RECT 76.17 4.345 77.12 4.365 ;
      RECT 76.17 4.285 77.08 4.365 ;
      RECT 76.17 3.295 77.06 3.465 ;
      RECT 77.23 3.795 77.56 4.215 ;
      RECT 77.23 3.305 77.45 4.215 ;
      RECT 77.15 7.165 77.36 7.765 ;
      RECT 77.01 7.165 77.36 7.365 ;
      RECT 75.73 4.765 76 5.465 ;
      RECT 75.95 3.255 76 5.465 ;
      RECT 75.83 4.065 76 5.465 ;
      RECT 75.83 3.255 76 4.055 ;
      RECT 75.74 3.255 76 3.735 ;
      RECT 73.87 4.425 74.12 4.965 ;
      RECT 74.84 4.425 75.56 4.895 ;
      RECT 73.87 4.425 75.66 4.595 ;
      RECT 75.43 4.065 75.66 4.595 ;
      RECT 74.43 3.305 74.68 4.595 ;
      RECT 75.43 3.995 75.49 4.895 ;
      RECT 75.43 3.995 75.66 4.055 ;
      RECT 73.89 3.305 74.68 3.575 ;
      RECT 74.85 7.115 75.53 7.365 ;
      RECT 75.26 6.755 75.53 7.365 ;
      RECT 75.01 7.535 75.34 8.085 ;
      RECT 73.95 7.535 75.34 7.725 ;
      RECT 73.95 6.695 74.12 7.725 ;
      RECT 73.83 7.115 74.12 7.445 ;
      RECT 73.95 6.695 74.89 6.865 ;
      RECT 74.59 6.145 74.89 6.865 ;
      RECT 74.85 3.725 75.26 4.245 ;
      RECT 74.85 3.305 75.05 4.245 ;
      RECT 73.46 3.485 73.63 5.465 ;
      RECT 73.46 3.995 74.26 4.245 ;
      RECT 73.46 3.485 73.71 4.245 ;
      RECT 73.38 3.485 73.71 3.905 ;
      RECT 73.41 7.895 73.97 8.185 ;
      RECT 73.41 5.975 73.66 8.185 ;
      RECT 73.41 5.975 73.87 6.525 ;
      RECT 70.24 7.3 70.41 10.59 ;
      RECT 70.24 9.6 70.645 9.93 ;
      RECT 70.24 8.76 70.645 9.09 ;
      RECT 68.245 3.035 68.415 4.225 ;
      RECT 68.245 3.035 68.715 3.205 ;
      RECT 68.245 9.255 68.715 9.425 ;
      RECT 68.245 8.235 68.415 9.425 ;
      RECT 67.255 3.035 67.425 4.225 ;
      RECT 67.255 3.035 67.725 3.205 ;
      RECT 67.255 9.255 67.725 9.425 ;
      RECT 67.255 8.235 67.425 9.425 ;
      RECT 65.405 3.93 65.575 5.16 ;
      RECT 65.46 2.15 65.63 4.1 ;
      RECT 65.405 1.87 65.575 2.32 ;
      RECT 65.405 10.14 65.575 10.59 ;
      RECT 65.46 8.36 65.63 10.31 ;
      RECT 65.405 7.3 65.575 8.53 ;
      RECT 64.885 1.87 65.055 5.16 ;
      RECT 64.885 3.37 65.29 3.7 ;
      RECT 64.885 2.53 65.29 2.86 ;
      RECT 64.885 7.3 65.055 10.59 ;
      RECT 64.885 9.6 65.29 9.93 ;
      RECT 64.885 8.76 65.29 9.09 ;
      RECT 60.14 7.935 61.45 8.185 ;
      RECT 60.14 7.615 60.32 8.185 ;
      RECT 59.59 7.615 60.32 7.785 ;
      RECT 59.59 6.775 59.76 7.785 ;
      RECT 60.43 6.815 62.17 6.995 ;
      RECT 61.84 5.975 62.17 6.995 ;
      RECT 59.59 6.775 60.65 6.945 ;
      RECT 61.84 6.145 62.66 6.315 ;
      RECT 61 5.975 61.33 6.185 ;
      RECT 61 5.975 62.17 6.145 ;
      RECT 61.9 4.495 62.23 5.455 ;
      RECT 61.9 4.495 62.58 4.665 ;
      RECT 62.41 3.255 62.58 4.665 ;
      RECT 62.32 3.255 62.65 3.895 ;
      RECT 61.45 4.765 61.72 5.465 ;
      RECT 61.55 3.255 61.72 5.465 ;
      RECT 61.89 4.075 62.24 4.325 ;
      RECT 61.55 4.105 62.24 4.275 ;
      RECT 61.46 3.255 61.72 3.735 ;
      RECT 60.79 6.405 61.67 6.645 ;
      RECT 61.44 6.315 61.67 6.645 ;
      RECT 60.14 6.405 61.67 6.605 ;
      RECT 61.06 6.355 61.67 6.645 ;
      RECT 60.14 6.275 60.31 6.605 ;
      RECT 61.03 7.165 61.28 7.765 ;
      RECT 61.03 7.165 61.5 7.365 ;
      RECT 60.52 4.385 61.28 4.885 ;
      RECT 59.59 4.195 59.85 4.815 ;
      RECT 60.51 4.325 60.52 4.635 ;
      RECT 60.49 4.315 60.51 4.605 ;
      RECT 61.15 3.995 61.38 4.595 ;
      RECT 60.47 4.265 60.49 4.575 ;
      RECT 60.45 4.385 61.38 4.565 ;
      RECT 60.42 4.385 61.38 4.555 ;
      RECT 60.35 4.385 61.38 4.545 ;
      RECT 60.33 4.385 61.38 4.515 ;
      RECT 60.31 3.295 60.48 4.485 ;
      RECT 60.28 4.385 61.38 4.455 ;
      RECT 60.25 4.385 61.38 4.425 ;
      RECT 60.22 4.375 60.58 4.395 ;
      RECT 60.22 4.365 60.57 4.395 ;
      RECT 59.59 4.195 60.48 4.365 ;
      RECT 59.59 4.355 60.55 4.365 ;
      RECT 59.59 4.345 60.54 4.365 ;
      RECT 59.59 4.285 60.5 4.365 ;
      RECT 59.59 3.295 60.48 3.465 ;
      RECT 60.65 3.795 60.98 4.215 ;
      RECT 60.65 3.305 60.87 4.215 ;
      RECT 60.57 7.165 60.78 7.765 ;
      RECT 60.43 7.165 60.78 7.365 ;
      RECT 59.15 4.765 59.42 5.465 ;
      RECT 59.37 3.255 59.42 5.465 ;
      RECT 59.25 4.065 59.42 5.465 ;
      RECT 59.25 3.255 59.42 4.055 ;
      RECT 59.16 3.255 59.42 3.735 ;
      RECT 57.29 4.425 57.54 4.965 ;
      RECT 58.26 4.425 58.98 4.895 ;
      RECT 57.29 4.425 59.08 4.595 ;
      RECT 58.85 4.065 59.08 4.595 ;
      RECT 57.85 3.305 58.1 4.595 ;
      RECT 58.85 3.995 58.91 4.895 ;
      RECT 58.85 3.995 59.08 4.055 ;
      RECT 57.31 3.305 58.1 3.575 ;
      RECT 58.27 7.115 58.95 7.365 ;
      RECT 58.68 6.755 58.95 7.365 ;
      RECT 58.43 7.535 58.76 8.085 ;
      RECT 57.37 7.535 58.76 7.725 ;
      RECT 57.37 6.695 57.54 7.725 ;
      RECT 57.25 7.115 57.54 7.445 ;
      RECT 57.37 6.695 58.31 6.865 ;
      RECT 58.01 6.145 58.31 6.865 ;
      RECT 58.27 3.725 58.68 4.245 ;
      RECT 58.27 3.305 58.47 4.245 ;
      RECT 56.88 3.485 57.05 5.465 ;
      RECT 56.88 3.995 57.68 4.245 ;
      RECT 56.88 3.485 57.13 4.245 ;
      RECT 56.8 3.485 57.13 3.905 ;
      RECT 56.83 7.895 57.39 8.185 ;
      RECT 56.83 5.975 57.08 8.185 ;
      RECT 56.83 5.975 57.29 6.525 ;
      RECT 53.66 7.3 53.83 10.59 ;
      RECT 53.66 9.6 54.065 9.93 ;
      RECT 53.66 8.76 54.065 9.09 ;
      RECT 51.66 3.035 51.83 4.225 ;
      RECT 51.66 3.035 52.13 3.205 ;
      RECT 51.66 9.255 52.13 9.425 ;
      RECT 51.66 8.235 51.83 9.425 ;
      RECT 50.67 3.035 50.84 4.225 ;
      RECT 50.67 3.035 51.14 3.205 ;
      RECT 50.67 9.255 51.14 9.425 ;
      RECT 50.67 8.235 50.84 9.425 ;
      RECT 48.82 3.93 48.99 5.16 ;
      RECT 48.875 2.15 49.045 4.1 ;
      RECT 48.82 1.87 48.99 2.32 ;
      RECT 48.82 10.14 48.99 10.59 ;
      RECT 48.875 8.36 49.045 10.31 ;
      RECT 48.82 7.3 48.99 8.53 ;
      RECT 48.3 1.87 48.47 5.16 ;
      RECT 48.3 3.37 48.705 3.7 ;
      RECT 48.3 2.53 48.705 2.86 ;
      RECT 48.3 7.3 48.47 10.59 ;
      RECT 48.3 9.6 48.705 9.93 ;
      RECT 48.3 8.76 48.705 9.09 ;
      RECT 43.555 7.935 44.865 8.185 ;
      RECT 43.555 7.615 43.735 8.185 ;
      RECT 43.005 7.615 43.735 7.785 ;
      RECT 43.005 6.775 43.175 7.785 ;
      RECT 43.845 6.815 45.585 6.995 ;
      RECT 45.255 5.975 45.585 6.995 ;
      RECT 43.005 6.775 44.065 6.945 ;
      RECT 45.255 6.145 46.075 6.315 ;
      RECT 44.415 5.975 44.745 6.185 ;
      RECT 44.415 5.975 45.585 6.145 ;
      RECT 45.315 4.495 45.645 5.455 ;
      RECT 45.315 4.495 45.995 4.665 ;
      RECT 45.825 3.255 45.995 4.665 ;
      RECT 45.735 3.255 46.065 3.895 ;
      RECT 44.865 4.765 45.135 5.465 ;
      RECT 44.965 3.255 45.135 5.465 ;
      RECT 45.305 4.075 45.655 4.325 ;
      RECT 44.965 4.105 45.655 4.275 ;
      RECT 44.875 3.255 45.135 3.735 ;
      RECT 44.205 6.405 45.085 6.645 ;
      RECT 44.855 6.315 45.085 6.645 ;
      RECT 43.555 6.405 45.085 6.605 ;
      RECT 44.475 6.355 45.085 6.645 ;
      RECT 43.555 6.275 43.725 6.605 ;
      RECT 44.445 7.165 44.695 7.765 ;
      RECT 44.445 7.165 44.915 7.365 ;
      RECT 43.935 4.385 44.695 4.885 ;
      RECT 43.005 4.195 43.265 4.815 ;
      RECT 43.925 4.325 43.935 4.635 ;
      RECT 43.905 4.315 43.925 4.605 ;
      RECT 44.565 3.995 44.795 4.595 ;
      RECT 43.885 4.265 43.905 4.575 ;
      RECT 43.865 4.385 44.795 4.565 ;
      RECT 43.835 4.385 44.795 4.555 ;
      RECT 43.765 4.385 44.795 4.545 ;
      RECT 43.745 4.385 44.795 4.515 ;
      RECT 43.725 3.295 43.895 4.485 ;
      RECT 43.695 4.385 44.795 4.455 ;
      RECT 43.665 4.385 44.795 4.425 ;
      RECT 43.635 4.375 43.995 4.395 ;
      RECT 43.635 4.365 43.985 4.395 ;
      RECT 43.005 4.195 43.895 4.365 ;
      RECT 43.005 4.355 43.965 4.365 ;
      RECT 43.005 4.345 43.955 4.365 ;
      RECT 43.005 4.285 43.915 4.365 ;
      RECT 43.005 3.295 43.895 3.465 ;
      RECT 44.065 3.795 44.395 4.215 ;
      RECT 44.065 3.305 44.285 4.215 ;
      RECT 43.985 7.165 44.195 7.765 ;
      RECT 43.845 7.165 44.195 7.365 ;
      RECT 42.565 4.765 42.835 5.465 ;
      RECT 42.785 3.255 42.835 5.465 ;
      RECT 42.665 4.065 42.835 5.465 ;
      RECT 42.665 3.255 42.835 4.055 ;
      RECT 42.575 3.255 42.835 3.735 ;
      RECT 40.705 4.425 40.955 4.965 ;
      RECT 41.675 4.425 42.395 4.895 ;
      RECT 40.705 4.425 42.495 4.595 ;
      RECT 42.265 4.065 42.495 4.595 ;
      RECT 41.265 3.305 41.515 4.595 ;
      RECT 42.265 3.995 42.325 4.895 ;
      RECT 42.265 3.995 42.495 4.055 ;
      RECT 40.725 3.305 41.515 3.575 ;
      RECT 41.685 7.115 42.365 7.365 ;
      RECT 42.095 6.755 42.365 7.365 ;
      RECT 41.845 7.535 42.175 8.085 ;
      RECT 40.785 7.535 42.175 7.725 ;
      RECT 40.785 6.695 40.955 7.725 ;
      RECT 40.665 7.115 40.955 7.445 ;
      RECT 40.785 6.695 41.725 6.865 ;
      RECT 41.425 6.145 41.725 6.865 ;
      RECT 41.685 3.725 42.095 4.245 ;
      RECT 41.685 3.305 41.885 4.245 ;
      RECT 40.295 3.485 40.465 5.465 ;
      RECT 40.295 3.995 41.095 4.245 ;
      RECT 40.295 3.485 40.545 4.245 ;
      RECT 40.215 3.485 40.545 3.905 ;
      RECT 40.245 7.895 40.805 8.185 ;
      RECT 40.245 5.975 40.495 8.185 ;
      RECT 40.245 5.975 40.705 6.525 ;
      RECT 37.075 7.3 37.245 10.59 ;
      RECT 37.075 9.6 37.48 9.93 ;
      RECT 37.075 8.76 37.48 9.09 ;
      RECT 35.075 3.035 35.245 4.225 ;
      RECT 35.075 3.035 35.545 3.205 ;
      RECT 35.075 9.255 35.545 9.425 ;
      RECT 35.075 8.235 35.245 9.425 ;
      RECT 34.085 3.035 34.255 4.225 ;
      RECT 34.085 3.035 34.555 3.205 ;
      RECT 34.085 9.255 34.555 9.425 ;
      RECT 34.085 8.235 34.255 9.425 ;
      RECT 32.235 3.93 32.405 5.16 ;
      RECT 32.29 2.15 32.46 4.1 ;
      RECT 32.235 1.87 32.405 2.32 ;
      RECT 32.235 10.14 32.405 10.59 ;
      RECT 32.29 8.36 32.46 10.31 ;
      RECT 32.235 7.3 32.405 8.53 ;
      RECT 31.715 1.87 31.885 5.16 ;
      RECT 31.715 3.37 32.12 3.7 ;
      RECT 31.715 2.53 32.12 2.86 ;
      RECT 31.715 7.3 31.885 10.59 ;
      RECT 31.715 9.6 32.12 9.93 ;
      RECT 31.715 8.76 32.12 9.09 ;
      RECT 26.97 7.935 28.28 8.185 ;
      RECT 26.97 7.615 27.15 8.185 ;
      RECT 26.42 7.615 27.15 7.785 ;
      RECT 26.42 6.775 26.59 7.785 ;
      RECT 27.26 6.815 29 6.995 ;
      RECT 28.67 5.975 29 6.995 ;
      RECT 26.42 6.775 27.48 6.945 ;
      RECT 28.67 6.145 29.49 6.315 ;
      RECT 27.83 5.975 28.16 6.185 ;
      RECT 27.83 5.975 29 6.145 ;
      RECT 28.73 4.495 29.06 5.455 ;
      RECT 28.73 4.495 29.41 4.665 ;
      RECT 29.24 3.255 29.41 4.665 ;
      RECT 29.15 3.255 29.48 3.895 ;
      RECT 28.28 4.765 28.55 5.465 ;
      RECT 28.38 3.255 28.55 5.465 ;
      RECT 28.72 4.075 29.07 4.325 ;
      RECT 28.38 4.105 29.07 4.275 ;
      RECT 28.29 3.255 28.55 3.735 ;
      RECT 27.62 6.405 28.5 6.645 ;
      RECT 28.27 6.315 28.5 6.645 ;
      RECT 26.97 6.405 28.5 6.605 ;
      RECT 27.89 6.355 28.5 6.645 ;
      RECT 26.97 6.275 27.14 6.605 ;
      RECT 27.86 7.165 28.11 7.765 ;
      RECT 27.86 7.165 28.33 7.365 ;
      RECT 27.35 4.385 28.11 4.885 ;
      RECT 26.42 4.195 26.68 4.815 ;
      RECT 27.34 4.325 27.35 4.635 ;
      RECT 27.32 4.315 27.34 4.605 ;
      RECT 27.98 3.995 28.21 4.595 ;
      RECT 27.3 4.265 27.32 4.575 ;
      RECT 27.28 4.385 28.21 4.565 ;
      RECT 27.25 4.385 28.21 4.555 ;
      RECT 27.18 4.385 28.21 4.545 ;
      RECT 27.16 4.385 28.21 4.515 ;
      RECT 27.14 3.295 27.31 4.485 ;
      RECT 27.11 4.385 28.21 4.455 ;
      RECT 27.08 4.385 28.21 4.425 ;
      RECT 27.05 4.375 27.41 4.395 ;
      RECT 27.05 4.365 27.4 4.395 ;
      RECT 26.42 4.195 27.31 4.365 ;
      RECT 26.42 4.355 27.38 4.365 ;
      RECT 26.42 4.345 27.37 4.365 ;
      RECT 26.42 4.285 27.33 4.365 ;
      RECT 26.42 3.295 27.31 3.465 ;
      RECT 27.48 3.795 27.81 4.215 ;
      RECT 27.48 3.305 27.7 4.215 ;
      RECT 27.4 7.165 27.61 7.765 ;
      RECT 27.26 7.165 27.61 7.365 ;
      RECT 25.98 4.765 26.25 5.465 ;
      RECT 26.2 3.255 26.25 5.465 ;
      RECT 26.08 4.065 26.25 5.465 ;
      RECT 26.08 3.255 26.25 4.055 ;
      RECT 25.99 3.255 26.25 3.735 ;
      RECT 24.12 4.425 24.37 4.965 ;
      RECT 25.09 4.425 25.81 4.895 ;
      RECT 24.12 4.425 25.91 4.595 ;
      RECT 25.68 4.065 25.91 4.595 ;
      RECT 24.68 3.305 24.93 4.595 ;
      RECT 25.68 3.995 25.74 4.895 ;
      RECT 25.68 3.995 25.91 4.055 ;
      RECT 24.14 3.305 24.93 3.575 ;
      RECT 25.1 7.115 25.78 7.365 ;
      RECT 25.51 6.755 25.78 7.365 ;
      RECT 25.26 7.535 25.59 8.085 ;
      RECT 24.2 7.535 25.59 7.725 ;
      RECT 24.2 6.695 24.37 7.725 ;
      RECT 24.08 7.115 24.37 7.445 ;
      RECT 24.2 6.695 25.14 6.865 ;
      RECT 24.84 6.145 25.14 6.865 ;
      RECT 25.1 3.725 25.51 4.245 ;
      RECT 25.1 3.305 25.3 4.245 ;
      RECT 23.71 3.485 23.88 5.465 ;
      RECT 23.71 3.995 24.51 4.245 ;
      RECT 23.71 3.485 23.96 4.245 ;
      RECT 23.63 3.485 23.96 3.905 ;
      RECT 23.66 7.895 24.22 8.185 ;
      RECT 23.66 5.975 23.91 8.185 ;
      RECT 23.66 5.975 24.12 6.525 ;
      RECT 20.49 7.3 20.66 10.59 ;
      RECT 20.49 9.6 20.895 9.93 ;
      RECT 20.49 8.76 20.895 9.09 ;
      RECT 18.49 3.035 18.66 4.225 ;
      RECT 18.49 3.035 18.96 3.205 ;
      RECT 18.49 9.255 18.96 9.425 ;
      RECT 18.49 8.235 18.66 9.425 ;
      RECT 17.5 3.035 17.67 4.225 ;
      RECT 17.5 3.035 17.97 3.205 ;
      RECT 17.5 9.255 17.97 9.425 ;
      RECT 17.5 8.235 17.67 9.425 ;
      RECT 15.65 3.93 15.82 5.16 ;
      RECT 15.705 2.15 15.875 4.1 ;
      RECT 15.65 1.87 15.82 2.32 ;
      RECT 15.65 10.14 15.82 10.59 ;
      RECT 15.705 8.36 15.875 10.31 ;
      RECT 15.65 7.3 15.82 8.53 ;
      RECT 15.13 1.87 15.3 5.16 ;
      RECT 15.13 3.37 15.535 3.7 ;
      RECT 15.13 2.53 15.535 2.86 ;
      RECT 15.13 7.3 15.3 10.59 ;
      RECT 15.13 9.6 15.535 9.93 ;
      RECT 15.13 8.76 15.535 9.09 ;
      RECT 10.385 7.935 11.695 8.185 ;
      RECT 10.385 7.615 10.565 8.185 ;
      RECT 9.835 7.615 10.565 7.785 ;
      RECT 9.835 6.775 10.005 7.785 ;
      RECT 10.675 6.815 12.415 6.995 ;
      RECT 12.085 5.975 12.415 6.995 ;
      RECT 9.835 6.775 10.895 6.945 ;
      RECT 12.085 6.145 12.905 6.315 ;
      RECT 11.245 5.975 11.575 6.185 ;
      RECT 11.245 5.975 12.415 6.145 ;
      RECT 12.145 4.495 12.475 5.455 ;
      RECT 12.145 4.495 12.825 4.665 ;
      RECT 12.655 3.255 12.825 4.665 ;
      RECT 12.565 3.255 12.895 3.895 ;
      RECT 11.695 4.765 11.965 5.465 ;
      RECT 11.795 3.255 11.965 5.465 ;
      RECT 12.135 4.075 12.485 4.325 ;
      RECT 11.795 4.105 12.485 4.275 ;
      RECT 11.705 3.255 11.965 3.735 ;
      RECT 11.035 6.405 11.915 6.645 ;
      RECT 11.685 6.315 11.915 6.645 ;
      RECT 10.385 6.405 11.915 6.605 ;
      RECT 11.305 6.355 11.915 6.645 ;
      RECT 10.385 6.275 10.555 6.605 ;
      RECT 11.275 7.165 11.525 7.765 ;
      RECT 11.275 7.165 11.745 7.365 ;
      RECT 10.765 4.385 11.525 4.885 ;
      RECT 9.835 4.195 10.095 4.815 ;
      RECT 10.755 4.325 10.765 4.635 ;
      RECT 10.735 4.315 10.755 4.605 ;
      RECT 11.395 3.995 11.625 4.595 ;
      RECT 10.715 4.265 10.735 4.575 ;
      RECT 10.695 4.385 11.625 4.565 ;
      RECT 10.665 4.385 11.625 4.555 ;
      RECT 10.595 4.385 11.625 4.545 ;
      RECT 10.575 4.385 11.625 4.515 ;
      RECT 10.555 3.295 10.725 4.485 ;
      RECT 10.525 4.385 11.625 4.455 ;
      RECT 10.495 4.385 11.625 4.425 ;
      RECT 10.465 4.375 10.825 4.395 ;
      RECT 10.465 4.365 10.815 4.395 ;
      RECT 9.835 4.195 10.725 4.365 ;
      RECT 9.835 4.355 10.795 4.365 ;
      RECT 9.835 4.345 10.785 4.365 ;
      RECT 9.835 4.285 10.745 4.365 ;
      RECT 9.835 3.295 10.725 3.465 ;
      RECT 10.895 3.795 11.225 4.215 ;
      RECT 10.895 3.305 11.115 4.215 ;
      RECT 10.815 7.165 11.025 7.765 ;
      RECT 10.675 7.165 11.025 7.365 ;
      RECT 9.395 4.765 9.665 5.465 ;
      RECT 9.615 3.255 9.665 5.465 ;
      RECT 9.495 4.065 9.665 5.465 ;
      RECT 9.495 3.255 9.665 4.055 ;
      RECT 9.405 3.255 9.665 3.735 ;
      RECT 7.535 4.425 7.785 4.965 ;
      RECT 8.505 4.425 9.225 4.895 ;
      RECT 7.535 4.425 9.325 4.595 ;
      RECT 9.095 4.065 9.325 4.595 ;
      RECT 8.095 3.305 8.345 4.595 ;
      RECT 9.095 3.995 9.155 4.895 ;
      RECT 9.095 3.995 9.325 4.055 ;
      RECT 7.555 3.305 8.345 3.575 ;
      RECT 8.515 7.115 9.195 7.365 ;
      RECT 8.925 6.755 9.195 7.365 ;
      RECT 8.675 7.535 9.005 8.085 ;
      RECT 7.615 7.535 9.005 7.725 ;
      RECT 7.615 6.695 7.785 7.725 ;
      RECT 7.495 7.115 7.785 7.445 ;
      RECT 7.615 6.695 8.555 6.865 ;
      RECT 8.255 6.145 8.555 6.865 ;
      RECT 8.515 3.725 8.925 4.245 ;
      RECT 8.515 3.305 8.715 4.245 ;
      RECT 7.125 3.485 7.295 5.465 ;
      RECT 7.125 3.995 7.925 4.245 ;
      RECT 7.125 3.485 7.375 4.245 ;
      RECT 7.045 3.485 7.375 3.905 ;
      RECT 7.075 7.895 7.635 8.185 ;
      RECT 7.075 5.975 7.325 8.185 ;
      RECT 7.075 5.975 7.535 6.525 ;
      RECT 3.905 7.3 4.075 10.59 ;
      RECT 3.905 9.6 4.31 9.93 ;
      RECT 3.905 8.76 4.31 9.09 ;
      RECT 1.195 10.135 1.365 10.585 ;
      RECT 1.25 8.355 1.42 10.305 ;
      RECT 1.195 7.295 1.365 8.525 ;
      RECT 0.675 7.295 0.845 10.585 ;
      RECT 0.675 9.595 1.08 9.925 ;
      RECT 0.675 8.755 1.08 9.085 ;
      RECT 85.195 7.305 85.365 8.775 ;
      RECT 85.195 10.085 85.365 10.595 ;
      RECT 84.205 1.865 84.375 2.375 ;
      RECT 84.205 3.685 84.375 5.155 ;
      RECT 84.205 7.305 84.375 8.775 ;
      RECT 84.205 10.085 84.375 10.595 ;
      RECT 82.845 1.87 83.015 5.16 ;
      RECT 82.845 7.3 83.015 10.59 ;
      RECT 82.415 1.87 82.585 2.38 ;
      RECT 82.415 2.95 82.585 5.16 ;
      RECT 82.415 7.3 82.585 9.51 ;
      RECT 82.415 10.08 82.585 10.59 ;
      RECT 79.33 4.075 79.68 4.325 ;
      RECT 78.27 7.165 78.72 7.675 ;
      RECT 76.95 5.125 77.43 5.465 ;
      RECT 76.51 7.115 76.84 7.445 ;
      RECT 76.17 3.635 76.72 4.025 ;
      RECT 74.66 5.125 75.13 5.465 ;
      RECT 74.29 7.115 74.63 7.365 ;
      RECT 72.95 4.075 73.29 4.955 ;
      RECT 71.62 7.3 71.79 10.59 ;
      RECT 71.19 7.3 71.36 9.51 ;
      RECT 71.19 10.08 71.36 10.59 ;
      RECT 68.615 7.305 68.785 8.775 ;
      RECT 68.615 10.085 68.785 10.595 ;
      RECT 67.625 1.865 67.795 2.375 ;
      RECT 67.625 3.685 67.795 5.155 ;
      RECT 67.625 7.305 67.795 8.775 ;
      RECT 67.625 10.085 67.795 10.595 ;
      RECT 66.265 1.87 66.435 5.16 ;
      RECT 66.265 7.3 66.435 10.59 ;
      RECT 65.835 1.87 66.005 2.38 ;
      RECT 65.835 2.95 66.005 5.16 ;
      RECT 65.835 7.3 66.005 9.51 ;
      RECT 65.835 10.08 66.005 10.59 ;
      RECT 62.75 4.075 63.1 4.325 ;
      RECT 61.69 7.165 62.14 7.675 ;
      RECT 60.37 5.125 60.85 5.465 ;
      RECT 59.93 7.115 60.26 7.445 ;
      RECT 59.59 3.635 60.14 4.025 ;
      RECT 58.08 5.125 58.55 5.465 ;
      RECT 57.71 7.115 58.05 7.365 ;
      RECT 56.37 4.075 56.71 4.955 ;
      RECT 55.04 7.3 55.21 10.59 ;
      RECT 54.61 7.3 54.78 9.51 ;
      RECT 54.61 10.08 54.78 10.59 ;
      RECT 52.03 7.305 52.2 8.775 ;
      RECT 52.03 10.085 52.2 10.595 ;
      RECT 51.04 1.865 51.21 2.375 ;
      RECT 51.04 3.685 51.21 5.155 ;
      RECT 51.04 7.305 51.21 8.775 ;
      RECT 51.04 10.085 51.21 10.595 ;
      RECT 49.68 1.87 49.85 5.16 ;
      RECT 49.68 7.3 49.85 10.59 ;
      RECT 49.25 1.87 49.42 2.38 ;
      RECT 49.25 2.95 49.42 5.16 ;
      RECT 49.25 7.3 49.42 9.51 ;
      RECT 49.25 10.08 49.42 10.59 ;
      RECT 46.165 4.075 46.515 4.325 ;
      RECT 45.105 7.165 45.555 7.675 ;
      RECT 43.785 5.125 44.265 5.465 ;
      RECT 43.345 7.115 43.675 7.445 ;
      RECT 43.005 3.635 43.555 4.025 ;
      RECT 41.495 5.125 41.965 5.465 ;
      RECT 41.125 7.115 41.465 7.365 ;
      RECT 39.785 4.075 40.125 4.955 ;
      RECT 38.455 7.3 38.625 10.59 ;
      RECT 38.025 7.3 38.195 9.51 ;
      RECT 38.025 10.08 38.195 10.59 ;
      RECT 35.445 7.305 35.615 8.775 ;
      RECT 35.445 10.085 35.615 10.595 ;
      RECT 34.455 1.865 34.625 2.375 ;
      RECT 34.455 3.685 34.625 5.155 ;
      RECT 34.455 7.305 34.625 8.775 ;
      RECT 34.455 10.085 34.625 10.595 ;
      RECT 33.095 1.87 33.265 5.16 ;
      RECT 33.095 7.3 33.265 10.59 ;
      RECT 32.665 1.87 32.835 2.38 ;
      RECT 32.665 2.95 32.835 5.16 ;
      RECT 32.665 7.3 32.835 9.51 ;
      RECT 32.665 10.08 32.835 10.59 ;
      RECT 29.58 4.075 29.93 4.325 ;
      RECT 28.52 7.165 28.97 7.675 ;
      RECT 27.2 5.125 27.68 5.465 ;
      RECT 26.76 7.115 27.09 7.445 ;
      RECT 26.42 3.635 26.97 4.025 ;
      RECT 24.91 5.125 25.38 5.465 ;
      RECT 24.54 7.115 24.88 7.365 ;
      RECT 23.2 4.075 23.54 4.955 ;
      RECT 21.87 7.3 22.04 10.59 ;
      RECT 21.44 7.3 21.61 9.51 ;
      RECT 21.44 10.08 21.61 10.59 ;
      RECT 18.86 7.305 19.03 8.775 ;
      RECT 18.86 10.085 19.03 10.595 ;
      RECT 17.87 1.865 18.04 2.375 ;
      RECT 17.87 3.685 18.04 5.155 ;
      RECT 17.87 7.305 18.04 8.775 ;
      RECT 17.87 10.085 18.04 10.595 ;
      RECT 16.51 1.87 16.68 5.16 ;
      RECT 16.51 7.3 16.68 10.59 ;
      RECT 16.08 1.87 16.25 2.38 ;
      RECT 16.08 2.95 16.25 5.16 ;
      RECT 16.08 7.3 16.25 9.51 ;
      RECT 16.08 10.08 16.25 10.59 ;
      RECT 12.995 4.075 13.345 4.325 ;
      RECT 11.935 7.165 12.385 7.675 ;
      RECT 10.615 5.125 11.095 5.465 ;
      RECT 10.175 7.115 10.505 7.445 ;
      RECT 9.835 3.635 10.385 4.025 ;
      RECT 8.325 5.125 8.795 5.465 ;
      RECT 7.955 7.115 8.295 7.365 ;
      RECT 6.615 4.075 6.955 4.955 ;
      RECT 5.285 7.3 5.455 10.59 ;
      RECT 4.855 7.3 5.025 9.51 ;
      RECT 4.855 10.08 5.025 10.59 ;
      RECT 1.625 7.295 1.795 9.505 ;
      RECT 1.625 10.075 1.795 10.585 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  ORIGIN -9.95 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r2 ;
  SIZE 86.085 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 29.155 1.87 29.325 2.38 ;
        RECT 29.155 3.69 29.325 5.16 ;
      LAYER met1 ;
        RECT 29.095 3.66 29.385 3.89 ;
        RECT 29.095 2.18 29.385 2.41 ;
        RECT 29.155 2.18 29.325 3.89 ;
      LAYER mcon ;
        RECT 29.155 3.69 29.325 3.86 ;
        RECT 29.155 2.21 29.325 2.38 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 45.74 1.87 45.91 2.38 ;
        RECT 45.74 3.69 45.91 5.16 ;
      LAYER met1 ;
        RECT 45.68 3.66 45.97 3.89 ;
        RECT 45.68 2.18 45.97 2.41 ;
        RECT 45.74 2.18 45.91 3.89 ;
      LAYER mcon ;
        RECT 45.74 3.69 45.91 3.86 ;
        RECT 45.74 2.21 45.91 2.38 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 62.325 1.87 62.495 2.38 ;
        RECT 62.325 3.69 62.495 5.16 ;
      LAYER met1 ;
        RECT 62.265 3.66 62.555 3.89 ;
        RECT 62.265 2.18 62.555 2.41 ;
        RECT 62.325 2.18 62.495 3.89 ;
      LAYER mcon ;
        RECT 62.325 3.69 62.495 3.86 ;
        RECT 62.325 2.21 62.495 2.38 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 78.91 1.87 79.08 2.38 ;
        RECT 78.91 3.69 79.08 5.16 ;
      LAYER met1 ;
        RECT 78.85 3.66 79.14 3.89 ;
        RECT 78.85 2.18 79.14 2.41 ;
        RECT 78.91 2.18 79.08 3.89 ;
      LAYER mcon ;
        RECT 78.91 3.69 79.08 3.86 ;
        RECT 78.91 2.21 79.08 2.38 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 95.49 1.87 95.66 2.38 ;
        RECT 95.49 3.69 95.66 5.16 ;
      LAYER met1 ;
        RECT 95.43 3.66 95.72 3.89 ;
        RECT 95.43 2.18 95.72 2.41 ;
        RECT 95.49 2.18 95.66 3.89 ;
      LAYER mcon ;
        RECT 95.49 3.69 95.66 3.86 ;
        RECT 95.49 2.21 95.66 2.38 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 25.005 2.955 25.175 4.23 ;
        RECT 25.005 8.23 25.175 9.505 ;
        RECT 13.78 8.23 13.95 9.505 ;
      LAYER met2 ;
        RECT 24.93 8.15 25.255 8.475 ;
        RECT 24.925 4.93 25.25 5.255 ;
        RECT 16.085 9.3 25.17 9.47 ;
        RECT 24.995 4.93 25.17 9.47 ;
        RECT 16.03 8.145 16.31 8.485 ;
        RECT 16.085 8.145 16.255 9.47 ;
      LAYER met1 ;
        RECT 24.945 4.06 25.405 4.23 ;
        RECT 24.925 4.93 25.25 5.255 ;
        RECT 24.945 4.03 25.235 4.26 ;
        RECT 25 4.03 25.18 5.255 ;
        RECT 24.93 8.23 25.405 8.4 ;
        RECT 24.93 8.15 25.255 8.475 ;
        RECT 16 8.175 16.34 8.455 ;
        RECT 13.72 8.23 16.34 8.4 ;
        RECT 13.72 8.2 14.01 8.43 ;
      LAYER via1 ;
        RECT 16.095 8.24 16.245 8.39 ;
        RECT 25.015 5.015 25.165 5.165 ;
        RECT 25.02 8.235 25.17 8.385 ;
      LAYER mcon ;
        RECT 13.78 8.23 13.95 8.4 ;
        RECT 25.005 8.23 25.175 8.4 ;
        RECT 25.005 4.06 25.175 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 41.59 2.955 41.76 4.23 ;
        RECT 41.59 8.23 41.76 9.505 ;
        RECT 30.365 8.23 30.535 9.505 ;
      LAYER met2 ;
        RECT 41.515 8.15 41.84 8.475 ;
        RECT 41.51 4.93 41.835 5.255 ;
        RECT 32.67 9.3 41.755 9.47 ;
        RECT 41.58 4.93 41.755 9.47 ;
        RECT 32.615 8.145 32.895 8.485 ;
        RECT 32.67 8.145 32.84 9.47 ;
      LAYER met1 ;
        RECT 41.53 4.06 41.99 4.23 ;
        RECT 41.51 4.93 41.835 5.255 ;
        RECT 41.53 4.03 41.82 4.26 ;
        RECT 41.585 4.03 41.765 5.255 ;
        RECT 41.515 8.23 41.99 8.4 ;
        RECT 41.515 8.15 41.84 8.475 ;
        RECT 32.585 8.175 32.925 8.455 ;
        RECT 30.305 8.23 32.925 8.4 ;
        RECT 30.305 8.2 30.595 8.43 ;
      LAYER via1 ;
        RECT 32.68 8.24 32.83 8.39 ;
        RECT 41.6 5.015 41.75 5.165 ;
        RECT 41.605 8.235 41.755 8.385 ;
      LAYER mcon ;
        RECT 30.365 8.23 30.535 8.4 ;
        RECT 41.59 8.23 41.76 8.4 ;
        RECT 41.59 4.06 41.76 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 58.175 2.955 58.345 4.23 ;
        RECT 58.175 8.23 58.345 9.505 ;
        RECT 46.95 8.23 47.12 9.505 ;
      LAYER met2 ;
        RECT 58.1 8.15 58.425 8.475 ;
        RECT 58.095 4.93 58.42 5.255 ;
        RECT 49.255 9.3 58.34 9.47 ;
        RECT 58.165 4.93 58.34 9.47 ;
        RECT 49.2 8.145 49.48 8.485 ;
        RECT 49.255 8.145 49.425 9.47 ;
      LAYER met1 ;
        RECT 58.115 4.06 58.575 4.23 ;
        RECT 58.095 4.93 58.42 5.255 ;
        RECT 58.115 4.03 58.405 4.26 ;
        RECT 58.17 4.03 58.35 5.255 ;
        RECT 58.1 8.23 58.575 8.4 ;
        RECT 58.1 8.15 58.425 8.475 ;
        RECT 49.17 8.175 49.51 8.455 ;
        RECT 46.89 8.23 49.51 8.4 ;
        RECT 46.89 8.2 47.18 8.43 ;
      LAYER via1 ;
        RECT 49.265 8.24 49.415 8.39 ;
        RECT 58.185 5.015 58.335 5.165 ;
        RECT 58.19 8.235 58.34 8.385 ;
      LAYER mcon ;
        RECT 46.95 8.23 47.12 8.4 ;
        RECT 58.175 8.23 58.345 8.4 ;
        RECT 58.175 4.06 58.345 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 74.76 2.955 74.93 4.23 ;
        RECT 74.76 8.23 74.93 9.505 ;
        RECT 63.535 8.23 63.705 9.505 ;
      LAYER met2 ;
        RECT 74.685 8.15 75.01 8.475 ;
        RECT 74.68 4.93 75.005 5.255 ;
        RECT 65.84 9.3 74.925 9.47 ;
        RECT 74.75 4.93 74.925 9.47 ;
        RECT 65.785 8.145 66.065 8.485 ;
        RECT 65.84 8.145 66.01 9.47 ;
      LAYER met1 ;
        RECT 74.7 4.06 75.16 4.23 ;
        RECT 74.68 4.93 75.005 5.255 ;
        RECT 74.7 4.03 74.99 4.26 ;
        RECT 74.755 4.03 74.935 5.255 ;
        RECT 74.685 8.23 75.16 8.4 ;
        RECT 74.685 8.15 75.01 8.475 ;
        RECT 65.755 8.175 66.095 8.455 ;
        RECT 63.475 8.23 66.095 8.4 ;
        RECT 63.475 8.2 63.765 8.43 ;
      LAYER via1 ;
        RECT 65.85 8.24 66 8.39 ;
        RECT 74.77 5.015 74.92 5.165 ;
        RECT 74.775 8.235 74.925 8.385 ;
      LAYER mcon ;
        RECT 63.535 8.23 63.705 8.4 ;
        RECT 74.76 8.23 74.93 8.4 ;
        RECT 74.76 4.06 74.93 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 91.34 2.955 91.51 4.23 ;
        RECT 91.34 8.23 91.51 9.505 ;
        RECT 80.115 8.23 80.285 9.505 ;
      LAYER met2 ;
        RECT 91.265 8.15 91.59 8.475 ;
        RECT 91.26 4.93 91.585 5.255 ;
        RECT 82.42 9.3 91.505 9.47 ;
        RECT 91.33 4.93 91.505 9.47 ;
        RECT 82.365 8.145 82.645 8.485 ;
        RECT 82.42 8.145 82.59 9.47 ;
      LAYER met1 ;
        RECT 91.28 4.06 91.74 4.23 ;
        RECT 91.26 4.93 91.585 5.255 ;
        RECT 91.28 4.03 91.57 4.26 ;
        RECT 91.335 4.03 91.515 5.255 ;
        RECT 91.265 8.23 91.74 8.4 ;
        RECT 91.265 8.15 91.59 8.475 ;
        RECT 82.335 8.175 82.675 8.455 ;
        RECT 80.055 8.23 82.675 8.4 ;
        RECT 80.055 8.2 80.345 8.43 ;
      LAYER via1 ;
        RECT 82.43 8.24 82.58 8.39 ;
        RECT 91.35 5.015 91.5 5.165 ;
        RECT 91.355 8.235 91.505 8.385 ;
      LAYER mcon ;
        RECT 80.115 8.23 80.285 8.4 ;
        RECT 91.34 8.23 91.51 8.4 ;
        RECT 91.34 4.06 91.51 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 10.55 8.23 10.72 9.505 ;
      LAYER met1 ;
        RECT 10.49 8.23 10.95 8.4 ;
        RECT 10.49 8.2 10.78 8.43 ;
      LAYER mcon ;
        RECT 10.55 8.23 10.72 8.4 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 90.095 5.43 96.035 7.04 ;
        RECT 95.06 4.7 95.23 7.765 ;
        RECT 94.07 4.7 94.24 7.765 ;
        RECT 91.33 4.7 91.5 7.76 ;
        RECT 89.965 5.43 96.035 5.965 ;
        RECT 89.635 4.495 89.965 5.805 ;
        RECT 10.155 5.635 96.035 5.805 ;
        RECT 87.895 5.095 88.155 5.805 ;
        RECT 87.335 5.635 87.705 6.185 ;
        RECT 86.895 4.715 87.225 4.955 ;
        RECT 86.895 4.715 87.085 5.085 ;
        RECT 86.465 4.985 87.075 5.805 ;
        RECT 86.515 4.985 86.785 6.585 ;
        RECT 85.595 5.095 85.815 5.805 ;
        RECT 85.355 5.635 85.635 6.475 ;
        RECT 84.585 4.765 84.915 4.955 ;
        RECT 84.165 5.135 84.785 5.805 ;
        RECT 84.585 4.765 84.785 5.805 ;
        RECT 84.355 5.135 84.685 6.525 ;
        RECT 83.245 5.125 83.505 5.805 ;
        RECT 73.515 5.43 83.28 7.03 ;
        RECT 79.45 5.425 83.025 7.03 ;
        RECT 80.105 5.425 80.275 7.76 ;
        RECT 73.515 5.43 79.455 7.04 ;
        RECT 78.48 4.7 78.65 7.765 ;
        RECT 77.49 4.7 77.66 7.765 ;
        RECT 74.75 4.7 74.92 7.76 ;
        RECT 73.385 5.43 83.28 5.965 ;
        RECT 73.055 4.495 73.385 5.805 ;
        RECT 71.315 5.095 71.575 5.805 ;
        RECT 70.755 5.635 71.125 6.185 ;
        RECT 70.315 4.715 70.645 4.955 ;
        RECT 70.315 4.715 70.505 5.085 ;
        RECT 69.885 4.985 70.495 5.805 ;
        RECT 69.935 4.985 70.205 6.585 ;
        RECT 69.015 5.095 69.235 5.805 ;
        RECT 68.775 5.635 69.055 6.475 ;
        RECT 68.005 4.765 68.335 4.955 ;
        RECT 67.585 5.135 68.205 5.805 ;
        RECT 68.005 4.765 68.205 5.805 ;
        RECT 67.775 5.135 68.105 6.525 ;
        RECT 66.665 5.125 66.925 5.805 ;
        RECT 56.93 5.43 66.695 7.03 ;
        RECT 62.87 5.425 66.445 7.03 ;
        RECT 63.525 5.425 63.695 7.76 ;
        RECT 56.93 5.43 62.87 7.04 ;
        RECT 61.895 4.7 62.065 7.765 ;
        RECT 60.905 4.7 61.075 7.765 ;
        RECT 58.165 4.7 58.335 7.76 ;
        RECT 56.8 5.43 66.695 5.965 ;
        RECT 56.47 4.495 56.8 5.805 ;
        RECT 54.73 5.095 54.99 5.805 ;
        RECT 54.17 5.635 54.54 6.185 ;
        RECT 53.73 4.715 54.06 4.955 ;
        RECT 53.73 4.715 53.92 5.085 ;
        RECT 53.3 4.985 53.91 5.805 ;
        RECT 53.35 4.985 53.62 6.585 ;
        RECT 52.43 5.095 52.65 5.805 ;
        RECT 52.19 5.635 52.47 6.475 ;
        RECT 51.42 4.765 51.75 4.955 ;
        RECT 51 5.135 51.62 5.805 ;
        RECT 51.42 4.765 51.62 5.805 ;
        RECT 51.19 5.135 51.52 6.525 ;
        RECT 50.08 5.125 50.34 5.805 ;
        RECT 40.345 5.43 50.11 7.03 ;
        RECT 46.285 5.425 49.86 7.03 ;
        RECT 46.94 5.425 47.11 7.76 ;
        RECT 40.345 5.43 46.285 7.04 ;
        RECT 45.31 4.7 45.48 7.765 ;
        RECT 44.32 4.7 44.49 7.765 ;
        RECT 41.58 4.7 41.75 7.76 ;
        RECT 40.215 5.43 50.11 5.965 ;
        RECT 39.885 4.495 40.215 5.805 ;
        RECT 38.145 5.095 38.405 5.805 ;
        RECT 37.585 5.635 37.955 6.185 ;
        RECT 37.145 4.715 37.475 4.955 ;
        RECT 37.145 4.715 37.335 5.085 ;
        RECT 36.715 4.985 37.325 5.805 ;
        RECT 36.765 4.985 37.035 6.585 ;
        RECT 35.845 5.095 36.065 5.805 ;
        RECT 35.605 5.635 35.885 6.475 ;
        RECT 34.835 4.765 35.165 4.955 ;
        RECT 34.415 5.135 35.035 5.805 ;
        RECT 34.835 4.765 35.035 5.805 ;
        RECT 34.605 5.135 34.935 6.525 ;
        RECT 33.495 5.125 33.755 5.805 ;
        RECT 23.76 5.43 33.525 7.03 ;
        RECT 29.7 5.425 33.275 7.03 ;
        RECT 30.355 5.425 30.525 7.76 ;
        RECT 23.76 5.43 29.7 7.04 ;
        RECT 28.725 4.7 28.895 7.765 ;
        RECT 27.735 4.7 27.905 7.765 ;
        RECT 24.995 4.7 25.165 7.76 ;
        RECT 23.63 5.43 33.525 5.965 ;
        RECT 23.3 4.495 23.63 5.805 ;
        RECT 21.56 5.095 21.82 5.805 ;
        RECT 21 5.635 21.37 6.185 ;
        RECT 20.56 4.715 20.89 4.955 ;
        RECT 20.56 4.715 20.75 5.085 ;
        RECT 20.13 4.985 20.74 5.805 ;
        RECT 20.18 4.985 20.45 6.585 ;
        RECT 19.26 5.095 19.48 5.805 ;
        RECT 19.02 5.635 19.3 6.475 ;
        RECT 18.25 4.765 18.58 4.955 ;
        RECT 17.83 5.135 18.45 5.805 ;
        RECT 18.25 4.765 18.45 5.805 ;
        RECT 18.02 5.135 18.35 6.525 ;
        RECT 16.91 5.125 17.17 5.805 ;
        RECT 10.155 5.425 16.915 7.025 ;
        RECT 10.155 5.425 16.345 7.03 ;
        RECT 13.77 5.425 13.94 7.76 ;
        RECT 12.35 5.425 12.52 10.59 ;
        RECT 10.54 5.425 10.71 7.76 ;
      LAYER met1 ;
        RECT 90.095 5.43 96.035 7.04 ;
        RECT 10.155 5.485 96.035 5.965 ;
        RECT 89.97 5.43 96.035 5.965 ;
        RECT 89.965 5.445 96.035 5.965 ;
        RECT 73.515 5.43 83.28 7.03 ;
        RECT 79.45 5.425 83.025 7.03 ;
        RECT 73.515 5.43 79.455 7.04 ;
        RECT 73.385 5.445 83.28 5.965 ;
        RECT 73.39 5.43 83.28 5.965 ;
        RECT 56.93 5.43 66.695 7.03 ;
        RECT 62.87 5.425 66.445 7.03 ;
        RECT 56.93 5.43 62.87 7.04 ;
        RECT 56.8 5.445 66.695 5.965 ;
        RECT 56.805 5.43 66.695 5.965 ;
        RECT 40.345 5.43 50.11 7.03 ;
        RECT 46.285 5.425 49.86 7.03 ;
        RECT 40.345 5.43 46.285 7.04 ;
        RECT 40.215 5.445 50.11 5.965 ;
        RECT 40.22 5.43 50.11 5.965 ;
        RECT 23.76 5.43 33.525 7.03 ;
        RECT 29.7 5.425 33.275 7.03 ;
        RECT 23.76 5.43 29.7 7.04 ;
        RECT 23.63 5.445 33.525 5.965 ;
        RECT 23.635 5.43 33.525 5.965 ;
        RECT 10.155 5.425 16.915 7.025 ;
        RECT 13.595 5.425 16.345 7.03 ;
        RECT 10.155 5.425 13.115 7.03 ;
        RECT 12.29 8.94 12.58 9.17 ;
        RECT 12.12 8.97 12.58 9.14 ;
      LAYER mcon ;
        RECT 12.35 8.97 12.52 9.14 ;
        RECT 12.66 6.83 12.83 7 ;
        RECT 15.89 6.83 16.06 7 ;
        RECT 16.97 5.635 17.14 5.805 ;
        RECT 17.43 5.635 17.6 5.805 ;
        RECT 17.89 5.635 18.06 5.805 ;
        RECT 18.35 5.635 18.52 5.805 ;
        RECT 18.81 5.635 18.98 5.805 ;
        RECT 19.27 5.635 19.44 5.805 ;
        RECT 19.73 5.635 19.9 5.805 ;
        RECT 20.19 5.635 20.36 5.805 ;
        RECT 20.65 5.635 20.82 5.805 ;
        RECT 21.11 5.635 21.28 5.805 ;
        RECT 21.57 5.635 21.74 5.805 ;
        RECT 22.03 5.635 22.2 5.805 ;
        RECT 22.49 5.635 22.66 5.805 ;
        RECT 22.95 5.635 23.12 5.805 ;
        RECT 23.41 5.635 23.58 5.805 ;
        RECT 27.115 6.83 27.285 7 ;
        RECT 27.115 5.46 27.285 5.63 ;
        RECT 27.815 6.835 27.985 7.005 ;
        RECT 27.815 5.46 27.985 5.63 ;
        RECT 28.805 6.835 28.975 7.005 ;
        RECT 28.805 5.46 28.975 5.63 ;
        RECT 32.475 6.83 32.645 7 ;
        RECT 33.555 5.635 33.725 5.805 ;
        RECT 34.015 5.635 34.185 5.805 ;
        RECT 34.475 5.635 34.645 5.805 ;
        RECT 34.935 5.635 35.105 5.805 ;
        RECT 35.395 5.635 35.565 5.805 ;
        RECT 35.855 5.635 36.025 5.805 ;
        RECT 36.315 5.635 36.485 5.805 ;
        RECT 36.775 5.635 36.945 5.805 ;
        RECT 37.235 5.635 37.405 5.805 ;
        RECT 37.695 5.635 37.865 5.805 ;
        RECT 38.155 5.635 38.325 5.805 ;
        RECT 38.615 5.635 38.785 5.805 ;
        RECT 39.075 5.635 39.245 5.805 ;
        RECT 39.535 5.635 39.705 5.805 ;
        RECT 39.995 5.635 40.165 5.805 ;
        RECT 43.7 6.83 43.87 7 ;
        RECT 43.7 5.46 43.87 5.63 ;
        RECT 44.4 6.835 44.57 7.005 ;
        RECT 44.4 5.46 44.57 5.63 ;
        RECT 45.39 6.835 45.56 7.005 ;
        RECT 45.39 5.46 45.56 5.63 ;
        RECT 49.06 6.83 49.23 7 ;
        RECT 50.14 5.635 50.31 5.805 ;
        RECT 50.6 5.635 50.77 5.805 ;
        RECT 51.06 5.635 51.23 5.805 ;
        RECT 51.52 5.635 51.69 5.805 ;
        RECT 51.98 5.635 52.15 5.805 ;
        RECT 52.44 5.635 52.61 5.805 ;
        RECT 52.9 5.635 53.07 5.805 ;
        RECT 53.36 5.635 53.53 5.805 ;
        RECT 53.82 5.635 53.99 5.805 ;
        RECT 54.28 5.635 54.45 5.805 ;
        RECT 54.74 5.635 54.91 5.805 ;
        RECT 55.2 5.635 55.37 5.805 ;
        RECT 55.66 5.635 55.83 5.805 ;
        RECT 56.12 5.635 56.29 5.805 ;
        RECT 56.58 5.635 56.75 5.805 ;
        RECT 60.285 6.83 60.455 7 ;
        RECT 60.285 5.46 60.455 5.63 ;
        RECT 60.985 6.835 61.155 7.005 ;
        RECT 60.985 5.46 61.155 5.63 ;
        RECT 61.975 6.835 62.145 7.005 ;
        RECT 61.975 5.46 62.145 5.63 ;
        RECT 65.645 6.83 65.815 7 ;
        RECT 66.725 5.635 66.895 5.805 ;
        RECT 67.185 5.635 67.355 5.805 ;
        RECT 67.645 5.635 67.815 5.805 ;
        RECT 68.105 5.635 68.275 5.805 ;
        RECT 68.565 5.635 68.735 5.805 ;
        RECT 69.025 5.635 69.195 5.805 ;
        RECT 69.485 5.635 69.655 5.805 ;
        RECT 69.945 5.635 70.115 5.805 ;
        RECT 70.405 5.635 70.575 5.805 ;
        RECT 70.865 5.635 71.035 5.805 ;
        RECT 71.325 5.635 71.495 5.805 ;
        RECT 71.785 5.635 71.955 5.805 ;
        RECT 72.245 5.635 72.415 5.805 ;
        RECT 72.705 5.635 72.875 5.805 ;
        RECT 73.165 5.635 73.335 5.805 ;
        RECT 76.87 6.83 77.04 7 ;
        RECT 76.87 5.46 77.04 5.63 ;
        RECT 77.57 6.835 77.74 7.005 ;
        RECT 77.57 5.46 77.74 5.63 ;
        RECT 78.56 6.835 78.73 7.005 ;
        RECT 78.56 5.46 78.73 5.63 ;
        RECT 82.225 6.83 82.395 7 ;
        RECT 83.305 5.635 83.475 5.805 ;
        RECT 83.765 5.635 83.935 5.805 ;
        RECT 84.225 5.635 84.395 5.805 ;
        RECT 84.685 5.635 84.855 5.805 ;
        RECT 85.145 5.635 85.315 5.805 ;
        RECT 85.605 5.635 85.775 5.805 ;
        RECT 86.065 5.635 86.235 5.805 ;
        RECT 86.525 5.635 86.695 5.805 ;
        RECT 86.985 5.635 87.155 5.805 ;
        RECT 87.445 5.635 87.615 5.805 ;
        RECT 87.905 5.635 88.075 5.805 ;
        RECT 88.365 5.635 88.535 5.805 ;
        RECT 88.825 5.635 88.995 5.805 ;
        RECT 89.285 5.635 89.455 5.805 ;
        RECT 89.745 5.635 89.915 5.805 ;
        RECT 93.45 6.83 93.62 7 ;
        RECT 93.45 5.46 93.62 5.63 ;
        RECT 94.15 6.835 94.32 7.005 ;
        RECT 94.15 5.46 94.32 5.63 ;
        RECT 95.14 6.835 95.31 7.005 ;
        RECT 95.14 5.46 95.31 5.63 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 85.535 7.765 85.865 8.095 ;
        RECT 85.505 7.785 85.805 8.195 ;
        RECT 85.065 7.785 85.865 8.085 ;
        RECT 68.955 7.765 69.285 8.095 ;
        RECT 68.925 7.785 69.225 8.195 ;
        RECT 68.485 7.785 69.285 8.085 ;
        RECT 52.37 7.765 52.7 8.095 ;
        RECT 52.34 7.785 52.64 8.195 ;
        RECT 51.9 7.785 52.7 8.085 ;
        RECT 35.785 7.765 36.115 8.095 ;
        RECT 35.755 7.785 36.055 8.195 ;
        RECT 35.315 7.785 36.115 8.085 ;
        RECT 19.2 7.765 19.53 8.095 ;
        RECT 19.17 7.785 19.47 8.195 ;
        RECT 18.73 7.785 19.53 8.085 ;
      LAYER li1 ;
        RECT 10.155 0 96.035 1.6 ;
        RECT 95.06 0 95.23 2.23 ;
        RECT 94.07 0 94.24 2.23 ;
        RECT 91.33 0 91.5 2.23 ;
        RECT 90.06 0 90.255 3.09 ;
        RECT 83.165 0 90.255 3.085 ;
        RECT 89.695 0 89.965 3.895 ;
        RECT 88.785 0 89.025 3.895 ;
        RECT 87.915 0 88.165 3.625 ;
        RECT 85.535 0 85.865 3.545 ;
        RECT 83.245 0 83.505 3.905 ;
        RECT 82.91 0 90.255 2.95 ;
        RECT 78.48 0 78.65 2.23 ;
        RECT 77.49 0 77.66 2.23 ;
        RECT 74.75 0 74.92 2.23 ;
        RECT 73.48 0 73.675 3.09 ;
        RECT 66.585 0 73.675 3.085 ;
        RECT 73.115 0 73.385 3.895 ;
        RECT 72.205 0 72.445 3.895 ;
        RECT 71.335 0 71.585 3.625 ;
        RECT 68.955 0 69.285 3.545 ;
        RECT 66.665 0 66.925 3.905 ;
        RECT 66.33 0 73.675 2.95 ;
        RECT 61.895 0 62.065 2.23 ;
        RECT 60.905 0 61.075 2.23 ;
        RECT 58.165 0 58.335 2.23 ;
        RECT 56.895 0 57.09 3.09 ;
        RECT 50 0 57.09 3.085 ;
        RECT 56.53 0 56.8 3.895 ;
        RECT 55.62 0 55.86 3.895 ;
        RECT 54.75 0 55 3.625 ;
        RECT 52.37 0 52.7 3.545 ;
        RECT 50.08 0 50.34 3.905 ;
        RECT 49.745 0 57.09 2.95 ;
        RECT 45.31 0 45.48 2.23 ;
        RECT 44.32 0 44.49 2.23 ;
        RECT 41.58 0 41.75 2.23 ;
        RECT 40.31 0 40.505 3.09 ;
        RECT 33.415 0 40.505 3.085 ;
        RECT 39.945 0 40.215 3.895 ;
        RECT 39.035 0 39.275 3.895 ;
        RECT 38.165 0 38.415 3.625 ;
        RECT 35.785 0 36.115 3.545 ;
        RECT 33.495 0 33.755 3.905 ;
        RECT 33.16 0 40.505 2.95 ;
        RECT 28.725 0 28.895 2.23 ;
        RECT 27.735 0 27.905 2.23 ;
        RECT 24.995 0 25.165 2.23 ;
        RECT 23.725 0 23.92 3.09 ;
        RECT 16.83 0 23.92 3.085 ;
        RECT 23.36 0 23.63 3.895 ;
        RECT 22.45 0 22.69 3.895 ;
        RECT 21.58 0 21.83 3.625 ;
        RECT 19.2 0 19.53 3.545 ;
        RECT 16.91 0 17.17 3.905 ;
        RECT 16.575 0 23.92 2.95 ;
        RECT 9.95 10.86 96.035 12.46 ;
        RECT 95.06 10.235 95.23 12.46 ;
        RECT 94.07 10.235 94.24 12.46 ;
        RECT 91.33 10.23 91.5 12.46 ;
        RECT 82.87 9.465 90.07 12.46 ;
        RECT 83.165 8.53 90.065 12.46 ;
        RECT 80.105 10.23 80.275 12.46 ;
        RECT 78.48 10.235 78.65 12.46 ;
        RECT 77.49 10.235 77.66 12.46 ;
        RECT 74.75 10.23 74.92 12.46 ;
        RECT 66.29 9.465 73.49 12.46 ;
        RECT 66.585 8.53 73.485 12.46 ;
        RECT 63.525 10.23 63.695 12.46 ;
        RECT 61.895 10.235 62.065 12.46 ;
        RECT 60.905 10.235 61.075 12.46 ;
        RECT 58.165 10.23 58.335 12.46 ;
        RECT 49.705 9.465 56.905 12.46 ;
        RECT 50 8.53 56.9 12.46 ;
        RECT 46.94 10.23 47.11 12.46 ;
        RECT 45.31 10.235 45.48 12.46 ;
        RECT 44.32 10.235 44.49 12.46 ;
        RECT 41.58 10.23 41.75 12.46 ;
        RECT 33.12 9.465 40.32 12.46 ;
        RECT 33.415 8.53 40.315 12.46 ;
        RECT 30.355 10.23 30.525 12.46 ;
        RECT 28.725 10.235 28.895 12.46 ;
        RECT 27.735 10.235 27.905 12.46 ;
        RECT 24.995 10.23 25.165 12.46 ;
        RECT 16.535 9.465 23.735 12.46 ;
        RECT 16.83 8.53 23.73 12.46 ;
        RECT 13.77 10.23 13.94 12.46 ;
        RECT 10.54 10.23 10.71 12.46 ;
        RECT 83.165 8.355 90.065 8.525 ;
        RECT 88.595 7.845 89.045 8.525 ;
        RECT 86.505 7.955 86.835 8.525 ;
        RECT 84.435 7.895 84.685 8.525 ;
        RECT 86.805 7.115 87.135 7.445 ;
        RECT 84.585 7.115 84.925 7.365 ;
        RECT 81.11 8.36 81.28 10.31 ;
        RECT 81.055 10.14 81.225 10.59 ;
        RECT 81.055 7.3 81.225 8.53 ;
        RECT 66.585 8.355 73.485 8.525 ;
        RECT 72.015 7.845 72.465 8.525 ;
        RECT 69.925 7.955 70.255 8.525 ;
        RECT 67.855 7.895 68.105 8.525 ;
        RECT 70.225 7.115 70.555 7.445 ;
        RECT 68.005 7.115 68.345 7.365 ;
        RECT 64.53 8.36 64.7 10.31 ;
        RECT 64.475 10.14 64.645 10.59 ;
        RECT 64.475 7.3 64.645 8.53 ;
        RECT 50 8.355 56.9 8.525 ;
        RECT 55.43 7.845 55.88 8.525 ;
        RECT 53.34 7.955 53.67 8.525 ;
        RECT 51.27 7.895 51.52 8.525 ;
        RECT 53.64 7.115 53.97 7.445 ;
        RECT 51.42 7.115 51.76 7.365 ;
        RECT 47.945 8.36 48.115 10.31 ;
        RECT 47.89 10.14 48.06 10.59 ;
        RECT 47.89 7.3 48.06 8.53 ;
        RECT 33.415 8.355 40.315 8.525 ;
        RECT 38.845 7.845 39.295 8.525 ;
        RECT 36.755 7.955 37.085 8.525 ;
        RECT 34.685 7.895 34.935 8.525 ;
        RECT 37.055 7.115 37.385 7.445 ;
        RECT 34.835 7.115 35.175 7.365 ;
        RECT 31.36 8.36 31.53 10.31 ;
        RECT 31.305 10.14 31.475 10.59 ;
        RECT 31.305 7.3 31.475 8.53 ;
        RECT 16.83 8.355 23.73 8.525 ;
        RECT 22.26 7.845 22.71 8.525 ;
        RECT 20.17 7.955 20.5 8.525 ;
        RECT 18.1 7.895 18.35 8.525 ;
        RECT 20.47 7.115 20.8 7.445 ;
        RECT 18.25 7.115 18.59 7.365 ;
        RECT 14.775 8.36 14.945 10.31 ;
        RECT 14.72 10.14 14.89 10.59 ;
        RECT 14.72 7.3 14.89 8.53 ;
      LAYER met2 ;
        RECT 85.565 7.745 85.845 8.115 ;
        RECT 68.985 7.745 69.265 8.115 ;
        RECT 52.4 7.745 52.68 8.115 ;
        RECT 35.815 7.745 36.095 8.115 ;
        RECT 19.23 7.745 19.51 8.115 ;
      LAYER met1 ;
        RECT 10.155 0 96.035 1.6 ;
        RECT 83.165 0 90.255 3.09 ;
        RECT 83.165 0 90.065 3.245 ;
        RECT 82.91 0 90.255 2.95 ;
        RECT 66.585 0 73.675 3.09 ;
        RECT 66.585 0 73.485 3.245 ;
        RECT 66.33 0 73.675 2.95 ;
        RECT 50 0 57.09 3.09 ;
        RECT 50 0 56.9 3.245 ;
        RECT 49.745 0 57.09 2.95 ;
        RECT 33.415 0 40.505 3.09 ;
        RECT 33.415 0 40.315 3.245 ;
        RECT 33.16 0 40.505 2.95 ;
        RECT 16.83 0 23.92 3.09 ;
        RECT 16.83 0 23.73 3.245 ;
        RECT 16.575 0 23.92 2.95 ;
        RECT 9.95 10.86 96.035 12.46 ;
        RECT 82.87 9.465 90.07 12.46 ;
        RECT 83.165 8.205 90.065 12.46 ;
        RECT 86.755 7.135 87.045 7.365 ;
        RECT 84.625 7.805 86.975 7.945 ;
        RECT 86.835 7.135 86.975 7.945 ;
        RECT 85.555 7.805 85.875 8.065 ;
        RECT 85.59 7.805 85.845 12.46 ;
        RECT 84.545 7.135 84.835 7.365 ;
        RECT 84.625 7.135 84.765 7.945 ;
        RECT 81.05 8.57 81.34 8.8 ;
        RECT 80.89 10.85 81.065 12.46 ;
        RECT 80.89 8.6 81.06 12.46 ;
        RECT 80.88 8.6 81.34 8.77 ;
        RECT 66.29 9.465 73.49 12.46 ;
        RECT 66.585 8.205 73.485 12.46 ;
        RECT 70.175 7.135 70.465 7.365 ;
        RECT 68.045 7.805 70.395 7.945 ;
        RECT 70.255 7.135 70.395 7.945 ;
        RECT 68.975 7.805 69.295 8.065 ;
        RECT 69.01 7.805 69.265 12.46 ;
        RECT 67.965 7.135 68.255 7.365 ;
        RECT 68.045 7.135 68.185 7.945 ;
        RECT 64.47 8.57 64.76 8.8 ;
        RECT 64.31 10.85 64.485 12.46 ;
        RECT 64.31 8.6 64.48 12.46 ;
        RECT 64.3 8.6 64.76 8.77 ;
        RECT 49.705 9.465 56.905 12.46 ;
        RECT 50 8.205 56.9 12.46 ;
        RECT 53.59 7.135 53.88 7.365 ;
        RECT 51.46 7.805 53.81 7.945 ;
        RECT 53.67 7.135 53.81 7.945 ;
        RECT 52.39 7.805 52.71 8.065 ;
        RECT 52.425 7.805 52.68 12.46 ;
        RECT 51.38 7.135 51.67 7.365 ;
        RECT 51.46 7.135 51.6 7.945 ;
        RECT 47.885 8.57 48.175 8.8 ;
        RECT 47.725 10.85 47.9 12.46 ;
        RECT 47.725 8.6 47.895 12.46 ;
        RECT 47.715 8.6 48.175 8.77 ;
        RECT 33.12 9.465 40.32 12.46 ;
        RECT 33.415 8.205 40.315 12.46 ;
        RECT 37.005 7.135 37.295 7.365 ;
        RECT 34.875 7.805 37.225 7.945 ;
        RECT 37.085 7.135 37.225 7.945 ;
        RECT 35.805 7.805 36.125 8.065 ;
        RECT 35.84 7.805 36.095 12.46 ;
        RECT 34.795 7.135 35.085 7.365 ;
        RECT 34.875 7.135 35.015 7.945 ;
        RECT 31.3 8.57 31.59 8.8 ;
        RECT 31.14 10.85 31.315 12.46 ;
        RECT 31.14 8.6 31.31 12.46 ;
        RECT 31.13 8.6 31.59 8.77 ;
        RECT 16.535 9.465 23.735 12.46 ;
        RECT 16.83 8.205 23.73 12.46 ;
        RECT 20.42 7.135 20.71 7.365 ;
        RECT 18.29 7.805 20.64 7.945 ;
        RECT 20.5 7.135 20.64 7.945 ;
        RECT 19.22 7.805 19.54 8.065 ;
        RECT 19.255 7.805 19.51 12.46 ;
        RECT 18.21 7.135 18.5 7.365 ;
        RECT 18.29 7.135 18.43 7.945 ;
        RECT 14.715 8.57 15.005 8.8 ;
        RECT 14.555 10.85 14.73 12.46 ;
        RECT 14.555 8.6 14.725 12.46 ;
        RECT 14.545 8.6 15.005 8.77 ;
      LAYER via2 ;
        RECT 19.27 7.835 19.47 8.035 ;
        RECT 35.855 7.835 36.055 8.035 ;
        RECT 52.44 7.835 52.64 8.035 ;
        RECT 69.025 7.835 69.225 8.035 ;
        RECT 85.605 7.835 85.805 8.035 ;
      LAYER via1 ;
        RECT 19.305 7.86 19.455 8.01 ;
        RECT 35.89 7.86 36.04 8.01 ;
        RECT 52.475 7.86 52.625 8.01 ;
        RECT 69.06 7.86 69.21 8.01 ;
        RECT 85.64 7.86 85.79 8.01 ;
      LAYER mcon ;
        RECT 10.62 10.89 10.79 11.06 ;
        RECT 11.3 10.89 11.47 11.06 ;
        RECT 11.98 10.89 12.15 11.06 ;
        RECT 12.66 10.89 12.83 11.06 ;
        RECT 13.85 10.89 14.02 11.06 ;
        RECT 14.53 10.89 14.7 11.06 ;
        RECT 14.775 8.6 14.945 8.77 ;
        RECT 15.21 10.89 15.38 11.06 ;
        RECT 15.89 10.89 16.06 11.06 ;
        RECT 16.97 8.355 17.14 8.525 ;
        RECT 17.43 8.355 17.6 8.525 ;
        RECT 17.89 8.355 18.06 8.525 ;
        RECT 18.27 7.165 18.44 7.335 ;
        RECT 18.35 8.355 18.52 8.525 ;
        RECT 18.81 8.355 18.98 8.525 ;
        RECT 19.27 8.355 19.44 8.525 ;
        RECT 19.73 8.355 19.9 8.525 ;
        RECT 20.19 8.355 20.36 8.525 ;
        RECT 20.48 7.165 20.65 7.335 ;
        RECT 20.65 8.355 20.82 8.525 ;
        RECT 21.11 8.355 21.28 8.525 ;
        RECT 21.57 8.355 21.74 8.525 ;
        RECT 22.03 8.355 22.2 8.525 ;
        RECT 22.49 8.355 22.66 8.525 ;
        RECT 22.95 8.355 23.12 8.525 ;
        RECT 23.41 8.355 23.58 8.525 ;
        RECT 25.075 10.89 25.245 11.06 ;
        RECT 25.075 1.4 25.245 1.57 ;
        RECT 25.755 10.89 25.925 11.06 ;
        RECT 25.755 1.4 25.925 1.57 ;
        RECT 26.435 10.89 26.605 11.06 ;
        RECT 26.435 1.4 26.605 1.57 ;
        RECT 27.115 10.89 27.285 11.06 ;
        RECT 27.115 1.4 27.285 1.57 ;
        RECT 27.815 10.895 27.985 11.065 ;
        RECT 27.815 1.4 27.985 1.57 ;
        RECT 28.805 10.895 28.975 11.065 ;
        RECT 28.805 1.4 28.975 1.57 ;
        RECT 30.435 10.89 30.605 11.06 ;
        RECT 31.115 10.89 31.285 11.06 ;
        RECT 31.36 8.6 31.53 8.77 ;
        RECT 31.795 10.89 31.965 11.06 ;
        RECT 32.475 10.89 32.645 11.06 ;
        RECT 33.555 8.355 33.725 8.525 ;
        RECT 34.015 8.355 34.185 8.525 ;
        RECT 34.475 8.355 34.645 8.525 ;
        RECT 34.855 7.165 35.025 7.335 ;
        RECT 34.935 8.355 35.105 8.525 ;
        RECT 35.395 8.355 35.565 8.525 ;
        RECT 35.855 8.355 36.025 8.525 ;
        RECT 36.315 8.355 36.485 8.525 ;
        RECT 36.775 8.355 36.945 8.525 ;
        RECT 37.065 7.165 37.235 7.335 ;
        RECT 37.235 8.355 37.405 8.525 ;
        RECT 37.695 8.355 37.865 8.525 ;
        RECT 38.155 8.355 38.325 8.525 ;
        RECT 38.615 8.355 38.785 8.525 ;
        RECT 39.075 8.355 39.245 8.525 ;
        RECT 39.535 8.355 39.705 8.525 ;
        RECT 39.995 8.355 40.165 8.525 ;
        RECT 41.66 10.89 41.83 11.06 ;
        RECT 41.66 1.4 41.83 1.57 ;
        RECT 42.34 10.89 42.51 11.06 ;
        RECT 42.34 1.4 42.51 1.57 ;
        RECT 43.02 10.89 43.19 11.06 ;
        RECT 43.02 1.4 43.19 1.57 ;
        RECT 43.7 10.89 43.87 11.06 ;
        RECT 43.7 1.4 43.87 1.57 ;
        RECT 44.4 10.895 44.57 11.065 ;
        RECT 44.4 1.4 44.57 1.57 ;
        RECT 45.39 10.895 45.56 11.065 ;
        RECT 45.39 1.4 45.56 1.57 ;
        RECT 47.02 10.89 47.19 11.06 ;
        RECT 47.7 10.89 47.87 11.06 ;
        RECT 47.945 8.6 48.115 8.77 ;
        RECT 48.38 10.89 48.55 11.06 ;
        RECT 49.06 10.89 49.23 11.06 ;
        RECT 50.14 8.355 50.31 8.525 ;
        RECT 50.6 8.355 50.77 8.525 ;
        RECT 51.06 8.355 51.23 8.525 ;
        RECT 51.44 7.165 51.61 7.335 ;
        RECT 51.52 8.355 51.69 8.525 ;
        RECT 51.98 8.355 52.15 8.525 ;
        RECT 52.44 8.355 52.61 8.525 ;
        RECT 52.9 8.355 53.07 8.525 ;
        RECT 53.36 8.355 53.53 8.525 ;
        RECT 53.65 7.165 53.82 7.335 ;
        RECT 53.82 8.355 53.99 8.525 ;
        RECT 54.28 8.355 54.45 8.525 ;
        RECT 54.74 8.355 54.91 8.525 ;
        RECT 55.2 8.355 55.37 8.525 ;
        RECT 55.66 8.355 55.83 8.525 ;
        RECT 56.12 8.355 56.29 8.525 ;
        RECT 56.58 8.355 56.75 8.525 ;
        RECT 58.245 10.89 58.415 11.06 ;
        RECT 58.245 1.4 58.415 1.57 ;
        RECT 58.925 10.89 59.095 11.06 ;
        RECT 58.925 1.4 59.095 1.57 ;
        RECT 59.605 10.89 59.775 11.06 ;
        RECT 59.605 1.4 59.775 1.57 ;
        RECT 60.285 10.89 60.455 11.06 ;
        RECT 60.285 1.4 60.455 1.57 ;
        RECT 60.985 10.895 61.155 11.065 ;
        RECT 60.985 1.4 61.155 1.57 ;
        RECT 61.975 10.895 62.145 11.065 ;
        RECT 61.975 1.4 62.145 1.57 ;
        RECT 63.605 10.89 63.775 11.06 ;
        RECT 64.285 10.89 64.455 11.06 ;
        RECT 64.53 8.6 64.7 8.77 ;
        RECT 64.965 10.89 65.135 11.06 ;
        RECT 65.645 10.89 65.815 11.06 ;
        RECT 66.725 8.355 66.895 8.525 ;
        RECT 67.185 8.355 67.355 8.525 ;
        RECT 67.645 8.355 67.815 8.525 ;
        RECT 68.025 7.165 68.195 7.335 ;
        RECT 68.105 8.355 68.275 8.525 ;
        RECT 68.565 8.355 68.735 8.525 ;
        RECT 69.025 8.355 69.195 8.525 ;
        RECT 69.485 8.355 69.655 8.525 ;
        RECT 69.945 8.355 70.115 8.525 ;
        RECT 70.235 7.165 70.405 7.335 ;
        RECT 70.405 8.355 70.575 8.525 ;
        RECT 70.865 8.355 71.035 8.525 ;
        RECT 71.325 8.355 71.495 8.525 ;
        RECT 71.785 8.355 71.955 8.525 ;
        RECT 72.245 8.355 72.415 8.525 ;
        RECT 72.705 8.355 72.875 8.525 ;
        RECT 73.165 8.355 73.335 8.525 ;
        RECT 74.83 10.89 75 11.06 ;
        RECT 74.83 1.4 75 1.57 ;
        RECT 75.51 10.89 75.68 11.06 ;
        RECT 75.51 1.4 75.68 1.57 ;
        RECT 76.19 10.89 76.36 11.06 ;
        RECT 76.19 1.4 76.36 1.57 ;
        RECT 76.87 10.89 77.04 11.06 ;
        RECT 76.87 1.4 77.04 1.57 ;
        RECT 77.57 10.895 77.74 11.065 ;
        RECT 77.57 1.4 77.74 1.57 ;
        RECT 78.56 10.895 78.73 11.065 ;
        RECT 78.56 1.4 78.73 1.57 ;
        RECT 80.185 10.89 80.355 11.06 ;
        RECT 80.865 10.89 81.035 11.06 ;
        RECT 81.11 8.6 81.28 8.77 ;
        RECT 81.545 10.89 81.715 11.06 ;
        RECT 82.225 10.89 82.395 11.06 ;
        RECT 83.305 8.355 83.475 8.525 ;
        RECT 83.765 8.355 83.935 8.525 ;
        RECT 84.225 8.355 84.395 8.525 ;
        RECT 84.605 7.165 84.775 7.335 ;
        RECT 84.685 8.355 84.855 8.525 ;
        RECT 85.145 8.355 85.315 8.525 ;
        RECT 85.605 8.355 85.775 8.525 ;
        RECT 86.065 8.355 86.235 8.525 ;
        RECT 86.525 8.355 86.695 8.525 ;
        RECT 86.815 7.165 86.985 7.335 ;
        RECT 86.985 8.355 87.155 8.525 ;
        RECT 87.445 8.355 87.615 8.525 ;
        RECT 87.905 8.355 88.075 8.525 ;
        RECT 88.365 8.355 88.535 8.525 ;
        RECT 88.825 8.355 88.995 8.525 ;
        RECT 89.285 8.355 89.455 8.525 ;
        RECT 89.745 8.355 89.915 8.525 ;
        RECT 91.41 10.89 91.58 11.06 ;
        RECT 91.41 1.4 91.58 1.57 ;
        RECT 92.09 10.89 92.26 11.06 ;
        RECT 92.09 1.4 92.26 1.57 ;
        RECT 92.77 10.89 92.94 11.06 ;
        RECT 92.77 1.4 92.94 1.57 ;
        RECT 93.45 10.89 93.62 11.06 ;
        RECT 93.45 1.4 93.62 1.57 ;
        RECT 94.15 10.895 94.32 11.065 ;
        RECT 94.15 1.4 94.32 1.57 ;
        RECT 95.14 10.895 95.31 11.065 ;
        RECT 95.14 1.4 95.31 1.57 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 87.96 4.025 88.26 4.36 ;
      RECT 87.935 4.025 88.265 4.355 ;
      RECT 87.935 4.045 88.735 4.345 ;
      RECT 81.385 9.28 81.755 9.65 ;
      RECT 81.385 9.315 86.54 9.615 ;
      RECT 86.235 7.085 86.535 9.615 ;
      RECT 85.61 7.09 86.545 7.42 ;
      RECT 86.215 7.085 86.545 7.42 ;
      RECT 87.255 7.085 87.585 7.415 ;
      RECT 85.61 7.105 88.055 7.405 ;
      RECT 85.61 7.09 87.585 7.405 ;
      RECT 85.61 5.06 85.94 7.42 ;
      RECT 85.61 5.06 87.905 5.39 ;
      RECT 85.61 5.06 88.26 5.38 ;
      RECT 87.935 5.045 88.265 5.375 ;
      RECT 85.61 5.065 88.735 5.365 ;
      RECT 87.945 4.995 88.245 5.38 ;
      RECT 87.235 4.365 87.565 4.695 ;
      RECT 87.265 4.355 87.565 4.695 ;
      RECT 86.765 4.385 87.565 4.685 ;
      RECT 86.58 6.065 86.615 6.4 ;
      RECT 86.575 6.065 86.905 6.395 ;
      RECT 86.575 6.085 87.375 6.385 ;
      RECT 86.575 6.08 86.91 6.385 ;
      RECT 85.895 3.685 86.225 4.015 ;
      RECT 85.425 3.705 85.785 4.005 ;
      RECT 85.785 3.695 86.225 3.995 ;
      RECT 71.38 4.025 71.68 4.36 ;
      RECT 71.355 4.025 71.685 4.355 ;
      RECT 71.355 4.045 72.155 4.345 ;
      RECT 64.805 9.28 65.175 9.65 ;
      RECT 64.805 9.315 69.96 9.615 ;
      RECT 69.655 7.085 69.955 9.615 ;
      RECT 69.03 7.09 69.965 7.42 ;
      RECT 69.635 7.085 69.965 7.42 ;
      RECT 70.675 7.085 71.005 7.415 ;
      RECT 69.03 7.105 71.475 7.405 ;
      RECT 69.03 7.09 71.005 7.405 ;
      RECT 69.03 5.06 69.36 7.42 ;
      RECT 69.03 5.06 71.325 5.39 ;
      RECT 69.03 5.06 71.68 5.38 ;
      RECT 71.355 5.045 71.685 5.375 ;
      RECT 69.03 5.065 72.155 5.365 ;
      RECT 71.365 4.995 71.665 5.38 ;
      RECT 70.655 4.365 70.985 4.695 ;
      RECT 70.685 4.355 70.985 4.695 ;
      RECT 70.185 4.385 70.985 4.685 ;
      RECT 70 6.065 70.035 6.4 ;
      RECT 69.995 6.065 70.325 6.395 ;
      RECT 69.995 6.085 70.795 6.385 ;
      RECT 69.995 6.08 70.33 6.385 ;
      RECT 69.315 3.685 69.645 4.015 ;
      RECT 68.845 3.705 69.205 4.005 ;
      RECT 69.205 3.695 69.645 3.995 ;
      RECT 54.795 4.025 55.095 4.36 ;
      RECT 54.77 4.025 55.1 4.355 ;
      RECT 54.77 4.045 55.57 4.345 ;
      RECT 48.22 9.28 48.59 9.65 ;
      RECT 48.22 9.315 53.375 9.615 ;
      RECT 53.07 7.085 53.37 9.615 ;
      RECT 52.445 7.09 53.38 7.42 ;
      RECT 53.05 7.085 53.38 7.42 ;
      RECT 54.09 7.085 54.42 7.415 ;
      RECT 52.445 7.105 54.89 7.405 ;
      RECT 52.445 7.09 54.42 7.405 ;
      RECT 52.445 5.06 52.775 7.42 ;
      RECT 52.445 5.06 54.74 5.39 ;
      RECT 52.445 5.06 55.095 5.38 ;
      RECT 54.77 5.045 55.1 5.375 ;
      RECT 52.445 5.065 55.57 5.365 ;
      RECT 54.78 4.995 55.08 5.38 ;
      RECT 54.07 4.365 54.4 4.695 ;
      RECT 54.1 4.355 54.4 4.695 ;
      RECT 53.6 4.385 54.4 4.685 ;
      RECT 53.415 6.065 53.45 6.4 ;
      RECT 53.41 6.065 53.74 6.395 ;
      RECT 53.41 6.085 54.21 6.385 ;
      RECT 53.41 6.08 53.745 6.385 ;
      RECT 52.73 3.685 53.06 4.015 ;
      RECT 52.26 3.705 52.62 4.005 ;
      RECT 52.62 3.695 53.06 3.995 ;
      RECT 38.21 4.025 38.51 4.36 ;
      RECT 38.185 4.025 38.515 4.355 ;
      RECT 38.185 4.045 38.985 4.345 ;
      RECT 31.635 9.28 32.005 9.65 ;
      RECT 31.635 9.315 36.79 9.615 ;
      RECT 36.485 7.085 36.785 9.615 ;
      RECT 35.86 7.09 36.795 7.42 ;
      RECT 36.465 7.085 36.795 7.42 ;
      RECT 37.505 7.085 37.835 7.415 ;
      RECT 35.86 7.105 38.305 7.405 ;
      RECT 35.86 7.09 37.835 7.405 ;
      RECT 35.86 5.06 36.19 7.42 ;
      RECT 35.86 5.06 38.155 5.39 ;
      RECT 35.86 5.06 38.51 5.38 ;
      RECT 38.185 5.045 38.515 5.375 ;
      RECT 35.86 5.065 38.985 5.365 ;
      RECT 38.195 4.995 38.495 5.38 ;
      RECT 37.485 4.365 37.815 4.695 ;
      RECT 37.515 4.355 37.815 4.695 ;
      RECT 37.015 4.385 37.815 4.685 ;
      RECT 36.83 6.065 36.865 6.4 ;
      RECT 36.825 6.065 37.155 6.395 ;
      RECT 36.825 6.085 37.625 6.385 ;
      RECT 36.825 6.08 37.16 6.385 ;
      RECT 36.145 3.685 36.475 4.015 ;
      RECT 35.675 3.705 36.035 4.005 ;
      RECT 36.035 3.695 36.475 3.995 ;
      RECT 21.625 4.025 21.925 4.36 ;
      RECT 21.6 4.025 21.93 4.355 ;
      RECT 21.6 4.045 22.4 4.345 ;
      RECT 15.05 9.28 15.42 9.65 ;
      RECT 15.05 9.315 20.205 9.615 ;
      RECT 19.9 7.085 20.2 9.615 ;
      RECT 19.275 7.09 20.21 7.42 ;
      RECT 19.88 7.085 20.21 7.42 ;
      RECT 20.92 7.085 21.25 7.415 ;
      RECT 19.275 7.105 21.72 7.405 ;
      RECT 19.275 7.09 21.25 7.405 ;
      RECT 19.275 5.06 19.605 7.42 ;
      RECT 19.275 5.06 21.57 5.39 ;
      RECT 19.275 5.06 21.925 5.38 ;
      RECT 21.6 5.045 21.93 5.375 ;
      RECT 19.275 5.065 22.4 5.365 ;
      RECT 21.61 4.995 21.91 5.38 ;
      RECT 20.9 4.365 21.23 4.695 ;
      RECT 20.93 4.355 21.23 4.695 ;
      RECT 20.43 4.385 21.23 4.685 ;
      RECT 20.245 6.065 20.28 6.4 ;
      RECT 20.24 6.065 20.57 6.395 ;
      RECT 20.24 6.085 21.04 6.385 ;
      RECT 20.24 6.08 20.575 6.385 ;
      RECT 19.56 3.685 19.89 4.015 ;
      RECT 19.09 3.705 19.45 4.005 ;
      RECT 19.45 3.695 19.89 3.995 ;
    LAYER via2 ;
      RECT 88.005 4.095 88.205 4.295 ;
      RECT 88.005 5.115 88.205 5.315 ;
      RECT 87.325 7.155 87.525 7.355 ;
      RECT 87.305 4.435 87.505 4.635 ;
      RECT 86.645 6.135 86.845 6.335 ;
      RECT 86.275 7.155 86.475 7.355 ;
      RECT 85.965 3.745 86.165 3.945 ;
      RECT 81.47 9.365 81.67 9.565 ;
      RECT 71.425 4.095 71.625 4.295 ;
      RECT 71.425 5.115 71.625 5.315 ;
      RECT 70.745 7.155 70.945 7.355 ;
      RECT 70.725 4.435 70.925 4.635 ;
      RECT 70.065 6.135 70.265 6.335 ;
      RECT 69.695 7.155 69.895 7.355 ;
      RECT 69.385 3.745 69.585 3.945 ;
      RECT 64.89 9.365 65.09 9.565 ;
      RECT 54.84 4.095 55.04 4.295 ;
      RECT 54.84 5.115 55.04 5.315 ;
      RECT 54.16 7.155 54.36 7.355 ;
      RECT 54.14 4.435 54.34 4.635 ;
      RECT 53.48 6.135 53.68 6.335 ;
      RECT 53.11 7.155 53.31 7.355 ;
      RECT 52.8 3.745 53 3.945 ;
      RECT 48.305 9.365 48.505 9.565 ;
      RECT 38.255 4.095 38.455 4.295 ;
      RECT 38.255 5.115 38.455 5.315 ;
      RECT 37.575 7.155 37.775 7.355 ;
      RECT 37.555 4.435 37.755 4.635 ;
      RECT 36.895 6.135 37.095 6.335 ;
      RECT 36.525 7.155 36.725 7.355 ;
      RECT 36.215 3.745 36.415 3.945 ;
      RECT 31.72 9.365 31.92 9.565 ;
      RECT 21.67 4.095 21.87 4.295 ;
      RECT 21.67 5.115 21.87 5.315 ;
      RECT 20.99 7.155 21.19 7.355 ;
      RECT 20.97 4.435 21.17 4.635 ;
      RECT 20.31 6.135 20.51 6.335 ;
      RECT 19.94 7.155 20.14 7.355 ;
      RECT 19.63 3.745 19.83 3.945 ;
      RECT 15.135 9.365 15.335 9.565 ;
    LAYER met2 ;
      RECT 11.525 10.065 95.665 10.235 ;
      RECT 95.495 9.585 95.665 10.235 ;
      RECT 11.525 8.54 11.695 10.235 ;
      RECT 95.46 9.585 95.785 9.91 ;
      RECT 11.485 8.54 11.765 8.88 ;
      RECT 92.305 8.565 92.625 8.89 ;
      RECT 92.335 7.98 92.505 8.89 ;
      RECT 92.335 7.98 92.51 8.33 ;
      RECT 92.335 7.98 93.31 8.155 ;
      RECT 93.135 3.26 93.31 8.155 ;
      RECT 93.08 3.26 93.43 3.61 ;
      RECT 81.97 9.705 92.15 9.875 ;
      RECT 91.99 3.69 92.15 9.875 ;
      RECT 81.97 8.885 82.14 9.875 ;
      RECT 93.105 8.94 93.43 9.265 ;
      RECT 78.915 8.94 79.24 9.265 ;
      RECT 81.915 8.885 82.195 9.225 ;
      RECT 91.99 9.03 93.43 9.2 ;
      RECT 78.915 8.97 82.195 9.14 ;
      RECT 92.305 3.66 92.625 3.98 ;
      RECT 91.99 3.69 92.625 3.86 ;
      RECT 85.925 3.665 86.205 4.035 ;
      RECT 85.97 2.9 86.14 4.035 ;
      RECT 90.635 3.29 90.96 3.615 ;
      RECT 90.71 2.9 90.88 3.615 ;
      RECT 85.97 2.9 90.88 3.07 ;
      RECT 89.665 6.075 89.925 6.395 ;
      RECT 89.725 4.035 89.865 6.395 ;
      RECT 89.665 4.035 89.925 4.355 ;
      RECT 88.645 7.095 88.905 7.415 ;
      RECT 88.025 7.185 88.905 7.325 ;
      RECT 88.025 5.025 88.165 7.325 ;
      RECT 87.965 5.025 88.245 5.395 ;
      RECT 87.285 7.065 87.565 7.435 ;
      RECT 87.345 5.145 87.485 7.435 ;
      RECT 87.345 5.145 87.825 5.285 ;
      RECT 87.685 3.355 87.825 5.285 ;
      RECT 87.625 3.355 87.885 3.675 ;
      RECT 86.605 6.045 86.885 6.415 ;
      RECT 86.665 3.695 86.805 6.415 ;
      RECT 86.605 3.695 86.865 4.015 ;
      RECT 86.235 7.065 86.515 7.435 ;
      RECT 86.235 7.095 86.525 7.415 ;
      RECT 81.385 9.28 81.755 9.65 ;
      RECT 81.385 9.28 81.76 9.29 ;
      RECT 75.725 8.565 76.045 8.89 ;
      RECT 75.755 7.98 75.925 8.89 ;
      RECT 75.755 7.98 75.93 8.33 ;
      RECT 75.755 7.98 76.73 8.155 ;
      RECT 76.555 3.26 76.73 8.155 ;
      RECT 76.5 3.26 76.85 3.61 ;
      RECT 65.39 9.705 75.57 9.875 ;
      RECT 75.41 3.69 75.57 9.875 ;
      RECT 65.39 8.885 65.56 9.875 ;
      RECT 76.525 8.94 76.85 9.265 ;
      RECT 62.33 8.94 62.655 9.265 ;
      RECT 65.335 8.885 65.615 9.225 ;
      RECT 75.41 9.03 76.85 9.2 ;
      RECT 62.33 8.97 65.615 9.14 ;
      RECT 75.725 3.66 76.045 3.98 ;
      RECT 75.41 3.69 76.045 3.86 ;
      RECT 69.345 3.665 69.625 4.035 ;
      RECT 69.39 2.9 69.56 4.035 ;
      RECT 74.055 3.29 74.38 3.615 ;
      RECT 74.13 2.9 74.3 3.615 ;
      RECT 69.39 2.9 74.3 3.07 ;
      RECT 73.085 6.075 73.345 6.395 ;
      RECT 73.145 4.035 73.285 6.395 ;
      RECT 73.085 4.035 73.345 4.355 ;
      RECT 72.065 7.095 72.325 7.415 ;
      RECT 71.445 7.185 72.325 7.325 ;
      RECT 71.445 5.025 71.585 7.325 ;
      RECT 71.385 5.025 71.665 5.395 ;
      RECT 70.705 7.065 70.985 7.435 ;
      RECT 70.765 5.145 70.905 7.435 ;
      RECT 70.765 5.145 71.245 5.285 ;
      RECT 71.105 3.355 71.245 5.285 ;
      RECT 71.045 3.355 71.305 3.675 ;
      RECT 70.025 6.045 70.305 6.415 ;
      RECT 70.085 3.695 70.225 6.415 ;
      RECT 70.025 3.695 70.285 4.015 ;
      RECT 69.655 7.065 69.935 7.435 ;
      RECT 69.655 7.095 69.945 7.415 ;
      RECT 59.14 8.565 59.46 8.89 ;
      RECT 59.17 7.98 59.34 8.89 ;
      RECT 59.17 7.98 59.345 8.33 ;
      RECT 59.17 7.98 60.145 8.155 ;
      RECT 59.97 3.26 60.145 8.155 ;
      RECT 59.915 3.26 60.265 3.61 ;
      RECT 48.805 9.705 58.985 9.875 ;
      RECT 58.825 3.69 58.985 9.875 ;
      RECT 48.805 8.885 48.975 9.875 ;
      RECT 59.94 8.94 60.265 9.265 ;
      RECT 45.745 8.94 46.07 9.265 ;
      RECT 48.75 8.885 49.03 9.225 ;
      RECT 58.825 9.03 60.265 9.2 ;
      RECT 45.745 8.97 49.03 9.14 ;
      RECT 59.14 3.66 59.46 3.98 ;
      RECT 58.825 3.69 59.46 3.86 ;
      RECT 52.76 3.665 53.04 4.035 ;
      RECT 52.805 2.9 52.975 4.035 ;
      RECT 57.47 3.29 57.795 3.615 ;
      RECT 57.545 2.9 57.715 3.615 ;
      RECT 52.805 2.9 57.715 3.07 ;
      RECT 56.5 6.075 56.76 6.395 ;
      RECT 56.56 4.035 56.7 6.395 ;
      RECT 56.5 4.035 56.76 4.355 ;
      RECT 55.48 7.095 55.74 7.415 ;
      RECT 54.86 7.185 55.74 7.325 ;
      RECT 54.86 5.025 55 7.325 ;
      RECT 54.8 5.025 55.08 5.395 ;
      RECT 54.12 7.065 54.4 7.435 ;
      RECT 54.18 5.145 54.32 7.435 ;
      RECT 54.18 5.145 54.66 5.285 ;
      RECT 54.52 3.355 54.66 5.285 ;
      RECT 54.46 3.355 54.72 3.675 ;
      RECT 53.44 6.045 53.72 6.415 ;
      RECT 53.5 3.695 53.64 6.415 ;
      RECT 53.44 3.695 53.7 4.015 ;
      RECT 53.07 7.065 53.35 7.435 ;
      RECT 53.07 7.095 53.36 7.415 ;
      RECT 42.555 8.565 42.875 8.89 ;
      RECT 42.585 7.98 42.755 8.89 ;
      RECT 42.585 7.98 42.76 8.33 ;
      RECT 42.585 7.98 43.56 8.155 ;
      RECT 43.385 3.26 43.56 8.155 ;
      RECT 43.33 3.26 43.68 3.61 ;
      RECT 32.22 9.705 42.4 9.875 ;
      RECT 42.24 3.69 42.4 9.875 ;
      RECT 32.22 8.885 32.39 9.875 ;
      RECT 43.355 8.94 43.68 9.265 ;
      RECT 29.16 8.94 29.485 9.265 ;
      RECT 32.165 8.885 32.445 9.225 ;
      RECT 42.24 9.03 43.68 9.2 ;
      RECT 29.16 8.97 32.445 9.14 ;
      RECT 42.555 3.66 42.875 3.98 ;
      RECT 42.24 3.69 42.875 3.86 ;
      RECT 36.175 3.665 36.455 4.035 ;
      RECT 36.22 2.9 36.39 4.035 ;
      RECT 40.885 3.29 41.21 3.615 ;
      RECT 40.96 2.9 41.13 3.615 ;
      RECT 36.22 2.9 41.13 3.07 ;
      RECT 39.915 6.075 40.175 6.395 ;
      RECT 39.975 4.035 40.115 6.395 ;
      RECT 39.915 4.035 40.175 4.355 ;
      RECT 38.895 7.095 39.155 7.415 ;
      RECT 38.275 7.185 39.155 7.325 ;
      RECT 38.275 5.025 38.415 7.325 ;
      RECT 38.215 5.025 38.495 5.395 ;
      RECT 37.535 7.065 37.815 7.435 ;
      RECT 37.595 5.145 37.735 7.435 ;
      RECT 37.595 5.145 38.075 5.285 ;
      RECT 37.935 3.355 38.075 5.285 ;
      RECT 37.875 3.355 38.135 3.675 ;
      RECT 36.855 6.045 37.135 6.415 ;
      RECT 36.915 3.695 37.055 6.415 ;
      RECT 36.855 3.695 37.115 4.015 ;
      RECT 36.485 7.065 36.765 7.435 ;
      RECT 36.485 7.095 36.775 7.415 ;
      RECT 25.97 8.565 26.29 8.89 ;
      RECT 26 7.98 26.17 8.89 ;
      RECT 26 7.98 26.175 8.33 ;
      RECT 26 7.98 26.975 8.155 ;
      RECT 26.8 3.26 26.975 8.155 ;
      RECT 26.745 3.26 27.095 3.61 ;
      RECT 15.635 9.705 25.815 9.875 ;
      RECT 25.655 3.69 25.815 9.875 ;
      RECT 15.635 8.885 15.805 9.875 ;
      RECT 11.87 9.28 12.15 9.62 ;
      RECT 11.87 9.345 13.06 9.515 ;
      RECT 12.89 8.97 13.06 9.515 ;
      RECT 26.77 8.94 27.095 9.265 ;
      RECT 15.58 8.885 15.86 9.225 ;
      RECT 25.655 9.03 27.095 9.2 ;
      RECT 12.89 8.97 15.86 9.14 ;
      RECT 25.97 3.66 26.29 3.98 ;
      RECT 25.655 3.69 26.29 3.86 ;
      RECT 19.59 3.665 19.87 4.035 ;
      RECT 19.635 2.9 19.805 4.035 ;
      RECT 24.3 3.29 24.625 3.615 ;
      RECT 24.375 2.9 24.545 3.615 ;
      RECT 19.635 2.9 24.545 3.07 ;
      RECT 23.33 6.075 23.59 6.395 ;
      RECT 23.39 4.035 23.53 6.395 ;
      RECT 23.33 4.035 23.59 4.355 ;
      RECT 22.31 7.095 22.57 7.415 ;
      RECT 21.69 7.185 22.57 7.325 ;
      RECT 21.69 5.025 21.83 7.325 ;
      RECT 21.63 5.025 21.91 5.395 ;
      RECT 20.95 7.065 21.23 7.435 ;
      RECT 21.01 5.145 21.15 7.435 ;
      RECT 21.01 5.145 21.49 5.285 ;
      RECT 21.35 3.355 21.49 5.285 ;
      RECT 21.29 3.355 21.55 3.675 ;
      RECT 20.27 6.045 20.55 6.415 ;
      RECT 20.33 3.695 20.47 6.415 ;
      RECT 20.27 3.695 20.53 4.015 ;
      RECT 19.9 7.065 20.18 7.435 ;
      RECT 19.9 7.095 20.19 7.415 ;
      RECT 87.965 4.005 88.245 4.375 ;
      RECT 87.265 4.345 87.545 4.715 ;
      RECT 71.385 4.005 71.665 4.375 ;
      RECT 70.685 4.345 70.965 4.715 ;
      RECT 64.805 9.28 65.175 9.65 ;
      RECT 54.8 4.005 55.08 4.375 ;
      RECT 54.1 4.345 54.38 4.715 ;
      RECT 48.22 9.28 48.59 9.65 ;
      RECT 38.215 4.005 38.495 4.375 ;
      RECT 37.515 4.345 37.795 4.715 ;
      RECT 31.635 9.28 32.005 9.65 ;
      RECT 21.63 4.005 21.91 4.375 ;
      RECT 20.93 4.345 21.21 4.715 ;
      RECT 15.05 9.28 15.42 9.65 ;
    LAYER via1 ;
      RECT 95.55 9.67 95.7 9.82 ;
      RECT 93.195 9.025 93.345 9.175 ;
      RECT 93.18 3.36 93.33 3.51 ;
      RECT 92.39 3.745 92.54 3.895 ;
      RECT 92.39 8.655 92.54 8.805 ;
      RECT 90.725 3.375 90.875 3.525 ;
      RECT 89.72 4.12 89.87 4.27 ;
      RECT 89.72 6.16 89.87 6.31 ;
      RECT 88.7 7.18 88.85 7.33 ;
      RECT 88.02 4.12 88.17 4.27 ;
      RECT 88.02 5.14 88.17 5.29 ;
      RECT 87.68 3.44 87.83 3.59 ;
      RECT 87.34 4.46 87.49 4.61 ;
      RECT 87.34 7.18 87.49 7.33 ;
      RECT 86.66 3.78 86.81 3.93 ;
      RECT 86.66 6.16 86.81 6.31 ;
      RECT 86.32 7.18 86.47 7.33 ;
      RECT 85.98 3.77 86.13 3.92 ;
      RECT 81.98 8.98 82.13 9.13 ;
      RECT 81.495 9.39 81.645 9.54 ;
      RECT 79.005 9.025 79.155 9.175 ;
      RECT 76.615 9.025 76.765 9.175 ;
      RECT 76.6 3.36 76.75 3.51 ;
      RECT 75.81 3.745 75.96 3.895 ;
      RECT 75.81 8.655 75.96 8.805 ;
      RECT 74.145 3.375 74.295 3.525 ;
      RECT 73.14 4.12 73.29 4.27 ;
      RECT 73.14 6.16 73.29 6.31 ;
      RECT 72.12 7.18 72.27 7.33 ;
      RECT 71.44 4.12 71.59 4.27 ;
      RECT 71.44 5.14 71.59 5.29 ;
      RECT 71.1 3.44 71.25 3.59 ;
      RECT 70.76 4.46 70.91 4.61 ;
      RECT 70.76 7.18 70.91 7.33 ;
      RECT 70.08 3.78 70.23 3.93 ;
      RECT 70.08 6.16 70.23 6.31 ;
      RECT 69.74 7.18 69.89 7.33 ;
      RECT 69.4 3.77 69.55 3.92 ;
      RECT 65.4 8.98 65.55 9.13 ;
      RECT 64.915 9.39 65.065 9.54 ;
      RECT 62.42 9.025 62.57 9.175 ;
      RECT 60.03 9.025 60.18 9.175 ;
      RECT 60.015 3.36 60.165 3.51 ;
      RECT 59.225 3.745 59.375 3.895 ;
      RECT 59.225 8.655 59.375 8.805 ;
      RECT 57.56 3.375 57.71 3.525 ;
      RECT 56.555 4.12 56.705 4.27 ;
      RECT 56.555 6.16 56.705 6.31 ;
      RECT 55.535 7.18 55.685 7.33 ;
      RECT 54.855 4.12 55.005 4.27 ;
      RECT 54.855 5.14 55.005 5.29 ;
      RECT 54.515 3.44 54.665 3.59 ;
      RECT 54.175 4.46 54.325 4.61 ;
      RECT 54.175 7.18 54.325 7.33 ;
      RECT 53.495 3.78 53.645 3.93 ;
      RECT 53.495 6.16 53.645 6.31 ;
      RECT 53.155 7.18 53.305 7.33 ;
      RECT 52.815 3.77 52.965 3.92 ;
      RECT 48.815 8.98 48.965 9.13 ;
      RECT 48.33 9.39 48.48 9.54 ;
      RECT 45.835 9.025 45.985 9.175 ;
      RECT 43.445 9.025 43.595 9.175 ;
      RECT 43.43 3.36 43.58 3.51 ;
      RECT 42.64 3.745 42.79 3.895 ;
      RECT 42.64 8.655 42.79 8.805 ;
      RECT 40.975 3.375 41.125 3.525 ;
      RECT 39.97 4.12 40.12 4.27 ;
      RECT 39.97 6.16 40.12 6.31 ;
      RECT 38.95 7.18 39.1 7.33 ;
      RECT 38.27 4.12 38.42 4.27 ;
      RECT 38.27 5.14 38.42 5.29 ;
      RECT 37.93 3.44 38.08 3.59 ;
      RECT 37.59 4.46 37.74 4.61 ;
      RECT 37.59 7.18 37.74 7.33 ;
      RECT 36.91 3.78 37.06 3.93 ;
      RECT 36.91 6.16 37.06 6.31 ;
      RECT 36.57 7.18 36.72 7.33 ;
      RECT 36.23 3.77 36.38 3.92 ;
      RECT 32.23 8.98 32.38 9.13 ;
      RECT 31.745 9.39 31.895 9.54 ;
      RECT 29.25 9.025 29.4 9.175 ;
      RECT 26.86 9.025 27.01 9.175 ;
      RECT 26.845 3.36 26.995 3.51 ;
      RECT 26.055 3.745 26.205 3.895 ;
      RECT 26.055 8.655 26.205 8.805 ;
      RECT 24.39 3.375 24.54 3.525 ;
      RECT 23.385 4.12 23.535 4.27 ;
      RECT 23.385 6.16 23.535 6.31 ;
      RECT 22.365 7.18 22.515 7.33 ;
      RECT 21.685 4.12 21.835 4.27 ;
      RECT 21.685 5.14 21.835 5.29 ;
      RECT 21.345 3.44 21.495 3.59 ;
      RECT 21.005 4.46 21.155 4.61 ;
      RECT 21.005 7.18 21.155 7.33 ;
      RECT 20.325 3.78 20.475 3.93 ;
      RECT 20.325 6.16 20.475 6.31 ;
      RECT 19.985 7.18 20.135 7.33 ;
      RECT 19.645 3.77 19.795 3.92 ;
      RECT 15.645 8.98 15.795 9.13 ;
      RECT 15.16 9.39 15.31 9.54 ;
      RECT 11.935 9.375 12.085 9.525 ;
      RECT 11.55 8.635 11.7 8.785 ;
    LAYER met1 ;
      RECT 95.43 10.055 95.72 10.285 ;
      RECT 95.49 8.575 95.66 10.285 ;
      RECT 95.46 9.585 95.785 9.91 ;
      RECT 95.43 8.575 95.72 8.805 ;
      RECT 95.025 4.03 95.35 4.26 ;
      RECT 95.025 4.06 95.52 4.23 ;
      RECT 95.025 3.69 95.215 4.26 ;
      RECT 94.44 3.66 94.73 3.89 ;
      RECT 94.44 3.69 95.215 3.86 ;
      RECT 94.5 2.18 94.67 3.89 ;
      RECT 94.44 2.18 94.73 2.41 ;
      RECT 94.44 10.055 94.73 10.285 ;
      RECT 94.5 8.575 94.67 10.285 ;
      RECT 94.44 8.575 94.73 8.805 ;
      RECT 94.44 8.61 95.295 8.77 ;
      RECT 95.125 8.205 95.295 8.77 ;
      RECT 94.44 8.605 94.835 8.77 ;
      RECT 95.06 8.205 95.35 8.435 ;
      RECT 95.06 8.235 95.52 8.405 ;
      RECT 94.07 4.03 94.36 4.26 ;
      RECT 94.07 4.06 94.53 4.23 ;
      RECT 94.135 2.95 94.3 4.26 ;
      RECT 92.65 2.92 92.94 3.15 ;
      RECT 92.65 2.95 94.3 3.12 ;
      RECT 92.71 2.18 92.88 3.15 ;
      RECT 92.65 2.18 92.94 2.41 ;
      RECT 92.65 10.05 92.94 10.28 ;
      RECT 92.71 9.31 92.88 10.28 ;
      RECT 92.71 9.405 94.3 9.575 ;
      RECT 94.13 8.205 94.3 9.575 ;
      RECT 92.65 9.31 92.94 9.54 ;
      RECT 94.07 8.205 94.36 8.435 ;
      RECT 94.07 8.235 94.53 8.405 ;
      RECT 90.635 3.29 90.96 3.615 ;
      RECT 93.08 3.26 93.43 3.61 ;
      RECT 90.635 3.32 93.43 3.49 ;
      RECT 93.105 8.94 93.43 9.265 ;
      RECT 93.08 8.94 93.43 9.17 ;
      RECT 92.91 8.97 93.43 9.14 ;
      RECT 92.305 3.66 92.625 3.98 ;
      RECT 92.275 3.66 92.625 3.89 ;
      RECT 91.99 3.69 92.625 3.86 ;
      RECT 92.305 8.565 92.625 8.89 ;
      RECT 92.275 8.57 92.625 8.8 ;
      RECT 92.105 8.6 92.625 8.77 ;
      RECT 89.635 4.065 89.955 4.325 ;
      RECT 89.355 4.125 89.955 4.265 ;
      RECT 87.255 4.405 87.575 4.665 ;
      RECT 89.225 4.415 89.515 4.645 ;
      RECT 87.255 4.465 89.52 4.605 ;
      RECT 88.615 7.125 88.935 7.385 ;
      RECT 88.615 7.185 89.205 7.325 ;
      RECT 87.935 4.065 88.255 4.325 ;
      RECT 83.195 4.075 83.485 4.305 ;
      RECT 83.195 4.125 88.255 4.265 ;
      RECT 88.025 3.785 88.165 4.325 ;
      RECT 88.025 3.785 88.505 3.925 ;
      RECT 88.365 3.395 88.505 3.925 ;
      RECT 88.285 3.395 88.575 3.625 ;
      RECT 87.935 5.085 88.255 5.345 ;
      RECT 87.265 5.095 87.555 5.325 ;
      RECT 85.055 5.095 85.345 5.325 ;
      RECT 85.055 5.145 88.255 5.285 ;
      RECT 86.235 7.125 86.555 7.385 ;
      RECT 87.945 7.135 88.235 7.365 ;
      RECT 85.565 7.135 85.855 7.365 ;
      RECT 85.565 7.185 86.555 7.325 ;
      RECT 88.025 6.845 88.165 7.365 ;
      RECT 86.325 6.845 86.465 7.385 ;
      RECT 86.325 6.845 88.165 6.985 ;
      RECT 85.225 3.735 85.515 3.965 ;
      RECT 85.305 3.445 85.445 3.965 ;
      RECT 87.595 3.385 87.915 3.645 ;
      RECT 87.495 3.395 87.915 3.625 ;
      RECT 85.305 3.445 87.915 3.585 ;
      RECT 86.575 3.725 86.895 3.985 ;
      RECT 86.575 3.785 87.165 3.925 ;
      RECT 86.575 6.105 86.895 6.365 ;
      RECT 83.865 6.115 84.155 6.345 ;
      RECT 83.865 6.165 86.895 6.305 ;
      RECT 85.895 3.685 86.225 4.015 ;
      RECT 85.895 3.735 86.355 3.965 ;
      RECT 85.895 3.785 86.375 3.925 ;
      RECT 85.775 3.785 85.785 3.925 ;
      RECT 85.785 3.775 86.355 3.915 ;
      RECT 81.885 8.915 82.225 9.195 ;
      RECT 81.855 8.94 82.225 9.17 ;
      RECT 81.685 8.97 82.225 9.14 ;
      RECT 81.425 10.05 81.715 10.28 ;
      RECT 81.485 9.28 81.655 10.28 ;
      RECT 81.385 9.28 81.755 9.65 ;
      RECT 78.85 10.055 79.14 10.285 ;
      RECT 78.91 8.575 79.08 10.285 ;
      RECT 78.91 8.94 79.24 9.265 ;
      RECT 78.85 8.575 79.14 8.805 ;
      RECT 78.445 4.03 78.77 4.26 ;
      RECT 78.445 4.06 78.94 4.23 ;
      RECT 78.445 3.69 78.635 4.26 ;
      RECT 77.86 3.66 78.15 3.89 ;
      RECT 77.86 3.69 78.635 3.86 ;
      RECT 77.92 2.18 78.09 3.89 ;
      RECT 77.86 2.18 78.15 2.41 ;
      RECT 77.86 10.055 78.15 10.285 ;
      RECT 77.92 8.575 78.09 10.285 ;
      RECT 77.86 8.575 78.15 8.805 ;
      RECT 77.86 8.61 78.715 8.77 ;
      RECT 78.545 8.205 78.715 8.77 ;
      RECT 77.86 8.605 78.255 8.77 ;
      RECT 78.48 8.205 78.77 8.435 ;
      RECT 78.48 8.235 78.94 8.405 ;
      RECT 77.49 4.03 77.78 4.26 ;
      RECT 77.49 4.06 77.95 4.23 ;
      RECT 77.555 2.95 77.72 4.26 ;
      RECT 76.07 2.92 76.36 3.15 ;
      RECT 76.07 2.95 77.72 3.12 ;
      RECT 76.13 2.18 76.3 3.15 ;
      RECT 76.07 2.18 76.36 2.41 ;
      RECT 76.07 10.05 76.36 10.28 ;
      RECT 76.13 9.31 76.3 10.28 ;
      RECT 76.13 9.405 77.72 9.575 ;
      RECT 77.55 8.205 77.72 9.575 ;
      RECT 76.07 9.31 76.36 9.54 ;
      RECT 77.49 8.205 77.78 8.435 ;
      RECT 77.49 8.235 77.95 8.405 ;
      RECT 74.055 3.29 74.38 3.615 ;
      RECT 76.5 3.26 76.85 3.61 ;
      RECT 74.055 3.32 76.85 3.49 ;
      RECT 76.525 8.94 76.85 9.265 ;
      RECT 76.5 8.94 76.85 9.17 ;
      RECT 76.33 8.97 76.85 9.14 ;
      RECT 75.725 3.66 76.045 3.98 ;
      RECT 75.695 3.66 76.045 3.89 ;
      RECT 75.41 3.69 76.045 3.86 ;
      RECT 75.725 8.565 76.045 8.89 ;
      RECT 75.695 8.57 76.045 8.8 ;
      RECT 75.525 8.6 76.045 8.77 ;
      RECT 73.055 4.065 73.375 4.325 ;
      RECT 72.775 4.125 73.375 4.265 ;
      RECT 70.675 4.405 70.995 4.665 ;
      RECT 72.645 4.415 72.935 4.645 ;
      RECT 70.675 4.465 72.94 4.605 ;
      RECT 72.035 7.125 72.355 7.385 ;
      RECT 72.035 7.185 72.625 7.325 ;
      RECT 71.355 4.065 71.675 4.325 ;
      RECT 66.615 4.075 66.905 4.305 ;
      RECT 66.615 4.125 71.675 4.265 ;
      RECT 71.445 3.785 71.585 4.325 ;
      RECT 71.445 3.785 71.925 3.925 ;
      RECT 71.785 3.395 71.925 3.925 ;
      RECT 71.705 3.395 71.995 3.625 ;
      RECT 71.355 5.085 71.675 5.345 ;
      RECT 70.685 5.095 70.975 5.325 ;
      RECT 68.475 5.095 68.765 5.325 ;
      RECT 68.475 5.145 71.675 5.285 ;
      RECT 69.655 7.125 69.975 7.385 ;
      RECT 71.365 7.135 71.655 7.365 ;
      RECT 68.985 7.135 69.275 7.365 ;
      RECT 68.985 7.185 69.975 7.325 ;
      RECT 71.445 6.845 71.585 7.365 ;
      RECT 69.745 6.845 69.885 7.385 ;
      RECT 69.745 6.845 71.585 6.985 ;
      RECT 68.645 3.735 68.935 3.965 ;
      RECT 68.725 3.445 68.865 3.965 ;
      RECT 71.015 3.385 71.335 3.645 ;
      RECT 70.915 3.395 71.335 3.625 ;
      RECT 68.725 3.445 71.335 3.585 ;
      RECT 69.995 3.725 70.315 3.985 ;
      RECT 69.995 3.785 70.585 3.925 ;
      RECT 69.995 6.105 70.315 6.365 ;
      RECT 67.285 6.115 67.575 6.345 ;
      RECT 67.285 6.165 70.315 6.305 ;
      RECT 69.315 3.685 69.645 4.015 ;
      RECT 69.315 3.735 69.775 3.965 ;
      RECT 69.315 3.785 69.795 3.925 ;
      RECT 69.195 3.785 69.205 3.925 ;
      RECT 69.205 3.775 69.775 3.915 ;
      RECT 65.305 8.915 65.645 9.195 ;
      RECT 65.275 8.94 65.645 9.17 ;
      RECT 65.105 8.97 65.645 9.14 ;
      RECT 64.845 10.05 65.135 10.28 ;
      RECT 64.905 9.28 65.075 10.28 ;
      RECT 64.805 9.28 65.175 9.65 ;
      RECT 62.265 10.055 62.555 10.285 ;
      RECT 62.325 8.575 62.495 10.285 ;
      RECT 62.325 8.94 62.655 9.265 ;
      RECT 62.265 8.575 62.555 8.805 ;
      RECT 61.86 4.03 62.185 4.26 ;
      RECT 61.86 4.06 62.355 4.23 ;
      RECT 61.86 3.69 62.05 4.26 ;
      RECT 61.275 3.66 61.565 3.89 ;
      RECT 61.275 3.69 62.05 3.86 ;
      RECT 61.335 2.18 61.505 3.89 ;
      RECT 61.275 2.18 61.565 2.41 ;
      RECT 61.275 10.055 61.565 10.285 ;
      RECT 61.335 8.575 61.505 10.285 ;
      RECT 61.275 8.575 61.565 8.805 ;
      RECT 61.275 8.61 62.13 8.77 ;
      RECT 61.96 8.205 62.13 8.77 ;
      RECT 61.275 8.605 61.67 8.77 ;
      RECT 61.895 8.205 62.185 8.435 ;
      RECT 61.895 8.235 62.355 8.405 ;
      RECT 60.905 4.03 61.195 4.26 ;
      RECT 60.905 4.06 61.365 4.23 ;
      RECT 60.97 2.95 61.135 4.26 ;
      RECT 59.485 2.92 59.775 3.15 ;
      RECT 59.485 2.95 61.135 3.12 ;
      RECT 59.545 2.18 59.715 3.15 ;
      RECT 59.485 2.18 59.775 2.41 ;
      RECT 59.485 10.05 59.775 10.28 ;
      RECT 59.545 9.31 59.715 10.28 ;
      RECT 59.545 9.405 61.135 9.575 ;
      RECT 60.965 8.205 61.135 9.575 ;
      RECT 59.485 9.31 59.775 9.54 ;
      RECT 60.905 8.205 61.195 8.435 ;
      RECT 60.905 8.235 61.365 8.405 ;
      RECT 57.47 3.29 57.795 3.615 ;
      RECT 59.915 3.26 60.265 3.61 ;
      RECT 57.47 3.32 60.265 3.49 ;
      RECT 59.94 8.94 60.265 9.265 ;
      RECT 59.915 8.94 60.265 9.17 ;
      RECT 59.745 8.97 60.265 9.14 ;
      RECT 59.14 3.66 59.46 3.98 ;
      RECT 59.11 3.66 59.46 3.89 ;
      RECT 58.825 3.69 59.46 3.86 ;
      RECT 59.14 8.565 59.46 8.89 ;
      RECT 59.11 8.57 59.46 8.8 ;
      RECT 58.94 8.6 59.46 8.77 ;
      RECT 56.47 4.065 56.79 4.325 ;
      RECT 56.19 4.125 56.79 4.265 ;
      RECT 54.09 4.405 54.41 4.665 ;
      RECT 56.06 4.415 56.35 4.645 ;
      RECT 54.09 4.465 56.355 4.605 ;
      RECT 55.45 7.125 55.77 7.385 ;
      RECT 55.45 7.185 56.04 7.325 ;
      RECT 54.77 4.065 55.09 4.325 ;
      RECT 50.03 4.075 50.32 4.305 ;
      RECT 50.03 4.125 55.09 4.265 ;
      RECT 54.86 3.785 55 4.325 ;
      RECT 54.86 3.785 55.34 3.925 ;
      RECT 55.2 3.395 55.34 3.925 ;
      RECT 55.12 3.395 55.41 3.625 ;
      RECT 54.77 5.085 55.09 5.345 ;
      RECT 54.1 5.095 54.39 5.325 ;
      RECT 51.89 5.095 52.18 5.325 ;
      RECT 51.89 5.145 55.09 5.285 ;
      RECT 53.07 7.125 53.39 7.385 ;
      RECT 54.78 7.135 55.07 7.365 ;
      RECT 52.4 7.135 52.69 7.365 ;
      RECT 52.4 7.185 53.39 7.325 ;
      RECT 54.86 6.845 55 7.365 ;
      RECT 53.16 6.845 53.3 7.385 ;
      RECT 53.16 6.845 55 6.985 ;
      RECT 52.06 3.735 52.35 3.965 ;
      RECT 52.14 3.445 52.28 3.965 ;
      RECT 54.43 3.385 54.75 3.645 ;
      RECT 54.33 3.395 54.75 3.625 ;
      RECT 52.14 3.445 54.75 3.585 ;
      RECT 53.41 3.725 53.73 3.985 ;
      RECT 53.41 3.785 54 3.925 ;
      RECT 53.41 6.105 53.73 6.365 ;
      RECT 50.7 6.115 50.99 6.345 ;
      RECT 50.7 6.165 53.73 6.305 ;
      RECT 52.73 3.685 53.06 4.015 ;
      RECT 52.73 3.735 53.19 3.965 ;
      RECT 52.73 3.785 53.21 3.925 ;
      RECT 52.61 3.785 52.62 3.925 ;
      RECT 52.62 3.775 53.19 3.915 ;
      RECT 48.72 8.915 49.06 9.195 ;
      RECT 48.69 8.94 49.06 9.17 ;
      RECT 48.52 8.97 49.06 9.14 ;
      RECT 48.26 10.05 48.55 10.28 ;
      RECT 48.32 9.28 48.49 10.28 ;
      RECT 48.22 9.28 48.59 9.65 ;
      RECT 45.68 10.055 45.97 10.285 ;
      RECT 45.74 8.575 45.91 10.285 ;
      RECT 45.74 8.94 46.07 9.265 ;
      RECT 45.68 8.575 45.97 8.805 ;
      RECT 45.275 4.03 45.6 4.26 ;
      RECT 45.275 4.06 45.77 4.23 ;
      RECT 45.275 3.69 45.465 4.26 ;
      RECT 44.69 3.66 44.98 3.89 ;
      RECT 44.69 3.69 45.465 3.86 ;
      RECT 44.75 2.18 44.92 3.89 ;
      RECT 44.69 2.18 44.98 2.41 ;
      RECT 44.69 10.055 44.98 10.285 ;
      RECT 44.75 8.575 44.92 10.285 ;
      RECT 44.69 8.575 44.98 8.805 ;
      RECT 44.69 8.61 45.545 8.77 ;
      RECT 45.375 8.205 45.545 8.77 ;
      RECT 44.69 8.605 45.085 8.77 ;
      RECT 45.31 8.205 45.6 8.435 ;
      RECT 45.31 8.235 45.77 8.405 ;
      RECT 44.32 4.03 44.61 4.26 ;
      RECT 44.32 4.06 44.78 4.23 ;
      RECT 44.385 2.95 44.55 4.26 ;
      RECT 42.9 2.92 43.19 3.15 ;
      RECT 42.9 2.95 44.55 3.12 ;
      RECT 42.96 2.18 43.13 3.15 ;
      RECT 42.9 2.18 43.19 2.41 ;
      RECT 42.9 10.05 43.19 10.28 ;
      RECT 42.96 9.31 43.13 10.28 ;
      RECT 42.96 9.405 44.55 9.575 ;
      RECT 44.38 8.205 44.55 9.575 ;
      RECT 42.9 9.31 43.19 9.54 ;
      RECT 44.32 8.205 44.61 8.435 ;
      RECT 44.32 8.235 44.78 8.405 ;
      RECT 40.885 3.29 41.21 3.615 ;
      RECT 43.33 3.26 43.68 3.61 ;
      RECT 40.885 3.32 43.68 3.49 ;
      RECT 43.355 8.94 43.68 9.265 ;
      RECT 43.33 8.94 43.68 9.17 ;
      RECT 43.16 8.97 43.68 9.14 ;
      RECT 42.555 3.66 42.875 3.98 ;
      RECT 42.525 3.66 42.875 3.89 ;
      RECT 42.24 3.69 42.875 3.86 ;
      RECT 42.555 8.565 42.875 8.89 ;
      RECT 42.525 8.57 42.875 8.8 ;
      RECT 42.355 8.6 42.875 8.77 ;
      RECT 39.885 4.065 40.205 4.325 ;
      RECT 39.605 4.125 40.205 4.265 ;
      RECT 37.505 4.405 37.825 4.665 ;
      RECT 39.475 4.415 39.765 4.645 ;
      RECT 37.505 4.465 39.77 4.605 ;
      RECT 38.865 7.125 39.185 7.385 ;
      RECT 38.865 7.185 39.455 7.325 ;
      RECT 38.185 4.065 38.505 4.325 ;
      RECT 33.445 4.075 33.735 4.305 ;
      RECT 33.445 4.125 38.505 4.265 ;
      RECT 38.275 3.785 38.415 4.325 ;
      RECT 38.275 3.785 38.755 3.925 ;
      RECT 38.615 3.395 38.755 3.925 ;
      RECT 38.535 3.395 38.825 3.625 ;
      RECT 38.185 5.085 38.505 5.345 ;
      RECT 37.515 5.095 37.805 5.325 ;
      RECT 35.305 5.095 35.595 5.325 ;
      RECT 35.305 5.145 38.505 5.285 ;
      RECT 36.485 7.125 36.805 7.385 ;
      RECT 38.195 7.135 38.485 7.365 ;
      RECT 35.815 7.135 36.105 7.365 ;
      RECT 35.815 7.185 36.805 7.325 ;
      RECT 38.275 6.845 38.415 7.365 ;
      RECT 36.575 6.845 36.715 7.385 ;
      RECT 36.575 6.845 38.415 6.985 ;
      RECT 35.475 3.735 35.765 3.965 ;
      RECT 35.555 3.445 35.695 3.965 ;
      RECT 37.845 3.385 38.165 3.645 ;
      RECT 37.745 3.395 38.165 3.625 ;
      RECT 35.555 3.445 38.165 3.585 ;
      RECT 36.825 3.725 37.145 3.985 ;
      RECT 36.825 3.785 37.415 3.925 ;
      RECT 36.825 6.105 37.145 6.365 ;
      RECT 34.115 6.115 34.405 6.345 ;
      RECT 34.115 6.165 37.145 6.305 ;
      RECT 36.145 3.685 36.475 4.015 ;
      RECT 36.145 3.735 36.605 3.965 ;
      RECT 36.145 3.785 36.625 3.925 ;
      RECT 36.025 3.785 36.035 3.925 ;
      RECT 36.035 3.775 36.605 3.915 ;
      RECT 32.135 8.915 32.475 9.195 ;
      RECT 32.105 8.94 32.475 9.17 ;
      RECT 31.935 8.97 32.475 9.14 ;
      RECT 31.675 10.05 31.965 10.28 ;
      RECT 31.735 9.28 31.905 10.28 ;
      RECT 31.635 9.28 32.005 9.65 ;
      RECT 29.095 10.055 29.385 10.285 ;
      RECT 29.155 8.575 29.325 10.285 ;
      RECT 29.155 8.94 29.485 9.265 ;
      RECT 29.095 8.575 29.385 8.805 ;
      RECT 28.69 4.03 29.015 4.26 ;
      RECT 28.69 4.06 29.185 4.23 ;
      RECT 28.69 3.69 28.88 4.26 ;
      RECT 28.105 3.66 28.395 3.89 ;
      RECT 28.105 3.69 28.88 3.86 ;
      RECT 28.165 2.18 28.335 3.89 ;
      RECT 28.105 2.18 28.395 2.41 ;
      RECT 28.105 10.055 28.395 10.285 ;
      RECT 28.165 8.575 28.335 10.285 ;
      RECT 28.105 8.575 28.395 8.805 ;
      RECT 28.105 8.61 28.96 8.77 ;
      RECT 28.79 8.205 28.96 8.77 ;
      RECT 28.105 8.605 28.5 8.77 ;
      RECT 28.725 8.205 29.015 8.435 ;
      RECT 28.725 8.235 29.185 8.405 ;
      RECT 27.735 4.03 28.025 4.26 ;
      RECT 27.735 4.06 28.195 4.23 ;
      RECT 27.8 2.95 27.965 4.26 ;
      RECT 26.315 2.92 26.605 3.15 ;
      RECT 26.315 2.95 27.965 3.12 ;
      RECT 26.375 2.18 26.545 3.15 ;
      RECT 26.315 2.18 26.605 2.41 ;
      RECT 26.315 10.05 26.605 10.28 ;
      RECT 26.375 9.31 26.545 10.28 ;
      RECT 26.375 9.405 27.965 9.575 ;
      RECT 27.795 8.205 27.965 9.575 ;
      RECT 26.315 9.31 26.605 9.54 ;
      RECT 27.735 8.205 28.025 8.435 ;
      RECT 27.735 8.235 28.195 8.405 ;
      RECT 24.3 3.29 24.625 3.615 ;
      RECT 26.745 3.26 27.095 3.61 ;
      RECT 24.3 3.32 27.095 3.49 ;
      RECT 26.77 8.94 27.095 9.265 ;
      RECT 26.745 8.94 27.095 9.17 ;
      RECT 26.575 8.97 27.095 9.14 ;
      RECT 25.97 3.66 26.29 3.98 ;
      RECT 25.94 3.66 26.29 3.89 ;
      RECT 25.655 3.69 26.29 3.86 ;
      RECT 25.97 8.565 26.29 8.89 ;
      RECT 25.94 8.57 26.29 8.8 ;
      RECT 25.77 8.6 26.29 8.77 ;
      RECT 23.3 4.065 23.62 4.325 ;
      RECT 23.02 4.125 23.62 4.265 ;
      RECT 20.92 4.405 21.24 4.665 ;
      RECT 22.89 4.415 23.18 4.645 ;
      RECT 20.92 4.465 23.185 4.605 ;
      RECT 22.28 7.125 22.6 7.385 ;
      RECT 22.28 7.185 22.87 7.325 ;
      RECT 21.6 4.065 21.92 4.325 ;
      RECT 16.86 4.075 17.15 4.305 ;
      RECT 16.86 4.125 21.92 4.265 ;
      RECT 21.69 3.785 21.83 4.325 ;
      RECT 21.69 3.785 22.17 3.925 ;
      RECT 22.03 3.395 22.17 3.925 ;
      RECT 21.95 3.395 22.24 3.625 ;
      RECT 21.6 5.085 21.92 5.345 ;
      RECT 20.93 5.095 21.22 5.325 ;
      RECT 18.72 5.095 19.01 5.325 ;
      RECT 18.72 5.145 21.92 5.285 ;
      RECT 19.9 7.125 20.22 7.385 ;
      RECT 21.61 7.135 21.9 7.365 ;
      RECT 19.23 7.135 19.52 7.365 ;
      RECT 19.23 7.185 20.22 7.325 ;
      RECT 21.69 6.845 21.83 7.365 ;
      RECT 19.99 6.845 20.13 7.385 ;
      RECT 19.99 6.845 21.83 6.985 ;
      RECT 18.89 3.735 19.18 3.965 ;
      RECT 18.97 3.445 19.11 3.965 ;
      RECT 21.26 3.385 21.58 3.645 ;
      RECT 21.16 3.395 21.58 3.625 ;
      RECT 18.97 3.445 21.58 3.585 ;
      RECT 20.24 3.725 20.56 3.985 ;
      RECT 20.24 3.785 20.83 3.925 ;
      RECT 20.24 6.105 20.56 6.365 ;
      RECT 17.53 6.115 17.82 6.345 ;
      RECT 17.53 6.165 20.56 6.305 ;
      RECT 19.56 3.685 19.89 4.015 ;
      RECT 19.56 3.735 20.02 3.965 ;
      RECT 19.56 3.785 20.04 3.925 ;
      RECT 19.44 3.785 19.45 3.925 ;
      RECT 19.45 3.775 20.02 3.915 ;
      RECT 15.55 8.915 15.89 9.195 ;
      RECT 15.52 8.94 15.89 9.17 ;
      RECT 15.35 8.97 15.89 9.14 ;
      RECT 15.09 10.05 15.38 10.28 ;
      RECT 15.15 9.28 15.32 10.28 ;
      RECT 15.05 9.28 15.42 9.65 ;
      RECT 11.86 10.05 12.15 10.28 ;
      RECT 11.92 9.31 12.09 10.28 ;
      RECT 11.84 9.31 12.18 9.59 ;
      RECT 11.455 8.57 11.795 8.85 ;
      RECT 11.315 8.6 11.795 8.77 ;
      RECT 89.305 6.105 89.955 6.365 ;
      RECT 87.255 7.125 87.575 7.385 ;
      RECT 72.725 6.105 73.375 6.365 ;
      RECT 70.675 7.125 70.995 7.385 ;
      RECT 56.14 6.105 56.79 6.365 ;
      RECT 54.09 7.125 54.41 7.385 ;
      RECT 39.555 6.105 40.205 6.365 ;
      RECT 37.505 7.125 37.825 7.385 ;
      RECT 22.97 6.105 23.62 6.365 ;
      RECT 20.92 7.125 21.24 7.385 ;
    LAYER mcon ;
      RECT 95.49 8.605 95.66 8.775 ;
      RECT 95.49 10.085 95.66 10.255 ;
      RECT 95.12 4.06 95.29 4.23 ;
      RECT 95.12 8.235 95.29 8.405 ;
      RECT 94.5 2.21 94.67 2.38 ;
      RECT 94.5 3.69 94.67 3.86 ;
      RECT 94.5 8.605 94.67 8.775 ;
      RECT 94.5 10.085 94.67 10.255 ;
      RECT 94.13 4.06 94.3 4.23 ;
      RECT 94.13 8.235 94.3 8.405 ;
      RECT 93.14 3.32 93.31 3.49 ;
      RECT 93.14 8.97 93.31 9.14 ;
      RECT 92.71 2.21 92.88 2.38 ;
      RECT 92.71 2.95 92.88 3.12 ;
      RECT 92.71 9.34 92.88 9.51 ;
      RECT 92.71 10.08 92.88 10.25 ;
      RECT 92.335 3.69 92.505 3.86 ;
      RECT 92.335 8.6 92.505 8.77 ;
      RECT 89.705 4.105 89.875 4.275 ;
      RECT 89.365 6.145 89.535 6.315 ;
      RECT 89.285 4.445 89.455 4.615 ;
      RECT 88.685 7.165 88.855 7.335 ;
      RECT 88.345 3.425 88.515 3.595 ;
      RECT 88.005 7.165 88.175 7.335 ;
      RECT 87.555 3.425 87.725 3.595 ;
      RECT 87.325 5.125 87.495 5.295 ;
      RECT 87.325 7.165 87.495 7.335 ;
      RECT 86.645 3.765 86.815 3.935 ;
      RECT 86.125 3.765 86.295 3.935 ;
      RECT 85.625 7.165 85.795 7.335 ;
      RECT 85.285 3.765 85.455 3.935 ;
      RECT 85.115 5.125 85.285 5.295 ;
      RECT 83.925 6.145 84.095 6.315 ;
      RECT 83.255 4.105 83.425 4.275 ;
      RECT 81.915 8.97 82.085 9.14 ;
      RECT 81.485 9.34 81.655 9.51 ;
      RECT 81.485 10.08 81.655 10.25 ;
      RECT 78.91 8.605 79.08 8.775 ;
      RECT 78.91 10.085 79.08 10.255 ;
      RECT 78.54 4.06 78.71 4.23 ;
      RECT 78.54 8.235 78.71 8.405 ;
      RECT 77.92 2.21 78.09 2.38 ;
      RECT 77.92 3.69 78.09 3.86 ;
      RECT 77.92 8.605 78.09 8.775 ;
      RECT 77.92 10.085 78.09 10.255 ;
      RECT 77.55 4.06 77.72 4.23 ;
      RECT 77.55 8.235 77.72 8.405 ;
      RECT 76.56 3.32 76.73 3.49 ;
      RECT 76.56 8.97 76.73 9.14 ;
      RECT 76.13 2.21 76.3 2.38 ;
      RECT 76.13 2.95 76.3 3.12 ;
      RECT 76.13 9.34 76.3 9.51 ;
      RECT 76.13 10.08 76.3 10.25 ;
      RECT 75.755 3.69 75.925 3.86 ;
      RECT 75.755 8.6 75.925 8.77 ;
      RECT 73.125 4.105 73.295 4.275 ;
      RECT 72.785 6.145 72.955 6.315 ;
      RECT 72.705 4.445 72.875 4.615 ;
      RECT 72.105 7.165 72.275 7.335 ;
      RECT 71.765 3.425 71.935 3.595 ;
      RECT 71.425 7.165 71.595 7.335 ;
      RECT 70.975 3.425 71.145 3.595 ;
      RECT 70.745 5.125 70.915 5.295 ;
      RECT 70.745 7.165 70.915 7.335 ;
      RECT 70.065 3.765 70.235 3.935 ;
      RECT 69.545 3.765 69.715 3.935 ;
      RECT 69.045 7.165 69.215 7.335 ;
      RECT 68.705 3.765 68.875 3.935 ;
      RECT 68.535 5.125 68.705 5.295 ;
      RECT 67.345 6.145 67.515 6.315 ;
      RECT 66.675 4.105 66.845 4.275 ;
      RECT 65.335 8.97 65.505 9.14 ;
      RECT 64.905 9.34 65.075 9.51 ;
      RECT 64.905 10.08 65.075 10.25 ;
      RECT 62.325 8.605 62.495 8.775 ;
      RECT 62.325 10.085 62.495 10.255 ;
      RECT 61.955 4.06 62.125 4.23 ;
      RECT 61.955 8.235 62.125 8.405 ;
      RECT 61.335 2.21 61.505 2.38 ;
      RECT 61.335 3.69 61.505 3.86 ;
      RECT 61.335 8.605 61.505 8.775 ;
      RECT 61.335 10.085 61.505 10.255 ;
      RECT 60.965 4.06 61.135 4.23 ;
      RECT 60.965 8.235 61.135 8.405 ;
      RECT 59.975 3.32 60.145 3.49 ;
      RECT 59.975 8.97 60.145 9.14 ;
      RECT 59.545 2.21 59.715 2.38 ;
      RECT 59.545 2.95 59.715 3.12 ;
      RECT 59.545 9.34 59.715 9.51 ;
      RECT 59.545 10.08 59.715 10.25 ;
      RECT 59.17 3.69 59.34 3.86 ;
      RECT 59.17 8.6 59.34 8.77 ;
      RECT 56.54 4.105 56.71 4.275 ;
      RECT 56.2 6.145 56.37 6.315 ;
      RECT 56.12 4.445 56.29 4.615 ;
      RECT 55.52 7.165 55.69 7.335 ;
      RECT 55.18 3.425 55.35 3.595 ;
      RECT 54.84 7.165 55.01 7.335 ;
      RECT 54.39 3.425 54.56 3.595 ;
      RECT 54.16 5.125 54.33 5.295 ;
      RECT 54.16 7.165 54.33 7.335 ;
      RECT 53.48 3.765 53.65 3.935 ;
      RECT 52.96 3.765 53.13 3.935 ;
      RECT 52.46 7.165 52.63 7.335 ;
      RECT 52.12 3.765 52.29 3.935 ;
      RECT 51.95 5.125 52.12 5.295 ;
      RECT 50.76 6.145 50.93 6.315 ;
      RECT 50.09 4.105 50.26 4.275 ;
      RECT 48.75 8.97 48.92 9.14 ;
      RECT 48.32 9.34 48.49 9.51 ;
      RECT 48.32 10.08 48.49 10.25 ;
      RECT 45.74 8.605 45.91 8.775 ;
      RECT 45.74 10.085 45.91 10.255 ;
      RECT 45.37 4.06 45.54 4.23 ;
      RECT 45.37 8.235 45.54 8.405 ;
      RECT 44.75 2.21 44.92 2.38 ;
      RECT 44.75 3.69 44.92 3.86 ;
      RECT 44.75 8.605 44.92 8.775 ;
      RECT 44.75 10.085 44.92 10.255 ;
      RECT 44.38 4.06 44.55 4.23 ;
      RECT 44.38 8.235 44.55 8.405 ;
      RECT 43.39 3.32 43.56 3.49 ;
      RECT 43.39 8.97 43.56 9.14 ;
      RECT 42.96 2.21 43.13 2.38 ;
      RECT 42.96 2.95 43.13 3.12 ;
      RECT 42.96 9.34 43.13 9.51 ;
      RECT 42.96 10.08 43.13 10.25 ;
      RECT 42.585 3.69 42.755 3.86 ;
      RECT 42.585 8.6 42.755 8.77 ;
      RECT 39.955 4.105 40.125 4.275 ;
      RECT 39.615 6.145 39.785 6.315 ;
      RECT 39.535 4.445 39.705 4.615 ;
      RECT 38.935 7.165 39.105 7.335 ;
      RECT 38.595 3.425 38.765 3.595 ;
      RECT 38.255 7.165 38.425 7.335 ;
      RECT 37.805 3.425 37.975 3.595 ;
      RECT 37.575 5.125 37.745 5.295 ;
      RECT 37.575 7.165 37.745 7.335 ;
      RECT 36.895 3.765 37.065 3.935 ;
      RECT 36.375 3.765 36.545 3.935 ;
      RECT 35.875 7.165 36.045 7.335 ;
      RECT 35.535 3.765 35.705 3.935 ;
      RECT 35.365 5.125 35.535 5.295 ;
      RECT 34.175 6.145 34.345 6.315 ;
      RECT 33.505 4.105 33.675 4.275 ;
      RECT 32.165 8.97 32.335 9.14 ;
      RECT 31.735 9.34 31.905 9.51 ;
      RECT 31.735 10.08 31.905 10.25 ;
      RECT 29.155 8.605 29.325 8.775 ;
      RECT 29.155 10.085 29.325 10.255 ;
      RECT 28.785 4.06 28.955 4.23 ;
      RECT 28.785 8.235 28.955 8.405 ;
      RECT 28.165 2.21 28.335 2.38 ;
      RECT 28.165 3.69 28.335 3.86 ;
      RECT 28.165 8.605 28.335 8.775 ;
      RECT 28.165 10.085 28.335 10.255 ;
      RECT 27.795 4.06 27.965 4.23 ;
      RECT 27.795 8.235 27.965 8.405 ;
      RECT 26.805 3.32 26.975 3.49 ;
      RECT 26.805 8.97 26.975 9.14 ;
      RECT 26.375 2.21 26.545 2.38 ;
      RECT 26.375 2.95 26.545 3.12 ;
      RECT 26.375 9.34 26.545 9.51 ;
      RECT 26.375 10.08 26.545 10.25 ;
      RECT 26 3.69 26.17 3.86 ;
      RECT 26 8.6 26.17 8.77 ;
      RECT 23.37 4.105 23.54 4.275 ;
      RECT 23.03 6.145 23.2 6.315 ;
      RECT 22.95 4.445 23.12 4.615 ;
      RECT 22.35 7.165 22.52 7.335 ;
      RECT 22.01 3.425 22.18 3.595 ;
      RECT 21.67 7.165 21.84 7.335 ;
      RECT 21.22 3.425 21.39 3.595 ;
      RECT 20.99 5.125 21.16 5.295 ;
      RECT 20.99 7.165 21.16 7.335 ;
      RECT 20.31 3.765 20.48 3.935 ;
      RECT 19.79 3.765 19.96 3.935 ;
      RECT 19.29 7.165 19.46 7.335 ;
      RECT 18.95 3.765 19.12 3.935 ;
      RECT 18.78 5.125 18.95 5.295 ;
      RECT 17.59 6.145 17.76 6.315 ;
      RECT 16.92 4.105 17.09 4.275 ;
      RECT 15.58 8.97 15.75 9.14 ;
      RECT 15.15 9.34 15.32 9.51 ;
      RECT 15.15 10.08 15.32 10.25 ;
      RECT 11.92 9.34 12.09 9.51 ;
      RECT 11.92 10.08 12.09 10.25 ;
      RECT 11.545 8.6 11.715 8.77 ;
    LAYER li1 ;
      RECT 95.12 3.04 95.29 4.23 ;
      RECT 95.12 3.04 95.59 3.21 ;
      RECT 95.12 9.255 95.59 9.425 ;
      RECT 95.12 8.235 95.29 9.425 ;
      RECT 94.13 3.04 94.3 4.23 ;
      RECT 94.13 3.04 94.6 3.21 ;
      RECT 94.13 9.255 94.6 9.425 ;
      RECT 94.13 8.235 94.3 9.425 ;
      RECT 92.28 3.93 92.45 5.16 ;
      RECT 92.335 2.15 92.505 4.1 ;
      RECT 92.28 1.87 92.45 2.32 ;
      RECT 92.28 10.14 92.45 10.59 ;
      RECT 92.335 8.36 92.505 10.31 ;
      RECT 92.28 7.3 92.45 8.53 ;
      RECT 91.76 1.87 91.93 5.16 ;
      RECT 91.76 3.37 92.165 3.7 ;
      RECT 91.76 2.53 92.165 2.86 ;
      RECT 91.76 7.3 91.93 10.59 ;
      RECT 91.76 9.6 92.165 9.93 ;
      RECT 91.76 8.76 92.165 9.09 ;
      RECT 87.015 7.935 88.325 8.185 ;
      RECT 87.015 7.615 87.195 8.185 ;
      RECT 86.465 7.615 87.195 7.785 ;
      RECT 86.465 6.775 86.635 7.785 ;
      RECT 87.305 6.815 89.045 6.995 ;
      RECT 88.715 5.975 89.045 6.995 ;
      RECT 86.465 6.775 87.525 6.945 ;
      RECT 88.715 6.145 89.535 6.315 ;
      RECT 87.875 5.975 88.205 6.185 ;
      RECT 87.875 5.975 89.045 6.145 ;
      RECT 88.775 4.495 89.105 5.455 ;
      RECT 88.775 4.495 89.455 4.665 ;
      RECT 89.285 3.255 89.455 4.665 ;
      RECT 89.195 3.255 89.525 3.895 ;
      RECT 88.325 4.765 88.595 5.465 ;
      RECT 88.425 3.255 88.595 5.465 ;
      RECT 88.765 4.075 89.115 4.325 ;
      RECT 88.425 4.105 89.115 4.275 ;
      RECT 88.335 3.255 88.595 3.735 ;
      RECT 87.665 6.405 88.545 6.645 ;
      RECT 88.315 6.315 88.545 6.645 ;
      RECT 87.015 6.405 88.545 6.605 ;
      RECT 87.935 6.355 88.545 6.645 ;
      RECT 87.015 6.275 87.185 6.605 ;
      RECT 87.905 7.165 88.155 7.765 ;
      RECT 87.905 7.165 88.375 7.365 ;
      RECT 87.395 4.385 88.155 4.885 ;
      RECT 86.465 4.195 86.725 4.815 ;
      RECT 87.385 4.325 87.395 4.635 ;
      RECT 87.365 4.315 87.385 4.605 ;
      RECT 88.025 3.995 88.255 4.595 ;
      RECT 87.345 4.265 87.365 4.575 ;
      RECT 87.325 4.385 88.255 4.565 ;
      RECT 87.295 4.385 88.255 4.555 ;
      RECT 87.225 4.385 88.255 4.545 ;
      RECT 87.205 4.385 88.255 4.515 ;
      RECT 87.185 3.295 87.355 4.485 ;
      RECT 87.155 4.385 88.255 4.455 ;
      RECT 87.125 4.385 88.255 4.425 ;
      RECT 87.095 4.375 87.455 4.395 ;
      RECT 87.095 4.365 87.445 4.395 ;
      RECT 86.465 4.195 87.355 4.365 ;
      RECT 86.465 4.355 87.425 4.365 ;
      RECT 86.465 4.345 87.415 4.365 ;
      RECT 86.465 4.285 87.375 4.365 ;
      RECT 86.465 3.295 87.355 3.465 ;
      RECT 87.525 3.795 87.855 4.215 ;
      RECT 87.525 3.305 87.745 4.215 ;
      RECT 87.445 7.165 87.655 7.765 ;
      RECT 87.305 7.165 87.655 7.365 ;
      RECT 86.025 4.765 86.295 5.465 ;
      RECT 86.245 3.255 86.295 5.465 ;
      RECT 86.125 4.065 86.295 5.465 ;
      RECT 86.125 3.255 86.295 4.055 ;
      RECT 86.035 3.255 86.295 3.735 ;
      RECT 84.165 4.425 84.415 4.965 ;
      RECT 85.135 4.425 85.855 4.895 ;
      RECT 84.165 4.425 85.955 4.595 ;
      RECT 85.725 4.065 85.955 4.595 ;
      RECT 84.725 3.305 84.975 4.595 ;
      RECT 85.725 3.995 85.785 4.895 ;
      RECT 85.725 3.995 85.955 4.055 ;
      RECT 84.185 3.305 84.975 3.575 ;
      RECT 85.145 7.115 85.825 7.365 ;
      RECT 85.555 6.755 85.825 7.365 ;
      RECT 85.305 7.535 85.635 8.085 ;
      RECT 84.245 7.535 85.635 7.725 ;
      RECT 84.245 6.695 84.415 7.725 ;
      RECT 84.125 7.115 84.415 7.445 ;
      RECT 84.245 6.695 85.185 6.865 ;
      RECT 84.885 6.145 85.185 6.865 ;
      RECT 85.145 3.725 85.555 4.245 ;
      RECT 85.145 3.305 85.345 4.245 ;
      RECT 83.755 3.485 83.925 5.465 ;
      RECT 83.755 3.995 84.555 4.245 ;
      RECT 83.755 3.485 84.005 4.245 ;
      RECT 83.675 3.485 84.005 3.905 ;
      RECT 83.705 7.895 84.265 8.185 ;
      RECT 83.705 5.975 83.955 8.185 ;
      RECT 83.705 5.975 84.165 6.525 ;
      RECT 80.535 7.3 80.705 10.59 ;
      RECT 80.535 9.6 80.94 9.93 ;
      RECT 80.535 8.76 80.94 9.09 ;
      RECT 78.54 3.04 78.71 4.23 ;
      RECT 78.54 3.04 79.01 3.21 ;
      RECT 78.54 9.255 79.01 9.425 ;
      RECT 78.54 8.235 78.71 9.425 ;
      RECT 77.55 3.04 77.72 4.23 ;
      RECT 77.55 3.04 78.02 3.21 ;
      RECT 77.55 9.255 78.02 9.425 ;
      RECT 77.55 8.235 77.72 9.425 ;
      RECT 75.7 3.93 75.87 5.16 ;
      RECT 75.755 2.15 75.925 4.1 ;
      RECT 75.7 1.87 75.87 2.32 ;
      RECT 75.7 10.14 75.87 10.59 ;
      RECT 75.755 8.36 75.925 10.31 ;
      RECT 75.7 7.3 75.87 8.53 ;
      RECT 75.18 1.87 75.35 5.16 ;
      RECT 75.18 3.37 75.585 3.7 ;
      RECT 75.18 2.53 75.585 2.86 ;
      RECT 75.18 7.3 75.35 10.59 ;
      RECT 75.18 9.6 75.585 9.93 ;
      RECT 75.18 8.76 75.585 9.09 ;
      RECT 70.435 7.935 71.745 8.185 ;
      RECT 70.435 7.615 70.615 8.185 ;
      RECT 69.885 7.615 70.615 7.785 ;
      RECT 69.885 6.775 70.055 7.785 ;
      RECT 70.725 6.815 72.465 6.995 ;
      RECT 72.135 5.975 72.465 6.995 ;
      RECT 69.885 6.775 70.945 6.945 ;
      RECT 72.135 6.145 72.955 6.315 ;
      RECT 71.295 5.975 71.625 6.185 ;
      RECT 71.295 5.975 72.465 6.145 ;
      RECT 72.195 4.495 72.525 5.455 ;
      RECT 72.195 4.495 72.875 4.665 ;
      RECT 72.705 3.255 72.875 4.665 ;
      RECT 72.615 3.255 72.945 3.895 ;
      RECT 71.745 4.765 72.015 5.465 ;
      RECT 71.845 3.255 72.015 5.465 ;
      RECT 72.185 4.075 72.535 4.325 ;
      RECT 71.845 4.105 72.535 4.275 ;
      RECT 71.755 3.255 72.015 3.735 ;
      RECT 71.085 6.405 71.965 6.645 ;
      RECT 71.735 6.315 71.965 6.645 ;
      RECT 70.435 6.405 71.965 6.605 ;
      RECT 71.355 6.355 71.965 6.645 ;
      RECT 70.435 6.275 70.605 6.605 ;
      RECT 71.325 7.165 71.575 7.765 ;
      RECT 71.325 7.165 71.795 7.365 ;
      RECT 70.815 4.385 71.575 4.885 ;
      RECT 69.885 4.195 70.145 4.815 ;
      RECT 70.805 4.325 70.815 4.635 ;
      RECT 70.785 4.315 70.805 4.605 ;
      RECT 71.445 3.995 71.675 4.595 ;
      RECT 70.765 4.265 70.785 4.575 ;
      RECT 70.745 4.385 71.675 4.565 ;
      RECT 70.715 4.385 71.675 4.555 ;
      RECT 70.645 4.385 71.675 4.545 ;
      RECT 70.625 4.385 71.675 4.515 ;
      RECT 70.605 3.295 70.775 4.485 ;
      RECT 70.575 4.385 71.675 4.455 ;
      RECT 70.545 4.385 71.675 4.425 ;
      RECT 70.515 4.375 70.875 4.395 ;
      RECT 70.515 4.365 70.865 4.395 ;
      RECT 69.885 4.195 70.775 4.365 ;
      RECT 69.885 4.355 70.845 4.365 ;
      RECT 69.885 4.345 70.835 4.365 ;
      RECT 69.885 4.285 70.795 4.365 ;
      RECT 69.885 3.295 70.775 3.465 ;
      RECT 70.945 3.795 71.275 4.215 ;
      RECT 70.945 3.305 71.165 4.215 ;
      RECT 70.865 7.165 71.075 7.765 ;
      RECT 70.725 7.165 71.075 7.365 ;
      RECT 69.445 4.765 69.715 5.465 ;
      RECT 69.665 3.255 69.715 5.465 ;
      RECT 69.545 4.065 69.715 5.465 ;
      RECT 69.545 3.255 69.715 4.055 ;
      RECT 69.455 3.255 69.715 3.735 ;
      RECT 67.585 4.425 67.835 4.965 ;
      RECT 68.555 4.425 69.275 4.895 ;
      RECT 67.585 4.425 69.375 4.595 ;
      RECT 69.145 4.065 69.375 4.595 ;
      RECT 68.145 3.305 68.395 4.595 ;
      RECT 69.145 3.995 69.205 4.895 ;
      RECT 69.145 3.995 69.375 4.055 ;
      RECT 67.605 3.305 68.395 3.575 ;
      RECT 68.565 7.115 69.245 7.365 ;
      RECT 68.975 6.755 69.245 7.365 ;
      RECT 68.725 7.535 69.055 8.085 ;
      RECT 67.665 7.535 69.055 7.725 ;
      RECT 67.665 6.695 67.835 7.725 ;
      RECT 67.545 7.115 67.835 7.445 ;
      RECT 67.665 6.695 68.605 6.865 ;
      RECT 68.305 6.145 68.605 6.865 ;
      RECT 68.565 3.725 68.975 4.245 ;
      RECT 68.565 3.305 68.765 4.245 ;
      RECT 67.175 3.485 67.345 5.465 ;
      RECT 67.175 3.995 67.975 4.245 ;
      RECT 67.175 3.485 67.425 4.245 ;
      RECT 67.095 3.485 67.425 3.905 ;
      RECT 67.125 7.895 67.685 8.185 ;
      RECT 67.125 5.975 67.375 8.185 ;
      RECT 67.125 5.975 67.585 6.525 ;
      RECT 63.955 7.3 64.125 10.59 ;
      RECT 63.955 9.6 64.36 9.93 ;
      RECT 63.955 8.76 64.36 9.09 ;
      RECT 61.955 3.04 62.125 4.23 ;
      RECT 61.955 3.04 62.425 3.21 ;
      RECT 61.955 9.255 62.425 9.425 ;
      RECT 61.955 8.235 62.125 9.425 ;
      RECT 60.965 3.04 61.135 4.23 ;
      RECT 60.965 3.04 61.435 3.21 ;
      RECT 60.965 9.255 61.435 9.425 ;
      RECT 60.965 8.235 61.135 9.425 ;
      RECT 59.115 3.93 59.285 5.16 ;
      RECT 59.17 2.15 59.34 4.1 ;
      RECT 59.115 1.87 59.285 2.32 ;
      RECT 59.115 10.14 59.285 10.59 ;
      RECT 59.17 8.36 59.34 10.31 ;
      RECT 59.115 7.3 59.285 8.53 ;
      RECT 58.595 1.87 58.765 5.16 ;
      RECT 58.595 3.37 59 3.7 ;
      RECT 58.595 2.53 59 2.86 ;
      RECT 58.595 7.3 58.765 10.59 ;
      RECT 58.595 9.6 59 9.93 ;
      RECT 58.595 8.76 59 9.09 ;
      RECT 53.85 7.935 55.16 8.185 ;
      RECT 53.85 7.615 54.03 8.185 ;
      RECT 53.3 7.615 54.03 7.785 ;
      RECT 53.3 6.775 53.47 7.785 ;
      RECT 54.14 6.815 55.88 6.995 ;
      RECT 55.55 5.975 55.88 6.995 ;
      RECT 53.3 6.775 54.36 6.945 ;
      RECT 55.55 6.145 56.37 6.315 ;
      RECT 54.71 5.975 55.04 6.185 ;
      RECT 54.71 5.975 55.88 6.145 ;
      RECT 55.61 4.495 55.94 5.455 ;
      RECT 55.61 4.495 56.29 4.665 ;
      RECT 56.12 3.255 56.29 4.665 ;
      RECT 56.03 3.255 56.36 3.895 ;
      RECT 55.16 4.765 55.43 5.465 ;
      RECT 55.26 3.255 55.43 5.465 ;
      RECT 55.6 4.075 55.95 4.325 ;
      RECT 55.26 4.105 55.95 4.275 ;
      RECT 55.17 3.255 55.43 3.735 ;
      RECT 54.5 6.405 55.38 6.645 ;
      RECT 55.15 6.315 55.38 6.645 ;
      RECT 53.85 6.405 55.38 6.605 ;
      RECT 54.77 6.355 55.38 6.645 ;
      RECT 53.85 6.275 54.02 6.605 ;
      RECT 54.74 7.165 54.99 7.765 ;
      RECT 54.74 7.165 55.21 7.365 ;
      RECT 54.23 4.385 54.99 4.885 ;
      RECT 53.3 4.195 53.56 4.815 ;
      RECT 54.22 4.325 54.23 4.635 ;
      RECT 54.2 4.315 54.22 4.605 ;
      RECT 54.86 3.995 55.09 4.595 ;
      RECT 54.18 4.265 54.2 4.575 ;
      RECT 54.16 4.385 55.09 4.565 ;
      RECT 54.13 4.385 55.09 4.555 ;
      RECT 54.06 4.385 55.09 4.545 ;
      RECT 54.04 4.385 55.09 4.515 ;
      RECT 54.02 3.295 54.19 4.485 ;
      RECT 53.99 4.385 55.09 4.455 ;
      RECT 53.96 4.385 55.09 4.425 ;
      RECT 53.93 4.375 54.29 4.395 ;
      RECT 53.93 4.365 54.28 4.395 ;
      RECT 53.3 4.195 54.19 4.365 ;
      RECT 53.3 4.355 54.26 4.365 ;
      RECT 53.3 4.345 54.25 4.365 ;
      RECT 53.3 4.285 54.21 4.365 ;
      RECT 53.3 3.295 54.19 3.465 ;
      RECT 54.36 3.795 54.69 4.215 ;
      RECT 54.36 3.305 54.58 4.215 ;
      RECT 54.28 7.165 54.49 7.765 ;
      RECT 54.14 7.165 54.49 7.365 ;
      RECT 52.86 4.765 53.13 5.465 ;
      RECT 53.08 3.255 53.13 5.465 ;
      RECT 52.96 4.065 53.13 5.465 ;
      RECT 52.96 3.255 53.13 4.055 ;
      RECT 52.87 3.255 53.13 3.735 ;
      RECT 51 4.425 51.25 4.965 ;
      RECT 51.97 4.425 52.69 4.895 ;
      RECT 51 4.425 52.79 4.595 ;
      RECT 52.56 4.065 52.79 4.595 ;
      RECT 51.56 3.305 51.81 4.595 ;
      RECT 52.56 3.995 52.62 4.895 ;
      RECT 52.56 3.995 52.79 4.055 ;
      RECT 51.02 3.305 51.81 3.575 ;
      RECT 51.98 7.115 52.66 7.365 ;
      RECT 52.39 6.755 52.66 7.365 ;
      RECT 52.14 7.535 52.47 8.085 ;
      RECT 51.08 7.535 52.47 7.725 ;
      RECT 51.08 6.695 51.25 7.725 ;
      RECT 50.96 7.115 51.25 7.445 ;
      RECT 51.08 6.695 52.02 6.865 ;
      RECT 51.72 6.145 52.02 6.865 ;
      RECT 51.98 3.725 52.39 4.245 ;
      RECT 51.98 3.305 52.18 4.245 ;
      RECT 50.59 3.485 50.76 5.465 ;
      RECT 50.59 3.995 51.39 4.245 ;
      RECT 50.59 3.485 50.84 4.245 ;
      RECT 50.51 3.485 50.84 3.905 ;
      RECT 50.54 7.895 51.1 8.185 ;
      RECT 50.54 5.975 50.79 8.185 ;
      RECT 50.54 5.975 51 6.525 ;
      RECT 47.37 7.3 47.54 10.59 ;
      RECT 47.37 9.6 47.775 9.93 ;
      RECT 47.37 8.76 47.775 9.09 ;
      RECT 45.37 3.04 45.54 4.23 ;
      RECT 45.37 3.04 45.84 3.21 ;
      RECT 45.37 9.255 45.84 9.425 ;
      RECT 45.37 8.235 45.54 9.425 ;
      RECT 44.38 3.04 44.55 4.23 ;
      RECT 44.38 3.04 44.85 3.21 ;
      RECT 44.38 9.255 44.85 9.425 ;
      RECT 44.38 8.235 44.55 9.425 ;
      RECT 42.53 3.93 42.7 5.16 ;
      RECT 42.585 2.15 42.755 4.1 ;
      RECT 42.53 1.87 42.7 2.32 ;
      RECT 42.53 10.14 42.7 10.59 ;
      RECT 42.585 8.36 42.755 10.31 ;
      RECT 42.53 7.3 42.7 8.53 ;
      RECT 42.01 1.87 42.18 5.16 ;
      RECT 42.01 3.37 42.415 3.7 ;
      RECT 42.01 2.53 42.415 2.86 ;
      RECT 42.01 7.3 42.18 10.59 ;
      RECT 42.01 9.6 42.415 9.93 ;
      RECT 42.01 8.76 42.415 9.09 ;
      RECT 37.265 7.935 38.575 8.185 ;
      RECT 37.265 7.615 37.445 8.185 ;
      RECT 36.715 7.615 37.445 7.785 ;
      RECT 36.715 6.775 36.885 7.785 ;
      RECT 37.555 6.815 39.295 6.995 ;
      RECT 38.965 5.975 39.295 6.995 ;
      RECT 36.715 6.775 37.775 6.945 ;
      RECT 38.965 6.145 39.785 6.315 ;
      RECT 38.125 5.975 38.455 6.185 ;
      RECT 38.125 5.975 39.295 6.145 ;
      RECT 39.025 4.495 39.355 5.455 ;
      RECT 39.025 4.495 39.705 4.665 ;
      RECT 39.535 3.255 39.705 4.665 ;
      RECT 39.445 3.255 39.775 3.895 ;
      RECT 38.575 4.765 38.845 5.465 ;
      RECT 38.675 3.255 38.845 5.465 ;
      RECT 39.015 4.075 39.365 4.325 ;
      RECT 38.675 4.105 39.365 4.275 ;
      RECT 38.585 3.255 38.845 3.735 ;
      RECT 37.915 6.405 38.795 6.645 ;
      RECT 38.565 6.315 38.795 6.645 ;
      RECT 37.265 6.405 38.795 6.605 ;
      RECT 38.185 6.355 38.795 6.645 ;
      RECT 37.265 6.275 37.435 6.605 ;
      RECT 38.155 7.165 38.405 7.765 ;
      RECT 38.155 7.165 38.625 7.365 ;
      RECT 37.645 4.385 38.405 4.885 ;
      RECT 36.715 4.195 36.975 4.815 ;
      RECT 37.635 4.325 37.645 4.635 ;
      RECT 37.615 4.315 37.635 4.605 ;
      RECT 38.275 3.995 38.505 4.595 ;
      RECT 37.595 4.265 37.615 4.575 ;
      RECT 37.575 4.385 38.505 4.565 ;
      RECT 37.545 4.385 38.505 4.555 ;
      RECT 37.475 4.385 38.505 4.545 ;
      RECT 37.455 4.385 38.505 4.515 ;
      RECT 37.435 3.295 37.605 4.485 ;
      RECT 37.405 4.385 38.505 4.455 ;
      RECT 37.375 4.385 38.505 4.425 ;
      RECT 37.345 4.375 37.705 4.395 ;
      RECT 37.345 4.365 37.695 4.395 ;
      RECT 36.715 4.195 37.605 4.365 ;
      RECT 36.715 4.355 37.675 4.365 ;
      RECT 36.715 4.345 37.665 4.365 ;
      RECT 36.715 4.285 37.625 4.365 ;
      RECT 36.715 3.295 37.605 3.465 ;
      RECT 37.775 3.795 38.105 4.215 ;
      RECT 37.775 3.305 37.995 4.215 ;
      RECT 37.695 7.165 37.905 7.765 ;
      RECT 37.555 7.165 37.905 7.365 ;
      RECT 36.275 4.765 36.545 5.465 ;
      RECT 36.495 3.255 36.545 5.465 ;
      RECT 36.375 4.065 36.545 5.465 ;
      RECT 36.375 3.255 36.545 4.055 ;
      RECT 36.285 3.255 36.545 3.735 ;
      RECT 34.415 4.425 34.665 4.965 ;
      RECT 35.385 4.425 36.105 4.895 ;
      RECT 34.415 4.425 36.205 4.595 ;
      RECT 35.975 4.065 36.205 4.595 ;
      RECT 34.975 3.305 35.225 4.595 ;
      RECT 35.975 3.995 36.035 4.895 ;
      RECT 35.975 3.995 36.205 4.055 ;
      RECT 34.435 3.305 35.225 3.575 ;
      RECT 35.395 7.115 36.075 7.365 ;
      RECT 35.805 6.755 36.075 7.365 ;
      RECT 35.555 7.535 35.885 8.085 ;
      RECT 34.495 7.535 35.885 7.725 ;
      RECT 34.495 6.695 34.665 7.725 ;
      RECT 34.375 7.115 34.665 7.445 ;
      RECT 34.495 6.695 35.435 6.865 ;
      RECT 35.135 6.145 35.435 6.865 ;
      RECT 35.395 3.725 35.805 4.245 ;
      RECT 35.395 3.305 35.595 4.245 ;
      RECT 34.005 3.485 34.175 5.465 ;
      RECT 34.005 3.995 34.805 4.245 ;
      RECT 34.005 3.485 34.255 4.245 ;
      RECT 33.925 3.485 34.255 3.905 ;
      RECT 33.955 7.895 34.515 8.185 ;
      RECT 33.955 5.975 34.205 8.185 ;
      RECT 33.955 5.975 34.415 6.525 ;
      RECT 30.785 7.3 30.955 10.59 ;
      RECT 30.785 9.6 31.19 9.93 ;
      RECT 30.785 8.76 31.19 9.09 ;
      RECT 28.785 3.04 28.955 4.23 ;
      RECT 28.785 3.04 29.255 3.21 ;
      RECT 28.785 9.255 29.255 9.425 ;
      RECT 28.785 8.235 28.955 9.425 ;
      RECT 27.795 3.04 27.965 4.23 ;
      RECT 27.795 3.04 28.265 3.21 ;
      RECT 27.795 9.255 28.265 9.425 ;
      RECT 27.795 8.235 27.965 9.425 ;
      RECT 25.945 3.93 26.115 5.16 ;
      RECT 26 2.15 26.17 4.1 ;
      RECT 25.945 1.87 26.115 2.32 ;
      RECT 25.945 10.14 26.115 10.59 ;
      RECT 26 8.36 26.17 10.31 ;
      RECT 25.945 7.3 26.115 8.53 ;
      RECT 25.425 1.87 25.595 5.16 ;
      RECT 25.425 3.37 25.83 3.7 ;
      RECT 25.425 2.53 25.83 2.86 ;
      RECT 25.425 7.3 25.595 10.59 ;
      RECT 25.425 9.6 25.83 9.93 ;
      RECT 25.425 8.76 25.83 9.09 ;
      RECT 20.68 7.935 21.99 8.185 ;
      RECT 20.68 7.615 20.86 8.185 ;
      RECT 20.13 7.615 20.86 7.785 ;
      RECT 20.13 6.775 20.3 7.785 ;
      RECT 20.97 6.815 22.71 6.995 ;
      RECT 22.38 5.975 22.71 6.995 ;
      RECT 20.13 6.775 21.19 6.945 ;
      RECT 22.38 6.145 23.2 6.315 ;
      RECT 21.54 5.975 21.87 6.185 ;
      RECT 21.54 5.975 22.71 6.145 ;
      RECT 22.44 4.495 22.77 5.455 ;
      RECT 22.44 4.495 23.12 4.665 ;
      RECT 22.95 3.255 23.12 4.665 ;
      RECT 22.86 3.255 23.19 3.895 ;
      RECT 21.99 4.765 22.26 5.465 ;
      RECT 22.09 3.255 22.26 5.465 ;
      RECT 22.43 4.075 22.78 4.325 ;
      RECT 22.09 4.105 22.78 4.275 ;
      RECT 22 3.255 22.26 3.735 ;
      RECT 21.33 6.405 22.21 6.645 ;
      RECT 21.98 6.315 22.21 6.645 ;
      RECT 20.68 6.405 22.21 6.605 ;
      RECT 21.6 6.355 22.21 6.645 ;
      RECT 20.68 6.275 20.85 6.605 ;
      RECT 21.57 7.165 21.82 7.765 ;
      RECT 21.57 7.165 22.04 7.365 ;
      RECT 21.06 4.385 21.82 4.885 ;
      RECT 20.13 4.195 20.39 4.815 ;
      RECT 21.05 4.325 21.06 4.635 ;
      RECT 21.03 4.315 21.05 4.605 ;
      RECT 21.69 3.995 21.92 4.595 ;
      RECT 21.01 4.265 21.03 4.575 ;
      RECT 20.99 4.385 21.92 4.565 ;
      RECT 20.96 4.385 21.92 4.555 ;
      RECT 20.89 4.385 21.92 4.545 ;
      RECT 20.87 4.385 21.92 4.515 ;
      RECT 20.85 3.295 21.02 4.485 ;
      RECT 20.82 4.385 21.92 4.455 ;
      RECT 20.79 4.385 21.92 4.425 ;
      RECT 20.76 4.375 21.12 4.395 ;
      RECT 20.76 4.365 21.11 4.395 ;
      RECT 20.13 4.195 21.02 4.365 ;
      RECT 20.13 4.355 21.09 4.365 ;
      RECT 20.13 4.345 21.08 4.365 ;
      RECT 20.13 4.285 21.04 4.365 ;
      RECT 20.13 3.295 21.02 3.465 ;
      RECT 21.19 3.795 21.52 4.215 ;
      RECT 21.19 3.305 21.41 4.215 ;
      RECT 21.11 7.165 21.32 7.765 ;
      RECT 20.97 7.165 21.32 7.365 ;
      RECT 19.69 4.765 19.96 5.465 ;
      RECT 19.91 3.255 19.96 5.465 ;
      RECT 19.79 4.065 19.96 5.465 ;
      RECT 19.79 3.255 19.96 4.055 ;
      RECT 19.7 3.255 19.96 3.735 ;
      RECT 17.83 4.425 18.08 4.965 ;
      RECT 18.8 4.425 19.52 4.895 ;
      RECT 17.83 4.425 19.62 4.595 ;
      RECT 19.39 4.065 19.62 4.595 ;
      RECT 18.39 3.305 18.64 4.595 ;
      RECT 19.39 3.995 19.45 4.895 ;
      RECT 19.39 3.995 19.62 4.055 ;
      RECT 17.85 3.305 18.64 3.575 ;
      RECT 18.81 7.115 19.49 7.365 ;
      RECT 19.22 6.755 19.49 7.365 ;
      RECT 18.97 7.535 19.3 8.085 ;
      RECT 17.91 7.535 19.3 7.725 ;
      RECT 17.91 6.695 18.08 7.725 ;
      RECT 17.79 7.115 18.08 7.445 ;
      RECT 17.91 6.695 18.85 6.865 ;
      RECT 18.55 6.145 18.85 6.865 ;
      RECT 18.81 3.725 19.22 4.245 ;
      RECT 18.81 3.305 19.01 4.245 ;
      RECT 17.42 3.485 17.59 5.465 ;
      RECT 17.42 3.995 18.22 4.245 ;
      RECT 17.42 3.485 17.67 4.245 ;
      RECT 17.34 3.485 17.67 3.905 ;
      RECT 17.37 7.895 17.93 8.185 ;
      RECT 17.37 5.975 17.62 8.185 ;
      RECT 17.37 5.975 17.83 6.525 ;
      RECT 14.2 7.3 14.37 10.59 ;
      RECT 14.2 9.6 14.605 9.93 ;
      RECT 14.2 8.76 14.605 9.09 ;
      RECT 11.49 10.14 11.66 10.59 ;
      RECT 11.545 8.36 11.715 10.31 ;
      RECT 11.49 7.3 11.66 8.53 ;
      RECT 10.97 7.3 11.14 10.59 ;
      RECT 10.97 9.6 11.375 9.93 ;
      RECT 10.97 8.76 11.375 9.09 ;
      RECT 95.49 7.305 95.66 8.775 ;
      RECT 95.49 10.085 95.66 10.595 ;
      RECT 94.5 1.87 94.67 2.38 ;
      RECT 94.5 3.69 94.67 5.16 ;
      RECT 94.5 7.305 94.67 8.775 ;
      RECT 94.5 10.085 94.67 10.595 ;
      RECT 93.14 1.87 93.31 5.16 ;
      RECT 93.14 7.3 93.31 10.59 ;
      RECT 92.71 1.87 92.88 2.38 ;
      RECT 92.71 2.95 92.88 5.16 ;
      RECT 92.71 7.3 92.88 9.51 ;
      RECT 92.71 10.08 92.88 10.59 ;
      RECT 89.625 4.075 89.975 4.325 ;
      RECT 88.565 7.165 89.015 7.675 ;
      RECT 87.245 5.125 87.725 5.465 ;
      RECT 86.465 3.635 87.015 4.025 ;
      RECT 84.955 5.125 85.425 5.465 ;
      RECT 83.245 4.075 83.585 4.955 ;
      RECT 81.915 7.3 82.085 10.59 ;
      RECT 81.485 7.3 81.655 9.51 ;
      RECT 81.485 10.08 81.655 10.59 ;
      RECT 78.91 7.305 79.08 8.775 ;
      RECT 78.91 10.085 79.08 10.595 ;
      RECT 77.92 1.87 78.09 2.38 ;
      RECT 77.92 3.69 78.09 5.16 ;
      RECT 77.92 7.305 78.09 8.775 ;
      RECT 77.92 10.085 78.09 10.595 ;
      RECT 76.56 1.87 76.73 5.16 ;
      RECT 76.56 7.3 76.73 10.59 ;
      RECT 76.13 1.87 76.3 2.38 ;
      RECT 76.13 2.95 76.3 5.16 ;
      RECT 76.13 7.3 76.3 9.51 ;
      RECT 76.13 10.08 76.3 10.59 ;
      RECT 73.045 4.075 73.395 4.325 ;
      RECT 71.985 7.165 72.435 7.675 ;
      RECT 70.665 5.125 71.145 5.465 ;
      RECT 69.885 3.635 70.435 4.025 ;
      RECT 68.375 5.125 68.845 5.465 ;
      RECT 66.665 4.075 67.005 4.955 ;
      RECT 65.335 7.3 65.505 10.59 ;
      RECT 64.905 7.3 65.075 9.51 ;
      RECT 64.905 10.08 65.075 10.59 ;
      RECT 62.325 7.305 62.495 8.775 ;
      RECT 62.325 10.085 62.495 10.595 ;
      RECT 61.335 1.87 61.505 2.38 ;
      RECT 61.335 3.69 61.505 5.16 ;
      RECT 61.335 7.305 61.505 8.775 ;
      RECT 61.335 10.085 61.505 10.595 ;
      RECT 59.975 1.87 60.145 5.16 ;
      RECT 59.975 7.3 60.145 10.59 ;
      RECT 59.545 1.87 59.715 2.38 ;
      RECT 59.545 2.95 59.715 5.16 ;
      RECT 59.545 7.3 59.715 9.51 ;
      RECT 59.545 10.08 59.715 10.59 ;
      RECT 56.46 4.075 56.81 4.325 ;
      RECT 55.4 7.165 55.85 7.675 ;
      RECT 54.08 5.125 54.56 5.465 ;
      RECT 53.3 3.635 53.85 4.025 ;
      RECT 51.79 5.125 52.26 5.465 ;
      RECT 50.08 4.075 50.42 4.955 ;
      RECT 48.75 7.3 48.92 10.59 ;
      RECT 48.32 7.3 48.49 9.51 ;
      RECT 48.32 10.08 48.49 10.59 ;
      RECT 45.74 7.305 45.91 8.775 ;
      RECT 45.74 10.085 45.91 10.595 ;
      RECT 44.75 1.87 44.92 2.38 ;
      RECT 44.75 3.69 44.92 5.16 ;
      RECT 44.75 7.305 44.92 8.775 ;
      RECT 44.75 10.085 44.92 10.595 ;
      RECT 43.39 1.87 43.56 5.16 ;
      RECT 43.39 7.3 43.56 10.59 ;
      RECT 42.96 1.87 43.13 2.38 ;
      RECT 42.96 2.95 43.13 5.16 ;
      RECT 42.96 7.3 43.13 9.51 ;
      RECT 42.96 10.08 43.13 10.59 ;
      RECT 39.875 4.075 40.225 4.325 ;
      RECT 38.815 7.165 39.265 7.675 ;
      RECT 37.495 5.125 37.975 5.465 ;
      RECT 36.715 3.635 37.265 4.025 ;
      RECT 35.205 5.125 35.675 5.465 ;
      RECT 33.495 4.075 33.835 4.955 ;
      RECT 32.165 7.3 32.335 10.59 ;
      RECT 31.735 7.3 31.905 9.51 ;
      RECT 31.735 10.08 31.905 10.59 ;
      RECT 29.155 7.305 29.325 8.775 ;
      RECT 29.155 10.085 29.325 10.595 ;
      RECT 28.165 1.87 28.335 2.38 ;
      RECT 28.165 3.69 28.335 5.16 ;
      RECT 28.165 7.305 28.335 8.775 ;
      RECT 28.165 10.085 28.335 10.595 ;
      RECT 26.805 1.87 26.975 5.16 ;
      RECT 26.805 7.3 26.975 10.59 ;
      RECT 26.375 1.87 26.545 2.38 ;
      RECT 26.375 2.95 26.545 5.16 ;
      RECT 26.375 7.3 26.545 9.51 ;
      RECT 26.375 10.08 26.545 10.59 ;
      RECT 23.29 4.075 23.64 4.325 ;
      RECT 22.23 7.165 22.68 7.675 ;
      RECT 20.91 5.125 21.39 5.465 ;
      RECT 20.13 3.635 20.68 4.025 ;
      RECT 18.62 5.125 19.09 5.465 ;
      RECT 16.91 4.075 17.25 4.955 ;
      RECT 15.58 7.3 15.75 10.59 ;
      RECT 15.15 7.3 15.32 9.51 ;
      RECT 15.15 10.08 15.32 10.59 ;
      RECT 11.92 7.3 12.09 9.51 ;
      RECT 11.92 10.08 12.09 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0.015 1.295 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r1 ;
  SIZE 88.925 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 19.485 0.57 19.655 1.08 ;
        RECT 19.485 2.39 19.655 3.86 ;
      LAYER met1 ;
        RECT 19.425 2.36 19.715 2.59 ;
        RECT 19.425 0.88 19.715 1.11 ;
        RECT 19.485 0.88 19.655 2.59 ;
      LAYER mcon ;
        RECT 19.485 2.39 19.655 2.56 ;
        RECT 19.485 0.91 19.655 1.08 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 36.705 0.57 36.875 1.08 ;
        RECT 36.705 2.39 36.875 3.86 ;
      LAYER met1 ;
        RECT 36.645 2.36 36.935 2.59 ;
        RECT 36.645 0.88 36.935 1.11 ;
        RECT 36.705 0.88 36.875 2.59 ;
      LAYER mcon ;
        RECT 36.705 2.39 36.875 2.56 ;
        RECT 36.705 0.91 36.875 1.08 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 53.925 0.57 54.095 1.08 ;
        RECT 53.925 2.39 54.095 3.86 ;
      LAYER met1 ;
        RECT 53.865 2.36 54.155 2.59 ;
        RECT 53.865 0.88 54.155 1.11 ;
        RECT 53.925 0.88 54.095 2.59 ;
      LAYER mcon ;
        RECT 53.925 2.39 54.095 2.56 ;
        RECT 53.925 0.91 54.095 1.08 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 71.145 0.57 71.315 1.08 ;
        RECT 71.145 2.39 71.315 3.86 ;
      LAYER met1 ;
        RECT 71.085 2.36 71.375 2.59 ;
        RECT 71.085 0.88 71.375 1.11 ;
        RECT 71.145 0.88 71.315 2.59 ;
      LAYER mcon ;
        RECT 71.145 2.39 71.315 2.56 ;
        RECT 71.145 0.91 71.315 1.08 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 88.365 0.57 88.535 1.08 ;
        RECT 88.365 2.39 88.535 3.86 ;
      LAYER met1 ;
        RECT 88.305 2.36 88.595 2.59 ;
        RECT 88.305 0.88 88.595 1.11 ;
        RECT 88.365 0.88 88.535 2.59 ;
      LAYER mcon ;
        RECT 88.365 2.39 88.535 2.56 ;
        RECT 88.365 0.91 88.535 1.08 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.335 1.66 15.505 2.935 ;
        RECT 15.335 6.93 15.505 8.21 ;
        RECT 15.325 6.93 15.505 7.17 ;
        RECT 3.65 6.935 3.82 8.21 ;
      LAYER met2 ;
        RECT 15.255 6.845 15.58 7.17 ;
        RECT 15.255 3.495 15.58 3.82 ;
        RECT 5.955 8.025 15.505 8.195 ;
        RECT 15.335 6.845 15.505 8.195 ;
        RECT 15.325 3.495 15.495 7.17 ;
        RECT 5.9 6.85 6.18 7.19 ;
        RECT 5.955 6.85 6.125 8.195 ;
      LAYER met1 ;
        RECT 15.275 2.765 15.735 2.935 ;
        RECT 15.255 3.495 15.58 3.82 ;
        RECT 15.275 2.735 15.565 2.965 ;
        RECT 15.335 2.735 15.505 3.82 ;
        RECT 15.255 6.935 15.735 7.105 ;
        RECT 15.255 6.845 15.58 7.17 ;
        RECT 5.87 6.88 6.21 7.16 ;
        RECT 3.59 6.935 6.21 7.105 ;
        RECT 3.59 6.905 3.88 7.135 ;
      LAYER via1 ;
        RECT 5.965 6.945 6.115 7.095 ;
        RECT 15.345 6.93 15.495 7.08 ;
        RECT 15.345 3.58 15.495 3.73 ;
      LAYER mcon ;
        RECT 3.65 6.935 3.82 7.105 ;
        RECT 15.335 6.935 15.505 7.105 ;
        RECT 15.335 2.765 15.505 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 32.555 1.66 32.725 2.935 ;
        RECT 32.555 6.93 32.725 8.21 ;
        RECT 32.545 6.93 32.725 7.17 ;
        RECT 20.87 6.935 21.04 8.21 ;
      LAYER met2 ;
        RECT 32.475 6.845 32.8 7.17 ;
        RECT 32.475 3.495 32.8 3.82 ;
        RECT 23.175 8.025 32.725 8.195 ;
        RECT 32.555 6.845 32.725 8.195 ;
        RECT 32.545 3.495 32.715 7.17 ;
        RECT 23.12 6.85 23.4 7.19 ;
        RECT 23.175 6.85 23.345 8.195 ;
      LAYER met1 ;
        RECT 32.495 2.765 32.955 2.935 ;
        RECT 32.475 3.495 32.8 3.82 ;
        RECT 32.495 2.735 32.785 2.965 ;
        RECT 32.555 2.735 32.725 3.82 ;
        RECT 32.475 6.935 32.955 7.105 ;
        RECT 32.475 6.845 32.8 7.17 ;
        RECT 23.09 6.88 23.43 7.16 ;
        RECT 20.81 6.935 23.43 7.105 ;
        RECT 20.81 6.905 21.1 7.135 ;
      LAYER via1 ;
        RECT 23.185 6.945 23.335 7.095 ;
        RECT 32.565 6.93 32.715 7.08 ;
        RECT 32.565 3.58 32.715 3.73 ;
      LAYER mcon ;
        RECT 20.87 6.935 21.04 7.105 ;
        RECT 32.555 6.935 32.725 7.105 ;
        RECT 32.555 2.765 32.725 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 49.775 1.66 49.945 2.935 ;
        RECT 49.775 6.93 49.945 8.21 ;
        RECT 49.765 6.93 49.945 7.17 ;
        RECT 38.09 6.935 38.26 8.21 ;
      LAYER met2 ;
        RECT 49.695 6.845 50.02 7.17 ;
        RECT 49.695 3.495 50.02 3.82 ;
        RECT 40.395 8.025 49.945 8.195 ;
        RECT 49.775 6.845 49.945 8.195 ;
        RECT 49.765 3.495 49.935 7.17 ;
        RECT 40.34 6.85 40.62 7.19 ;
        RECT 40.395 6.85 40.565 8.195 ;
      LAYER met1 ;
        RECT 49.715 2.765 50.175 2.935 ;
        RECT 49.695 3.495 50.02 3.82 ;
        RECT 49.715 2.735 50.005 2.965 ;
        RECT 49.775 2.735 49.945 3.82 ;
        RECT 49.695 6.935 50.175 7.105 ;
        RECT 49.695 6.845 50.02 7.17 ;
        RECT 40.31 6.88 40.65 7.16 ;
        RECT 38.03 6.935 40.65 7.105 ;
        RECT 38.03 6.905 38.32 7.135 ;
      LAYER via1 ;
        RECT 40.405 6.945 40.555 7.095 ;
        RECT 49.785 6.93 49.935 7.08 ;
        RECT 49.785 3.58 49.935 3.73 ;
      LAYER mcon ;
        RECT 38.09 6.935 38.26 7.105 ;
        RECT 49.775 6.935 49.945 7.105 ;
        RECT 49.775 2.765 49.945 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 66.995 1.66 67.165 2.935 ;
        RECT 66.995 6.93 67.165 8.21 ;
        RECT 66.985 6.93 67.165 7.17 ;
        RECT 55.31 6.935 55.48 8.21 ;
      LAYER met2 ;
        RECT 66.915 6.845 67.24 7.17 ;
        RECT 66.915 3.495 67.24 3.82 ;
        RECT 57.615 8.025 67.165 8.195 ;
        RECT 66.995 6.845 67.165 8.195 ;
        RECT 66.985 3.495 67.155 7.17 ;
        RECT 57.56 6.85 57.84 7.19 ;
        RECT 57.615 6.85 57.785 8.195 ;
      LAYER met1 ;
        RECT 66.935 2.765 67.395 2.935 ;
        RECT 66.915 3.495 67.24 3.82 ;
        RECT 66.935 2.735 67.225 2.965 ;
        RECT 66.995 2.735 67.165 3.82 ;
        RECT 66.915 6.935 67.395 7.105 ;
        RECT 66.915 6.845 67.24 7.17 ;
        RECT 57.53 6.88 57.87 7.16 ;
        RECT 55.25 6.935 57.87 7.105 ;
        RECT 55.25 6.905 55.54 7.135 ;
      LAYER via1 ;
        RECT 57.625 6.945 57.775 7.095 ;
        RECT 67.005 6.93 67.155 7.08 ;
        RECT 67.005 3.58 67.155 3.73 ;
      LAYER mcon ;
        RECT 55.31 6.935 55.48 7.105 ;
        RECT 66.995 6.935 67.165 7.105 ;
        RECT 66.995 2.765 67.165 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 84.215 1.66 84.385 2.935 ;
        RECT 84.215 6.93 84.385 8.21 ;
        RECT 84.205 6.93 84.385 7.17 ;
        RECT 72.53 6.935 72.7 8.21 ;
      LAYER met2 ;
        RECT 84.135 6.845 84.46 7.17 ;
        RECT 84.135 3.495 84.46 3.82 ;
        RECT 74.835 8.025 84.385 8.195 ;
        RECT 84.215 6.845 84.385 8.195 ;
        RECT 84.205 3.495 84.375 7.17 ;
        RECT 74.78 6.85 75.06 7.19 ;
        RECT 74.835 6.85 75.005 8.195 ;
      LAYER met1 ;
        RECT 84.155 2.765 84.615 2.935 ;
        RECT 84.135 3.495 84.46 3.82 ;
        RECT 84.155 2.735 84.445 2.965 ;
        RECT 84.215 2.735 84.385 3.82 ;
        RECT 84.135 6.935 84.615 7.105 ;
        RECT 84.135 6.845 84.46 7.17 ;
        RECT 74.75 6.88 75.09 7.16 ;
        RECT 72.47 6.935 75.09 7.105 ;
        RECT 72.47 6.905 72.76 7.135 ;
      LAYER via1 ;
        RECT 74.845 6.945 74.995 7.095 ;
        RECT 84.225 6.93 84.375 7.08 ;
        RECT 84.225 3.58 84.375 3.73 ;
      LAYER mcon ;
        RECT 72.53 6.935 72.7 7.105 ;
        RECT 84.215 6.935 84.385 7.105 ;
        RECT 84.215 2.765 84.385 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.24 6.935 0.41 8.21 ;
      LAYER met1 ;
        RECT 0.18 6.935 0.64 7.105 ;
        RECT 0.18 6.905 0.47 7.135 ;
      LAYER mcon ;
        RECT 0.24 6.935 0.41 7.105 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 82.825 4.345 88.91 5.735 ;
        RECT 82.92 4.135 88.91 5.735 ;
        RECT 86.775 4.13 88.755 5.74 ;
        RECT 87.935 3.4 88.105 6.47 ;
        RECT 86.945 3.4 87.115 6.47 ;
        RECT 84.205 3.405 84.375 6.465 ;
        RECT 0 4.345 88.91 4.515 ;
        RECT 82.01 4.345 82.29 5.655 ;
        RECT 81.61 3.495 81.78 4.515 ;
        RECT 81.08 4.345 81.34 5.655 ;
        RECT 80.77 3.835 80.94 4.515 ;
        RECT 80.63 4.345 80.91 5.655 ;
        RECT 79.7 4.345 79.96 5.655 ;
        RECT 79.27 4.345 79.53 5.655 ;
        RECT 79.19 3.205 79.52 4.515 ;
        RECT 78.32 4.345 78.6 5.655 ;
        RECT 76.95 3.205 77.28 4.515 ;
        RECT 76.97 3.205 77.23 5.655 ;
        RECT 76.5 3.205 76.73 4.515 ;
        RECT 76.02 4.345 76.3 5.655 ;
        RECT 65.7 4.135 75.83 4.515 ;
        RECT 75.62 3.205 75.83 4.515 ;
        RECT 71.685 4.13 75.83 4.515 ;
        RECT 65.605 4.345 75.49 5.705 ;
        RECT 72.345 4.13 75.36 5.735 ;
        RECT 72.52 4.13 72.69 6.465 ;
        RECT 65.605 4.345 75.36 5.73 ;
        RECT 65.605 4.345 71.69 5.735 ;
        RECT 69.555 4.13 71.535 5.74 ;
        RECT 70.715 3.4 70.885 6.47 ;
        RECT 69.725 3.4 69.895 6.47 ;
        RECT 66.985 3.405 67.155 6.465 ;
        RECT 64.79 4.345 65.07 5.655 ;
        RECT 64.39 3.495 64.56 4.515 ;
        RECT 63.86 4.345 64.12 5.655 ;
        RECT 63.55 3.835 63.72 4.515 ;
        RECT 63.41 4.345 63.69 5.655 ;
        RECT 62.48 4.345 62.74 5.655 ;
        RECT 62.05 4.345 62.31 5.655 ;
        RECT 61.97 3.205 62.3 4.515 ;
        RECT 61.1 4.345 61.38 5.655 ;
        RECT 59.73 3.205 60.06 4.515 ;
        RECT 59.75 3.205 60.01 5.655 ;
        RECT 59.28 3.205 59.51 4.515 ;
        RECT 58.8 4.345 59.08 5.655 ;
        RECT 48.48 4.135 58.61 4.515 ;
        RECT 58.4 3.205 58.61 4.515 ;
        RECT 54.465 4.13 58.61 4.515 ;
        RECT 48.385 4.345 58.27 5.705 ;
        RECT 55.125 4.13 58.14 5.735 ;
        RECT 55.3 4.13 55.47 6.465 ;
        RECT 48.385 4.345 58.14 5.73 ;
        RECT 48.385 4.345 54.47 5.735 ;
        RECT 52.335 4.13 54.315 5.74 ;
        RECT 53.495 3.4 53.665 6.47 ;
        RECT 52.505 3.4 52.675 6.47 ;
        RECT 49.765 3.405 49.935 6.465 ;
        RECT 47.57 4.345 47.85 5.655 ;
        RECT 47.17 3.495 47.34 4.515 ;
        RECT 46.64 4.345 46.9 5.655 ;
        RECT 46.33 3.835 46.5 4.515 ;
        RECT 46.19 4.345 46.47 5.655 ;
        RECT 45.26 4.345 45.52 5.655 ;
        RECT 44.83 4.345 45.09 5.655 ;
        RECT 44.75 3.205 45.08 4.515 ;
        RECT 43.88 4.345 44.16 5.655 ;
        RECT 42.51 3.205 42.84 4.515 ;
        RECT 42.53 3.205 42.79 5.655 ;
        RECT 42.06 3.205 42.29 4.515 ;
        RECT 41.58 4.345 41.86 5.655 ;
        RECT 31.26 4.135 41.39 4.515 ;
        RECT 41.18 3.205 41.39 4.515 ;
        RECT 37.245 4.13 41.39 4.515 ;
        RECT 31.165 4.345 41.05 5.705 ;
        RECT 31.165 4.345 40.92 5.735 ;
        RECT 38.08 4.13 38.25 6.465 ;
        RECT 35.115 4.13 37.095 5.74 ;
        RECT 36.275 3.4 36.445 6.47 ;
        RECT 35.285 3.4 35.455 6.47 ;
        RECT 32.545 3.405 32.715 6.465 ;
        RECT 30.35 4.345 30.63 5.655 ;
        RECT 29.95 3.495 30.12 4.515 ;
        RECT 29.42 4.345 29.68 5.655 ;
        RECT 29.11 3.835 29.28 4.515 ;
        RECT 28.97 4.345 29.25 5.655 ;
        RECT 28.04 4.345 28.3 5.655 ;
        RECT 27.61 4.345 27.87 5.655 ;
        RECT 27.53 3.205 27.86 4.515 ;
        RECT 26.66 4.345 26.94 5.655 ;
        RECT 25.29 3.205 25.62 4.515 ;
        RECT 25.31 3.205 25.57 5.655 ;
        RECT 24.84 3.205 25.07 4.515 ;
        RECT 24.36 4.345 24.64 5.655 ;
        RECT 14.04 4.135 24.17 4.515 ;
        RECT 23.96 3.205 24.17 4.515 ;
        RECT 20.025 4.13 24.17 4.515 ;
        RECT 13.945 4.345 23.83 5.705 ;
        RECT 20.685 4.13 23.7 5.735 ;
        RECT 20.86 4.13 21.03 6.465 ;
        RECT 13.945 4.345 23.7 5.73 ;
        RECT 13.945 4.345 20.03 5.735 ;
        RECT 17.895 4.13 19.875 5.74 ;
        RECT 19.055 3.4 19.225 6.47 ;
        RECT 18.065 3.4 18.235 6.47 ;
        RECT 15.325 3.405 15.495 6.465 ;
        RECT 13.13 4.345 13.41 5.655 ;
        RECT 12.73 3.495 12.9 4.515 ;
        RECT 12.2 4.345 12.46 5.655 ;
        RECT 11.89 3.835 12.06 4.515 ;
        RECT 11.75 4.345 12.03 5.655 ;
        RECT 10.82 4.345 11.08 5.655 ;
        RECT 10.39 4.345 10.65 5.655 ;
        RECT 10.31 3.205 10.64 4.515 ;
        RECT 9.44 4.345 9.72 5.655 ;
        RECT 8.07 3.205 8.4 4.515 ;
        RECT 8.09 3.205 8.35 5.655 ;
        RECT 7.62 3.205 7.85 4.515 ;
        RECT 7.14 4.345 7.42 5.655 ;
        RECT 0 4.13 6.95 4.515 ;
        RECT 6.74 3.205 6.95 4.515 ;
        RECT 0 4.13 6.61 5.705 ;
        RECT 0 4.13 6.485 5.73 ;
        RECT 3.465 4.13 6.48 5.735 ;
        RECT 3.64 4.13 3.81 6.465 ;
        RECT 0.055 4.13 2.805 5.735 ;
        RECT 2.04 4.13 2.21 9.295 ;
        RECT 0.23 4.13 0.4 6.465 ;
      LAYER met1 ;
        RECT 82.825 4.19 88.91 5.735 ;
        RECT 82.92 4.135 88.91 5.735 ;
        RECT 86.775 4.13 88.755 5.74 ;
        RECT 0 4.19 88.91 4.67 ;
        RECT 65.7 4.135 75.65 4.67 ;
        RECT 71.685 4.13 75.65 4.67 ;
        RECT 65.605 4.19 75.49 5.705 ;
        RECT 65.605 4.19 75.36 5.735 ;
        RECT 69.555 4.13 71.535 5.74 ;
        RECT 48.48 4.135 58.43 4.67 ;
        RECT 54.465 4.13 58.43 4.67 ;
        RECT 48.385 4.19 58.27 5.705 ;
        RECT 48.385 4.19 58.14 5.735 ;
        RECT 52.335 4.13 54.315 5.74 ;
        RECT 31.26 4.135 41.21 4.67 ;
        RECT 37.245 4.13 41.21 4.67 ;
        RECT 31.165 4.19 41.05 5.705 ;
        RECT 31.165 4.19 40.92 5.735 ;
        RECT 35.115 4.13 37.095 5.74 ;
        RECT 14.04 4.135 23.99 4.67 ;
        RECT 20.025 4.13 23.99 4.67 ;
        RECT 13.945 4.19 23.83 5.705 ;
        RECT 13.945 4.19 23.7 5.735 ;
        RECT 17.895 4.13 19.875 5.74 ;
        RECT 0 4.13 6.77 4.67 ;
        RECT 0 4.13 6.61 5.705 ;
        RECT 0 4.13 6.485 5.73 ;
        RECT 3.465 4.13 6.48 5.735 ;
        RECT 0.055 4.13 2.805 5.735 ;
        RECT 1.98 7.645 2.27 7.875 ;
        RECT 1.81 7.675 2.27 7.845 ;
      LAYER mcon ;
        RECT 2.04 7.675 2.21 7.845 ;
        RECT 2.35 5.535 2.52 5.705 ;
        RECT 5.76 5.535 5.93 5.705 ;
        RECT 6.74 4.345 6.91 4.515 ;
        RECT 7.2 4.345 7.37 4.515 ;
        RECT 7.66 4.345 7.83 4.515 ;
        RECT 8.12 4.345 8.29 4.515 ;
        RECT 8.58 4.345 8.75 4.515 ;
        RECT 9.04 4.345 9.21 4.515 ;
        RECT 9.5 4.345 9.67 4.515 ;
        RECT 9.96 4.345 10.13 4.515 ;
        RECT 10.42 4.345 10.59 4.515 ;
        RECT 10.88 4.345 11.05 4.515 ;
        RECT 11.34 4.345 11.51 4.515 ;
        RECT 11.8 4.345 11.97 4.515 ;
        RECT 12.26 4.345 12.43 4.515 ;
        RECT 12.72 4.345 12.89 4.515 ;
        RECT 13.18 4.345 13.35 4.515 ;
        RECT 13.64 4.345 13.81 4.515 ;
        RECT 17.445 5.535 17.615 5.705 ;
        RECT 17.445 4.165 17.615 4.335 ;
        RECT 18.145 5.54 18.315 5.71 ;
        RECT 18.145 4.16 18.315 4.33 ;
        RECT 19.135 5.54 19.305 5.71 ;
        RECT 19.135 4.16 19.305 4.33 ;
        RECT 22.98 5.535 23.15 5.705 ;
        RECT 23.96 4.345 24.13 4.515 ;
        RECT 24.42 4.345 24.59 4.515 ;
        RECT 24.88 4.345 25.05 4.515 ;
        RECT 25.34 4.345 25.51 4.515 ;
        RECT 25.8 4.345 25.97 4.515 ;
        RECT 26.26 4.345 26.43 4.515 ;
        RECT 26.72 4.345 26.89 4.515 ;
        RECT 27.18 4.345 27.35 4.515 ;
        RECT 27.64 4.345 27.81 4.515 ;
        RECT 28.1 4.345 28.27 4.515 ;
        RECT 28.56 4.345 28.73 4.515 ;
        RECT 29.02 4.345 29.19 4.515 ;
        RECT 29.48 4.345 29.65 4.515 ;
        RECT 29.94 4.345 30.11 4.515 ;
        RECT 30.4 4.345 30.57 4.515 ;
        RECT 30.86 4.345 31.03 4.515 ;
        RECT 34.665 5.535 34.835 5.705 ;
        RECT 34.665 4.165 34.835 4.335 ;
        RECT 35.365 5.54 35.535 5.71 ;
        RECT 35.365 4.16 35.535 4.33 ;
        RECT 36.355 5.54 36.525 5.71 ;
        RECT 36.355 4.16 36.525 4.33 ;
        RECT 40.2 5.535 40.37 5.705 ;
        RECT 41.18 4.345 41.35 4.515 ;
        RECT 41.64 4.345 41.81 4.515 ;
        RECT 42.1 4.345 42.27 4.515 ;
        RECT 42.56 4.345 42.73 4.515 ;
        RECT 43.02 4.345 43.19 4.515 ;
        RECT 43.48 4.345 43.65 4.515 ;
        RECT 43.94 4.345 44.11 4.515 ;
        RECT 44.4 4.345 44.57 4.515 ;
        RECT 44.86 4.345 45.03 4.515 ;
        RECT 45.32 4.345 45.49 4.515 ;
        RECT 45.78 4.345 45.95 4.515 ;
        RECT 46.24 4.345 46.41 4.515 ;
        RECT 46.7 4.345 46.87 4.515 ;
        RECT 47.16 4.345 47.33 4.515 ;
        RECT 47.62 4.345 47.79 4.515 ;
        RECT 48.08 4.345 48.25 4.515 ;
        RECT 51.885 5.535 52.055 5.705 ;
        RECT 51.885 4.165 52.055 4.335 ;
        RECT 52.585 5.54 52.755 5.71 ;
        RECT 52.585 4.16 52.755 4.33 ;
        RECT 53.575 5.54 53.745 5.71 ;
        RECT 53.575 4.16 53.745 4.33 ;
        RECT 57.42 5.535 57.59 5.705 ;
        RECT 58.4 4.345 58.57 4.515 ;
        RECT 58.86 4.345 59.03 4.515 ;
        RECT 59.32 4.345 59.49 4.515 ;
        RECT 59.78 4.345 59.95 4.515 ;
        RECT 60.24 4.345 60.41 4.515 ;
        RECT 60.7 4.345 60.87 4.515 ;
        RECT 61.16 4.345 61.33 4.515 ;
        RECT 61.62 4.345 61.79 4.515 ;
        RECT 62.08 4.345 62.25 4.515 ;
        RECT 62.54 4.345 62.71 4.515 ;
        RECT 63 4.345 63.17 4.515 ;
        RECT 63.46 4.345 63.63 4.515 ;
        RECT 63.92 4.345 64.09 4.515 ;
        RECT 64.38 4.345 64.55 4.515 ;
        RECT 64.84 4.345 65.01 4.515 ;
        RECT 65.3 4.345 65.47 4.515 ;
        RECT 69.105 5.535 69.275 5.705 ;
        RECT 69.105 4.165 69.275 4.335 ;
        RECT 69.805 5.54 69.975 5.71 ;
        RECT 69.805 4.16 69.975 4.33 ;
        RECT 70.795 5.54 70.965 5.71 ;
        RECT 70.795 4.16 70.965 4.33 ;
        RECT 74.64 5.535 74.81 5.705 ;
        RECT 75.62 4.345 75.79 4.515 ;
        RECT 76.08 4.345 76.25 4.515 ;
        RECT 76.54 4.345 76.71 4.515 ;
        RECT 77 4.345 77.17 4.515 ;
        RECT 77.46 4.345 77.63 4.515 ;
        RECT 77.92 4.345 78.09 4.515 ;
        RECT 78.38 4.345 78.55 4.515 ;
        RECT 78.84 4.345 79.01 4.515 ;
        RECT 79.3 4.345 79.47 4.515 ;
        RECT 79.76 4.345 79.93 4.515 ;
        RECT 80.22 4.345 80.39 4.515 ;
        RECT 80.68 4.345 80.85 4.515 ;
        RECT 81.14 4.345 81.31 4.515 ;
        RECT 81.6 4.345 81.77 4.515 ;
        RECT 82.06 4.345 82.23 4.515 ;
        RECT 82.52 4.345 82.69 4.515 ;
        RECT 86.325 5.535 86.495 5.705 ;
        RECT 86.325 4.165 86.495 4.335 ;
        RECT 87.025 5.54 87.195 5.71 ;
        RECT 87.025 4.16 87.195 4.33 ;
        RECT 88.015 5.54 88.185 5.71 ;
        RECT 88.015 4.16 88.185 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.86 5.79 78.19 6.12 ;
        RECT 77.39 5.805 78.19 6.105 ;
        RECT 60.64 5.79 60.97 6.12 ;
        RECT 60.17 5.805 60.97 6.105 ;
        RECT 43.42 5.79 43.75 6.12 ;
        RECT 42.95 5.805 43.75 6.105 ;
        RECT 26.2 5.79 26.53 6.12 ;
        RECT 25.73 5.805 26.53 6.105 ;
        RECT 8.98 5.79 9.31 6.12 ;
        RECT 8.51 5.805 9.31 6.105 ;
      LAYER li1 ;
        RECT 0 -1.295 88.91 0.305 ;
        RECT 87.935 -1.295 88.105 0.93 ;
        RECT 86.945 -1.295 87.115 0.93 ;
        RECT 84.205 -1.295 84.375 0.935 ;
        RECT 75.475 -1.295 83.13 1.795 ;
        RECT 82.37 -1.295 82.7 2.185 ;
        RECT 81.53 -1.295 81.86 2.185 ;
        RECT 79.7 -1.295 79.99 2.63 ;
        RECT 79.25 -1.295 79.52 2.605 ;
        RECT 78.34 -1.295 78.58 2.605 ;
        RECT 77.89 -1.295 78.13 2.605 ;
        RECT 76.95 -1.295 77.22 2.605 ;
        RECT 76.5 -1.295 76.73 2.615 ;
        RECT 75.62 -1.295 75.83 2.615 ;
        RECT 75.47 -1.295 83.13 1.635 ;
        RECT 70.715 -1.295 70.885 0.93 ;
        RECT 69.725 -1.295 69.895 0.93 ;
        RECT 66.985 -1.295 67.155 0.935 ;
        RECT 58.255 -1.295 65.91 1.795 ;
        RECT 65.15 -1.295 65.48 2.185 ;
        RECT 64.31 -1.295 64.64 2.185 ;
        RECT 62.48 -1.295 62.77 2.63 ;
        RECT 62.03 -1.295 62.3 2.605 ;
        RECT 61.12 -1.295 61.36 2.605 ;
        RECT 60.67 -1.295 60.91 2.605 ;
        RECT 59.73 -1.295 60 2.605 ;
        RECT 59.28 -1.295 59.51 2.615 ;
        RECT 58.4 -1.295 58.61 2.615 ;
        RECT 58.25 -1.295 65.91 1.635 ;
        RECT 53.495 -1.295 53.665 0.93 ;
        RECT 52.505 -1.295 52.675 0.93 ;
        RECT 49.765 -1.295 49.935 0.935 ;
        RECT 41.035 -1.295 48.69 1.795 ;
        RECT 47.93 -1.295 48.26 2.185 ;
        RECT 47.09 -1.295 47.42 2.185 ;
        RECT 45.26 -1.295 45.55 2.63 ;
        RECT 44.81 -1.295 45.08 2.605 ;
        RECT 43.9 -1.295 44.14 2.605 ;
        RECT 43.45 -1.295 43.69 2.605 ;
        RECT 42.51 -1.295 42.78 2.605 ;
        RECT 42.06 -1.295 42.29 2.615 ;
        RECT 41.18 -1.295 41.39 2.615 ;
        RECT 41.03 -1.295 48.69 1.635 ;
        RECT 36.275 -1.295 36.445 0.93 ;
        RECT 35.285 -1.295 35.455 0.93 ;
        RECT 32.545 -1.295 32.715 0.935 ;
        RECT 23.815 -1.295 31.47 1.795 ;
        RECT 30.71 -1.295 31.04 2.185 ;
        RECT 29.87 -1.295 30.2 2.185 ;
        RECT 28.04 -1.295 28.33 2.63 ;
        RECT 27.59 -1.295 27.86 2.605 ;
        RECT 26.68 -1.295 26.92 2.605 ;
        RECT 26.23 -1.295 26.47 2.605 ;
        RECT 25.29 -1.295 25.56 2.605 ;
        RECT 24.84 -1.295 25.07 2.615 ;
        RECT 23.96 -1.295 24.17 2.615 ;
        RECT 23.81 -1.295 31.47 1.635 ;
        RECT 19.055 -1.295 19.225 0.93 ;
        RECT 18.065 -1.295 18.235 0.93 ;
        RECT 15.325 -1.295 15.495 0.935 ;
        RECT 6.595 -1.295 14.25 1.795 ;
        RECT 13.49 -1.295 13.82 2.185 ;
        RECT 12.65 -1.295 12.98 2.185 ;
        RECT 10.82 -1.295 11.11 2.63 ;
        RECT 10.37 -1.295 10.64 2.605 ;
        RECT 9.46 -1.295 9.7 2.605 ;
        RECT 9.01 -1.295 9.25 2.605 ;
        RECT 8.07 -1.295 8.34 2.605 ;
        RECT 7.62 -1.295 7.85 2.615 ;
        RECT 6.74 -1.295 6.95 2.615 ;
        RECT 6.59 -1.295 14.25 1.635 ;
        RECT -0.015 9.565 88.91 11.165 ;
        RECT 87.935 8.94 88.105 11.165 ;
        RECT 86.945 8.94 87.115 11.165 ;
        RECT 84.205 8.935 84.375 11.165 ;
        RECT 75.475 9.56 82.945 11.165 ;
        RECT 75.475 7.065 82.835 11.165 ;
        RECT 81.98 6.265 82.29 11.165 ;
        RECT 80.6 6.265 80.91 11.165 ;
        RECT 78.33 5.825 78.665 6.095 ;
        RECT 78.32 6.265 78.63 11.165 ;
        RECT 77.94 5.875 78.665 6.045 ;
        RECT 77.95 5.875 78.12 11.165 ;
        RECT 76.02 6.265 76.33 11.165 ;
        RECT 72.52 8.935 72.69 11.165 ;
        RECT 70.715 8.94 70.885 11.165 ;
        RECT 69.725 8.94 69.895 11.165 ;
        RECT 66.985 8.935 67.155 11.165 ;
        RECT 58.255 9.56 65.725 11.165 ;
        RECT 58.255 7.065 65.615 11.165 ;
        RECT 64.76 6.265 65.07 11.165 ;
        RECT 63.38 6.265 63.69 11.165 ;
        RECT 61.11 5.825 61.445 6.095 ;
        RECT 61.1 6.265 61.41 11.165 ;
        RECT 60.72 5.875 61.445 6.045 ;
        RECT 60.73 5.875 60.9 11.165 ;
        RECT 58.8 6.265 59.11 11.165 ;
        RECT 55.3 8.935 55.47 11.165 ;
        RECT 53.495 8.94 53.665 11.165 ;
        RECT 52.505 8.94 52.675 11.165 ;
        RECT 49.765 8.935 49.935 11.165 ;
        RECT 41.035 9.56 48.505 11.165 ;
        RECT 41.035 7.065 48.395 11.165 ;
        RECT 47.54 6.265 47.85 11.165 ;
        RECT 46.16 6.265 46.47 11.165 ;
        RECT 43.89 5.825 44.225 6.095 ;
        RECT 43.88 6.265 44.19 11.165 ;
        RECT 43.5 5.875 44.225 6.045 ;
        RECT 43.51 5.875 43.68 11.165 ;
        RECT 41.58 6.265 41.89 11.165 ;
        RECT 38.08 8.935 38.25 11.165 ;
        RECT 36.275 8.94 36.445 11.165 ;
        RECT 35.285 8.94 35.455 11.165 ;
        RECT 32.545 8.935 32.715 11.165 ;
        RECT 23.815 9.56 31.285 11.165 ;
        RECT 23.815 7.065 31.175 11.165 ;
        RECT 30.32 6.265 30.63 11.165 ;
        RECT 28.94 6.265 29.25 11.165 ;
        RECT 26.67 5.825 27.005 6.095 ;
        RECT 26.66 6.265 26.97 11.165 ;
        RECT 26.28 5.875 27.005 6.045 ;
        RECT 26.29 5.875 26.46 11.165 ;
        RECT 24.36 6.265 24.67 11.165 ;
        RECT 20.86 8.935 21.03 11.165 ;
        RECT 19.055 8.94 19.225 11.165 ;
        RECT 18.065 8.94 18.235 11.165 ;
        RECT 15.325 8.935 15.495 11.165 ;
        RECT 6.595 9.56 14.065 11.165 ;
        RECT 6.595 7.065 13.955 11.165 ;
        RECT 13.1 6.265 13.41 11.165 ;
        RECT 11.72 6.265 12.03 11.165 ;
        RECT 9.45 5.825 9.785 6.095 ;
        RECT 9.44 6.265 9.75 11.165 ;
        RECT 9.06 5.875 9.785 6.045 ;
        RECT 9.07 5.875 9.24 11.165 ;
        RECT 7.14 6.265 7.45 11.165 ;
        RECT 3.64 8.935 3.81 11.165 ;
        RECT 0.23 8.935 0.4 11.165 ;
        RECT 76.03 5.825 76.365 6.095 ;
        RECT 75.56 5.875 76.365 6.045 ;
        RECT 73.525 7.065 73.695 9.015 ;
        RECT 73.47 8.845 73.64 9.295 ;
        RECT 73.47 6.005 73.64 7.235 ;
        RECT 58.81 5.825 59.145 6.095 ;
        RECT 58.34 5.875 59.145 6.045 ;
        RECT 56.305 7.065 56.475 9.015 ;
        RECT 56.25 8.845 56.42 9.295 ;
        RECT 56.25 6.005 56.42 7.235 ;
        RECT 41.59 5.825 41.925 6.095 ;
        RECT 41.12 5.875 41.925 6.045 ;
        RECT 39.085 7.065 39.255 9.015 ;
        RECT 39.03 8.845 39.2 9.295 ;
        RECT 39.03 6.005 39.2 7.235 ;
        RECT 24.37 5.825 24.705 6.095 ;
        RECT 23.9 5.875 24.705 6.045 ;
        RECT 21.865 7.065 22.035 9.015 ;
        RECT 21.81 8.845 21.98 9.295 ;
        RECT 21.81 6.005 21.98 7.235 ;
        RECT 7.15 5.825 7.485 6.095 ;
        RECT 6.68 5.875 7.485 6.045 ;
        RECT 4.645 7.065 4.815 9.015 ;
        RECT 4.59 8.845 4.76 9.295 ;
        RECT 4.59 6.005 4.76 7.235 ;
      LAYER met2 ;
        RECT 77.885 5.77 78.165 6.14 ;
        RECT 60.665 5.77 60.945 6.14 ;
        RECT 43.445 5.77 43.725 6.14 ;
        RECT 26.225 5.77 26.505 6.14 ;
        RECT 9.005 5.77 9.285 6.14 ;
      LAYER met1 ;
        RECT 0 -1.295 88.91 0.305 ;
        RECT 75.475 -1.295 83.13 1.795 ;
        RECT 75.475 -1.295 82.835 1.95 ;
        RECT 75.47 -1.295 83.13 1.635 ;
        RECT 58.255 -1.295 65.91 1.795 ;
        RECT 58.255 -1.295 65.615 1.95 ;
        RECT 58.25 -1.295 65.91 1.635 ;
        RECT 41.035 -1.295 48.69 1.795 ;
        RECT 41.035 -1.295 48.395 1.95 ;
        RECT 41.03 -1.295 48.69 1.635 ;
        RECT 23.815 -1.295 31.47 1.795 ;
        RECT 23.815 -1.295 31.175 1.95 ;
        RECT 23.81 -1.295 31.47 1.635 ;
        RECT 6.595 -1.295 14.25 1.795 ;
        RECT 6.595 -1.295 13.955 1.95 ;
        RECT 6.59 -1.295 14.25 1.635 ;
        RECT -0.015 9.565 88.91 11.165 ;
        RECT 75.475 9.56 82.945 11.165 ;
        RECT 75.475 6.91 82.835 11.165 ;
        RECT 73.465 7.275 73.755 7.505 ;
        RECT 73.065 7.305 73.755 7.475 ;
        RECT 73.065 7.305 73.235 11.165 ;
        RECT 58.255 9.56 65.725 11.165 ;
        RECT 58.255 6.91 65.615 11.165 ;
        RECT 56.245 7.275 56.535 7.505 ;
        RECT 55.845 7.305 56.535 7.475 ;
        RECT 55.845 7.305 56.015 11.165 ;
        RECT 41.035 9.56 48.505 11.165 ;
        RECT 41.035 6.91 48.395 11.165 ;
        RECT 39.025 7.275 39.315 7.505 ;
        RECT 38.625 7.305 39.315 7.475 ;
        RECT 38.625 7.305 38.795 11.165 ;
        RECT 23.815 9.56 31.285 11.165 ;
        RECT 23.815 6.91 31.175 11.165 ;
        RECT 21.805 7.275 22.095 7.505 ;
        RECT 21.405 7.305 22.095 7.475 ;
        RECT 21.405 7.305 21.575 11.165 ;
        RECT 6.595 9.56 14.065 11.165 ;
        RECT 6.595 6.91 13.955 11.165 ;
        RECT 4.585 7.275 4.875 7.505 ;
        RECT 4.185 7.305 4.875 7.475 ;
        RECT 4.185 7.305 4.355 11.165 ;
        RECT 77.865 5.83 78.185 6.09 ;
        RECT 75.5 5.89 78.185 6.03 ;
        RECT 75.5 5.845 75.79 6.075 ;
        RECT 60.645 5.83 60.965 6.09 ;
        RECT 58.28 5.89 60.965 6.03 ;
        RECT 58.28 5.845 58.57 6.075 ;
        RECT 43.425 5.83 43.745 6.09 ;
        RECT 41.06 5.89 43.745 6.03 ;
        RECT 41.06 5.845 41.35 6.075 ;
        RECT 26.205 5.83 26.525 6.09 ;
        RECT 23.84 5.89 26.525 6.03 ;
        RECT 23.84 5.845 24.13 6.075 ;
        RECT 8.985 5.83 9.305 6.09 ;
        RECT 6.62 5.89 9.305 6.03 ;
        RECT 6.62 5.845 6.91 6.075 ;
      LAYER via2 ;
        RECT 9.045 5.855 9.245 6.055 ;
        RECT 26.265 5.855 26.465 6.055 ;
        RECT 43.485 5.855 43.685 6.055 ;
        RECT 60.705 5.855 60.905 6.055 ;
        RECT 77.925 5.855 78.125 6.055 ;
      LAYER via1 ;
        RECT 9.07 5.885 9.22 6.035 ;
        RECT 26.29 5.885 26.44 6.035 ;
        RECT 43.51 5.885 43.66 6.035 ;
        RECT 60.73 5.885 60.88 6.035 ;
        RECT 77.95 5.885 78.1 6.035 ;
      LAYER mcon ;
        RECT 0.31 9.595 0.48 9.765 ;
        RECT 0.99 9.595 1.16 9.765 ;
        RECT 1.67 9.595 1.84 9.765 ;
        RECT 2.35 9.595 2.52 9.765 ;
        RECT 3.72 9.595 3.89 9.765 ;
        RECT 4.4 9.595 4.57 9.765 ;
        RECT 4.645 7.305 4.815 7.475 ;
        RECT 5.08 9.595 5.25 9.765 ;
        RECT 5.76 9.595 5.93 9.765 ;
        RECT 6.68 5.875 6.85 6.045 ;
        RECT 6.74 7.065 6.91 7.235 ;
        RECT 6.74 1.625 6.91 1.795 ;
        RECT 7.2 7.065 7.37 7.235 ;
        RECT 7.2 1.625 7.37 1.795 ;
        RECT 7.66 7.065 7.83 7.235 ;
        RECT 7.66 1.625 7.83 1.795 ;
        RECT 8.12 7.065 8.29 7.235 ;
        RECT 8.12 1.625 8.29 1.795 ;
        RECT 8.58 7.065 8.75 7.235 ;
        RECT 8.58 1.625 8.75 1.795 ;
        RECT 9.04 7.065 9.21 7.235 ;
        RECT 9.04 1.625 9.21 1.795 ;
        RECT 9.06 5.875 9.23 6.045 ;
        RECT 9.5 7.065 9.67 7.235 ;
        RECT 9.5 1.625 9.67 1.795 ;
        RECT 9.96 7.065 10.13 7.235 ;
        RECT 9.96 1.625 10.13 1.795 ;
        RECT 10.42 7.065 10.59 7.235 ;
        RECT 10.42 1.625 10.59 1.795 ;
        RECT 10.88 7.065 11.05 7.235 ;
        RECT 10.88 1.625 11.05 1.795 ;
        RECT 11.34 7.065 11.51 7.235 ;
        RECT 11.34 1.625 11.51 1.795 ;
        RECT 11.8 7.065 11.97 7.235 ;
        RECT 11.8 1.625 11.97 1.795 ;
        RECT 12.26 7.065 12.43 7.235 ;
        RECT 12.26 1.625 12.43 1.795 ;
        RECT 12.72 7.065 12.89 7.235 ;
        RECT 12.72 1.625 12.89 1.795 ;
        RECT 13.18 7.065 13.35 7.235 ;
        RECT 13.18 1.625 13.35 1.795 ;
        RECT 13.64 7.065 13.81 7.235 ;
        RECT 13.64 1.625 13.81 1.795 ;
        RECT 15.405 9.595 15.575 9.765 ;
        RECT 15.405 0.105 15.575 0.275 ;
        RECT 16.085 9.595 16.255 9.765 ;
        RECT 16.085 0.105 16.255 0.275 ;
        RECT 16.765 9.595 16.935 9.765 ;
        RECT 16.765 0.105 16.935 0.275 ;
        RECT 17.445 9.595 17.615 9.765 ;
        RECT 17.445 0.105 17.615 0.275 ;
        RECT 18.145 9.6 18.315 9.77 ;
        RECT 18.145 0.1 18.315 0.27 ;
        RECT 19.135 9.6 19.305 9.77 ;
        RECT 19.135 0.1 19.305 0.27 ;
        RECT 20.94 9.595 21.11 9.765 ;
        RECT 21.62 9.595 21.79 9.765 ;
        RECT 21.865 7.305 22.035 7.475 ;
        RECT 22.3 9.595 22.47 9.765 ;
        RECT 22.98 9.595 23.15 9.765 ;
        RECT 23.9 5.875 24.07 6.045 ;
        RECT 23.96 7.065 24.13 7.235 ;
        RECT 23.96 1.625 24.13 1.795 ;
        RECT 24.42 7.065 24.59 7.235 ;
        RECT 24.42 1.625 24.59 1.795 ;
        RECT 24.88 7.065 25.05 7.235 ;
        RECT 24.88 1.625 25.05 1.795 ;
        RECT 25.34 7.065 25.51 7.235 ;
        RECT 25.34 1.625 25.51 1.795 ;
        RECT 25.8 7.065 25.97 7.235 ;
        RECT 25.8 1.625 25.97 1.795 ;
        RECT 26.26 7.065 26.43 7.235 ;
        RECT 26.26 1.625 26.43 1.795 ;
        RECT 26.28 5.875 26.45 6.045 ;
        RECT 26.72 7.065 26.89 7.235 ;
        RECT 26.72 1.625 26.89 1.795 ;
        RECT 27.18 7.065 27.35 7.235 ;
        RECT 27.18 1.625 27.35 1.795 ;
        RECT 27.64 7.065 27.81 7.235 ;
        RECT 27.64 1.625 27.81 1.795 ;
        RECT 28.1 7.065 28.27 7.235 ;
        RECT 28.1 1.625 28.27 1.795 ;
        RECT 28.56 7.065 28.73 7.235 ;
        RECT 28.56 1.625 28.73 1.795 ;
        RECT 29.02 7.065 29.19 7.235 ;
        RECT 29.02 1.625 29.19 1.795 ;
        RECT 29.48 7.065 29.65 7.235 ;
        RECT 29.48 1.625 29.65 1.795 ;
        RECT 29.94 7.065 30.11 7.235 ;
        RECT 29.94 1.625 30.11 1.795 ;
        RECT 30.4 7.065 30.57 7.235 ;
        RECT 30.4 1.625 30.57 1.795 ;
        RECT 30.86 7.065 31.03 7.235 ;
        RECT 30.86 1.625 31.03 1.795 ;
        RECT 32.625 9.595 32.795 9.765 ;
        RECT 32.625 0.105 32.795 0.275 ;
        RECT 33.305 9.595 33.475 9.765 ;
        RECT 33.305 0.105 33.475 0.275 ;
        RECT 33.985 9.595 34.155 9.765 ;
        RECT 33.985 0.105 34.155 0.275 ;
        RECT 34.665 9.595 34.835 9.765 ;
        RECT 34.665 0.105 34.835 0.275 ;
        RECT 35.365 9.6 35.535 9.77 ;
        RECT 35.365 0.1 35.535 0.27 ;
        RECT 36.355 9.6 36.525 9.77 ;
        RECT 36.355 0.1 36.525 0.27 ;
        RECT 38.16 9.595 38.33 9.765 ;
        RECT 38.84 9.595 39.01 9.765 ;
        RECT 39.085 7.305 39.255 7.475 ;
        RECT 39.52 9.595 39.69 9.765 ;
        RECT 40.2 9.595 40.37 9.765 ;
        RECT 41.12 5.875 41.29 6.045 ;
        RECT 41.18 7.065 41.35 7.235 ;
        RECT 41.18 1.625 41.35 1.795 ;
        RECT 41.64 7.065 41.81 7.235 ;
        RECT 41.64 1.625 41.81 1.795 ;
        RECT 42.1 7.065 42.27 7.235 ;
        RECT 42.1 1.625 42.27 1.795 ;
        RECT 42.56 7.065 42.73 7.235 ;
        RECT 42.56 1.625 42.73 1.795 ;
        RECT 43.02 7.065 43.19 7.235 ;
        RECT 43.02 1.625 43.19 1.795 ;
        RECT 43.48 7.065 43.65 7.235 ;
        RECT 43.48 1.625 43.65 1.795 ;
        RECT 43.5 5.875 43.67 6.045 ;
        RECT 43.94 7.065 44.11 7.235 ;
        RECT 43.94 1.625 44.11 1.795 ;
        RECT 44.4 7.065 44.57 7.235 ;
        RECT 44.4 1.625 44.57 1.795 ;
        RECT 44.86 7.065 45.03 7.235 ;
        RECT 44.86 1.625 45.03 1.795 ;
        RECT 45.32 7.065 45.49 7.235 ;
        RECT 45.32 1.625 45.49 1.795 ;
        RECT 45.78 7.065 45.95 7.235 ;
        RECT 45.78 1.625 45.95 1.795 ;
        RECT 46.24 7.065 46.41 7.235 ;
        RECT 46.24 1.625 46.41 1.795 ;
        RECT 46.7 7.065 46.87 7.235 ;
        RECT 46.7 1.625 46.87 1.795 ;
        RECT 47.16 7.065 47.33 7.235 ;
        RECT 47.16 1.625 47.33 1.795 ;
        RECT 47.62 7.065 47.79 7.235 ;
        RECT 47.62 1.625 47.79 1.795 ;
        RECT 48.08 7.065 48.25 7.235 ;
        RECT 48.08 1.625 48.25 1.795 ;
        RECT 49.845 9.595 50.015 9.765 ;
        RECT 49.845 0.105 50.015 0.275 ;
        RECT 50.525 9.595 50.695 9.765 ;
        RECT 50.525 0.105 50.695 0.275 ;
        RECT 51.205 9.595 51.375 9.765 ;
        RECT 51.205 0.105 51.375 0.275 ;
        RECT 51.885 9.595 52.055 9.765 ;
        RECT 51.885 0.105 52.055 0.275 ;
        RECT 52.585 9.6 52.755 9.77 ;
        RECT 52.585 0.1 52.755 0.27 ;
        RECT 53.575 9.6 53.745 9.77 ;
        RECT 53.575 0.1 53.745 0.27 ;
        RECT 55.38 9.595 55.55 9.765 ;
        RECT 56.06 9.595 56.23 9.765 ;
        RECT 56.305 7.305 56.475 7.475 ;
        RECT 56.74 9.595 56.91 9.765 ;
        RECT 57.42 9.595 57.59 9.765 ;
        RECT 58.34 5.875 58.51 6.045 ;
        RECT 58.4 7.065 58.57 7.235 ;
        RECT 58.4 1.625 58.57 1.795 ;
        RECT 58.86 7.065 59.03 7.235 ;
        RECT 58.86 1.625 59.03 1.795 ;
        RECT 59.32 7.065 59.49 7.235 ;
        RECT 59.32 1.625 59.49 1.795 ;
        RECT 59.78 7.065 59.95 7.235 ;
        RECT 59.78 1.625 59.95 1.795 ;
        RECT 60.24 7.065 60.41 7.235 ;
        RECT 60.24 1.625 60.41 1.795 ;
        RECT 60.7 7.065 60.87 7.235 ;
        RECT 60.7 1.625 60.87 1.795 ;
        RECT 60.72 5.875 60.89 6.045 ;
        RECT 61.16 7.065 61.33 7.235 ;
        RECT 61.16 1.625 61.33 1.795 ;
        RECT 61.62 7.065 61.79 7.235 ;
        RECT 61.62 1.625 61.79 1.795 ;
        RECT 62.08 7.065 62.25 7.235 ;
        RECT 62.08 1.625 62.25 1.795 ;
        RECT 62.54 7.065 62.71 7.235 ;
        RECT 62.54 1.625 62.71 1.795 ;
        RECT 63 7.065 63.17 7.235 ;
        RECT 63 1.625 63.17 1.795 ;
        RECT 63.46 7.065 63.63 7.235 ;
        RECT 63.46 1.625 63.63 1.795 ;
        RECT 63.92 7.065 64.09 7.235 ;
        RECT 63.92 1.625 64.09 1.795 ;
        RECT 64.38 7.065 64.55 7.235 ;
        RECT 64.38 1.625 64.55 1.795 ;
        RECT 64.84 7.065 65.01 7.235 ;
        RECT 64.84 1.625 65.01 1.795 ;
        RECT 65.3 7.065 65.47 7.235 ;
        RECT 65.3 1.625 65.47 1.795 ;
        RECT 67.065 9.595 67.235 9.765 ;
        RECT 67.065 0.105 67.235 0.275 ;
        RECT 67.745 9.595 67.915 9.765 ;
        RECT 67.745 0.105 67.915 0.275 ;
        RECT 68.425 9.595 68.595 9.765 ;
        RECT 68.425 0.105 68.595 0.275 ;
        RECT 69.105 9.595 69.275 9.765 ;
        RECT 69.105 0.105 69.275 0.275 ;
        RECT 69.805 9.6 69.975 9.77 ;
        RECT 69.805 0.1 69.975 0.27 ;
        RECT 70.795 9.6 70.965 9.77 ;
        RECT 70.795 0.1 70.965 0.27 ;
        RECT 72.6 9.595 72.77 9.765 ;
        RECT 73.28 9.595 73.45 9.765 ;
        RECT 73.525 7.305 73.695 7.475 ;
        RECT 73.96 9.595 74.13 9.765 ;
        RECT 74.64 9.595 74.81 9.765 ;
        RECT 75.56 5.875 75.73 6.045 ;
        RECT 75.62 7.065 75.79 7.235 ;
        RECT 75.62 1.625 75.79 1.795 ;
        RECT 76.08 7.065 76.25 7.235 ;
        RECT 76.08 1.625 76.25 1.795 ;
        RECT 76.54 7.065 76.71 7.235 ;
        RECT 76.54 1.625 76.71 1.795 ;
        RECT 77 7.065 77.17 7.235 ;
        RECT 77 1.625 77.17 1.795 ;
        RECT 77.46 7.065 77.63 7.235 ;
        RECT 77.46 1.625 77.63 1.795 ;
        RECT 77.92 7.065 78.09 7.235 ;
        RECT 77.92 1.625 78.09 1.795 ;
        RECT 77.94 5.875 78.11 6.045 ;
        RECT 78.38 7.065 78.55 7.235 ;
        RECT 78.38 1.625 78.55 1.795 ;
        RECT 78.84 7.065 79.01 7.235 ;
        RECT 78.84 1.625 79.01 1.795 ;
        RECT 79.3 7.065 79.47 7.235 ;
        RECT 79.3 1.625 79.47 1.795 ;
        RECT 79.76 7.065 79.93 7.235 ;
        RECT 79.76 1.625 79.93 1.795 ;
        RECT 80.22 7.065 80.39 7.235 ;
        RECT 80.22 1.625 80.39 1.795 ;
        RECT 80.68 7.065 80.85 7.235 ;
        RECT 80.68 1.625 80.85 1.795 ;
        RECT 81.14 7.065 81.31 7.235 ;
        RECT 81.14 1.625 81.31 1.795 ;
        RECT 81.6 7.065 81.77 7.235 ;
        RECT 81.6 1.625 81.77 1.795 ;
        RECT 82.06 7.065 82.23 7.235 ;
        RECT 82.06 1.625 82.23 1.795 ;
        RECT 82.52 7.065 82.69 7.235 ;
        RECT 82.52 1.625 82.69 1.795 ;
        RECT 84.285 9.595 84.455 9.765 ;
        RECT 84.285 0.105 84.455 0.275 ;
        RECT 84.965 9.595 85.135 9.765 ;
        RECT 84.965 0.105 85.135 0.275 ;
        RECT 85.645 9.595 85.815 9.765 ;
        RECT 85.645 0.105 85.815 0.275 ;
        RECT 86.325 9.595 86.495 9.765 ;
        RECT 86.325 0.105 86.495 0.275 ;
        RECT 87.025 9.6 87.195 9.77 ;
        RECT 87.025 0.1 87.195 0.27 ;
        RECT 88.015 9.6 88.185 9.77 ;
        RECT 88.015 0.1 88.185 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 73.805 7.99 74.175 8.36 ;
      RECT 73.805 8.025 80.955 8.325 ;
      RECT 80.655 5.805 80.955 8.325 ;
      RECT 79.6 5.785 79.9 8.325 ;
      RECT 78.57 6.48 78.87 8.325 ;
      RECT 78.54 6.48 78.87 6.81 ;
      RECT 78.07 6.495 78.87 6.795 ;
      RECT 78.45 6.455 78.75 6.795 ;
      RECT 80.58 5.805 80.955 6.17 ;
      RECT 80.645 5.765 80.945 6.17 ;
      RECT 79.56 5.785 79.9 6.135 ;
      RECT 79.575 5.745 79.875 6.135 ;
      RECT 79.55 5.79 79.9 6.12 ;
      RECT 80.58 5.805 81.39 6.105 ;
      RECT 79.08 5.805 79.9 6.105 ;
      RECT 80.59 5.79 80.945 6.17 ;
      RECT 80.24 3.755 80.57 4.085 ;
      RECT 80.24 3.77 81.04 4.07 ;
      RECT 80.255 3.725 80.555 4.085 ;
      RECT 79.9 3.075 80.23 3.405 ;
      RECT 79.9 3.09 80.7 3.39 ;
      RECT 79.985 3.065 80.285 3.39 ;
      RECT 79.22 4.155 79.55 4.485 ;
      RECT 77.18 4.155 77.51 4.485 ;
      RECT 77.18 4.17 79.55 4.47 ;
      RECT 78.87 3.415 79.2 3.745 ;
      RECT 78.41 3.43 79.21 3.73 ;
      RECT 78.54 2.225 78.87 2.555 ;
      RECT 78.07 2.24 78.87 2.54 ;
      RECT 78.53 2.235 78.87 2.54 ;
      RECT 56.585 7.99 56.955 8.36 ;
      RECT 56.585 8.025 63.735 8.325 ;
      RECT 63.435 5.805 63.735 8.325 ;
      RECT 62.38 5.785 62.68 8.325 ;
      RECT 61.35 6.48 61.65 8.325 ;
      RECT 61.32 6.48 61.65 6.81 ;
      RECT 60.85 6.495 61.65 6.795 ;
      RECT 61.23 6.455 61.53 6.795 ;
      RECT 63.36 5.805 63.735 6.17 ;
      RECT 63.425 5.765 63.725 6.17 ;
      RECT 62.34 5.785 62.68 6.135 ;
      RECT 62.355 5.745 62.655 6.135 ;
      RECT 62.33 5.79 62.68 6.12 ;
      RECT 63.36 5.805 64.17 6.105 ;
      RECT 61.86 5.805 62.68 6.105 ;
      RECT 63.37 5.79 63.725 6.17 ;
      RECT 63.02 3.755 63.35 4.085 ;
      RECT 63.02 3.77 63.82 4.07 ;
      RECT 63.035 3.725 63.335 4.085 ;
      RECT 62.68 3.075 63.01 3.405 ;
      RECT 62.68 3.09 63.48 3.39 ;
      RECT 62.765 3.065 63.065 3.39 ;
      RECT 62 4.155 62.33 4.485 ;
      RECT 59.96 4.155 60.29 4.485 ;
      RECT 59.96 4.17 62.33 4.47 ;
      RECT 61.65 3.415 61.98 3.745 ;
      RECT 61.19 3.43 61.99 3.73 ;
      RECT 61.32 2.225 61.65 2.555 ;
      RECT 60.85 2.24 61.65 2.54 ;
      RECT 61.31 2.235 61.65 2.54 ;
      RECT 39.365 7.99 39.735 8.36 ;
      RECT 39.365 8.025 46.515 8.325 ;
      RECT 46.215 5.805 46.515 8.325 ;
      RECT 45.16 5.785 45.46 8.325 ;
      RECT 44.13 6.48 44.43 8.325 ;
      RECT 44.1 6.48 44.43 6.81 ;
      RECT 43.63 6.495 44.43 6.795 ;
      RECT 44.01 6.455 44.31 6.795 ;
      RECT 46.14 5.805 46.515 6.17 ;
      RECT 46.205 5.765 46.505 6.17 ;
      RECT 45.12 5.785 45.46 6.135 ;
      RECT 45.135 5.745 45.435 6.135 ;
      RECT 45.11 5.79 45.46 6.12 ;
      RECT 46.14 5.805 46.95 6.105 ;
      RECT 44.64 5.805 45.46 6.105 ;
      RECT 46.15 5.79 46.505 6.17 ;
      RECT 45.8 3.755 46.13 4.085 ;
      RECT 45.8 3.77 46.6 4.07 ;
      RECT 45.815 3.725 46.115 4.085 ;
      RECT 45.46 3.075 45.79 3.405 ;
      RECT 45.46 3.09 46.26 3.39 ;
      RECT 45.545 3.065 45.845 3.39 ;
      RECT 44.78 4.155 45.11 4.485 ;
      RECT 42.74 4.155 43.07 4.485 ;
      RECT 42.74 4.17 45.11 4.47 ;
      RECT 44.43 3.415 44.76 3.745 ;
      RECT 43.97 3.43 44.77 3.73 ;
      RECT 44.1 2.225 44.43 2.555 ;
      RECT 43.63 2.24 44.43 2.54 ;
      RECT 44.09 2.235 44.43 2.54 ;
      RECT 22.145 7.99 22.515 8.36 ;
      RECT 22.145 8.025 29.295 8.325 ;
      RECT 28.995 5.805 29.295 8.325 ;
      RECT 27.94 5.785 28.24 8.325 ;
      RECT 26.91 6.48 27.21 8.325 ;
      RECT 26.88 6.48 27.21 6.81 ;
      RECT 26.41 6.495 27.21 6.795 ;
      RECT 26.79 6.455 27.09 6.795 ;
      RECT 28.92 5.805 29.295 6.17 ;
      RECT 28.985 5.765 29.285 6.17 ;
      RECT 27.9 5.785 28.24 6.135 ;
      RECT 27.915 5.745 28.215 6.135 ;
      RECT 27.89 5.79 28.24 6.12 ;
      RECT 28.92 5.805 29.73 6.105 ;
      RECT 27.42 5.805 28.24 6.105 ;
      RECT 28.93 5.79 29.285 6.17 ;
      RECT 28.58 3.755 28.91 4.085 ;
      RECT 28.58 3.77 29.38 4.07 ;
      RECT 28.595 3.725 28.895 4.085 ;
      RECT 28.24 3.075 28.57 3.405 ;
      RECT 28.24 3.09 29.04 3.39 ;
      RECT 28.325 3.065 28.625 3.39 ;
      RECT 27.56 4.155 27.89 4.485 ;
      RECT 25.52 4.155 25.85 4.485 ;
      RECT 25.52 4.17 27.89 4.47 ;
      RECT 27.21 3.415 27.54 3.745 ;
      RECT 26.75 3.43 27.55 3.73 ;
      RECT 26.88 2.225 27.21 2.555 ;
      RECT 26.41 2.24 27.21 2.54 ;
      RECT 26.87 2.235 27.21 2.54 ;
      RECT 4.925 7.99 5.295 8.36 ;
      RECT 4.925 8.025 12.075 8.325 ;
      RECT 11.775 5.805 12.075 8.325 ;
      RECT 10.72 5.785 11.02 8.325 ;
      RECT 9.69 6.48 9.99 8.325 ;
      RECT 9.66 6.48 9.99 6.81 ;
      RECT 9.19 6.495 9.99 6.795 ;
      RECT 9.57 6.455 9.87 6.795 ;
      RECT 11.7 5.805 12.075 6.17 ;
      RECT 11.765 5.765 12.065 6.17 ;
      RECT 10.68 5.785 11.02 6.135 ;
      RECT 10.695 5.745 10.995 6.135 ;
      RECT 10.67 5.79 11.02 6.12 ;
      RECT 11.7 5.805 12.51 6.105 ;
      RECT 10.2 5.805 11.02 6.105 ;
      RECT 11.71 5.79 12.065 6.17 ;
      RECT 11.36 3.755 11.69 4.085 ;
      RECT 11.36 3.77 12.16 4.07 ;
      RECT 11.375 3.725 11.675 4.085 ;
      RECT 11.02 3.075 11.35 3.405 ;
      RECT 11.02 3.09 11.82 3.39 ;
      RECT 11.105 3.065 11.405 3.39 ;
      RECT 10.34 4.155 10.67 4.485 ;
      RECT 8.3 4.155 8.63 4.485 ;
      RECT 8.3 4.17 10.67 4.47 ;
      RECT 9.99 3.415 10.32 3.745 ;
      RECT 9.53 3.43 10.33 3.73 ;
      RECT 9.66 2.225 9.99 2.555 ;
      RECT 9.19 2.24 9.99 2.54 ;
      RECT 9.65 2.235 9.99 2.54 ;
    LAYER via2 ;
      RECT 80.655 5.855 80.855 6.055 ;
      RECT 80.305 3.82 80.505 4.02 ;
      RECT 79.965 3.14 80.165 3.34 ;
      RECT 79.615 5.855 79.815 6.055 ;
      RECT 79.285 4.22 79.485 4.42 ;
      RECT 78.935 3.48 79.135 3.68 ;
      RECT 78.605 2.29 78.805 2.49 ;
      RECT 78.605 6.545 78.805 6.745 ;
      RECT 77.245 4.22 77.445 4.42 ;
      RECT 73.89 8.075 74.09 8.275 ;
      RECT 63.435 5.855 63.635 6.055 ;
      RECT 63.085 3.82 63.285 4.02 ;
      RECT 62.745 3.14 62.945 3.34 ;
      RECT 62.395 5.855 62.595 6.055 ;
      RECT 62.065 4.22 62.265 4.42 ;
      RECT 61.715 3.48 61.915 3.68 ;
      RECT 61.385 2.29 61.585 2.49 ;
      RECT 61.385 6.545 61.585 6.745 ;
      RECT 60.025 4.22 60.225 4.42 ;
      RECT 56.67 8.075 56.87 8.275 ;
      RECT 46.215 5.855 46.415 6.055 ;
      RECT 45.865 3.82 46.065 4.02 ;
      RECT 45.525 3.14 45.725 3.34 ;
      RECT 45.175 5.855 45.375 6.055 ;
      RECT 44.845 4.22 45.045 4.42 ;
      RECT 44.495 3.48 44.695 3.68 ;
      RECT 44.165 2.29 44.365 2.49 ;
      RECT 44.165 6.545 44.365 6.745 ;
      RECT 42.805 4.22 43.005 4.42 ;
      RECT 39.45 8.075 39.65 8.275 ;
      RECT 28.995 5.855 29.195 6.055 ;
      RECT 28.645 3.82 28.845 4.02 ;
      RECT 28.305 3.14 28.505 3.34 ;
      RECT 27.955 5.855 28.155 6.055 ;
      RECT 27.625 4.22 27.825 4.42 ;
      RECT 27.275 3.48 27.475 3.68 ;
      RECT 26.945 2.29 27.145 2.49 ;
      RECT 26.945 6.545 27.145 6.745 ;
      RECT 25.585 4.22 25.785 4.42 ;
      RECT 22.23 8.075 22.43 8.275 ;
      RECT 11.775 5.855 11.975 6.055 ;
      RECT 11.425 3.82 11.625 4.02 ;
      RECT 11.085 3.14 11.285 3.34 ;
      RECT 10.735 5.855 10.935 6.055 ;
      RECT 10.405 4.22 10.605 4.42 ;
      RECT 10.055 3.48 10.255 3.68 ;
      RECT 9.725 2.29 9.925 2.49 ;
      RECT 9.725 6.545 9.925 6.745 ;
      RECT 8.365 4.22 8.565 4.42 ;
      RECT 5.01 8.075 5.21 8.275 ;
    LAYER met2 ;
      RECT 1.23 8.77 88.54 8.94 ;
      RECT 88.37 8.29 88.54 8.94 ;
      RECT 1.23 7.245 1.4 8.94 ;
      RECT 88.335 8.29 88.66 8.615 ;
      RECT 1.175 7.245 1.455 7.585 ;
      RECT 85.18 7.27 85.5 7.595 ;
      RECT 85.21 6.685 85.38 7.595 ;
      RECT 85.21 6.685 85.385 7.035 ;
      RECT 85.21 6.685 86.185 6.86 ;
      RECT 86.01 1.965 86.185 6.86 ;
      RECT 79.925 3.055 80.205 3.425 ;
      RECT 79.995 2.345 80.17 3.425 ;
      RECT 79.995 2.345 83.215 2.52 ;
      RECT 83.04 2.025 83.215 2.52 ;
      RECT 83.51 1.995 83.835 2.32 ;
      RECT 85.955 1.965 86.305 2.315 ;
      RECT 83.04 2.025 86.305 2.195 ;
      RECT 74.33 8.355 85.025 8.525 ;
      RECT 84.865 2.395 85.025 8.525 ;
      RECT 74.33 7.535 74.5 8.525 ;
      RECT 85.98 7.645 86.305 7.97 ;
      RECT 71.15 7.645 71.475 7.97 ;
      RECT 84.865 7.735 86.305 7.905 ;
      RECT 74.28 7.535 74.56 7.875 ;
      RECT 71.15 7.675 74.56 7.845 ;
      RECT 85.18 2.365 85.5 2.685 ;
      RECT 84.865 2.395 85.5 2.565 ;
      RECT 81.635 6.48 81.895 6.8 ;
      RECT 81.695 2.74 81.835 6.8 ;
      RECT 81.635 2.74 81.895 3.06 ;
      RECT 80.955 4.78 81.215 5.1 ;
      RECT 81.015 3.76 81.155 5.1 ;
      RECT 80.955 3.76 81.215 4.08 ;
      RECT 79.935 6.48 80.195 6.8 ;
      RECT 79.995 5.21 80.135 6.8 ;
      RECT 79.315 5.21 80.135 5.35 ;
      RECT 79.315 2.74 79.455 5.35 ;
      RECT 79.245 4.135 79.525 4.505 ;
      RECT 79.255 2.74 79.515 3.06 ;
      RECT 77.205 4.135 77.485 4.505 ;
      RECT 77.275 2.4 77.415 4.505 ;
      RECT 77.215 2.4 77.475 2.72 ;
      RECT 76.535 4.78 76.795 5.1 ;
      RECT 76.595 2.74 76.735 5.1 ;
      RECT 76.535 2.74 76.795 3.06 ;
      RECT 67.96 7.27 68.28 7.595 ;
      RECT 67.99 6.685 68.16 7.595 ;
      RECT 67.99 6.685 68.165 7.035 ;
      RECT 67.99 6.685 68.965 6.86 ;
      RECT 68.79 1.965 68.965 6.86 ;
      RECT 62.705 3.055 62.985 3.425 ;
      RECT 62.775 2.345 62.95 3.425 ;
      RECT 62.775 2.345 65.995 2.52 ;
      RECT 65.82 2.025 65.995 2.52 ;
      RECT 66.29 1.995 66.615 2.32 ;
      RECT 68.735 1.965 69.085 2.315 ;
      RECT 65.82 2.025 69.085 2.195 ;
      RECT 57.11 8.355 67.805 8.525 ;
      RECT 67.645 2.395 67.805 8.525 ;
      RECT 57.11 7.535 57.28 8.525 ;
      RECT 68.76 7.645 69.085 7.97 ;
      RECT 53.93 7.645 54.255 7.97 ;
      RECT 67.645 7.735 69.085 7.905 ;
      RECT 57.06 7.535 57.34 7.875 ;
      RECT 53.93 7.675 57.34 7.845 ;
      RECT 67.96 2.365 68.28 2.685 ;
      RECT 67.645 2.395 68.28 2.565 ;
      RECT 64.415 6.48 64.675 6.8 ;
      RECT 64.475 2.74 64.615 6.8 ;
      RECT 64.415 2.74 64.675 3.06 ;
      RECT 63.735 4.78 63.995 5.1 ;
      RECT 63.795 3.76 63.935 5.1 ;
      RECT 63.735 3.76 63.995 4.08 ;
      RECT 62.715 6.48 62.975 6.8 ;
      RECT 62.775 5.21 62.915 6.8 ;
      RECT 62.095 5.21 62.915 5.35 ;
      RECT 62.095 2.74 62.235 5.35 ;
      RECT 62.025 4.135 62.305 4.505 ;
      RECT 62.035 2.74 62.295 3.06 ;
      RECT 59.985 4.135 60.265 4.505 ;
      RECT 60.055 2.4 60.195 4.505 ;
      RECT 59.995 2.4 60.255 2.72 ;
      RECT 59.315 4.78 59.575 5.1 ;
      RECT 59.375 2.74 59.515 5.1 ;
      RECT 59.315 2.74 59.575 3.06 ;
      RECT 50.74 7.27 51.06 7.595 ;
      RECT 50.77 6.685 50.94 7.595 ;
      RECT 50.77 6.685 50.945 7.035 ;
      RECT 50.77 6.685 51.745 6.86 ;
      RECT 51.57 1.965 51.745 6.86 ;
      RECT 45.485 3.055 45.765 3.425 ;
      RECT 45.555 2.345 45.73 3.425 ;
      RECT 45.555 2.345 48.775 2.52 ;
      RECT 48.6 2.025 48.775 2.52 ;
      RECT 49.07 1.995 49.395 2.32 ;
      RECT 51.515 1.965 51.865 2.315 ;
      RECT 48.6 2.025 51.865 2.195 ;
      RECT 39.89 8.355 50.585 8.525 ;
      RECT 50.425 2.395 50.585 8.525 ;
      RECT 39.89 7.535 40.06 8.525 ;
      RECT 51.54 7.645 51.865 7.97 ;
      RECT 36.71 7.645 37.035 7.97 ;
      RECT 50.425 7.735 51.865 7.905 ;
      RECT 39.84 7.535 40.12 7.875 ;
      RECT 36.71 7.675 40.13 7.845 ;
      RECT 50.74 2.365 51.06 2.685 ;
      RECT 50.425 2.395 51.06 2.565 ;
      RECT 47.195 6.48 47.455 6.8 ;
      RECT 47.255 2.74 47.395 6.8 ;
      RECT 47.195 2.74 47.455 3.06 ;
      RECT 46.515 4.78 46.775 5.1 ;
      RECT 46.575 3.76 46.715 5.1 ;
      RECT 46.515 3.76 46.775 4.08 ;
      RECT 45.495 6.48 45.755 6.8 ;
      RECT 45.555 5.21 45.695 6.8 ;
      RECT 44.875 5.21 45.695 5.35 ;
      RECT 44.875 2.74 45.015 5.35 ;
      RECT 44.805 4.135 45.085 4.505 ;
      RECT 44.815 2.74 45.075 3.06 ;
      RECT 42.765 4.135 43.045 4.505 ;
      RECT 42.835 2.4 42.975 4.505 ;
      RECT 42.775 2.4 43.035 2.72 ;
      RECT 42.095 4.78 42.355 5.1 ;
      RECT 42.155 2.74 42.295 5.1 ;
      RECT 42.095 2.74 42.355 3.06 ;
      RECT 33.52 7.27 33.84 7.595 ;
      RECT 33.55 6.685 33.72 7.595 ;
      RECT 33.55 6.685 33.725 7.035 ;
      RECT 33.55 6.685 34.525 6.86 ;
      RECT 34.35 1.965 34.525 6.86 ;
      RECT 28.265 3.055 28.545 3.425 ;
      RECT 28.335 2.345 28.51 3.425 ;
      RECT 28.335 2.345 31.555 2.52 ;
      RECT 31.38 2.025 31.555 2.52 ;
      RECT 31.85 1.995 32.175 2.32 ;
      RECT 34.295 1.965 34.645 2.315 ;
      RECT 31.38 2.025 34.645 2.195 ;
      RECT 22.67 8.355 33.365 8.525 ;
      RECT 33.205 2.395 33.365 8.525 ;
      RECT 22.67 7.535 22.84 8.525 ;
      RECT 34.32 7.645 34.645 7.97 ;
      RECT 19.49 7.645 19.815 7.97 ;
      RECT 33.205 7.735 34.645 7.905 ;
      RECT 22.62 7.535 22.9 7.875 ;
      RECT 19.49 7.675 22.9 7.845 ;
      RECT 33.52 2.365 33.84 2.685 ;
      RECT 33.205 2.395 33.84 2.565 ;
      RECT 29.975 6.48 30.235 6.8 ;
      RECT 30.035 2.74 30.175 6.8 ;
      RECT 29.975 2.74 30.235 3.06 ;
      RECT 29.295 4.78 29.555 5.1 ;
      RECT 29.355 3.76 29.495 5.1 ;
      RECT 29.295 3.76 29.555 4.08 ;
      RECT 28.275 6.48 28.535 6.8 ;
      RECT 28.335 5.21 28.475 6.8 ;
      RECT 27.655 5.21 28.475 5.35 ;
      RECT 27.655 2.74 27.795 5.35 ;
      RECT 27.585 4.135 27.865 4.505 ;
      RECT 27.595 2.74 27.855 3.06 ;
      RECT 25.545 4.135 25.825 4.505 ;
      RECT 25.615 2.4 25.755 4.505 ;
      RECT 25.555 2.4 25.815 2.72 ;
      RECT 24.875 4.78 25.135 5.1 ;
      RECT 24.935 2.74 25.075 5.1 ;
      RECT 24.875 2.74 25.135 3.06 ;
      RECT 16.3 7.27 16.62 7.595 ;
      RECT 16.33 6.685 16.5 7.595 ;
      RECT 16.33 6.685 16.505 7.035 ;
      RECT 16.33 6.685 17.305 6.86 ;
      RECT 17.13 1.965 17.305 6.86 ;
      RECT 11.045 3.055 11.325 3.425 ;
      RECT 11.115 2.345 11.29 3.425 ;
      RECT 11.115 2.345 14.335 2.52 ;
      RECT 14.16 2.025 14.335 2.52 ;
      RECT 14.63 1.995 14.955 2.32 ;
      RECT 17.075 1.965 17.425 2.315 ;
      RECT 14.16 2.025 17.425 2.195 ;
      RECT 5.45 8.355 16.145 8.525 ;
      RECT 15.985 2.395 16.145 8.525 ;
      RECT 5.45 7.535 5.62 8.525 ;
      RECT 1.55 7.985 1.83 8.325 ;
      RECT 1.55 8.05 2.76 8.22 ;
      RECT 2.59 7.675 2.76 8.22 ;
      RECT 17.1 7.645 17.425 7.97 ;
      RECT 15.985 7.735 17.425 7.905 ;
      RECT 5.4 7.535 5.68 7.875 ;
      RECT 2.59 7.675 5.68 7.845 ;
      RECT 16.3 2.365 16.62 2.685 ;
      RECT 15.985 2.395 16.62 2.565 ;
      RECT 12.755 6.48 13.015 6.8 ;
      RECT 12.815 2.74 12.955 6.8 ;
      RECT 12.755 2.74 13.015 3.06 ;
      RECT 12.075 4.78 12.335 5.1 ;
      RECT 12.135 3.76 12.275 5.1 ;
      RECT 12.075 3.76 12.335 4.08 ;
      RECT 11.055 6.48 11.315 6.8 ;
      RECT 11.115 5.21 11.255 6.8 ;
      RECT 10.435 5.21 11.255 5.35 ;
      RECT 10.435 2.74 10.575 5.35 ;
      RECT 10.365 4.135 10.645 4.505 ;
      RECT 10.375 2.74 10.635 3.06 ;
      RECT 8.325 4.135 8.605 4.505 ;
      RECT 8.395 2.4 8.535 4.505 ;
      RECT 8.335 2.4 8.595 2.72 ;
      RECT 7.655 4.78 7.915 5.1 ;
      RECT 7.715 2.74 7.855 5.1 ;
      RECT 7.655 2.74 7.915 3.06 ;
      RECT 80.615 5.77 80.895 6.14 ;
      RECT 80.265 3.735 80.545 4.105 ;
      RECT 79.575 5.77 79.855 6.14 ;
      RECT 78.895 3.395 79.175 3.765 ;
      RECT 78.565 2.205 78.845 2.575 ;
      RECT 78.565 6.46 78.845 6.83 ;
      RECT 73.805 7.99 74.175 8.36 ;
      RECT 63.395 5.77 63.675 6.14 ;
      RECT 63.045 3.735 63.325 4.105 ;
      RECT 62.355 5.77 62.635 6.14 ;
      RECT 61.675 3.395 61.955 3.765 ;
      RECT 61.345 2.205 61.625 2.575 ;
      RECT 61.345 6.46 61.625 6.83 ;
      RECT 56.585 7.99 56.955 8.36 ;
      RECT 46.175 5.77 46.455 6.14 ;
      RECT 45.825 3.735 46.105 4.105 ;
      RECT 45.135 5.77 45.415 6.14 ;
      RECT 44.455 3.395 44.735 3.765 ;
      RECT 44.125 2.205 44.405 2.575 ;
      RECT 44.125 6.46 44.405 6.83 ;
      RECT 39.365 7.99 39.735 8.36 ;
      RECT 28.955 5.77 29.235 6.14 ;
      RECT 28.605 3.735 28.885 4.105 ;
      RECT 27.915 5.77 28.195 6.14 ;
      RECT 27.235 3.395 27.515 3.765 ;
      RECT 26.905 2.205 27.185 2.575 ;
      RECT 26.905 6.46 27.185 6.83 ;
      RECT 22.145 7.99 22.515 8.36 ;
      RECT 11.735 5.77 12.015 6.14 ;
      RECT 11.385 3.735 11.665 4.105 ;
      RECT 10.695 5.77 10.975 6.14 ;
      RECT 10.015 3.395 10.295 3.765 ;
      RECT 9.685 2.205 9.965 2.575 ;
      RECT 9.685 6.46 9.965 6.83 ;
      RECT 4.925 7.99 5.295 8.36 ;
    LAYER via1 ;
      RECT 88.425 8.375 88.575 8.525 ;
      RECT 86.07 7.73 86.22 7.88 ;
      RECT 86.055 2.065 86.205 2.215 ;
      RECT 85.265 2.45 85.415 2.6 ;
      RECT 85.265 7.36 85.415 7.51 ;
      RECT 83.6 2.08 83.75 2.23 ;
      RECT 81.69 2.825 81.84 2.975 ;
      RECT 81.69 6.565 81.84 6.715 ;
      RECT 81.01 3.845 81.16 3.995 ;
      RECT 81.01 4.865 81.16 5.015 ;
      RECT 80.67 5.885 80.82 6.035 ;
      RECT 80.33 3.845 80.48 3.995 ;
      RECT 79.99 3.165 80.14 3.315 ;
      RECT 79.99 6.565 80.14 6.715 ;
      RECT 79.64 5.885 79.79 6.035 ;
      RECT 79.31 2.825 79.46 2.975 ;
      RECT 78.97 3.505 79.12 3.655 ;
      RECT 78.63 2.315 78.78 2.465 ;
      RECT 78.63 6.565 78.78 6.715 ;
      RECT 77.27 2.485 77.42 2.635 ;
      RECT 76.59 2.825 76.74 2.975 ;
      RECT 76.59 4.865 76.74 5.015 ;
      RECT 74.345 7.63 74.495 7.78 ;
      RECT 73.915 8.1 74.065 8.25 ;
      RECT 71.24 7.73 71.39 7.88 ;
      RECT 68.85 7.73 69 7.88 ;
      RECT 68.835 2.065 68.985 2.215 ;
      RECT 68.045 2.45 68.195 2.6 ;
      RECT 68.045 7.36 68.195 7.51 ;
      RECT 66.38 2.08 66.53 2.23 ;
      RECT 64.47 2.825 64.62 2.975 ;
      RECT 64.47 6.565 64.62 6.715 ;
      RECT 63.79 3.845 63.94 3.995 ;
      RECT 63.79 4.865 63.94 5.015 ;
      RECT 63.45 5.885 63.6 6.035 ;
      RECT 63.11 3.845 63.26 3.995 ;
      RECT 62.77 3.165 62.92 3.315 ;
      RECT 62.77 6.565 62.92 6.715 ;
      RECT 62.42 5.885 62.57 6.035 ;
      RECT 62.09 2.825 62.24 2.975 ;
      RECT 61.75 3.505 61.9 3.655 ;
      RECT 61.41 2.315 61.56 2.465 ;
      RECT 61.41 6.565 61.56 6.715 ;
      RECT 60.05 2.485 60.2 2.635 ;
      RECT 59.37 2.825 59.52 2.975 ;
      RECT 59.37 4.865 59.52 5.015 ;
      RECT 57.125 7.63 57.275 7.78 ;
      RECT 56.695 8.1 56.845 8.25 ;
      RECT 54.02 7.73 54.17 7.88 ;
      RECT 51.63 7.73 51.78 7.88 ;
      RECT 51.615 2.065 51.765 2.215 ;
      RECT 50.825 2.45 50.975 2.6 ;
      RECT 50.825 7.36 50.975 7.51 ;
      RECT 49.16 2.08 49.31 2.23 ;
      RECT 47.25 2.825 47.4 2.975 ;
      RECT 47.25 6.565 47.4 6.715 ;
      RECT 46.57 3.845 46.72 3.995 ;
      RECT 46.57 4.865 46.72 5.015 ;
      RECT 46.23 5.885 46.38 6.035 ;
      RECT 45.89 3.845 46.04 3.995 ;
      RECT 45.55 3.165 45.7 3.315 ;
      RECT 45.55 6.565 45.7 6.715 ;
      RECT 45.2 5.885 45.35 6.035 ;
      RECT 44.87 2.825 45.02 2.975 ;
      RECT 44.53 3.505 44.68 3.655 ;
      RECT 44.19 2.315 44.34 2.465 ;
      RECT 44.19 6.565 44.34 6.715 ;
      RECT 42.83 2.485 42.98 2.635 ;
      RECT 42.15 2.825 42.3 2.975 ;
      RECT 42.15 4.865 42.3 5.015 ;
      RECT 39.905 7.63 40.055 7.78 ;
      RECT 39.475 8.1 39.625 8.25 ;
      RECT 36.8 7.73 36.95 7.88 ;
      RECT 34.41 7.73 34.56 7.88 ;
      RECT 34.395 2.065 34.545 2.215 ;
      RECT 33.605 2.45 33.755 2.6 ;
      RECT 33.605 7.36 33.755 7.51 ;
      RECT 31.94 2.08 32.09 2.23 ;
      RECT 30.03 2.825 30.18 2.975 ;
      RECT 30.03 6.565 30.18 6.715 ;
      RECT 29.35 3.845 29.5 3.995 ;
      RECT 29.35 4.865 29.5 5.015 ;
      RECT 29.01 5.885 29.16 6.035 ;
      RECT 28.67 3.845 28.82 3.995 ;
      RECT 28.33 3.165 28.48 3.315 ;
      RECT 28.33 6.565 28.48 6.715 ;
      RECT 27.98 5.885 28.13 6.035 ;
      RECT 27.65 2.825 27.8 2.975 ;
      RECT 27.31 3.505 27.46 3.655 ;
      RECT 26.97 2.315 27.12 2.465 ;
      RECT 26.97 6.565 27.12 6.715 ;
      RECT 25.61 2.485 25.76 2.635 ;
      RECT 24.93 2.825 25.08 2.975 ;
      RECT 24.93 4.865 25.08 5.015 ;
      RECT 22.685 7.63 22.835 7.78 ;
      RECT 22.255 8.1 22.405 8.25 ;
      RECT 19.58 7.73 19.73 7.88 ;
      RECT 17.19 7.73 17.34 7.88 ;
      RECT 17.175 2.065 17.325 2.215 ;
      RECT 16.385 2.45 16.535 2.6 ;
      RECT 16.385 7.36 16.535 7.51 ;
      RECT 14.72 2.08 14.87 2.23 ;
      RECT 12.81 2.825 12.96 2.975 ;
      RECT 12.81 6.565 12.96 6.715 ;
      RECT 12.13 3.845 12.28 3.995 ;
      RECT 12.13 4.865 12.28 5.015 ;
      RECT 11.79 5.885 11.94 6.035 ;
      RECT 11.45 3.845 11.6 3.995 ;
      RECT 11.11 3.165 11.26 3.315 ;
      RECT 11.11 6.565 11.26 6.715 ;
      RECT 10.76 5.885 10.91 6.035 ;
      RECT 10.43 2.825 10.58 2.975 ;
      RECT 10.09 3.505 10.24 3.655 ;
      RECT 9.75 2.315 9.9 2.465 ;
      RECT 9.75 6.565 9.9 6.715 ;
      RECT 8.39 2.485 8.54 2.635 ;
      RECT 7.71 2.825 7.86 2.975 ;
      RECT 7.71 4.865 7.86 5.015 ;
      RECT 5.465 7.63 5.615 7.78 ;
      RECT 5.035 8.1 5.185 8.25 ;
      RECT 1.615 8.08 1.765 8.23 ;
      RECT 1.24 7.34 1.39 7.49 ;
    LAYER met1 ;
      RECT 88.305 8.76 88.595 8.99 ;
      RECT 88.365 7.28 88.535 8.99 ;
      RECT 88.335 8.29 88.66 8.615 ;
      RECT 88.305 7.28 88.595 7.51 ;
      RECT 87.9 2.395 88.005 2.965 ;
      RECT 87.9 2.73 88.225 2.96 ;
      RECT 87.9 2.76 88.395 2.93 ;
      RECT 87.9 2.395 88.09 2.96 ;
      RECT 87.315 2.36 87.605 2.59 ;
      RECT 87.315 2.395 88.09 2.565 ;
      RECT 87.375 0.88 87.545 2.59 ;
      RECT 87.315 0.88 87.605 1.11 ;
      RECT 87.315 8.76 87.605 8.99 ;
      RECT 87.375 7.28 87.545 8.99 ;
      RECT 87.315 7.28 87.605 7.51 ;
      RECT 87.315 7.315 88.17 7.475 ;
      RECT 88 6.91 88.17 7.475 ;
      RECT 87.315 7.31 87.71 7.475 ;
      RECT 87.935 6.91 88.225 7.14 ;
      RECT 87.935 6.94 88.395 7.11 ;
      RECT 86.945 2.73 87.235 2.96 ;
      RECT 86.945 2.76 87.405 2.93 ;
      RECT 87.01 1.655 87.175 2.96 ;
      RECT 85.525 1.625 85.815 1.855 ;
      RECT 85.525 1.655 87.175 1.825 ;
      RECT 85.585 0.885 85.755 1.855 ;
      RECT 85.525 0.885 85.815 1.115 ;
      RECT 85.525 8.755 85.815 8.985 ;
      RECT 85.585 8.015 85.755 8.985 ;
      RECT 85.585 8.11 87.175 8.28 ;
      RECT 87.005 6.91 87.175 8.28 ;
      RECT 85.525 8.015 85.815 8.245 ;
      RECT 86.945 6.91 87.235 7.14 ;
      RECT 86.945 6.94 87.405 7.11 ;
      RECT 85.955 1.965 86.305 2.315 ;
      RECT 85.785 2.025 86.305 2.195 ;
      RECT 85.98 7.645 86.305 7.97 ;
      RECT 85.955 7.645 86.305 7.875 ;
      RECT 85.785 7.675 86.305 7.845 ;
      RECT 85.18 2.365 85.5 2.685 ;
      RECT 85.15 2.365 85.5 2.595 ;
      RECT 84.865 2.395 85.5 2.565 ;
      RECT 85.18 7.27 85.5 7.595 ;
      RECT 85.15 7.275 85.5 7.505 ;
      RECT 84.98 7.305 85.5 7.475 ;
      RECT 80.925 3.79 81.245 4.05 ;
      RECT 81.96 3.805 82.25 4.035 ;
      RECT 80.925 3.85 82.25 3.99 ;
      RECT 80.585 5.83 80.905 6.09 ;
      RECT 81.96 5.845 82.25 6.075 ;
      RECT 82.035 5.55 82.175 6.075 ;
      RECT 80.675 5.55 80.815 6.09 ;
      RECT 80.675 5.55 82.175 5.69 ;
      RECT 81.605 2.77 81.925 3.03 ;
      RECT 81.33 2.83 81.925 2.97 ;
      RECT 78.545 6.51 78.865 6.77 ;
      RECT 77.54 6.525 77.83 6.755 ;
      RECT 77.54 6.57 79.455 6.71 ;
      RECT 79.315 6.23 79.455 6.71 ;
      RECT 79.315 6.23 81.325 6.37 ;
      RECT 81.185 5.845 81.325 6.37 ;
      RECT 81.11 5.845 81.4 6.075 ;
      RECT 80.925 4.81 81.245 5.07 ;
      RECT 78.78 4.825 79.07 5.055 ;
      RECT 78.78 4.87 81.245 5.01 ;
      RECT 80.245 3.79 80.565 4.05 ;
      RECT 77.88 3.805 78.17 4.035 ;
      RECT 77.88 3.85 80.565 3.99 ;
      RECT 79.905 6.51 80.225 6.77 ;
      RECT 79.905 6.57 80.5 6.71 ;
      RECT 79.905 3.11 80.225 3.37 ;
      RECT 79.63 3.17 80.225 3.31 ;
      RECT 79.225 2.77 79.545 3.03 ;
      RECT 78.95 2.83 79.545 2.97 ;
      RECT 78.885 3.45 79.205 3.71 ;
      RECT 76.01 3.465 76.3 3.695 ;
      RECT 76.01 3.51 79.205 3.65 ;
      RECT 78.465 2.79 78.605 3.65 ;
      RECT 78.39 2.79 78.68 3.02 ;
      RECT 78.545 2.26 78.865 2.52 ;
      RECT 78.545 2.275 79.05 2.505 ;
      RECT 78.455 2.32 79.05 2.46 ;
      RECT 77.88 2.79 78.17 3.02 ;
      RECT 77.275 2.835 78.17 2.975 ;
      RECT 77.275 2.43 77.415 2.975 ;
      RECT 77.185 2.43 77.505 2.69 ;
      RECT 76.505 2.77 76.825 3.03 ;
      RECT 76.23 2.83 76.825 2.97 ;
      RECT 76.505 4.81 76.825 5.07 ;
      RECT 76.23 4.87 76.825 5.01 ;
      RECT 74.27 7.565 74.56 7.875 ;
      RECT 74.1 7.675 74.59 7.845 ;
      RECT 74.25 7.565 74.59 7.845 ;
      RECT 73.84 8.755 74.13 8.985 ;
      RECT 73.9 7.985 74.07 8.985 ;
      RECT 73.805 7.985 74.175 8.36 ;
      RECT 71.085 8.76 71.375 8.99 ;
      RECT 71.145 7.28 71.315 8.99 ;
      RECT 71.145 7.645 71.475 7.97 ;
      RECT 71.085 7.28 71.375 7.51 ;
      RECT 70.68 2.395 70.785 2.965 ;
      RECT 70.68 2.73 71.005 2.96 ;
      RECT 70.68 2.76 71.175 2.93 ;
      RECT 70.68 2.395 70.87 2.96 ;
      RECT 70.095 2.36 70.385 2.59 ;
      RECT 70.095 2.395 70.87 2.565 ;
      RECT 70.155 0.88 70.325 2.59 ;
      RECT 70.095 0.88 70.385 1.11 ;
      RECT 70.095 8.76 70.385 8.99 ;
      RECT 70.155 7.28 70.325 8.99 ;
      RECT 70.095 7.28 70.385 7.51 ;
      RECT 70.095 7.315 70.95 7.475 ;
      RECT 70.78 6.91 70.95 7.475 ;
      RECT 70.095 7.31 70.49 7.475 ;
      RECT 70.715 6.91 71.005 7.14 ;
      RECT 70.715 6.94 71.175 7.11 ;
      RECT 69.725 2.73 70.015 2.96 ;
      RECT 69.725 2.76 70.185 2.93 ;
      RECT 69.79 1.655 69.955 2.96 ;
      RECT 68.305 1.625 68.595 1.855 ;
      RECT 68.305 1.655 69.955 1.825 ;
      RECT 68.365 0.885 68.535 1.855 ;
      RECT 68.305 0.885 68.595 1.115 ;
      RECT 68.305 8.755 68.595 8.985 ;
      RECT 68.365 8.015 68.535 8.985 ;
      RECT 68.365 8.11 69.955 8.28 ;
      RECT 69.785 6.91 69.955 8.28 ;
      RECT 68.305 8.015 68.595 8.245 ;
      RECT 69.725 6.91 70.015 7.14 ;
      RECT 69.725 6.94 70.185 7.11 ;
      RECT 68.735 1.965 69.085 2.315 ;
      RECT 68.565 2.025 69.085 2.195 ;
      RECT 68.76 7.645 69.085 7.97 ;
      RECT 68.735 7.645 69.085 7.875 ;
      RECT 68.565 7.675 69.085 7.845 ;
      RECT 67.96 2.365 68.28 2.685 ;
      RECT 67.93 2.365 68.28 2.595 ;
      RECT 67.645 2.395 68.28 2.565 ;
      RECT 67.96 7.27 68.28 7.595 ;
      RECT 67.93 7.275 68.28 7.505 ;
      RECT 67.76 7.305 68.28 7.475 ;
      RECT 63.705 3.79 64.025 4.05 ;
      RECT 64.74 3.805 65.03 4.035 ;
      RECT 63.705 3.85 65.03 3.99 ;
      RECT 63.365 5.83 63.685 6.09 ;
      RECT 64.74 5.845 65.03 6.075 ;
      RECT 64.815 5.55 64.955 6.075 ;
      RECT 63.455 5.55 63.595 6.09 ;
      RECT 63.455 5.55 64.955 5.69 ;
      RECT 64.385 2.77 64.705 3.03 ;
      RECT 64.11 2.83 64.705 2.97 ;
      RECT 61.325 6.51 61.645 6.77 ;
      RECT 60.32 6.525 60.61 6.755 ;
      RECT 60.32 6.57 62.235 6.71 ;
      RECT 62.095 6.23 62.235 6.71 ;
      RECT 62.095 6.23 64.105 6.37 ;
      RECT 63.965 5.845 64.105 6.37 ;
      RECT 63.89 5.845 64.18 6.075 ;
      RECT 63.705 4.81 64.025 5.07 ;
      RECT 61.56 4.825 61.85 5.055 ;
      RECT 61.56 4.87 64.025 5.01 ;
      RECT 63.025 3.79 63.345 4.05 ;
      RECT 60.66 3.805 60.95 4.035 ;
      RECT 60.66 3.85 63.345 3.99 ;
      RECT 62.685 6.51 63.005 6.77 ;
      RECT 62.685 6.57 63.28 6.71 ;
      RECT 62.685 3.11 63.005 3.37 ;
      RECT 62.41 3.17 63.005 3.31 ;
      RECT 62.005 2.77 62.325 3.03 ;
      RECT 61.73 2.83 62.325 2.97 ;
      RECT 61.665 3.45 61.985 3.71 ;
      RECT 58.79 3.465 59.08 3.695 ;
      RECT 58.79 3.51 61.985 3.65 ;
      RECT 61.245 2.79 61.385 3.65 ;
      RECT 61.17 2.79 61.46 3.02 ;
      RECT 61.325 2.26 61.645 2.52 ;
      RECT 61.325 2.275 61.83 2.505 ;
      RECT 61.235 2.32 61.83 2.46 ;
      RECT 60.66 2.79 60.95 3.02 ;
      RECT 60.055 2.835 60.95 2.975 ;
      RECT 60.055 2.43 60.195 2.975 ;
      RECT 59.965 2.43 60.285 2.69 ;
      RECT 59.285 2.77 59.605 3.03 ;
      RECT 59.01 2.83 59.605 2.97 ;
      RECT 59.285 4.81 59.605 5.07 ;
      RECT 59.01 4.87 59.605 5.01 ;
      RECT 57.05 7.565 57.34 7.875 ;
      RECT 56.88 7.675 57.37 7.845 ;
      RECT 57.03 7.565 57.37 7.845 ;
      RECT 56.62 8.755 56.91 8.985 ;
      RECT 56.68 7.985 56.85 8.985 ;
      RECT 56.585 7.985 56.955 8.36 ;
      RECT 53.865 8.76 54.155 8.99 ;
      RECT 53.925 7.28 54.095 8.99 ;
      RECT 53.925 7.645 54.255 7.97 ;
      RECT 53.865 7.28 54.155 7.51 ;
      RECT 53.46 2.395 53.565 2.965 ;
      RECT 53.46 2.73 53.785 2.96 ;
      RECT 53.46 2.76 53.955 2.93 ;
      RECT 53.46 2.395 53.65 2.96 ;
      RECT 52.875 2.36 53.165 2.59 ;
      RECT 52.875 2.395 53.65 2.565 ;
      RECT 52.935 0.88 53.105 2.59 ;
      RECT 52.875 0.88 53.165 1.11 ;
      RECT 52.875 8.76 53.165 8.99 ;
      RECT 52.935 7.28 53.105 8.99 ;
      RECT 52.875 7.28 53.165 7.51 ;
      RECT 52.875 7.315 53.73 7.475 ;
      RECT 53.56 6.91 53.73 7.475 ;
      RECT 52.875 7.31 53.27 7.475 ;
      RECT 53.495 6.91 53.785 7.14 ;
      RECT 53.495 6.94 53.955 7.11 ;
      RECT 52.505 2.73 52.795 2.96 ;
      RECT 52.505 2.76 52.965 2.93 ;
      RECT 52.57 1.655 52.735 2.96 ;
      RECT 51.085 1.625 51.375 1.855 ;
      RECT 51.085 1.655 52.735 1.825 ;
      RECT 51.145 0.885 51.315 1.855 ;
      RECT 51.085 0.885 51.375 1.115 ;
      RECT 51.085 8.755 51.375 8.985 ;
      RECT 51.145 8.015 51.315 8.985 ;
      RECT 51.145 8.11 52.735 8.28 ;
      RECT 52.565 6.91 52.735 8.28 ;
      RECT 51.085 8.015 51.375 8.245 ;
      RECT 52.505 6.91 52.795 7.14 ;
      RECT 52.505 6.94 52.965 7.11 ;
      RECT 51.515 1.965 51.865 2.315 ;
      RECT 51.345 2.025 51.865 2.195 ;
      RECT 51.54 7.645 51.865 7.97 ;
      RECT 51.515 7.645 51.865 7.875 ;
      RECT 51.345 7.675 51.865 7.845 ;
      RECT 50.74 2.365 51.06 2.685 ;
      RECT 50.71 2.365 51.06 2.595 ;
      RECT 50.425 2.395 51.06 2.565 ;
      RECT 50.74 7.27 51.06 7.595 ;
      RECT 50.71 7.275 51.06 7.505 ;
      RECT 50.54 7.305 51.06 7.475 ;
      RECT 46.485 3.79 46.805 4.05 ;
      RECT 47.52 3.805 47.81 4.035 ;
      RECT 46.485 3.85 47.81 3.99 ;
      RECT 46.145 5.83 46.465 6.09 ;
      RECT 47.52 5.845 47.81 6.075 ;
      RECT 47.595 5.55 47.735 6.075 ;
      RECT 46.235 5.55 46.375 6.09 ;
      RECT 46.235 5.55 47.735 5.69 ;
      RECT 47.165 2.77 47.485 3.03 ;
      RECT 46.89 2.83 47.485 2.97 ;
      RECT 44.105 6.51 44.425 6.77 ;
      RECT 43.1 6.525 43.39 6.755 ;
      RECT 43.1 6.57 45.015 6.71 ;
      RECT 44.875 6.23 45.015 6.71 ;
      RECT 44.875 6.23 46.885 6.37 ;
      RECT 46.745 5.845 46.885 6.37 ;
      RECT 46.67 5.845 46.96 6.075 ;
      RECT 46.485 4.81 46.805 5.07 ;
      RECT 44.34 4.825 44.63 5.055 ;
      RECT 44.34 4.87 46.805 5.01 ;
      RECT 45.805 3.79 46.125 4.05 ;
      RECT 43.44 3.805 43.73 4.035 ;
      RECT 43.44 3.85 46.125 3.99 ;
      RECT 45.465 6.51 45.785 6.77 ;
      RECT 45.465 6.57 46.06 6.71 ;
      RECT 45.465 3.11 45.785 3.37 ;
      RECT 45.19 3.17 45.785 3.31 ;
      RECT 44.785 2.77 45.105 3.03 ;
      RECT 44.51 2.83 45.105 2.97 ;
      RECT 44.445 3.45 44.765 3.71 ;
      RECT 41.57 3.465 41.86 3.695 ;
      RECT 41.57 3.51 44.765 3.65 ;
      RECT 44.025 2.79 44.165 3.65 ;
      RECT 43.95 2.79 44.24 3.02 ;
      RECT 44.105 2.26 44.425 2.52 ;
      RECT 44.105 2.275 44.61 2.505 ;
      RECT 44.015 2.32 44.61 2.46 ;
      RECT 43.44 2.79 43.73 3.02 ;
      RECT 42.835 2.835 43.73 2.975 ;
      RECT 42.835 2.43 42.975 2.975 ;
      RECT 42.745 2.43 43.065 2.69 ;
      RECT 42.065 2.77 42.385 3.03 ;
      RECT 41.79 2.83 42.385 2.97 ;
      RECT 42.065 4.81 42.385 5.07 ;
      RECT 41.79 4.87 42.385 5.01 ;
      RECT 39.83 7.565 40.12 7.875 ;
      RECT 39.66 7.675 40.15 7.845 ;
      RECT 39.81 7.565 40.15 7.845 ;
      RECT 39.4 8.755 39.69 8.985 ;
      RECT 39.46 7.985 39.63 8.985 ;
      RECT 39.365 7.985 39.735 8.36 ;
      RECT 36.645 8.76 36.935 8.99 ;
      RECT 36.705 7.28 36.875 8.99 ;
      RECT 36.705 7.645 37.035 7.97 ;
      RECT 36.645 7.28 36.935 7.51 ;
      RECT 36.24 2.395 36.345 2.965 ;
      RECT 36.24 2.73 36.565 2.96 ;
      RECT 36.24 2.76 36.735 2.93 ;
      RECT 36.24 2.395 36.43 2.96 ;
      RECT 35.655 2.36 35.945 2.59 ;
      RECT 35.655 2.395 36.43 2.565 ;
      RECT 35.715 0.88 35.885 2.59 ;
      RECT 35.655 0.88 35.945 1.11 ;
      RECT 35.655 8.76 35.945 8.99 ;
      RECT 35.715 7.28 35.885 8.99 ;
      RECT 35.655 7.28 35.945 7.51 ;
      RECT 35.655 7.315 36.51 7.475 ;
      RECT 36.34 6.91 36.51 7.475 ;
      RECT 35.655 7.31 36.05 7.475 ;
      RECT 36.275 6.91 36.565 7.14 ;
      RECT 36.275 6.94 36.735 7.11 ;
      RECT 35.285 2.73 35.575 2.96 ;
      RECT 35.285 2.76 35.745 2.93 ;
      RECT 35.35 1.655 35.515 2.96 ;
      RECT 33.865 1.625 34.155 1.855 ;
      RECT 33.865 1.655 35.515 1.825 ;
      RECT 33.925 0.885 34.095 1.855 ;
      RECT 33.865 0.885 34.155 1.115 ;
      RECT 33.865 8.755 34.155 8.985 ;
      RECT 33.925 8.015 34.095 8.985 ;
      RECT 33.925 8.11 35.515 8.28 ;
      RECT 35.345 6.91 35.515 8.28 ;
      RECT 33.865 8.015 34.155 8.245 ;
      RECT 35.285 6.91 35.575 7.14 ;
      RECT 35.285 6.94 35.745 7.11 ;
      RECT 34.295 1.965 34.645 2.315 ;
      RECT 34.125 2.025 34.645 2.195 ;
      RECT 34.32 7.645 34.645 7.97 ;
      RECT 34.295 7.645 34.645 7.875 ;
      RECT 34.125 7.675 34.645 7.845 ;
      RECT 33.52 2.365 33.84 2.685 ;
      RECT 33.49 2.365 33.84 2.595 ;
      RECT 33.205 2.395 33.84 2.565 ;
      RECT 33.52 7.27 33.84 7.595 ;
      RECT 33.49 7.275 33.84 7.505 ;
      RECT 33.32 7.305 33.84 7.475 ;
      RECT 29.265 3.79 29.585 4.05 ;
      RECT 30.3 3.805 30.59 4.035 ;
      RECT 29.265 3.85 30.59 3.99 ;
      RECT 28.925 5.83 29.245 6.09 ;
      RECT 30.3 5.845 30.59 6.075 ;
      RECT 30.375 5.55 30.515 6.075 ;
      RECT 29.015 5.55 29.155 6.09 ;
      RECT 29.015 5.55 30.515 5.69 ;
      RECT 29.945 2.77 30.265 3.03 ;
      RECT 29.67 2.83 30.265 2.97 ;
      RECT 26.885 6.51 27.205 6.77 ;
      RECT 25.88 6.525 26.17 6.755 ;
      RECT 25.88 6.57 27.795 6.71 ;
      RECT 27.655 6.23 27.795 6.71 ;
      RECT 27.655 6.23 29.665 6.37 ;
      RECT 29.525 5.845 29.665 6.37 ;
      RECT 29.45 5.845 29.74 6.075 ;
      RECT 29.265 4.81 29.585 5.07 ;
      RECT 27.12 4.825 27.41 5.055 ;
      RECT 27.12 4.87 29.585 5.01 ;
      RECT 28.585 3.79 28.905 4.05 ;
      RECT 26.22 3.805 26.51 4.035 ;
      RECT 26.22 3.85 28.905 3.99 ;
      RECT 28.245 6.51 28.565 6.77 ;
      RECT 28.245 6.57 28.84 6.71 ;
      RECT 28.245 3.11 28.565 3.37 ;
      RECT 27.97 3.17 28.565 3.31 ;
      RECT 27.565 2.77 27.885 3.03 ;
      RECT 27.29 2.83 27.885 2.97 ;
      RECT 27.225 3.45 27.545 3.71 ;
      RECT 24.35 3.465 24.64 3.695 ;
      RECT 24.35 3.51 27.545 3.65 ;
      RECT 26.805 2.79 26.945 3.65 ;
      RECT 26.73 2.79 27.02 3.02 ;
      RECT 26.885 2.26 27.205 2.52 ;
      RECT 26.885 2.275 27.39 2.505 ;
      RECT 26.795 2.32 27.39 2.46 ;
      RECT 26.22 2.79 26.51 3.02 ;
      RECT 25.615 2.835 26.51 2.975 ;
      RECT 25.615 2.43 25.755 2.975 ;
      RECT 25.525 2.43 25.845 2.69 ;
      RECT 24.845 2.77 25.165 3.03 ;
      RECT 24.57 2.83 25.165 2.97 ;
      RECT 24.845 4.81 25.165 5.07 ;
      RECT 24.57 4.87 25.165 5.01 ;
      RECT 22.61 7.565 22.9 7.875 ;
      RECT 22.44 7.675 22.93 7.845 ;
      RECT 22.59 7.565 22.93 7.845 ;
      RECT 22.18 8.755 22.47 8.985 ;
      RECT 22.24 7.985 22.41 8.985 ;
      RECT 22.145 7.985 22.515 8.36 ;
      RECT 19.425 8.76 19.715 8.99 ;
      RECT 19.485 7.28 19.655 8.99 ;
      RECT 19.485 7.645 19.815 7.97 ;
      RECT 19.425 7.28 19.715 7.51 ;
      RECT 19.02 2.395 19.125 2.965 ;
      RECT 19.02 2.73 19.345 2.96 ;
      RECT 19.02 2.76 19.515 2.93 ;
      RECT 19.02 2.395 19.21 2.96 ;
      RECT 18.435 2.36 18.725 2.59 ;
      RECT 18.435 2.395 19.21 2.565 ;
      RECT 18.495 0.88 18.665 2.59 ;
      RECT 18.435 0.88 18.725 1.11 ;
      RECT 18.435 8.76 18.725 8.99 ;
      RECT 18.495 7.28 18.665 8.99 ;
      RECT 18.435 7.28 18.725 7.51 ;
      RECT 18.435 7.315 19.29 7.475 ;
      RECT 19.12 6.91 19.29 7.475 ;
      RECT 18.435 7.31 18.83 7.475 ;
      RECT 19.055 6.91 19.345 7.14 ;
      RECT 19.055 6.94 19.515 7.11 ;
      RECT 18.065 2.73 18.355 2.96 ;
      RECT 18.065 2.76 18.525 2.93 ;
      RECT 18.13 1.655 18.295 2.96 ;
      RECT 16.645 1.625 16.935 1.855 ;
      RECT 16.645 1.655 18.295 1.825 ;
      RECT 16.705 0.885 16.875 1.855 ;
      RECT 16.645 0.885 16.935 1.115 ;
      RECT 16.645 8.755 16.935 8.985 ;
      RECT 16.705 8.015 16.875 8.985 ;
      RECT 16.705 8.11 18.295 8.28 ;
      RECT 18.125 6.91 18.295 8.28 ;
      RECT 16.645 8.015 16.935 8.245 ;
      RECT 18.065 6.91 18.355 7.14 ;
      RECT 18.065 6.94 18.525 7.11 ;
      RECT 17.075 1.965 17.425 2.315 ;
      RECT 16.905 2.025 17.425 2.195 ;
      RECT 17.1 7.645 17.425 7.97 ;
      RECT 17.075 7.645 17.425 7.875 ;
      RECT 16.905 7.675 17.425 7.845 ;
      RECT 16.3 2.365 16.62 2.685 ;
      RECT 16.27 2.365 16.62 2.595 ;
      RECT 15.985 2.395 16.62 2.565 ;
      RECT 16.3 7.27 16.62 7.595 ;
      RECT 16.27 7.275 16.62 7.505 ;
      RECT 16.1 7.305 16.62 7.475 ;
      RECT 12.045 3.79 12.365 4.05 ;
      RECT 13.08 3.805 13.37 4.035 ;
      RECT 12.045 3.85 13.37 3.99 ;
      RECT 11.705 5.83 12.025 6.09 ;
      RECT 13.08 5.845 13.37 6.075 ;
      RECT 13.155 5.55 13.295 6.075 ;
      RECT 11.795 5.55 11.935 6.09 ;
      RECT 11.795 5.55 13.295 5.69 ;
      RECT 12.725 2.77 13.045 3.03 ;
      RECT 12.45 2.83 13.045 2.97 ;
      RECT 9.665 6.51 9.985 6.77 ;
      RECT 8.66 6.525 8.95 6.755 ;
      RECT 8.66 6.57 10.575 6.71 ;
      RECT 10.435 6.23 10.575 6.71 ;
      RECT 10.435 6.23 12.445 6.37 ;
      RECT 12.305 5.845 12.445 6.37 ;
      RECT 12.23 5.845 12.52 6.075 ;
      RECT 12.045 4.81 12.365 5.07 ;
      RECT 9.9 4.825 10.19 5.055 ;
      RECT 9.9 4.87 12.365 5.01 ;
      RECT 11.365 3.79 11.685 4.05 ;
      RECT 9 3.805 9.29 4.035 ;
      RECT 9 3.85 11.685 3.99 ;
      RECT 11.025 6.51 11.345 6.77 ;
      RECT 11.025 6.57 11.62 6.71 ;
      RECT 11.025 3.11 11.345 3.37 ;
      RECT 10.75 3.17 11.345 3.31 ;
      RECT 10.345 2.77 10.665 3.03 ;
      RECT 10.07 2.83 10.665 2.97 ;
      RECT 10.005 3.45 10.325 3.71 ;
      RECT 7.13 3.465 7.42 3.695 ;
      RECT 7.13 3.51 10.325 3.65 ;
      RECT 9.585 2.79 9.725 3.65 ;
      RECT 9.51 2.79 9.8 3.02 ;
      RECT 9.665 2.26 9.985 2.52 ;
      RECT 9.665 2.275 10.17 2.505 ;
      RECT 9.575 2.32 10.17 2.46 ;
      RECT 9 2.79 9.29 3.02 ;
      RECT 8.395 2.835 9.29 2.975 ;
      RECT 8.395 2.43 8.535 2.975 ;
      RECT 8.305 2.43 8.625 2.69 ;
      RECT 7.625 2.77 7.945 3.03 ;
      RECT 7.35 2.83 7.945 2.97 ;
      RECT 7.625 4.81 7.945 5.07 ;
      RECT 7.35 4.87 7.945 5.01 ;
      RECT 5.39 7.565 5.68 7.875 ;
      RECT 5.22 7.675 5.71 7.845 ;
      RECT 5.37 7.565 5.71 7.845 ;
      RECT 4.96 8.755 5.25 8.985 ;
      RECT 5.02 7.985 5.19 8.985 ;
      RECT 4.925 7.985 5.295 8.36 ;
      RECT 1.55 8.755 1.84 8.985 ;
      RECT 1.61 8.015 1.78 8.985 ;
      RECT 1.52 8.015 1.86 8.295 ;
      RECT 1.145 7.275 1.485 7.555 ;
      RECT 1.005 7.305 1.485 7.475 ;
      RECT 83.51 1.995 83.835 2.32 ;
      RECT 81.28 6.51 81.925 6.77 ;
      RECT 79.23 5.83 79.875 6.09 ;
      RECT 66.29 1.995 66.615 2.32 ;
      RECT 64.06 6.51 64.705 6.77 ;
      RECT 62.01 5.83 62.655 6.09 ;
      RECT 49.07 1.995 49.395 2.32 ;
      RECT 46.84 6.51 47.485 6.77 ;
      RECT 44.79 5.83 45.435 6.09 ;
      RECT 31.85 1.995 32.175 2.32 ;
      RECT 29.62 6.51 30.265 6.77 ;
      RECT 27.57 5.83 28.215 6.09 ;
      RECT 14.63 1.995 14.955 2.32 ;
      RECT 12.4 6.51 13.045 6.77 ;
      RECT 10.35 5.83 10.995 6.09 ;
    LAYER mcon ;
      RECT 88.365 7.31 88.535 7.48 ;
      RECT 88.365 8.79 88.535 8.96 ;
      RECT 87.995 2.76 88.165 2.93 ;
      RECT 87.995 6.94 88.165 7.11 ;
      RECT 87.375 0.91 87.545 1.08 ;
      RECT 87.375 2.39 87.545 2.56 ;
      RECT 87.375 7.31 87.545 7.48 ;
      RECT 87.375 8.79 87.545 8.96 ;
      RECT 87.005 2.76 87.175 2.93 ;
      RECT 87.005 6.94 87.175 7.11 ;
      RECT 86.015 2.025 86.185 2.195 ;
      RECT 86.015 7.675 86.185 7.845 ;
      RECT 85.585 0.915 85.755 1.085 ;
      RECT 85.585 1.655 85.755 1.825 ;
      RECT 85.585 8.045 85.755 8.215 ;
      RECT 85.585 8.785 85.755 8.955 ;
      RECT 85.21 2.395 85.38 2.565 ;
      RECT 85.21 7.305 85.38 7.475 ;
      RECT 82.02 3.835 82.19 4.005 ;
      RECT 82.02 5.875 82.19 6.045 ;
      RECT 81.68 2.815 81.85 2.985 ;
      RECT 81.34 6.555 81.51 6.725 ;
      RECT 81.17 5.875 81.34 6.045 ;
      RECT 80.66 5.875 80.83 6.045 ;
      RECT 79.98 3.155 80.15 3.325 ;
      RECT 79.98 6.555 80.15 6.725 ;
      RECT 79.3 2.815 79.47 2.985 ;
      RECT 79.29 5.875 79.46 6.045 ;
      RECT 78.84 4.855 79.01 5.025 ;
      RECT 78.82 2.305 78.99 2.475 ;
      RECT 78.45 2.82 78.62 2.99 ;
      RECT 77.94 2.82 78.11 2.99 ;
      RECT 77.94 3.835 78.11 4.005 ;
      RECT 77.6 6.555 77.77 6.725 ;
      RECT 76.58 2.815 76.75 2.985 ;
      RECT 76.58 4.855 76.75 5.025 ;
      RECT 76.07 3.495 76.24 3.665 ;
      RECT 74.33 7.675 74.5 7.845 ;
      RECT 73.9 8.045 74.07 8.215 ;
      RECT 73.9 8.785 74.07 8.955 ;
      RECT 71.145 7.31 71.315 7.48 ;
      RECT 71.145 8.79 71.315 8.96 ;
      RECT 70.775 2.76 70.945 2.93 ;
      RECT 70.775 6.94 70.945 7.11 ;
      RECT 70.155 0.91 70.325 1.08 ;
      RECT 70.155 2.39 70.325 2.56 ;
      RECT 70.155 7.31 70.325 7.48 ;
      RECT 70.155 8.79 70.325 8.96 ;
      RECT 69.785 2.76 69.955 2.93 ;
      RECT 69.785 6.94 69.955 7.11 ;
      RECT 68.795 2.025 68.965 2.195 ;
      RECT 68.795 7.675 68.965 7.845 ;
      RECT 68.365 0.915 68.535 1.085 ;
      RECT 68.365 1.655 68.535 1.825 ;
      RECT 68.365 8.045 68.535 8.215 ;
      RECT 68.365 8.785 68.535 8.955 ;
      RECT 67.99 2.395 68.16 2.565 ;
      RECT 67.99 7.305 68.16 7.475 ;
      RECT 64.8 3.835 64.97 4.005 ;
      RECT 64.8 5.875 64.97 6.045 ;
      RECT 64.46 2.815 64.63 2.985 ;
      RECT 64.12 6.555 64.29 6.725 ;
      RECT 63.95 5.875 64.12 6.045 ;
      RECT 63.44 5.875 63.61 6.045 ;
      RECT 62.76 3.155 62.93 3.325 ;
      RECT 62.76 6.555 62.93 6.725 ;
      RECT 62.08 2.815 62.25 2.985 ;
      RECT 62.07 5.875 62.24 6.045 ;
      RECT 61.62 4.855 61.79 5.025 ;
      RECT 61.6 2.305 61.77 2.475 ;
      RECT 61.23 2.82 61.4 2.99 ;
      RECT 60.72 2.82 60.89 2.99 ;
      RECT 60.72 3.835 60.89 4.005 ;
      RECT 60.38 6.555 60.55 6.725 ;
      RECT 59.36 2.815 59.53 2.985 ;
      RECT 59.36 4.855 59.53 5.025 ;
      RECT 58.85 3.495 59.02 3.665 ;
      RECT 57.11 7.675 57.28 7.845 ;
      RECT 56.68 8.045 56.85 8.215 ;
      RECT 56.68 8.785 56.85 8.955 ;
      RECT 53.925 7.31 54.095 7.48 ;
      RECT 53.925 8.79 54.095 8.96 ;
      RECT 53.555 2.76 53.725 2.93 ;
      RECT 53.555 6.94 53.725 7.11 ;
      RECT 52.935 0.91 53.105 1.08 ;
      RECT 52.935 2.39 53.105 2.56 ;
      RECT 52.935 7.31 53.105 7.48 ;
      RECT 52.935 8.79 53.105 8.96 ;
      RECT 52.565 2.76 52.735 2.93 ;
      RECT 52.565 6.94 52.735 7.11 ;
      RECT 51.575 2.025 51.745 2.195 ;
      RECT 51.575 7.675 51.745 7.845 ;
      RECT 51.145 0.915 51.315 1.085 ;
      RECT 51.145 1.655 51.315 1.825 ;
      RECT 51.145 8.045 51.315 8.215 ;
      RECT 51.145 8.785 51.315 8.955 ;
      RECT 50.77 2.395 50.94 2.565 ;
      RECT 50.77 7.305 50.94 7.475 ;
      RECT 47.58 3.835 47.75 4.005 ;
      RECT 47.58 5.875 47.75 6.045 ;
      RECT 47.24 2.815 47.41 2.985 ;
      RECT 46.9 6.555 47.07 6.725 ;
      RECT 46.73 5.875 46.9 6.045 ;
      RECT 46.22 5.875 46.39 6.045 ;
      RECT 45.54 3.155 45.71 3.325 ;
      RECT 45.54 6.555 45.71 6.725 ;
      RECT 44.86 2.815 45.03 2.985 ;
      RECT 44.85 5.875 45.02 6.045 ;
      RECT 44.4 4.855 44.57 5.025 ;
      RECT 44.38 2.305 44.55 2.475 ;
      RECT 44.01 2.82 44.18 2.99 ;
      RECT 43.5 2.82 43.67 2.99 ;
      RECT 43.5 3.835 43.67 4.005 ;
      RECT 43.16 6.555 43.33 6.725 ;
      RECT 42.14 2.815 42.31 2.985 ;
      RECT 42.14 4.855 42.31 5.025 ;
      RECT 41.63 3.495 41.8 3.665 ;
      RECT 39.89 7.675 40.06 7.845 ;
      RECT 39.46 8.045 39.63 8.215 ;
      RECT 39.46 8.785 39.63 8.955 ;
      RECT 36.705 7.31 36.875 7.48 ;
      RECT 36.705 8.79 36.875 8.96 ;
      RECT 36.335 2.76 36.505 2.93 ;
      RECT 36.335 6.94 36.505 7.11 ;
      RECT 35.715 0.91 35.885 1.08 ;
      RECT 35.715 2.39 35.885 2.56 ;
      RECT 35.715 7.31 35.885 7.48 ;
      RECT 35.715 8.79 35.885 8.96 ;
      RECT 35.345 2.76 35.515 2.93 ;
      RECT 35.345 6.94 35.515 7.11 ;
      RECT 34.355 2.025 34.525 2.195 ;
      RECT 34.355 7.675 34.525 7.845 ;
      RECT 33.925 0.915 34.095 1.085 ;
      RECT 33.925 1.655 34.095 1.825 ;
      RECT 33.925 8.045 34.095 8.215 ;
      RECT 33.925 8.785 34.095 8.955 ;
      RECT 33.55 2.395 33.72 2.565 ;
      RECT 33.55 7.305 33.72 7.475 ;
      RECT 30.36 3.835 30.53 4.005 ;
      RECT 30.36 5.875 30.53 6.045 ;
      RECT 30.02 2.815 30.19 2.985 ;
      RECT 29.68 6.555 29.85 6.725 ;
      RECT 29.51 5.875 29.68 6.045 ;
      RECT 29 5.875 29.17 6.045 ;
      RECT 28.32 3.155 28.49 3.325 ;
      RECT 28.32 6.555 28.49 6.725 ;
      RECT 27.64 2.815 27.81 2.985 ;
      RECT 27.63 5.875 27.8 6.045 ;
      RECT 27.18 4.855 27.35 5.025 ;
      RECT 27.16 2.305 27.33 2.475 ;
      RECT 26.79 2.82 26.96 2.99 ;
      RECT 26.28 2.82 26.45 2.99 ;
      RECT 26.28 3.835 26.45 4.005 ;
      RECT 25.94 6.555 26.11 6.725 ;
      RECT 24.92 2.815 25.09 2.985 ;
      RECT 24.92 4.855 25.09 5.025 ;
      RECT 24.41 3.495 24.58 3.665 ;
      RECT 22.67 7.675 22.84 7.845 ;
      RECT 22.24 8.045 22.41 8.215 ;
      RECT 22.24 8.785 22.41 8.955 ;
      RECT 19.485 7.31 19.655 7.48 ;
      RECT 19.485 8.79 19.655 8.96 ;
      RECT 19.115 2.76 19.285 2.93 ;
      RECT 19.115 6.94 19.285 7.11 ;
      RECT 18.495 0.91 18.665 1.08 ;
      RECT 18.495 2.39 18.665 2.56 ;
      RECT 18.495 7.31 18.665 7.48 ;
      RECT 18.495 8.79 18.665 8.96 ;
      RECT 18.125 2.76 18.295 2.93 ;
      RECT 18.125 6.94 18.295 7.11 ;
      RECT 17.135 2.025 17.305 2.195 ;
      RECT 17.135 7.675 17.305 7.845 ;
      RECT 16.705 0.915 16.875 1.085 ;
      RECT 16.705 1.655 16.875 1.825 ;
      RECT 16.705 8.045 16.875 8.215 ;
      RECT 16.705 8.785 16.875 8.955 ;
      RECT 16.33 2.395 16.5 2.565 ;
      RECT 16.33 7.305 16.5 7.475 ;
      RECT 13.14 3.835 13.31 4.005 ;
      RECT 13.14 5.875 13.31 6.045 ;
      RECT 12.8 2.815 12.97 2.985 ;
      RECT 12.46 6.555 12.63 6.725 ;
      RECT 12.29 5.875 12.46 6.045 ;
      RECT 11.78 5.875 11.95 6.045 ;
      RECT 11.1 3.155 11.27 3.325 ;
      RECT 11.1 6.555 11.27 6.725 ;
      RECT 10.42 2.815 10.59 2.985 ;
      RECT 10.41 5.875 10.58 6.045 ;
      RECT 9.96 4.855 10.13 5.025 ;
      RECT 9.94 2.305 10.11 2.475 ;
      RECT 9.57 2.82 9.74 2.99 ;
      RECT 9.06 2.82 9.23 2.99 ;
      RECT 9.06 3.835 9.23 4.005 ;
      RECT 8.72 6.555 8.89 6.725 ;
      RECT 7.7 2.815 7.87 2.985 ;
      RECT 7.7 4.855 7.87 5.025 ;
      RECT 7.19 3.495 7.36 3.665 ;
      RECT 5.45 7.675 5.62 7.845 ;
      RECT 5.02 8.045 5.19 8.215 ;
      RECT 5.02 8.785 5.19 8.955 ;
      RECT 1.61 8.045 1.78 8.215 ;
      RECT 1.61 8.785 1.78 8.955 ;
      RECT 1.235 7.305 1.405 7.475 ;
    LAYER li1 ;
      RECT 87.995 1.74 88.165 2.93 ;
      RECT 87.995 1.74 88.465 1.91 ;
      RECT 87.995 7.96 88.465 8.13 ;
      RECT 87.995 6.94 88.165 8.13 ;
      RECT 87.005 1.74 87.175 2.93 ;
      RECT 87.005 1.74 87.475 1.91 ;
      RECT 87.005 7.96 87.475 8.13 ;
      RECT 87.005 6.94 87.175 8.13 ;
      RECT 85.155 2.635 85.325 3.865 ;
      RECT 85.21 0.855 85.38 2.805 ;
      RECT 85.155 0.575 85.325 1.025 ;
      RECT 85.155 8.845 85.325 9.295 ;
      RECT 85.21 7.065 85.38 9.015 ;
      RECT 85.155 6.005 85.325 7.235 ;
      RECT 84.635 0.575 84.805 3.865 ;
      RECT 84.635 2.075 85.04 2.405 ;
      RECT 84.635 1.235 85.04 1.565 ;
      RECT 84.635 6.005 84.805 9.295 ;
      RECT 84.635 8.305 85.04 8.635 ;
      RECT 84.635 7.465 85.04 7.795 ;
      RECT 82.37 3.495 82.75 4.175 ;
      RECT 82.58 2.365 82.75 4.175 ;
      RECT 80.5 2.365 80.73 3.035 ;
      RECT 80.5 2.365 82.75 2.535 ;
      RECT 82.03 2.045 82.2 2.535 ;
      RECT 82.02 3.155 82.19 4.005 ;
      RECT 81.105 3.155 82.41 3.325 ;
      RECT 82.165 2.705 82.41 3.325 ;
      RECT 81.105 2.785 81.275 3.325 ;
      RECT 80.9 2.785 81.275 2.955 ;
      RECT 81.08 6.265 81.775 6.895 ;
      RECT 81.605 4.685 81.775 6.895 ;
      RECT 81.51 4.685 81.84 5.665 ;
      RECT 81.11 3.495 81.44 4.175 ;
      RECT 80.2 3.495 80.6 4.175 ;
      RECT 80.2 3.495 81.44 3.665 ;
      RECT 79.7 3.075 80.02 4.175 ;
      RECT 79.7 3.075 80.15 3.325 ;
      RECT 79.7 3.075 80.33 3.245 ;
      RECT 80.16 2.025 80.33 3.245 ;
      RECT 80.16 2.025 81.115 2.195 ;
      RECT 79.7 6.265 80.395 6.895 ;
      RECT 80.225 4.685 80.395 6.895 ;
      RECT 80.13 4.685 80.46 5.665 ;
      RECT 79.72 5.825 80.055 6.075 ;
      RECT 79.175 5.825 79.51 6.075 ;
      RECT 79.175 5.875 80.055 6.045 ;
      RECT 78.835 6.265 79.53 6.895 ;
      RECT 78.835 4.685 79.005 6.895 ;
      RECT 78.77 4.685 79.1 5.665 ;
      RECT 78.33 3.205 78.66 4.16 ;
      RECT 78.33 3.205 79.01 3.375 ;
      RECT 78.84 1.965 79.01 3.375 ;
      RECT 78.75 1.965 79.08 2.605 ;
      RECT 77.81 3.205 78.14 4.16 ;
      RECT 77.46 3.205 78.14 3.375 ;
      RECT 77.46 1.965 77.63 3.375 ;
      RECT 77.39 1.965 77.72 2.605 ;
      RECT 77.6 5.875 77.77 6.725 ;
      RECT 76.875 5.825 77.21 6.075 ;
      RECT 76.875 5.875 77.77 6.045 ;
      RECT 76.94 2.785 77.29 3.035 ;
      RECT 76.42 2.785 76.75 3.035 ;
      RECT 76.42 2.815 77.29 2.985 ;
      RECT 76.535 6.265 77.23 6.895 ;
      RECT 76.535 4.685 76.705 6.895 ;
      RECT 76.47 4.685 76.8 5.665 ;
      RECT 76 3.195 76.33 4.175 ;
      RECT 76 1.965 76.25 4.175 ;
      RECT 76 1.965 76.33 2.595 ;
      RECT 72.95 6.005 73.12 9.295 ;
      RECT 72.95 8.305 73.355 8.635 ;
      RECT 72.95 7.465 73.355 7.795 ;
      RECT 70.775 1.74 70.945 2.93 ;
      RECT 70.775 1.74 71.245 1.91 ;
      RECT 70.775 7.96 71.245 8.13 ;
      RECT 70.775 6.94 70.945 8.13 ;
      RECT 69.785 1.74 69.955 2.93 ;
      RECT 69.785 1.74 70.255 1.91 ;
      RECT 69.785 7.96 70.255 8.13 ;
      RECT 69.785 6.94 69.955 8.13 ;
      RECT 67.935 2.635 68.105 3.865 ;
      RECT 67.99 0.855 68.16 2.805 ;
      RECT 67.935 0.575 68.105 1.025 ;
      RECT 67.935 8.845 68.105 9.295 ;
      RECT 67.99 7.065 68.16 9.015 ;
      RECT 67.935 6.005 68.105 7.235 ;
      RECT 67.415 0.575 67.585 3.865 ;
      RECT 67.415 2.075 67.82 2.405 ;
      RECT 67.415 1.235 67.82 1.565 ;
      RECT 67.415 6.005 67.585 9.295 ;
      RECT 67.415 8.305 67.82 8.635 ;
      RECT 67.415 7.465 67.82 7.795 ;
      RECT 65.15 3.495 65.53 4.175 ;
      RECT 65.36 2.365 65.53 4.175 ;
      RECT 63.28 2.365 63.51 3.035 ;
      RECT 63.28 2.365 65.53 2.535 ;
      RECT 64.81 2.045 64.98 2.535 ;
      RECT 64.8 3.155 64.97 4.005 ;
      RECT 63.885 3.155 65.19 3.325 ;
      RECT 64.945 2.705 65.19 3.325 ;
      RECT 63.885 2.785 64.055 3.325 ;
      RECT 63.68 2.785 64.055 2.955 ;
      RECT 63.86 6.265 64.555 6.895 ;
      RECT 64.385 4.685 64.555 6.895 ;
      RECT 64.29 4.685 64.62 5.665 ;
      RECT 63.89 3.495 64.22 4.175 ;
      RECT 62.98 3.495 63.38 4.175 ;
      RECT 62.98 3.495 64.22 3.665 ;
      RECT 62.48 3.075 62.8 4.175 ;
      RECT 62.48 3.075 62.93 3.325 ;
      RECT 62.48 3.075 63.11 3.245 ;
      RECT 62.94 2.025 63.11 3.245 ;
      RECT 62.94 2.025 63.895 2.195 ;
      RECT 62.48 6.265 63.175 6.895 ;
      RECT 63.005 4.685 63.175 6.895 ;
      RECT 62.91 4.685 63.24 5.665 ;
      RECT 62.5 5.825 62.835 6.075 ;
      RECT 61.955 5.825 62.29 6.075 ;
      RECT 61.955 5.875 62.835 6.045 ;
      RECT 61.615 6.265 62.31 6.895 ;
      RECT 61.615 4.685 61.785 6.895 ;
      RECT 61.55 4.685 61.88 5.665 ;
      RECT 61.11 3.205 61.44 4.16 ;
      RECT 61.11 3.205 61.79 3.375 ;
      RECT 61.62 1.965 61.79 3.375 ;
      RECT 61.53 1.965 61.86 2.605 ;
      RECT 60.59 3.205 60.92 4.16 ;
      RECT 60.24 3.205 60.92 3.375 ;
      RECT 60.24 1.965 60.41 3.375 ;
      RECT 60.17 1.965 60.5 2.605 ;
      RECT 60.38 5.875 60.55 6.725 ;
      RECT 59.655 5.825 59.99 6.075 ;
      RECT 59.655 5.875 60.55 6.045 ;
      RECT 59.72 2.785 60.07 3.035 ;
      RECT 59.2 2.785 59.53 3.035 ;
      RECT 59.2 2.815 60.07 2.985 ;
      RECT 59.315 6.265 60.01 6.895 ;
      RECT 59.315 4.685 59.485 6.895 ;
      RECT 59.25 4.685 59.58 5.665 ;
      RECT 58.78 3.195 59.11 4.175 ;
      RECT 58.78 1.965 59.03 4.175 ;
      RECT 58.78 1.965 59.11 2.595 ;
      RECT 55.73 6.005 55.9 9.295 ;
      RECT 55.73 8.305 56.135 8.635 ;
      RECT 55.73 7.465 56.135 7.795 ;
      RECT 53.555 1.74 53.725 2.93 ;
      RECT 53.555 1.74 54.025 1.91 ;
      RECT 53.555 7.96 54.025 8.13 ;
      RECT 53.555 6.94 53.725 8.13 ;
      RECT 52.565 1.74 52.735 2.93 ;
      RECT 52.565 1.74 53.035 1.91 ;
      RECT 52.565 7.96 53.035 8.13 ;
      RECT 52.565 6.94 52.735 8.13 ;
      RECT 50.715 2.635 50.885 3.865 ;
      RECT 50.77 0.855 50.94 2.805 ;
      RECT 50.715 0.575 50.885 1.025 ;
      RECT 50.715 8.845 50.885 9.295 ;
      RECT 50.77 7.065 50.94 9.015 ;
      RECT 50.715 6.005 50.885 7.235 ;
      RECT 50.195 0.575 50.365 3.865 ;
      RECT 50.195 2.075 50.6 2.405 ;
      RECT 50.195 1.235 50.6 1.565 ;
      RECT 50.195 6.005 50.365 9.295 ;
      RECT 50.195 8.305 50.6 8.635 ;
      RECT 50.195 7.465 50.6 7.795 ;
      RECT 47.93 3.495 48.31 4.175 ;
      RECT 48.14 2.365 48.31 4.175 ;
      RECT 46.06 2.365 46.29 3.035 ;
      RECT 46.06 2.365 48.31 2.535 ;
      RECT 47.59 2.045 47.76 2.535 ;
      RECT 47.58 3.155 47.75 4.005 ;
      RECT 46.665 3.155 47.97 3.325 ;
      RECT 47.725 2.705 47.97 3.325 ;
      RECT 46.665 2.785 46.835 3.325 ;
      RECT 46.46 2.785 46.835 2.955 ;
      RECT 46.64 6.265 47.335 6.895 ;
      RECT 47.165 4.685 47.335 6.895 ;
      RECT 47.07 4.685 47.4 5.665 ;
      RECT 46.67 3.495 47 4.175 ;
      RECT 45.76 3.495 46.16 4.175 ;
      RECT 45.76 3.495 47 3.665 ;
      RECT 45.26 3.075 45.58 4.175 ;
      RECT 45.26 3.075 45.71 3.325 ;
      RECT 45.26 3.075 45.89 3.245 ;
      RECT 45.72 2.025 45.89 3.245 ;
      RECT 45.72 2.025 46.675 2.195 ;
      RECT 45.26 6.265 45.955 6.895 ;
      RECT 45.785 4.685 45.955 6.895 ;
      RECT 45.69 4.685 46.02 5.665 ;
      RECT 45.28 5.825 45.615 6.075 ;
      RECT 44.735 5.825 45.07 6.075 ;
      RECT 44.735 5.875 45.615 6.045 ;
      RECT 44.395 6.265 45.09 6.895 ;
      RECT 44.395 4.685 44.565 6.895 ;
      RECT 44.33 4.685 44.66 5.665 ;
      RECT 43.89 3.205 44.22 4.16 ;
      RECT 43.89 3.205 44.57 3.375 ;
      RECT 44.4 1.965 44.57 3.375 ;
      RECT 44.31 1.965 44.64 2.605 ;
      RECT 43.37 3.205 43.7 4.16 ;
      RECT 43.02 3.205 43.7 3.375 ;
      RECT 43.02 1.965 43.19 3.375 ;
      RECT 42.95 1.965 43.28 2.605 ;
      RECT 43.16 5.875 43.33 6.725 ;
      RECT 42.435 5.825 42.77 6.075 ;
      RECT 42.435 5.875 43.33 6.045 ;
      RECT 42.5 2.785 42.85 3.035 ;
      RECT 41.98 2.785 42.31 3.035 ;
      RECT 41.98 2.815 42.85 2.985 ;
      RECT 42.095 6.265 42.79 6.895 ;
      RECT 42.095 4.685 42.265 6.895 ;
      RECT 42.03 4.685 42.36 5.665 ;
      RECT 41.56 3.195 41.89 4.175 ;
      RECT 41.56 1.965 41.81 4.175 ;
      RECT 41.56 1.965 41.89 2.595 ;
      RECT 38.51 6.005 38.68 9.295 ;
      RECT 38.51 8.305 38.915 8.635 ;
      RECT 38.51 7.465 38.915 7.795 ;
      RECT 36.335 1.74 36.505 2.93 ;
      RECT 36.335 1.74 36.805 1.91 ;
      RECT 36.335 7.96 36.805 8.13 ;
      RECT 36.335 6.94 36.505 8.13 ;
      RECT 35.345 1.74 35.515 2.93 ;
      RECT 35.345 1.74 35.815 1.91 ;
      RECT 35.345 7.96 35.815 8.13 ;
      RECT 35.345 6.94 35.515 8.13 ;
      RECT 33.495 2.635 33.665 3.865 ;
      RECT 33.55 0.855 33.72 2.805 ;
      RECT 33.495 0.575 33.665 1.025 ;
      RECT 33.495 8.845 33.665 9.295 ;
      RECT 33.55 7.065 33.72 9.015 ;
      RECT 33.495 6.005 33.665 7.235 ;
      RECT 32.975 0.575 33.145 3.865 ;
      RECT 32.975 2.075 33.38 2.405 ;
      RECT 32.975 1.235 33.38 1.565 ;
      RECT 32.975 6.005 33.145 9.295 ;
      RECT 32.975 8.305 33.38 8.635 ;
      RECT 32.975 7.465 33.38 7.795 ;
      RECT 30.71 3.495 31.09 4.175 ;
      RECT 30.92 2.365 31.09 4.175 ;
      RECT 28.84 2.365 29.07 3.035 ;
      RECT 28.84 2.365 31.09 2.535 ;
      RECT 30.37 2.045 30.54 2.535 ;
      RECT 30.36 3.155 30.53 4.005 ;
      RECT 29.445 3.155 30.75 3.325 ;
      RECT 30.505 2.705 30.75 3.325 ;
      RECT 29.445 2.785 29.615 3.325 ;
      RECT 29.24 2.785 29.615 2.955 ;
      RECT 29.42 6.265 30.115 6.895 ;
      RECT 29.945 4.685 30.115 6.895 ;
      RECT 29.85 4.685 30.18 5.665 ;
      RECT 29.45 3.495 29.78 4.175 ;
      RECT 28.54 3.495 28.94 4.175 ;
      RECT 28.54 3.495 29.78 3.665 ;
      RECT 28.04 3.075 28.36 4.175 ;
      RECT 28.04 3.075 28.49 3.325 ;
      RECT 28.04 3.075 28.67 3.245 ;
      RECT 28.5 2.025 28.67 3.245 ;
      RECT 28.5 2.025 29.455 2.195 ;
      RECT 28.04 6.265 28.735 6.895 ;
      RECT 28.565 4.685 28.735 6.895 ;
      RECT 28.47 4.685 28.8 5.665 ;
      RECT 28.06 5.825 28.395 6.075 ;
      RECT 27.515 5.825 27.85 6.075 ;
      RECT 27.515 5.875 28.395 6.045 ;
      RECT 27.175 6.265 27.87 6.895 ;
      RECT 27.175 4.685 27.345 6.895 ;
      RECT 27.11 4.685 27.44 5.665 ;
      RECT 26.67 3.205 27 4.16 ;
      RECT 26.67 3.205 27.35 3.375 ;
      RECT 27.18 1.965 27.35 3.375 ;
      RECT 27.09 1.965 27.42 2.605 ;
      RECT 26.15 3.205 26.48 4.16 ;
      RECT 25.8 3.205 26.48 3.375 ;
      RECT 25.8 1.965 25.97 3.375 ;
      RECT 25.73 1.965 26.06 2.605 ;
      RECT 25.94 5.875 26.11 6.725 ;
      RECT 25.215 5.825 25.55 6.075 ;
      RECT 25.215 5.875 26.11 6.045 ;
      RECT 25.28 2.785 25.63 3.035 ;
      RECT 24.76 2.785 25.09 3.035 ;
      RECT 24.76 2.815 25.63 2.985 ;
      RECT 24.875 6.265 25.57 6.895 ;
      RECT 24.875 4.685 25.045 6.895 ;
      RECT 24.81 4.685 25.14 5.665 ;
      RECT 24.34 3.195 24.67 4.175 ;
      RECT 24.34 1.965 24.59 4.175 ;
      RECT 24.34 1.965 24.67 2.595 ;
      RECT 21.29 6.005 21.46 9.295 ;
      RECT 21.29 8.305 21.695 8.635 ;
      RECT 21.29 7.465 21.695 7.795 ;
      RECT 19.115 1.74 19.285 2.93 ;
      RECT 19.115 1.74 19.585 1.91 ;
      RECT 19.115 7.96 19.585 8.13 ;
      RECT 19.115 6.94 19.285 8.13 ;
      RECT 18.125 1.74 18.295 2.93 ;
      RECT 18.125 1.74 18.595 1.91 ;
      RECT 18.125 7.96 18.595 8.13 ;
      RECT 18.125 6.94 18.295 8.13 ;
      RECT 16.275 2.635 16.445 3.865 ;
      RECT 16.33 0.855 16.5 2.805 ;
      RECT 16.275 0.575 16.445 1.025 ;
      RECT 16.275 8.845 16.445 9.295 ;
      RECT 16.33 7.065 16.5 9.015 ;
      RECT 16.275 6.005 16.445 7.235 ;
      RECT 15.755 0.575 15.925 3.865 ;
      RECT 15.755 2.075 16.16 2.405 ;
      RECT 15.755 1.235 16.16 1.565 ;
      RECT 15.755 6.005 15.925 9.295 ;
      RECT 15.755 8.305 16.16 8.635 ;
      RECT 15.755 7.465 16.16 7.795 ;
      RECT 13.49 3.495 13.87 4.175 ;
      RECT 13.7 2.365 13.87 4.175 ;
      RECT 11.62 2.365 11.85 3.035 ;
      RECT 11.62 2.365 13.87 2.535 ;
      RECT 13.15 2.045 13.32 2.535 ;
      RECT 13.14 3.155 13.31 4.005 ;
      RECT 12.225 3.155 13.53 3.325 ;
      RECT 13.285 2.705 13.53 3.325 ;
      RECT 12.225 2.785 12.395 3.325 ;
      RECT 12.02 2.785 12.395 2.955 ;
      RECT 12.2 6.265 12.895 6.895 ;
      RECT 12.725 4.685 12.895 6.895 ;
      RECT 12.63 4.685 12.96 5.665 ;
      RECT 12.23 3.495 12.56 4.175 ;
      RECT 11.32 3.495 11.72 4.175 ;
      RECT 11.32 3.495 12.56 3.665 ;
      RECT 10.82 3.075 11.14 4.175 ;
      RECT 10.82 3.075 11.27 3.325 ;
      RECT 10.82 3.075 11.45 3.245 ;
      RECT 11.28 2.025 11.45 3.245 ;
      RECT 11.28 2.025 12.235 2.195 ;
      RECT 10.82 6.265 11.515 6.895 ;
      RECT 11.345 4.685 11.515 6.895 ;
      RECT 11.25 4.685 11.58 5.665 ;
      RECT 10.84 5.825 11.175 6.075 ;
      RECT 10.295 5.825 10.63 6.075 ;
      RECT 10.295 5.875 11.175 6.045 ;
      RECT 9.955 6.265 10.65 6.895 ;
      RECT 9.955 4.685 10.125 6.895 ;
      RECT 9.89 4.685 10.22 5.665 ;
      RECT 9.45 3.205 9.78 4.16 ;
      RECT 9.45 3.205 10.13 3.375 ;
      RECT 9.96 1.965 10.13 3.375 ;
      RECT 9.87 1.965 10.2 2.605 ;
      RECT 8.93 3.205 9.26 4.16 ;
      RECT 8.58 3.205 9.26 3.375 ;
      RECT 8.58 1.965 8.75 3.375 ;
      RECT 8.51 1.965 8.84 2.605 ;
      RECT 8.72 5.875 8.89 6.725 ;
      RECT 7.995 5.825 8.33 6.075 ;
      RECT 7.995 5.875 8.89 6.045 ;
      RECT 8.06 2.785 8.41 3.035 ;
      RECT 7.54 2.785 7.87 3.035 ;
      RECT 7.54 2.815 8.41 2.985 ;
      RECT 7.655 6.265 8.35 6.895 ;
      RECT 7.655 4.685 7.825 6.895 ;
      RECT 7.59 4.685 7.92 5.665 ;
      RECT 7.12 3.195 7.45 4.175 ;
      RECT 7.12 1.965 7.37 4.175 ;
      RECT 7.12 1.965 7.45 2.595 ;
      RECT 4.07 6.005 4.24 9.295 ;
      RECT 4.07 8.305 4.475 8.635 ;
      RECT 4.07 7.465 4.475 7.795 ;
      RECT 1.18 8.845 1.35 9.295 ;
      RECT 1.235 7.065 1.405 9.015 ;
      RECT 1.18 6.005 1.35 7.235 ;
      RECT 0.66 6.005 0.83 9.295 ;
      RECT 0.66 8.305 1.065 8.635 ;
      RECT 0.66 7.465 1.065 7.795 ;
      RECT 88.365 6.01 88.535 7.48 ;
      RECT 88.365 8.79 88.535 9.3 ;
      RECT 87.375 0.57 87.545 1.08 ;
      RECT 87.375 2.39 87.545 3.86 ;
      RECT 87.375 6.01 87.545 7.48 ;
      RECT 87.375 8.79 87.545 9.3 ;
      RECT 86.015 0.575 86.185 3.865 ;
      RECT 86.015 6.005 86.185 9.295 ;
      RECT 85.585 0.575 85.755 1.085 ;
      RECT 85.585 1.655 85.755 3.865 ;
      RECT 85.585 6.005 85.755 8.215 ;
      RECT 85.585 8.785 85.755 9.295 ;
      RECT 81.945 5.825 82.28 6.095 ;
      RECT 81.445 2.785 81.995 2.985 ;
      RECT 81.1 5.825 81.435 6.075 ;
      RECT 80.565 5.825 80.9 6.095 ;
      RECT 79.18 2.785 79.53 3.035 ;
      RECT 78.32 2.785 78.67 3.035 ;
      RECT 77.8 2.785 78.15 3.035 ;
      RECT 74.33 6.005 74.5 9.295 ;
      RECT 73.9 6.005 74.07 8.215 ;
      RECT 73.9 8.785 74.07 9.295 ;
      RECT 71.145 6.01 71.315 7.48 ;
      RECT 71.145 8.79 71.315 9.3 ;
      RECT 70.155 0.57 70.325 1.08 ;
      RECT 70.155 2.39 70.325 3.86 ;
      RECT 70.155 6.01 70.325 7.48 ;
      RECT 70.155 8.79 70.325 9.3 ;
      RECT 68.795 0.575 68.965 3.865 ;
      RECT 68.795 6.005 68.965 9.295 ;
      RECT 68.365 0.575 68.535 1.085 ;
      RECT 68.365 1.655 68.535 3.865 ;
      RECT 68.365 6.005 68.535 8.215 ;
      RECT 68.365 8.785 68.535 9.295 ;
      RECT 64.725 5.825 65.06 6.095 ;
      RECT 64.225 2.785 64.775 2.985 ;
      RECT 63.88 5.825 64.215 6.075 ;
      RECT 63.345 5.825 63.68 6.095 ;
      RECT 61.96 2.785 62.31 3.035 ;
      RECT 61.1 2.785 61.45 3.035 ;
      RECT 60.58 2.785 60.93 3.035 ;
      RECT 57.11 6.005 57.28 9.295 ;
      RECT 56.68 6.005 56.85 8.215 ;
      RECT 56.68 8.785 56.85 9.295 ;
      RECT 53.925 6.01 54.095 7.48 ;
      RECT 53.925 8.79 54.095 9.3 ;
      RECT 52.935 0.57 53.105 1.08 ;
      RECT 52.935 2.39 53.105 3.86 ;
      RECT 52.935 6.01 53.105 7.48 ;
      RECT 52.935 8.79 53.105 9.3 ;
      RECT 51.575 0.575 51.745 3.865 ;
      RECT 51.575 6.005 51.745 9.295 ;
      RECT 51.145 0.575 51.315 1.085 ;
      RECT 51.145 1.655 51.315 3.865 ;
      RECT 51.145 6.005 51.315 8.215 ;
      RECT 51.145 8.785 51.315 9.295 ;
      RECT 47.505 5.825 47.84 6.095 ;
      RECT 47.005 2.785 47.555 2.985 ;
      RECT 46.66 5.825 46.995 6.075 ;
      RECT 46.125 5.825 46.46 6.095 ;
      RECT 44.74 2.785 45.09 3.035 ;
      RECT 43.88 2.785 44.23 3.035 ;
      RECT 43.36 2.785 43.71 3.035 ;
      RECT 39.89 6.005 40.06 9.295 ;
      RECT 39.46 6.005 39.63 8.215 ;
      RECT 39.46 8.785 39.63 9.295 ;
      RECT 36.705 6.01 36.875 7.48 ;
      RECT 36.705 8.79 36.875 9.3 ;
      RECT 35.715 0.57 35.885 1.08 ;
      RECT 35.715 2.39 35.885 3.86 ;
      RECT 35.715 6.01 35.885 7.48 ;
      RECT 35.715 8.79 35.885 9.3 ;
      RECT 34.355 0.575 34.525 3.865 ;
      RECT 34.355 6.005 34.525 9.295 ;
      RECT 33.925 0.575 34.095 1.085 ;
      RECT 33.925 1.655 34.095 3.865 ;
      RECT 33.925 6.005 34.095 8.215 ;
      RECT 33.925 8.785 34.095 9.295 ;
      RECT 30.285 5.825 30.62 6.095 ;
      RECT 29.785 2.785 30.335 2.985 ;
      RECT 29.44 5.825 29.775 6.075 ;
      RECT 28.905 5.825 29.24 6.095 ;
      RECT 27.52 2.785 27.87 3.035 ;
      RECT 26.66 2.785 27.01 3.035 ;
      RECT 26.14 2.785 26.49 3.035 ;
      RECT 22.67 6.005 22.84 9.295 ;
      RECT 22.24 6.005 22.41 8.215 ;
      RECT 22.24 8.785 22.41 9.295 ;
      RECT 19.485 6.01 19.655 7.48 ;
      RECT 19.485 8.79 19.655 9.3 ;
      RECT 18.495 0.57 18.665 1.08 ;
      RECT 18.495 2.39 18.665 3.86 ;
      RECT 18.495 6.01 18.665 7.48 ;
      RECT 18.495 8.79 18.665 9.3 ;
      RECT 17.135 0.575 17.305 3.865 ;
      RECT 17.135 6.005 17.305 9.295 ;
      RECT 16.705 0.575 16.875 1.085 ;
      RECT 16.705 1.655 16.875 3.865 ;
      RECT 16.705 6.005 16.875 8.215 ;
      RECT 16.705 8.785 16.875 9.295 ;
      RECT 13.065 5.825 13.4 6.095 ;
      RECT 12.565 2.785 13.115 2.985 ;
      RECT 12.22 5.825 12.555 6.075 ;
      RECT 11.685 5.825 12.02 6.095 ;
      RECT 10.3 2.785 10.65 3.035 ;
      RECT 9.44 2.785 9.79 3.035 ;
      RECT 8.92 2.785 9.27 3.035 ;
      RECT 5.45 6.005 5.62 9.295 ;
      RECT 5.02 6.005 5.19 8.215 ;
      RECT 5.02 8.785 5.19 9.295 ;
      RECT 1.61 6.005 1.78 8.215 ;
      RECT 1.61 8.785 1.78 9.295 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r2 ;
  SIZE 88.92 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 19.48 1.865 19.65 2.375 ;
        RECT 19.48 3.685 19.65 5.155 ;
      LAYER met1 ;
        RECT 19.42 3.655 19.71 3.885 ;
        RECT 19.42 2.175 19.71 2.405 ;
        RECT 19.48 2.175 19.65 3.885 ;
      LAYER mcon ;
        RECT 19.48 3.685 19.65 3.855 ;
        RECT 19.48 2.205 19.65 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 36.7 1.865 36.87 2.375 ;
        RECT 36.7 3.685 36.87 5.155 ;
      LAYER met1 ;
        RECT 36.64 3.655 36.93 3.885 ;
        RECT 36.64 2.175 36.93 2.405 ;
        RECT 36.7 2.175 36.87 3.885 ;
      LAYER mcon ;
        RECT 36.7 3.685 36.87 3.855 ;
        RECT 36.7 2.205 36.87 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 53.92 1.865 54.09 2.375 ;
        RECT 53.92 3.685 54.09 5.155 ;
      LAYER met1 ;
        RECT 53.86 3.655 54.15 3.885 ;
        RECT 53.86 2.175 54.15 2.405 ;
        RECT 53.92 2.175 54.09 3.885 ;
      LAYER mcon ;
        RECT 53.92 3.685 54.09 3.855 ;
        RECT 53.92 2.205 54.09 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 71.14 1.865 71.31 2.375 ;
        RECT 71.14 3.685 71.31 5.155 ;
      LAYER met1 ;
        RECT 71.08 3.655 71.37 3.885 ;
        RECT 71.08 2.175 71.37 2.405 ;
        RECT 71.14 3.2 71.315 3.37 ;
        RECT 71.14 2.175 71.31 3.885 ;
      LAYER mcon ;
        RECT 71.14 3.685 71.31 3.855 ;
        RECT 71.14 2.205 71.31 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 88.36 1.865 88.53 2.375 ;
        RECT 88.36 3.685 88.53 5.155 ;
      LAYER met1 ;
        RECT 88.3 3.655 88.59 3.885 ;
        RECT 88.3 2.175 88.59 2.405 ;
        RECT 88.36 2.175 88.53 3.885 ;
      LAYER mcon ;
        RECT 88.36 3.685 88.53 3.855 ;
        RECT 88.36 2.205 88.53 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.33 2.955 15.5 4.23 ;
        RECT 15.33 8.225 15.5 9.505 ;
        RECT 15.32 8.225 15.5 8.465 ;
        RECT 3.645 8.23 3.815 9.505 ;
      LAYER met2 ;
        RECT 15.25 8.14 15.575 8.465 ;
        RECT 15.25 4.79 15.575 5.115 ;
        RECT 5.95 9.24 15.5 9.41 ;
        RECT 15.33 8.14 15.5 9.41 ;
        RECT 15.32 4.79 15.49 8.465 ;
        RECT 5.895 8.145 6.175 8.485 ;
        RECT 5.95 8.145 6.12 9.41 ;
      LAYER met1 ;
        RECT 15.27 4.06 15.73 4.23 ;
        RECT 15.25 4.79 15.575 5.115 ;
        RECT 15.27 4.03 15.56 4.26 ;
        RECT 15.33 4.03 15.5 5.115 ;
        RECT 15.25 8.23 15.73 8.4 ;
        RECT 15.25 8.14 15.575 8.465 ;
        RECT 5.865 8.175 6.205 8.455 ;
        RECT 3.585 8.23 6.205 8.4 ;
        RECT 3.585 8.2 3.875 8.43 ;
      LAYER via1 ;
        RECT 5.96 8.24 6.11 8.39 ;
        RECT 15.34 8.225 15.49 8.375 ;
        RECT 15.34 4.875 15.49 5.025 ;
      LAYER mcon ;
        RECT 3.645 8.23 3.815 8.4 ;
        RECT 15.33 8.23 15.5 8.4 ;
        RECT 15.33 4.06 15.5 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 32.55 2.955 32.72 4.23 ;
        RECT 32.55 8.225 32.72 9.505 ;
        RECT 32.54 8.225 32.72 8.465 ;
        RECT 20.865 8.23 21.035 9.505 ;
      LAYER met2 ;
        RECT 32.47 8.14 32.795 8.465 ;
        RECT 32.47 4.79 32.795 5.115 ;
        RECT 23.17 9.24 32.72 9.41 ;
        RECT 32.55 8.14 32.72 9.41 ;
        RECT 32.54 4.79 32.71 8.465 ;
        RECT 23.115 8.145 23.395 8.485 ;
        RECT 23.17 8.145 23.34 9.41 ;
      LAYER met1 ;
        RECT 32.49 4.06 32.95 4.23 ;
        RECT 32.47 4.79 32.795 5.115 ;
        RECT 32.49 4.03 32.78 4.26 ;
        RECT 32.55 4.03 32.72 5.115 ;
        RECT 32.47 8.23 32.95 8.4 ;
        RECT 32.47 8.14 32.795 8.465 ;
        RECT 23.085 8.175 23.425 8.455 ;
        RECT 20.805 8.23 23.425 8.4 ;
        RECT 20.805 8.2 21.095 8.43 ;
      LAYER via1 ;
        RECT 23.18 8.24 23.33 8.39 ;
        RECT 32.56 8.225 32.71 8.375 ;
        RECT 32.56 4.875 32.71 5.025 ;
      LAYER mcon ;
        RECT 20.865 8.23 21.035 8.4 ;
        RECT 32.55 8.23 32.72 8.4 ;
        RECT 32.55 4.06 32.72 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 49.77 2.955 49.94 4.23 ;
        RECT 49.77 8.225 49.94 9.505 ;
        RECT 49.76 8.225 49.94 8.465 ;
        RECT 38.085 8.23 38.255 9.505 ;
      LAYER met2 ;
        RECT 49.69 8.14 50.015 8.465 ;
        RECT 49.69 4.79 50.015 5.115 ;
        RECT 40.39 9.24 49.94 9.41 ;
        RECT 49.77 8.14 49.94 9.41 ;
        RECT 49.76 4.79 49.93 8.465 ;
        RECT 40.335 8.145 40.615 8.485 ;
        RECT 40.39 8.145 40.56 9.41 ;
      LAYER met1 ;
        RECT 49.71 4.06 50.17 4.23 ;
        RECT 49.69 4.79 50.015 5.115 ;
        RECT 49.71 4.03 50 4.26 ;
        RECT 49.77 4.03 49.94 5.115 ;
        RECT 49.69 8.23 50.17 8.4 ;
        RECT 49.69 8.14 50.015 8.465 ;
        RECT 40.305 8.175 40.645 8.455 ;
        RECT 38.025 8.23 40.645 8.4 ;
        RECT 38.025 8.2 38.315 8.43 ;
      LAYER via1 ;
        RECT 40.4 8.24 40.55 8.39 ;
        RECT 49.78 8.225 49.93 8.375 ;
        RECT 49.78 4.875 49.93 5.025 ;
      LAYER mcon ;
        RECT 38.085 8.23 38.255 8.4 ;
        RECT 49.77 8.23 49.94 8.4 ;
        RECT 49.77 4.06 49.94 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 66.99 2.955 67.16 4.23 ;
        RECT 66.99 8.225 67.16 9.505 ;
        RECT 66.98 8.225 67.16 8.465 ;
        RECT 55.305 8.23 55.475 9.505 ;
      LAYER met2 ;
        RECT 66.91 8.14 67.235 8.465 ;
        RECT 66.91 4.79 67.235 5.115 ;
        RECT 57.61 9.24 67.16 9.41 ;
        RECT 66.99 8.14 67.16 9.41 ;
        RECT 66.98 4.79 67.15 8.465 ;
        RECT 57.555 8.145 57.835 8.485 ;
        RECT 57.61 8.145 57.78 9.41 ;
      LAYER met1 ;
        RECT 66.93 4.06 67.39 4.23 ;
        RECT 66.91 4.79 67.235 5.115 ;
        RECT 66.93 4.03 67.22 4.26 ;
        RECT 66.99 4.03 67.16 5.115 ;
        RECT 66.91 8.23 67.39 8.4 ;
        RECT 66.91 8.14 67.235 8.465 ;
        RECT 57.525 8.175 57.865 8.455 ;
        RECT 55.245 8.23 57.865 8.4 ;
        RECT 55.245 8.2 55.535 8.43 ;
      LAYER via1 ;
        RECT 57.62 8.24 57.77 8.39 ;
        RECT 67 8.225 67.15 8.375 ;
        RECT 67 4.875 67.15 5.025 ;
      LAYER mcon ;
        RECT 55.305 8.23 55.475 8.4 ;
        RECT 66.99 8.23 67.16 8.4 ;
        RECT 66.99 4.06 67.16 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 84.21 2.955 84.38 4.23 ;
        RECT 84.21 8.225 84.38 9.505 ;
        RECT 84.2 8.225 84.38 8.465 ;
        RECT 72.525 8.23 72.695 9.505 ;
      LAYER met2 ;
        RECT 84.13 8.14 84.455 8.465 ;
        RECT 84.13 4.79 84.455 5.115 ;
        RECT 74.83 9.24 84.38 9.41 ;
        RECT 84.21 8.14 84.38 9.41 ;
        RECT 84.2 4.79 84.37 8.465 ;
        RECT 74.775 8.145 75.055 8.485 ;
        RECT 74.83 8.145 75 9.41 ;
      LAYER met1 ;
        RECT 84.15 4.06 84.61 4.23 ;
        RECT 84.13 4.79 84.455 5.115 ;
        RECT 84.15 4.03 84.44 4.26 ;
        RECT 84.21 4.03 84.38 5.115 ;
        RECT 84.13 8.23 84.61 8.4 ;
        RECT 84.13 8.14 84.455 8.465 ;
        RECT 74.745 8.175 75.085 8.455 ;
        RECT 72.465 8.23 75.085 8.4 ;
        RECT 72.465 8.2 72.755 8.43 ;
      LAYER via1 ;
        RECT 74.84 8.24 74.99 8.39 ;
        RECT 84.22 8.225 84.37 8.375 ;
        RECT 84.22 4.875 84.37 5.025 ;
      LAYER mcon ;
        RECT 72.525 8.23 72.695 8.4 ;
        RECT 84.21 8.23 84.38 8.4 ;
        RECT 84.21 4.06 84.38 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.235 8.23 0.405 9.505 ;
      LAYER met1 ;
        RECT 0.175 8.23 0.635 8.4 ;
        RECT 0.175 8.2 0.465 8.43 ;
      LAYER mcon ;
        RECT 0.235 8.23 0.405 8.4 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 82.92 5.43 88.905 7.03 ;
        RECT 86.77 5.425 88.75 7.035 ;
        RECT 87.93 4.695 88.1 7.765 ;
        RECT 86.94 4.695 87.11 7.765 ;
        RECT 84.2 4.7 84.37 7.76 ;
        RECT 82.82 5.64 88.905 6.8 ;
        RECT 82.915 5.43 88.905 6.8 ;
        RECT 0.005 5.64 88.905 5.81 ;
        RECT 82.005 5.64 82.285 6.95 ;
        RECT 81.605 4.79 81.775 5.81 ;
        RECT 81.075 5.64 81.335 6.95 ;
        RECT 80.765 5.13 80.935 5.81 ;
        RECT 80.625 5.64 80.905 6.95 ;
        RECT 79.695 5.64 79.955 6.95 ;
        RECT 79.265 5.64 79.525 6.95 ;
        RECT 79.185 4.5 79.515 5.81 ;
        RECT 78.315 5.64 78.595 6.95 ;
        RECT 76.945 4.5 77.275 5.81 ;
        RECT 76.965 4.5 77.225 6.95 ;
        RECT 76.495 4.5 76.725 5.81 ;
        RECT 76.015 5.64 76.295 6.95 ;
        RECT 65.6 5.64 75.83 6.8 ;
        RECT 65.695 5.43 75.825 6.8 ;
        RECT 75.615 4.5 75.825 6.8 ;
        RECT 71.68 5.425 75.825 6.8 ;
        RECT 65.7 5.43 75.25 7.03 ;
        RECT 72.515 5.425 72.685 7.76 ;
        RECT 69.55 5.425 71.53 7.035 ;
        RECT 70.71 4.695 70.88 7.765 ;
        RECT 69.72 4.695 69.89 7.765 ;
        RECT 66.98 4.7 67.15 7.76 ;
        RECT 64.785 5.64 65.065 6.95 ;
        RECT 64.385 4.79 64.555 5.81 ;
        RECT 63.855 5.64 64.115 6.95 ;
        RECT 63.545 5.13 63.715 5.81 ;
        RECT 63.405 5.64 63.685 6.95 ;
        RECT 62.475 5.64 62.735 6.95 ;
        RECT 62.045 5.64 62.305 6.95 ;
        RECT 61.965 4.5 62.295 5.81 ;
        RECT 61.095 5.64 61.375 6.95 ;
        RECT 59.725 4.5 60.055 5.81 ;
        RECT 59.745 4.5 60.005 6.95 ;
        RECT 59.275 4.5 59.505 5.81 ;
        RECT 58.795 5.64 59.075 6.95 ;
        RECT 48.38 5.64 58.61 6.8 ;
        RECT 48.475 5.43 58.605 6.8 ;
        RECT 58.395 4.5 58.605 6.8 ;
        RECT 54.46 5.425 58.605 6.8 ;
        RECT 48.48 5.43 58.03 7.03 ;
        RECT 55.295 5.425 55.465 7.76 ;
        RECT 52.33 5.425 54.31 7.035 ;
        RECT 53.49 4.695 53.66 7.765 ;
        RECT 52.5 4.695 52.67 7.765 ;
        RECT 49.76 4.7 49.93 7.76 ;
        RECT 47.565 5.64 47.845 6.95 ;
        RECT 47.165 4.79 47.335 5.81 ;
        RECT 46.635 5.64 46.895 6.95 ;
        RECT 46.325 5.13 46.495 5.81 ;
        RECT 46.185 5.64 46.465 6.95 ;
        RECT 45.255 5.64 45.515 6.95 ;
        RECT 44.825 5.64 45.085 6.95 ;
        RECT 44.745 4.5 45.075 5.81 ;
        RECT 43.875 5.64 44.155 6.95 ;
        RECT 42.505 4.5 42.835 5.81 ;
        RECT 42.525 4.5 42.785 6.95 ;
        RECT 42.055 4.5 42.285 5.81 ;
        RECT 41.575 5.64 41.855 6.95 ;
        RECT 31.16 5.64 41.39 6.8 ;
        RECT 31.255 5.43 41.385 6.8 ;
        RECT 41.175 4.5 41.385 6.8 ;
        RECT 37.24 5.425 41.385 6.8 ;
        RECT 31.26 5.43 40.81 7.03 ;
        RECT 38.075 5.425 38.245 7.76 ;
        RECT 35.11 5.425 37.09 7.035 ;
        RECT 36.27 4.695 36.44 7.765 ;
        RECT 35.28 4.695 35.45 7.765 ;
        RECT 32.54 4.7 32.71 7.76 ;
        RECT 30.345 5.64 30.625 6.95 ;
        RECT 29.945 4.79 30.115 5.81 ;
        RECT 29.415 5.64 29.675 6.95 ;
        RECT 29.105 5.13 29.275 5.81 ;
        RECT 28.965 5.64 29.245 6.95 ;
        RECT 28.035 5.64 28.295 6.95 ;
        RECT 27.605 5.64 27.865 6.95 ;
        RECT 27.525 4.5 27.855 5.81 ;
        RECT 26.655 5.64 26.935 6.95 ;
        RECT 25.285 4.5 25.615 5.81 ;
        RECT 25.305 4.5 25.565 6.95 ;
        RECT 24.835 4.5 25.065 5.81 ;
        RECT 24.355 5.64 24.635 6.95 ;
        RECT 13.94 5.64 24.17 6.8 ;
        RECT 14.035 5.43 24.165 6.8 ;
        RECT 23.955 4.5 24.165 6.8 ;
        RECT 20.02 5.425 24.165 6.8 ;
        RECT 14.04 5.43 23.59 7.005 ;
        RECT 14.04 5.43 23.585 7.03 ;
        RECT 20.855 5.425 21.025 7.76 ;
        RECT 17.89 5.425 19.87 7.035 ;
        RECT 19.05 4.695 19.22 7.765 ;
        RECT 18.06 4.695 18.23 7.765 ;
        RECT 15.32 4.7 15.49 7.76 ;
        RECT 13.125 5.64 13.405 6.95 ;
        RECT 12.725 4.79 12.895 5.81 ;
        RECT 12.195 5.64 12.455 6.95 ;
        RECT 11.885 5.13 12.055 5.81 ;
        RECT 11.745 5.64 12.025 6.95 ;
        RECT 10.815 5.64 11.075 6.95 ;
        RECT 10.385 5.64 10.645 6.95 ;
        RECT 10.305 4.5 10.635 5.81 ;
        RECT 9.435 5.64 9.715 6.95 ;
        RECT 8.065 4.5 8.395 5.81 ;
        RECT 8.085 4.5 8.345 6.95 ;
        RECT 7.615 4.5 7.845 5.81 ;
        RECT 7.135 5.64 7.415 6.95 ;
        RECT 0.005 5.64 6.95 6.8 ;
        RECT 0.005 5.425 6.945 7 ;
        RECT 6.735 4.5 6.945 7 ;
        RECT 0.005 5.425 6.475 7.025 ;
        RECT 3.46 5.425 6.21 7.03 ;
        RECT 3.635 5.425 3.805 7.76 ;
        RECT 0.05 5.425 2.8 7.03 ;
        RECT 2.035 5.425 2.205 10.59 ;
        RECT 0.225 5.425 0.395 7.76 ;
      LAYER met1 ;
        RECT 82.92 5.43 88.905 7.03 ;
        RECT 86.77 5.425 88.75 7.035 ;
        RECT 82.83 5.485 88.905 6.955 ;
        RECT 82.915 5.43 88.905 6.955 ;
        RECT 82.82 5.485 88.905 6.8 ;
        RECT 0.005 5.485 88.905 5.965 ;
        RECT 65.6 5.485 75.83 6.8 ;
        RECT 65.695 5.43 75.825 6.8 ;
        RECT 71.68 5.425 75.825 6.8 ;
        RECT 65.7 5.43 75.25 7.03 ;
        RECT 69.55 5.425 71.53 7.035 ;
        RECT 65.61 5.485 75.25 6.955 ;
        RECT 48.38 5.485 58.61 6.8 ;
        RECT 48.475 5.43 58.605 6.8 ;
        RECT 54.46 5.425 58.605 6.8 ;
        RECT 48.48 5.43 58.03 7.03 ;
        RECT 52.33 5.425 54.31 7.035 ;
        RECT 48.39 5.485 58.03 6.955 ;
        RECT 31.16 5.485 41.39 6.8 ;
        RECT 31.255 5.43 41.385 6.8 ;
        RECT 37.24 5.425 41.385 6.8 ;
        RECT 31.26 5.43 40.81 7.03 ;
        RECT 35.11 5.425 37.09 7.035 ;
        RECT 31.17 5.485 40.81 6.955 ;
        RECT 13.94 5.485 24.17 6.8 ;
        RECT 14.035 5.43 24.165 6.8 ;
        RECT 20.02 5.425 24.165 6.8 ;
        RECT 14.04 5.43 23.59 7.005 ;
        RECT 14.04 5.43 23.585 7.03 ;
        RECT 17.89 5.425 19.87 7.035 ;
        RECT 13.95 5.485 23.59 6.955 ;
        RECT 0.005 5.485 6.95 6.8 ;
        RECT 0.005 5.425 6.945 7 ;
        RECT 0.005 5.425 6.475 7.025 ;
        RECT 3.46 5.425 6.21 7.03 ;
        RECT 0.05 5.425 2.8 7.03 ;
        RECT 1.975 8.94 2.265 9.17 ;
        RECT 1.805 8.97 2.265 9.14 ;
      LAYER mcon ;
        RECT 2.035 8.97 2.205 9.14 ;
        RECT 2.345 6.83 2.515 7 ;
        RECT 5.755 6.83 5.925 7 ;
        RECT 6.735 5.64 6.905 5.81 ;
        RECT 7.195 5.64 7.365 5.81 ;
        RECT 7.655 5.64 7.825 5.81 ;
        RECT 8.115 5.64 8.285 5.81 ;
        RECT 8.575 5.64 8.745 5.81 ;
        RECT 9.035 5.64 9.205 5.81 ;
        RECT 9.495 5.64 9.665 5.81 ;
        RECT 9.955 5.64 10.125 5.81 ;
        RECT 10.415 5.64 10.585 5.81 ;
        RECT 10.875 5.64 11.045 5.81 ;
        RECT 11.335 5.64 11.505 5.81 ;
        RECT 11.795 5.64 11.965 5.81 ;
        RECT 12.255 5.64 12.425 5.81 ;
        RECT 12.715 5.64 12.885 5.81 ;
        RECT 13.175 5.64 13.345 5.81 ;
        RECT 13.635 5.64 13.805 5.81 ;
        RECT 17.44 6.83 17.61 7 ;
        RECT 17.44 5.46 17.61 5.63 ;
        RECT 18.14 6.835 18.31 7.005 ;
        RECT 18.14 5.455 18.31 5.625 ;
        RECT 19.13 6.835 19.3 7.005 ;
        RECT 19.13 5.455 19.3 5.625 ;
        RECT 22.975 6.83 23.145 7 ;
        RECT 23.955 5.64 24.125 5.81 ;
        RECT 24.415 5.64 24.585 5.81 ;
        RECT 24.875 5.64 25.045 5.81 ;
        RECT 25.335 5.64 25.505 5.81 ;
        RECT 25.795 5.64 25.965 5.81 ;
        RECT 26.255 5.64 26.425 5.81 ;
        RECT 26.715 5.64 26.885 5.81 ;
        RECT 27.175 5.64 27.345 5.81 ;
        RECT 27.635 5.64 27.805 5.81 ;
        RECT 28.095 5.64 28.265 5.81 ;
        RECT 28.555 5.64 28.725 5.81 ;
        RECT 29.015 5.64 29.185 5.81 ;
        RECT 29.475 5.64 29.645 5.81 ;
        RECT 29.935 5.64 30.105 5.81 ;
        RECT 30.395 5.64 30.565 5.81 ;
        RECT 30.855 5.64 31.025 5.81 ;
        RECT 34.66 6.83 34.83 7 ;
        RECT 34.66 5.46 34.83 5.63 ;
        RECT 35.36 6.835 35.53 7.005 ;
        RECT 35.36 5.455 35.53 5.625 ;
        RECT 36.35 6.835 36.52 7.005 ;
        RECT 36.35 5.455 36.52 5.625 ;
        RECT 40.195 6.83 40.365 7 ;
        RECT 41.175 5.64 41.345 5.81 ;
        RECT 41.635 5.64 41.805 5.81 ;
        RECT 42.095 5.64 42.265 5.81 ;
        RECT 42.555 5.64 42.725 5.81 ;
        RECT 43.015 5.64 43.185 5.81 ;
        RECT 43.475 5.64 43.645 5.81 ;
        RECT 43.935 5.64 44.105 5.81 ;
        RECT 44.395 5.64 44.565 5.81 ;
        RECT 44.855 5.64 45.025 5.81 ;
        RECT 45.315 5.64 45.485 5.81 ;
        RECT 45.775 5.64 45.945 5.81 ;
        RECT 46.235 5.64 46.405 5.81 ;
        RECT 46.695 5.64 46.865 5.81 ;
        RECT 47.155 5.64 47.325 5.81 ;
        RECT 47.615 5.64 47.785 5.81 ;
        RECT 48.075 5.64 48.245 5.81 ;
        RECT 51.88 6.83 52.05 7 ;
        RECT 51.88 5.46 52.05 5.63 ;
        RECT 52.58 6.835 52.75 7.005 ;
        RECT 52.58 5.455 52.75 5.625 ;
        RECT 53.57 6.835 53.74 7.005 ;
        RECT 53.57 5.455 53.74 5.625 ;
        RECT 57.415 6.83 57.585 7 ;
        RECT 58.395 5.64 58.565 5.81 ;
        RECT 58.855 5.64 59.025 5.81 ;
        RECT 59.315 5.64 59.485 5.81 ;
        RECT 59.775 5.64 59.945 5.81 ;
        RECT 60.235 5.64 60.405 5.81 ;
        RECT 60.695 5.64 60.865 5.81 ;
        RECT 61.155 5.64 61.325 5.81 ;
        RECT 61.615 5.64 61.785 5.81 ;
        RECT 62.075 5.64 62.245 5.81 ;
        RECT 62.535 5.64 62.705 5.81 ;
        RECT 62.995 5.64 63.165 5.81 ;
        RECT 63.455 5.64 63.625 5.81 ;
        RECT 63.915 5.64 64.085 5.81 ;
        RECT 64.375 5.64 64.545 5.81 ;
        RECT 64.835 5.64 65.005 5.81 ;
        RECT 65.295 5.64 65.465 5.81 ;
        RECT 69.1 6.83 69.27 7 ;
        RECT 69.1 5.46 69.27 5.63 ;
        RECT 69.8 6.835 69.97 7.005 ;
        RECT 69.8 5.455 69.97 5.625 ;
        RECT 70.79 6.835 70.96 7.005 ;
        RECT 70.79 5.455 70.96 5.625 ;
        RECT 74.635 6.83 74.805 7 ;
        RECT 75.615 5.64 75.785 5.81 ;
        RECT 76.075 5.64 76.245 5.81 ;
        RECT 76.535 5.64 76.705 5.81 ;
        RECT 76.995 5.64 77.165 5.81 ;
        RECT 77.455 5.64 77.625 5.81 ;
        RECT 77.915 5.64 78.085 5.81 ;
        RECT 78.375 5.64 78.545 5.81 ;
        RECT 78.835 5.64 79.005 5.81 ;
        RECT 79.295 5.64 79.465 5.81 ;
        RECT 79.755 5.64 79.925 5.81 ;
        RECT 80.215 5.64 80.385 5.81 ;
        RECT 80.675 5.64 80.845 5.81 ;
        RECT 81.135 5.64 81.305 5.81 ;
        RECT 81.595 5.64 81.765 5.81 ;
        RECT 82.055 5.64 82.225 5.81 ;
        RECT 82.515 5.64 82.685 5.81 ;
        RECT 86.32 6.83 86.49 7 ;
        RECT 86.32 5.46 86.49 5.63 ;
        RECT 87.02 6.835 87.19 7.005 ;
        RECT 87.02 5.455 87.19 5.625 ;
        RECT 88.01 6.835 88.18 7.005 ;
        RECT 88.01 5.455 88.18 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 77.855 7.085 78.185 7.415 ;
        RECT 77.385 7.1 78.185 7.4 ;
        RECT 60.635 7.085 60.965 7.415 ;
        RECT 60.165 7.1 60.965 7.4 ;
        RECT 43.415 7.085 43.745 7.415 ;
        RECT 42.945 7.1 43.745 7.4 ;
        RECT 26.195 7.085 26.525 7.415 ;
        RECT 25.725 7.1 26.525 7.4 ;
        RECT 8.975 7.085 9.305 7.415 ;
        RECT 8.505 7.1 9.305 7.4 ;
      LAYER li1 ;
        RECT 0.05 0 88.92 1.6 ;
        RECT 87.93 0 88.1 2.225 ;
        RECT 86.94 0 87.11 2.225 ;
        RECT 84.2 0 84.37 2.23 ;
        RECT 75.47 0 83.125 3.09 ;
        RECT 82.365 0 82.695 3.48 ;
        RECT 81.525 0 81.855 3.48 ;
        RECT 79.695 0 79.985 3.925 ;
        RECT 79.245 0 79.515 3.9 ;
        RECT 78.335 0 78.575 3.9 ;
        RECT 77.885 0 78.125 3.9 ;
        RECT 76.945 0 77.215 3.9 ;
        RECT 76.495 0 76.725 3.91 ;
        RECT 75.615 0 75.825 3.91 ;
        RECT 75.465 0 83.125 2.93 ;
        RECT 70.71 0 70.88 2.225 ;
        RECT 69.72 0 69.89 2.225 ;
        RECT 66.98 0 67.15 2.23 ;
        RECT 58.25 0 65.905 3.09 ;
        RECT 65.145 0 65.475 3.48 ;
        RECT 64.305 0 64.635 3.48 ;
        RECT 62.475 0 62.765 3.925 ;
        RECT 62.025 0 62.295 3.9 ;
        RECT 61.115 0 61.355 3.9 ;
        RECT 60.665 0 60.905 3.9 ;
        RECT 59.725 0 59.995 3.9 ;
        RECT 59.275 0 59.505 3.91 ;
        RECT 58.395 0 58.605 3.91 ;
        RECT 58.245 0 65.905 2.93 ;
        RECT 53.49 0 53.66 2.225 ;
        RECT 52.5 0 52.67 2.225 ;
        RECT 49.76 0 49.93 2.23 ;
        RECT 41.03 0 48.685 3.09 ;
        RECT 47.925 0 48.255 3.48 ;
        RECT 47.085 0 47.415 3.48 ;
        RECT 45.255 0 45.545 3.925 ;
        RECT 44.805 0 45.075 3.9 ;
        RECT 43.895 0 44.135 3.9 ;
        RECT 43.445 0 43.685 3.9 ;
        RECT 42.505 0 42.775 3.9 ;
        RECT 42.055 0 42.285 3.91 ;
        RECT 41.175 0 41.385 3.91 ;
        RECT 41.025 0 48.685 2.93 ;
        RECT 36.27 0 36.44 2.225 ;
        RECT 35.28 0 35.45 2.225 ;
        RECT 32.54 0 32.71 2.23 ;
        RECT 23.81 0 31.465 3.09 ;
        RECT 30.705 0 31.035 3.48 ;
        RECT 29.865 0 30.195 3.48 ;
        RECT 28.035 0 28.325 3.925 ;
        RECT 27.585 0 27.855 3.9 ;
        RECT 26.675 0 26.915 3.9 ;
        RECT 26.225 0 26.465 3.9 ;
        RECT 25.285 0 25.555 3.9 ;
        RECT 24.835 0 25.065 3.91 ;
        RECT 23.955 0 24.165 3.91 ;
        RECT 23.805 0 31.465 2.93 ;
        RECT 19.05 0 19.22 2.225 ;
        RECT 18.06 0 18.23 2.225 ;
        RECT 15.32 0 15.49 2.23 ;
        RECT 6.59 0 14.245 3.09 ;
        RECT 13.485 0 13.815 3.48 ;
        RECT 12.645 0 12.975 3.48 ;
        RECT 10.815 0 11.105 3.925 ;
        RECT 10.365 0 10.635 3.9 ;
        RECT 9.455 0 9.695 3.9 ;
        RECT 9.005 0 9.245 3.9 ;
        RECT 8.065 0 8.335 3.9 ;
        RECT 7.615 0 7.845 3.91 ;
        RECT 6.735 0 6.945 3.91 ;
        RECT 6.585 0 14.245 2.93 ;
        RECT 0.05 10.86 88.92 12.46 ;
        RECT 87.93 10.235 88.1 12.46 ;
        RECT 86.94 10.235 87.11 12.46 ;
        RECT 84.2 10.23 84.37 12.46 ;
        RECT 75.47 8.36 82.83 12.46 ;
        RECT 81.975 7.56 82.285 12.46 ;
        RECT 80.595 7.56 80.905 12.46 ;
        RECT 78.325 7.12 78.66 7.39 ;
        RECT 78.315 7.56 78.625 12.46 ;
        RECT 77.935 7.17 78.66 7.34 ;
        RECT 77.945 7.17 78.115 12.46 ;
        RECT 76.015 7.56 76.325 12.46 ;
        RECT 72.515 10.23 72.685 12.46 ;
        RECT 70.71 10.235 70.88 12.46 ;
        RECT 69.72 10.235 69.89 12.46 ;
        RECT 66.98 10.23 67.15 12.46 ;
        RECT 58.25 8.36 65.61 12.46 ;
        RECT 64.755 7.56 65.065 12.46 ;
        RECT 63.375 7.56 63.685 12.46 ;
        RECT 61.105 7.12 61.44 7.39 ;
        RECT 61.095 7.56 61.405 12.46 ;
        RECT 60.715 7.17 61.44 7.34 ;
        RECT 60.725 7.17 60.895 12.46 ;
        RECT 58.795 7.56 59.105 12.46 ;
        RECT 55.295 10.23 55.465 12.46 ;
        RECT 53.49 10.235 53.66 12.46 ;
        RECT 52.5 10.235 52.67 12.46 ;
        RECT 49.76 10.23 49.93 12.46 ;
        RECT 41.03 8.36 48.39 12.46 ;
        RECT 47.535 7.56 47.845 12.46 ;
        RECT 46.155 7.56 46.465 12.46 ;
        RECT 43.885 7.12 44.22 7.39 ;
        RECT 43.875 7.56 44.185 12.46 ;
        RECT 43.495 7.17 44.22 7.34 ;
        RECT 43.505 7.17 43.675 12.46 ;
        RECT 41.575 7.56 41.885 12.46 ;
        RECT 38.075 10.23 38.245 12.46 ;
        RECT 36.27 10.235 36.44 12.46 ;
        RECT 35.28 10.235 35.45 12.46 ;
        RECT 32.54 10.23 32.71 12.46 ;
        RECT 23.81 8.36 31.17 12.46 ;
        RECT 30.315 7.56 30.625 12.46 ;
        RECT 28.935 7.56 29.245 12.46 ;
        RECT 26.665 7.12 27 7.39 ;
        RECT 26.655 7.56 26.965 12.46 ;
        RECT 26.275 7.17 27 7.34 ;
        RECT 26.285 7.17 26.455 12.46 ;
        RECT 24.355 7.56 24.665 12.46 ;
        RECT 20.855 10.23 21.025 12.46 ;
        RECT 19.05 10.235 19.22 12.46 ;
        RECT 18.06 10.235 18.23 12.46 ;
        RECT 15.32 10.23 15.49 12.46 ;
        RECT 6.59 8.36 13.95 12.46 ;
        RECT 13.095 7.56 13.405 12.46 ;
        RECT 11.715 7.56 12.025 12.46 ;
        RECT 9.445 7.12 9.78 7.39 ;
        RECT 9.435 7.56 9.745 12.46 ;
        RECT 9.055 7.17 9.78 7.34 ;
        RECT 9.065 7.17 9.235 12.46 ;
        RECT 7.135 7.56 7.445 12.46 ;
        RECT 3.635 10.23 3.805 12.46 ;
        RECT 0.225 10.23 0.395 12.46 ;
        RECT 76.025 7.12 76.36 7.39 ;
        RECT 75.555 7.17 76.36 7.34 ;
        RECT 73.52 8.36 73.69 10.31 ;
        RECT 73.465 10.14 73.635 10.59 ;
        RECT 73.465 7.3 73.635 8.53 ;
        RECT 58.805 7.12 59.14 7.39 ;
        RECT 58.335 7.17 59.14 7.34 ;
        RECT 56.3 8.36 56.47 10.31 ;
        RECT 56.245 10.14 56.415 10.59 ;
        RECT 56.245 7.3 56.415 8.53 ;
        RECT 41.585 7.12 41.92 7.39 ;
        RECT 41.115 7.17 41.92 7.34 ;
        RECT 39.08 8.36 39.25 10.31 ;
        RECT 39.025 10.14 39.195 10.59 ;
        RECT 39.025 7.3 39.195 8.53 ;
        RECT 24.365 7.12 24.7 7.39 ;
        RECT 23.895 7.17 24.7 7.34 ;
        RECT 21.86 8.36 22.03 10.31 ;
        RECT 21.805 10.14 21.975 10.59 ;
        RECT 21.805 7.3 21.975 8.53 ;
        RECT 7.145 7.12 7.48 7.39 ;
        RECT 6.675 7.17 7.48 7.34 ;
        RECT 4.64 8.36 4.81 10.31 ;
        RECT 4.585 10.14 4.755 10.59 ;
        RECT 4.585 7.3 4.755 8.53 ;
      LAYER met2 ;
        RECT 77.88 7.065 78.16 7.435 ;
        RECT 60.66 7.065 60.94 7.435 ;
        RECT 43.44 7.065 43.72 7.435 ;
        RECT 26.22 7.065 26.5 7.435 ;
        RECT 9 7.065 9.28 7.435 ;
      LAYER met1 ;
        RECT 0.05 0 88.92 1.6 ;
        RECT 75.47 0 83.125 3.09 ;
        RECT 75.47 0 82.83 3.245 ;
        RECT 75.465 0 83.125 2.93 ;
        RECT 58.25 0 65.905 3.09 ;
        RECT 58.25 0 65.61 3.245 ;
        RECT 58.245 0 65.905 2.93 ;
        RECT 41.03 0 48.685 3.09 ;
        RECT 41.03 0 48.39 3.245 ;
        RECT 41.025 0 48.685 2.93 ;
        RECT 23.81 0 31.465 3.09 ;
        RECT 23.81 0 31.17 3.245 ;
        RECT 23.805 0 31.465 2.93 ;
        RECT 6.59 0 14.245 3.09 ;
        RECT 6.59 0 13.95 3.245 ;
        RECT 6.585 0 14.245 2.93 ;
        RECT 0.05 10.86 88.92 12.46 ;
        RECT 75.47 8.205 82.83 12.46 ;
        RECT 73.46 8.57 73.75 8.8 ;
        RECT 73.06 8.6 73.75 8.77 ;
        RECT 73.06 8.6 73.23 12.46 ;
        RECT 58.25 8.205 65.61 12.46 ;
        RECT 56.24 8.57 56.53 8.8 ;
        RECT 55.84 8.6 56.53 8.77 ;
        RECT 55.84 8.6 56.01 12.46 ;
        RECT 41.03 8.205 48.39 12.46 ;
        RECT 39.02 8.57 39.31 8.8 ;
        RECT 38.62 8.6 39.31 8.77 ;
        RECT 38.62 8.6 38.79 12.46 ;
        RECT 23.81 8.205 31.17 12.46 ;
        RECT 21.8 8.57 22.09 8.8 ;
        RECT 21.4 8.6 22.09 8.77 ;
        RECT 21.4 8.6 21.57 12.46 ;
        RECT 6.59 8.205 13.95 12.46 ;
        RECT 4.58 8.57 4.87 8.8 ;
        RECT 4.18 8.6 4.87 8.77 ;
        RECT 4.18 8.6 4.35 12.46 ;
        RECT 77.86 7.125 78.18 7.385 ;
        RECT 75.495 7.185 78.18 7.325 ;
        RECT 75.495 7.14 75.785 7.37 ;
        RECT 60.64 7.125 60.96 7.385 ;
        RECT 58.275 7.185 60.96 7.325 ;
        RECT 58.275 7.14 58.565 7.37 ;
        RECT 43.42 7.125 43.74 7.385 ;
        RECT 41.055 7.185 43.74 7.325 ;
        RECT 41.055 7.14 41.345 7.37 ;
        RECT 26.2 7.125 26.52 7.385 ;
        RECT 23.835 7.185 26.52 7.325 ;
        RECT 23.835 7.14 24.125 7.37 ;
        RECT 8.98 7.125 9.3 7.385 ;
        RECT 6.615 7.185 9.3 7.325 ;
        RECT 6.615 7.14 6.905 7.37 ;
      LAYER via2 ;
        RECT 9.04 7.15 9.24 7.35 ;
        RECT 26.26 7.15 26.46 7.35 ;
        RECT 43.48 7.15 43.68 7.35 ;
        RECT 60.7 7.15 60.9 7.35 ;
        RECT 77.92 7.15 78.12 7.35 ;
      LAYER via1 ;
        RECT 9.065 7.18 9.215 7.33 ;
        RECT 26.285 7.18 26.435 7.33 ;
        RECT 43.505 7.18 43.655 7.33 ;
        RECT 60.725 7.18 60.875 7.33 ;
        RECT 77.945 7.18 78.095 7.33 ;
      LAYER mcon ;
        RECT 0.305 10.89 0.475 11.06 ;
        RECT 0.985 10.89 1.155 11.06 ;
        RECT 1.665 10.89 1.835 11.06 ;
        RECT 2.345 10.89 2.515 11.06 ;
        RECT 3.715 10.89 3.885 11.06 ;
        RECT 4.395 10.89 4.565 11.06 ;
        RECT 4.64 8.6 4.81 8.77 ;
        RECT 5.075 10.89 5.245 11.06 ;
        RECT 5.755 10.89 5.925 11.06 ;
        RECT 6.675 7.17 6.845 7.34 ;
        RECT 6.735 8.36 6.905 8.53 ;
        RECT 6.735 2.92 6.905 3.09 ;
        RECT 7.195 8.36 7.365 8.53 ;
        RECT 7.195 2.92 7.365 3.09 ;
        RECT 7.655 8.36 7.825 8.53 ;
        RECT 7.655 2.92 7.825 3.09 ;
        RECT 8.115 8.36 8.285 8.53 ;
        RECT 8.115 2.92 8.285 3.09 ;
        RECT 8.575 8.36 8.745 8.53 ;
        RECT 8.575 2.92 8.745 3.09 ;
        RECT 9.035 8.36 9.205 8.53 ;
        RECT 9.035 2.92 9.205 3.09 ;
        RECT 9.055 7.17 9.225 7.34 ;
        RECT 9.495 8.36 9.665 8.53 ;
        RECT 9.495 2.92 9.665 3.09 ;
        RECT 9.955 8.36 10.125 8.53 ;
        RECT 9.955 2.92 10.125 3.09 ;
        RECT 10.415 8.36 10.585 8.53 ;
        RECT 10.415 2.92 10.585 3.09 ;
        RECT 10.875 8.36 11.045 8.53 ;
        RECT 10.875 2.92 11.045 3.09 ;
        RECT 11.335 8.36 11.505 8.53 ;
        RECT 11.335 2.92 11.505 3.09 ;
        RECT 11.795 8.36 11.965 8.53 ;
        RECT 11.795 2.92 11.965 3.09 ;
        RECT 12.255 8.36 12.425 8.53 ;
        RECT 12.255 2.92 12.425 3.09 ;
        RECT 12.715 8.36 12.885 8.53 ;
        RECT 12.715 2.92 12.885 3.09 ;
        RECT 13.175 8.36 13.345 8.53 ;
        RECT 13.175 2.92 13.345 3.09 ;
        RECT 13.635 8.36 13.805 8.53 ;
        RECT 13.635 2.92 13.805 3.09 ;
        RECT 15.4 10.89 15.57 11.06 ;
        RECT 15.4 1.4 15.57 1.57 ;
        RECT 16.08 10.89 16.25 11.06 ;
        RECT 16.08 1.4 16.25 1.57 ;
        RECT 16.76 10.89 16.93 11.06 ;
        RECT 16.76 1.4 16.93 1.57 ;
        RECT 17.44 10.89 17.61 11.06 ;
        RECT 17.44 1.4 17.61 1.57 ;
        RECT 18.14 10.895 18.31 11.065 ;
        RECT 18.14 1.395 18.31 1.565 ;
        RECT 19.13 10.895 19.3 11.065 ;
        RECT 19.13 1.395 19.3 1.565 ;
        RECT 20.935 10.89 21.105 11.06 ;
        RECT 21.615 10.89 21.785 11.06 ;
        RECT 21.86 8.6 22.03 8.77 ;
        RECT 22.295 10.89 22.465 11.06 ;
        RECT 22.975 10.89 23.145 11.06 ;
        RECT 23.895 7.17 24.065 7.34 ;
        RECT 23.955 8.36 24.125 8.53 ;
        RECT 23.955 2.92 24.125 3.09 ;
        RECT 24.415 8.36 24.585 8.53 ;
        RECT 24.415 2.92 24.585 3.09 ;
        RECT 24.875 8.36 25.045 8.53 ;
        RECT 24.875 2.92 25.045 3.09 ;
        RECT 25.335 8.36 25.505 8.53 ;
        RECT 25.335 2.92 25.505 3.09 ;
        RECT 25.795 8.36 25.965 8.53 ;
        RECT 25.795 2.92 25.965 3.09 ;
        RECT 26.255 8.36 26.425 8.53 ;
        RECT 26.255 2.92 26.425 3.09 ;
        RECT 26.275 7.17 26.445 7.34 ;
        RECT 26.715 8.36 26.885 8.53 ;
        RECT 26.715 2.92 26.885 3.09 ;
        RECT 27.175 8.36 27.345 8.53 ;
        RECT 27.175 2.92 27.345 3.09 ;
        RECT 27.635 8.36 27.805 8.53 ;
        RECT 27.635 2.92 27.805 3.09 ;
        RECT 28.095 8.36 28.265 8.53 ;
        RECT 28.095 2.92 28.265 3.09 ;
        RECT 28.555 8.36 28.725 8.53 ;
        RECT 28.555 2.92 28.725 3.09 ;
        RECT 29.015 8.36 29.185 8.53 ;
        RECT 29.015 2.92 29.185 3.09 ;
        RECT 29.475 8.36 29.645 8.53 ;
        RECT 29.475 2.92 29.645 3.09 ;
        RECT 29.935 8.36 30.105 8.53 ;
        RECT 29.935 2.92 30.105 3.09 ;
        RECT 30.395 8.36 30.565 8.53 ;
        RECT 30.395 2.92 30.565 3.09 ;
        RECT 30.855 8.36 31.025 8.53 ;
        RECT 30.855 2.92 31.025 3.09 ;
        RECT 32.62 10.89 32.79 11.06 ;
        RECT 32.62 1.4 32.79 1.57 ;
        RECT 33.3 10.89 33.47 11.06 ;
        RECT 33.3 1.4 33.47 1.57 ;
        RECT 33.98 10.89 34.15 11.06 ;
        RECT 33.98 1.4 34.15 1.57 ;
        RECT 34.66 10.89 34.83 11.06 ;
        RECT 34.66 1.4 34.83 1.57 ;
        RECT 35.36 10.895 35.53 11.065 ;
        RECT 35.36 1.395 35.53 1.565 ;
        RECT 36.35 10.895 36.52 11.065 ;
        RECT 36.35 1.395 36.52 1.565 ;
        RECT 38.155 10.89 38.325 11.06 ;
        RECT 38.835 10.89 39.005 11.06 ;
        RECT 39.08 8.6 39.25 8.77 ;
        RECT 39.515 10.89 39.685 11.06 ;
        RECT 40.195 10.89 40.365 11.06 ;
        RECT 41.115 7.17 41.285 7.34 ;
        RECT 41.175 8.36 41.345 8.53 ;
        RECT 41.175 2.92 41.345 3.09 ;
        RECT 41.635 8.36 41.805 8.53 ;
        RECT 41.635 2.92 41.805 3.09 ;
        RECT 42.095 8.36 42.265 8.53 ;
        RECT 42.095 2.92 42.265 3.09 ;
        RECT 42.555 8.36 42.725 8.53 ;
        RECT 42.555 2.92 42.725 3.09 ;
        RECT 43.015 8.36 43.185 8.53 ;
        RECT 43.015 2.92 43.185 3.09 ;
        RECT 43.475 8.36 43.645 8.53 ;
        RECT 43.475 2.92 43.645 3.09 ;
        RECT 43.495 7.17 43.665 7.34 ;
        RECT 43.935 8.36 44.105 8.53 ;
        RECT 43.935 2.92 44.105 3.09 ;
        RECT 44.395 8.36 44.565 8.53 ;
        RECT 44.395 2.92 44.565 3.09 ;
        RECT 44.855 8.36 45.025 8.53 ;
        RECT 44.855 2.92 45.025 3.09 ;
        RECT 45.315 8.36 45.485 8.53 ;
        RECT 45.315 2.92 45.485 3.09 ;
        RECT 45.775 8.36 45.945 8.53 ;
        RECT 45.775 2.92 45.945 3.09 ;
        RECT 46.235 8.36 46.405 8.53 ;
        RECT 46.235 2.92 46.405 3.09 ;
        RECT 46.695 8.36 46.865 8.53 ;
        RECT 46.695 2.92 46.865 3.09 ;
        RECT 47.155 8.36 47.325 8.53 ;
        RECT 47.155 2.92 47.325 3.09 ;
        RECT 47.615 8.36 47.785 8.53 ;
        RECT 47.615 2.92 47.785 3.09 ;
        RECT 48.075 8.36 48.245 8.53 ;
        RECT 48.075 2.92 48.245 3.09 ;
        RECT 49.84 10.89 50.01 11.06 ;
        RECT 49.84 1.4 50.01 1.57 ;
        RECT 50.52 10.89 50.69 11.06 ;
        RECT 50.52 1.4 50.69 1.57 ;
        RECT 51.2 10.89 51.37 11.06 ;
        RECT 51.2 1.4 51.37 1.57 ;
        RECT 51.88 10.89 52.05 11.06 ;
        RECT 51.88 1.4 52.05 1.57 ;
        RECT 52.58 10.895 52.75 11.065 ;
        RECT 52.58 1.395 52.75 1.565 ;
        RECT 53.57 10.895 53.74 11.065 ;
        RECT 53.57 1.395 53.74 1.565 ;
        RECT 55.375 10.89 55.545 11.06 ;
        RECT 56.055 10.89 56.225 11.06 ;
        RECT 56.3 8.6 56.47 8.77 ;
        RECT 56.735 10.89 56.905 11.06 ;
        RECT 57.415 10.89 57.585 11.06 ;
        RECT 58.335 7.17 58.505 7.34 ;
        RECT 58.395 8.36 58.565 8.53 ;
        RECT 58.395 2.92 58.565 3.09 ;
        RECT 58.855 8.36 59.025 8.53 ;
        RECT 58.855 2.92 59.025 3.09 ;
        RECT 59.315 8.36 59.485 8.53 ;
        RECT 59.315 2.92 59.485 3.09 ;
        RECT 59.775 8.36 59.945 8.53 ;
        RECT 59.775 2.92 59.945 3.09 ;
        RECT 60.235 8.36 60.405 8.53 ;
        RECT 60.235 2.92 60.405 3.09 ;
        RECT 60.695 8.36 60.865 8.53 ;
        RECT 60.695 2.92 60.865 3.09 ;
        RECT 60.715 7.17 60.885 7.34 ;
        RECT 61.155 8.36 61.325 8.53 ;
        RECT 61.155 2.92 61.325 3.09 ;
        RECT 61.615 8.36 61.785 8.53 ;
        RECT 61.615 2.92 61.785 3.09 ;
        RECT 62.075 8.36 62.245 8.53 ;
        RECT 62.075 2.92 62.245 3.09 ;
        RECT 62.535 8.36 62.705 8.53 ;
        RECT 62.535 2.92 62.705 3.09 ;
        RECT 62.995 8.36 63.165 8.53 ;
        RECT 62.995 2.92 63.165 3.09 ;
        RECT 63.455 8.36 63.625 8.53 ;
        RECT 63.455 2.92 63.625 3.09 ;
        RECT 63.915 8.36 64.085 8.53 ;
        RECT 63.915 2.92 64.085 3.09 ;
        RECT 64.375 8.36 64.545 8.53 ;
        RECT 64.375 2.92 64.545 3.09 ;
        RECT 64.835 8.36 65.005 8.53 ;
        RECT 64.835 2.92 65.005 3.09 ;
        RECT 65.295 8.36 65.465 8.53 ;
        RECT 65.295 2.92 65.465 3.09 ;
        RECT 67.06 10.89 67.23 11.06 ;
        RECT 67.06 1.4 67.23 1.57 ;
        RECT 67.74 10.89 67.91 11.06 ;
        RECT 67.74 1.4 67.91 1.57 ;
        RECT 68.42 10.89 68.59 11.06 ;
        RECT 68.42 1.4 68.59 1.57 ;
        RECT 69.1 10.89 69.27 11.06 ;
        RECT 69.1 1.4 69.27 1.57 ;
        RECT 69.8 10.895 69.97 11.065 ;
        RECT 69.8 1.395 69.97 1.565 ;
        RECT 70.79 10.895 70.96 11.065 ;
        RECT 70.79 1.395 70.96 1.565 ;
        RECT 72.595 10.89 72.765 11.06 ;
        RECT 73.275 10.89 73.445 11.06 ;
        RECT 73.52 8.6 73.69 8.77 ;
        RECT 73.955 10.89 74.125 11.06 ;
        RECT 74.635 10.89 74.805 11.06 ;
        RECT 75.555 7.17 75.725 7.34 ;
        RECT 75.615 8.36 75.785 8.53 ;
        RECT 75.615 2.92 75.785 3.09 ;
        RECT 76.075 8.36 76.245 8.53 ;
        RECT 76.075 2.92 76.245 3.09 ;
        RECT 76.535 8.36 76.705 8.53 ;
        RECT 76.535 2.92 76.705 3.09 ;
        RECT 76.995 8.36 77.165 8.53 ;
        RECT 76.995 2.92 77.165 3.09 ;
        RECT 77.455 8.36 77.625 8.53 ;
        RECT 77.455 2.92 77.625 3.09 ;
        RECT 77.915 8.36 78.085 8.53 ;
        RECT 77.915 2.92 78.085 3.09 ;
        RECT 77.935 7.17 78.105 7.34 ;
        RECT 78.375 8.36 78.545 8.53 ;
        RECT 78.375 2.92 78.545 3.09 ;
        RECT 78.835 8.36 79.005 8.53 ;
        RECT 78.835 2.92 79.005 3.09 ;
        RECT 79.295 8.36 79.465 8.53 ;
        RECT 79.295 2.92 79.465 3.09 ;
        RECT 79.755 8.36 79.925 8.53 ;
        RECT 79.755 2.92 79.925 3.09 ;
        RECT 80.215 8.36 80.385 8.53 ;
        RECT 80.215 2.92 80.385 3.09 ;
        RECT 80.675 8.36 80.845 8.53 ;
        RECT 80.675 2.92 80.845 3.09 ;
        RECT 81.135 8.36 81.305 8.53 ;
        RECT 81.135 2.92 81.305 3.09 ;
        RECT 81.595 8.36 81.765 8.53 ;
        RECT 81.595 2.92 81.765 3.09 ;
        RECT 82.055 8.36 82.225 8.53 ;
        RECT 82.055 2.92 82.225 3.09 ;
        RECT 82.515 8.36 82.685 8.53 ;
        RECT 82.515 2.92 82.685 3.09 ;
        RECT 84.28 10.89 84.45 11.06 ;
        RECT 84.28 1.4 84.45 1.57 ;
        RECT 84.96 10.89 85.13 11.06 ;
        RECT 84.96 1.4 85.13 1.57 ;
        RECT 85.64 10.89 85.81 11.06 ;
        RECT 85.64 1.4 85.81 1.57 ;
        RECT 86.32 10.89 86.49 11.06 ;
        RECT 86.32 1.4 86.49 1.57 ;
        RECT 87.02 10.895 87.19 11.065 ;
        RECT 87.02 1.395 87.19 1.565 ;
        RECT 88.01 10.895 88.18 11.065 ;
        RECT 88.01 1.395 88.18 1.565 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 73.8 9.285 74.17 9.655 ;
      RECT 73.8 9.32 80.95 9.62 ;
      RECT 80.65 7.1 80.95 9.62 ;
      RECT 79.595 7.08 79.895 9.62 ;
      RECT 78.565 7.775 78.865 9.62 ;
      RECT 78.535 7.775 78.865 8.105 ;
      RECT 78.065 7.79 78.865 8.09 ;
      RECT 78.445 7.75 78.745 8.09 ;
      RECT 80.575 7.1 80.95 7.465 ;
      RECT 80.64 7.06 80.94 7.465 ;
      RECT 79.555 7.08 79.895 7.43 ;
      RECT 79.57 7.04 79.87 7.43 ;
      RECT 79.545 7.085 79.895 7.415 ;
      RECT 80.575 7.1 81.385 7.4 ;
      RECT 79.075 7.1 79.895 7.4 ;
      RECT 80.585 7.085 80.94 7.465 ;
      RECT 80.235 5.05 80.565 5.38 ;
      RECT 80.235 5.065 81.035 5.365 ;
      RECT 80.25 5.02 80.55 5.38 ;
      RECT 79.895 4.37 80.225 4.7 ;
      RECT 79.895 4.385 80.695 4.685 ;
      RECT 79.98 4.36 80.28 4.685 ;
      RECT 79.215 5.45 79.545 5.78 ;
      RECT 77.175 5.45 77.505 5.78 ;
      RECT 77.175 5.465 79.545 5.765 ;
      RECT 78.865 4.71 79.195 5.04 ;
      RECT 78.405 4.725 79.205 5.025 ;
      RECT 78.535 3.52 78.865 3.85 ;
      RECT 78.065 3.535 78.865 3.835 ;
      RECT 78.525 3.53 78.865 3.835 ;
      RECT 56.58 9.285 56.95 9.655 ;
      RECT 56.58 9.32 63.73 9.62 ;
      RECT 63.43 7.1 63.73 9.62 ;
      RECT 62.375 7.08 62.675 9.62 ;
      RECT 61.345 7.775 61.645 9.62 ;
      RECT 61.315 7.775 61.645 8.105 ;
      RECT 60.845 7.79 61.645 8.09 ;
      RECT 61.225 7.75 61.525 8.09 ;
      RECT 63.355 7.1 63.73 7.465 ;
      RECT 63.42 7.06 63.72 7.465 ;
      RECT 62.335 7.08 62.675 7.43 ;
      RECT 62.35 7.04 62.65 7.43 ;
      RECT 62.325 7.085 62.675 7.415 ;
      RECT 63.355 7.1 64.165 7.4 ;
      RECT 61.855 7.1 62.675 7.4 ;
      RECT 63.365 7.085 63.72 7.465 ;
      RECT 63.015 5.05 63.345 5.38 ;
      RECT 63.015 5.065 63.815 5.365 ;
      RECT 63.03 5.02 63.33 5.38 ;
      RECT 62.675 4.37 63.005 4.7 ;
      RECT 62.675 4.385 63.475 4.685 ;
      RECT 62.76 4.36 63.06 4.685 ;
      RECT 61.995 5.45 62.325 5.78 ;
      RECT 59.955 5.45 60.285 5.78 ;
      RECT 59.955 5.465 62.325 5.765 ;
      RECT 61.645 4.71 61.975 5.04 ;
      RECT 61.185 4.725 61.985 5.025 ;
      RECT 61.315 3.52 61.645 3.85 ;
      RECT 60.845 3.535 61.645 3.835 ;
      RECT 61.305 3.53 61.645 3.835 ;
      RECT 39.36 9.285 39.73 9.655 ;
      RECT 39.36 9.32 46.51 9.62 ;
      RECT 46.21 7.1 46.51 9.62 ;
      RECT 45.155 7.08 45.455 9.62 ;
      RECT 44.125 7.775 44.425 9.62 ;
      RECT 44.095 7.775 44.425 8.105 ;
      RECT 43.625 7.79 44.425 8.09 ;
      RECT 44.005 7.75 44.305 8.09 ;
      RECT 46.135 7.1 46.51 7.465 ;
      RECT 46.2 7.06 46.5 7.465 ;
      RECT 45.115 7.08 45.455 7.43 ;
      RECT 45.13 7.04 45.43 7.43 ;
      RECT 45.105 7.085 45.455 7.415 ;
      RECT 46.135 7.1 46.945 7.4 ;
      RECT 44.635 7.1 45.455 7.4 ;
      RECT 46.145 7.085 46.5 7.465 ;
      RECT 45.795 5.05 46.125 5.38 ;
      RECT 45.795 5.065 46.595 5.365 ;
      RECT 45.81 5.02 46.11 5.38 ;
      RECT 45.455 4.37 45.785 4.7 ;
      RECT 45.455 4.385 46.255 4.685 ;
      RECT 45.54 4.36 45.84 4.685 ;
      RECT 44.775 5.45 45.105 5.78 ;
      RECT 42.735 5.45 43.065 5.78 ;
      RECT 42.735 5.465 45.105 5.765 ;
      RECT 44.425 4.71 44.755 5.04 ;
      RECT 43.965 4.725 44.765 5.025 ;
      RECT 44.095 3.52 44.425 3.85 ;
      RECT 43.625 3.535 44.425 3.835 ;
      RECT 44.085 3.53 44.425 3.835 ;
      RECT 22.14 9.285 22.51 9.655 ;
      RECT 22.14 9.32 29.29 9.62 ;
      RECT 28.99 7.1 29.29 9.62 ;
      RECT 27.935 7.08 28.235 9.62 ;
      RECT 26.905 7.775 27.205 9.62 ;
      RECT 26.875 7.775 27.205 8.105 ;
      RECT 26.405 7.79 27.205 8.09 ;
      RECT 26.785 7.75 27.085 8.09 ;
      RECT 28.915 7.1 29.29 7.465 ;
      RECT 28.98 7.06 29.28 7.465 ;
      RECT 27.895 7.08 28.235 7.43 ;
      RECT 27.91 7.04 28.21 7.43 ;
      RECT 27.885 7.085 28.235 7.415 ;
      RECT 28.915 7.1 29.725 7.4 ;
      RECT 27.415 7.1 28.235 7.4 ;
      RECT 28.925 7.085 29.28 7.465 ;
      RECT 28.575 5.05 28.905 5.38 ;
      RECT 28.575 5.065 29.375 5.365 ;
      RECT 28.59 5.02 28.89 5.38 ;
      RECT 28.235 4.37 28.565 4.7 ;
      RECT 28.235 4.385 29.035 4.685 ;
      RECT 28.32 4.36 28.62 4.685 ;
      RECT 27.555 5.45 27.885 5.78 ;
      RECT 25.515 5.45 25.845 5.78 ;
      RECT 25.515 5.465 27.885 5.765 ;
      RECT 27.205 4.71 27.535 5.04 ;
      RECT 26.745 4.725 27.545 5.025 ;
      RECT 26.875 3.52 27.205 3.85 ;
      RECT 26.405 3.535 27.205 3.835 ;
      RECT 26.865 3.53 27.205 3.835 ;
      RECT 4.92 9.285 5.29 9.655 ;
      RECT 4.92 9.32 12.07 9.62 ;
      RECT 11.77 7.1 12.07 9.62 ;
      RECT 10.715 7.08 11.015 9.62 ;
      RECT 9.685 7.775 9.985 9.62 ;
      RECT 9.655 7.775 9.985 8.105 ;
      RECT 9.185 7.79 9.985 8.09 ;
      RECT 9.565 7.75 9.865 8.09 ;
      RECT 11.695 7.1 12.07 7.465 ;
      RECT 11.76 7.06 12.06 7.465 ;
      RECT 10.675 7.08 11.015 7.43 ;
      RECT 10.69 7.04 10.99 7.43 ;
      RECT 10.665 7.085 11.015 7.415 ;
      RECT 11.695 7.1 12.505 7.4 ;
      RECT 10.195 7.1 11.015 7.4 ;
      RECT 11.705 7.085 12.06 7.465 ;
      RECT 11.355 5.05 11.685 5.38 ;
      RECT 11.355 5.065 12.155 5.365 ;
      RECT 11.37 5.02 11.67 5.38 ;
      RECT 11.015 4.37 11.345 4.7 ;
      RECT 11.015 4.385 11.815 4.685 ;
      RECT 11.1 4.36 11.4 4.685 ;
      RECT 10.335 5.45 10.665 5.78 ;
      RECT 8.295 5.45 8.625 5.78 ;
      RECT 8.295 5.465 10.665 5.765 ;
      RECT 9.985 4.71 10.315 5.04 ;
      RECT 9.525 4.725 10.325 5.025 ;
      RECT 9.655 3.52 9.985 3.85 ;
      RECT 9.185 3.535 9.985 3.835 ;
      RECT 9.645 3.53 9.985 3.835 ;
    LAYER via2 ;
      RECT 80.65 7.15 80.85 7.35 ;
      RECT 80.3 5.115 80.5 5.315 ;
      RECT 79.96 4.435 80.16 4.635 ;
      RECT 79.61 7.15 79.81 7.35 ;
      RECT 79.28 5.515 79.48 5.715 ;
      RECT 78.93 4.775 79.13 4.975 ;
      RECT 78.6 3.585 78.8 3.785 ;
      RECT 78.6 7.84 78.8 8.04 ;
      RECT 77.24 5.515 77.44 5.715 ;
      RECT 73.885 9.37 74.085 9.57 ;
      RECT 63.43 7.15 63.63 7.35 ;
      RECT 63.08 5.115 63.28 5.315 ;
      RECT 62.74 4.435 62.94 4.635 ;
      RECT 62.39 7.15 62.59 7.35 ;
      RECT 62.06 5.515 62.26 5.715 ;
      RECT 61.71 4.775 61.91 4.975 ;
      RECT 61.38 3.585 61.58 3.785 ;
      RECT 61.38 7.84 61.58 8.04 ;
      RECT 60.02 5.515 60.22 5.715 ;
      RECT 56.665 9.37 56.865 9.57 ;
      RECT 46.21 7.15 46.41 7.35 ;
      RECT 45.86 5.115 46.06 5.315 ;
      RECT 45.52 4.435 45.72 4.635 ;
      RECT 45.17 7.15 45.37 7.35 ;
      RECT 44.84 5.515 45.04 5.715 ;
      RECT 44.49 4.775 44.69 4.975 ;
      RECT 44.16 3.585 44.36 3.785 ;
      RECT 44.16 7.84 44.36 8.04 ;
      RECT 42.8 5.515 43 5.715 ;
      RECT 39.445 9.37 39.645 9.57 ;
      RECT 28.99 7.15 29.19 7.35 ;
      RECT 28.64 5.115 28.84 5.315 ;
      RECT 28.3 4.435 28.5 4.635 ;
      RECT 27.95 7.15 28.15 7.35 ;
      RECT 27.62 5.515 27.82 5.715 ;
      RECT 27.27 4.775 27.47 4.975 ;
      RECT 26.94 3.585 27.14 3.785 ;
      RECT 26.94 7.84 27.14 8.04 ;
      RECT 25.58 5.515 25.78 5.715 ;
      RECT 22.225 9.37 22.425 9.57 ;
      RECT 11.77 7.15 11.97 7.35 ;
      RECT 11.42 5.115 11.62 5.315 ;
      RECT 11.08 4.435 11.28 4.635 ;
      RECT 10.73 7.15 10.93 7.35 ;
      RECT 10.4 5.515 10.6 5.715 ;
      RECT 10.05 4.775 10.25 4.975 ;
      RECT 9.72 3.585 9.92 3.785 ;
      RECT 9.72 7.84 9.92 8.04 ;
      RECT 8.36 5.515 8.56 5.715 ;
      RECT 5.005 9.37 5.205 9.57 ;
    LAYER met2 ;
      RECT 1.215 10.055 88.535 10.225 ;
      RECT 88.365 9.585 88.535 10.225 ;
      RECT 1.215 8.54 1.385 10.225 ;
      RECT 88.33 9.585 88.655 9.91 ;
      RECT 1.17 8.54 1.45 8.88 ;
      RECT 85.175 8.565 85.495 8.89 ;
      RECT 85.205 7.98 85.375 8.89 ;
      RECT 85.205 7.98 85.38 8.33 ;
      RECT 85.205 7.98 86.18 8.155 ;
      RECT 86.005 3.26 86.18 8.155 ;
      RECT 78.56 3.5 78.84 3.87 ;
      RECT 78.56 3.64 83.21 3.815 ;
      RECT 83.035 3.32 83.21 3.815 ;
      RECT 83.505 3.29 83.83 3.615 ;
      RECT 85.95 3.26 86.3 3.61 ;
      RECT 83.035 3.32 86.3 3.49 ;
      RECT 74.325 9.55 85.02 9.72 ;
      RECT 84.86 3.69 85.02 9.72 ;
      RECT 74.325 8.83 74.495 9.72 ;
      RECT 85.975 8.94 86.3 9.265 ;
      RECT 71.145 8.94 71.47 9.265 ;
      RECT 84.86 9.03 86.3 9.2 ;
      RECT 74.275 8.83 74.555 9.17 ;
      RECT 71.145 8.97 74.555 9.14 ;
      RECT 85.175 3.66 85.495 3.98 ;
      RECT 84.86 3.69 85.495 3.86 ;
      RECT 81.63 7.775 81.89 8.095 ;
      RECT 81.69 4.035 81.83 8.095 ;
      RECT 81.63 4.035 81.89 4.355 ;
      RECT 80.95 6.075 81.21 6.395 ;
      RECT 81.01 5.055 81.15 6.395 ;
      RECT 80.95 5.055 81.21 5.375 ;
      RECT 79.93 7.775 80.19 8.095 ;
      RECT 79.99 6.505 80.13 8.095 ;
      RECT 79.31 6.505 80.13 6.645 ;
      RECT 79.31 4.035 79.45 6.645 ;
      RECT 79.24 5.43 79.52 5.8 ;
      RECT 79.25 4.035 79.51 4.355 ;
      RECT 77.2 5.43 77.48 5.8 ;
      RECT 77.27 3.695 77.41 5.8 ;
      RECT 77.21 3.695 77.47 4.015 ;
      RECT 76.53 6.075 76.79 6.395 ;
      RECT 76.59 4.035 76.73 6.395 ;
      RECT 76.53 4.035 76.79 4.355 ;
      RECT 67.955 8.565 68.275 8.89 ;
      RECT 67.985 7.98 68.155 8.89 ;
      RECT 67.985 7.98 68.16 8.33 ;
      RECT 67.985 7.98 68.96 8.155 ;
      RECT 68.785 3.26 68.96 8.155 ;
      RECT 61.34 3.5 61.62 3.87 ;
      RECT 61.34 3.64 65.99 3.815 ;
      RECT 65.815 3.32 65.99 3.815 ;
      RECT 66.285 3.29 66.61 3.615 ;
      RECT 68.73 3.26 69.08 3.61 ;
      RECT 65.815 3.32 69.08 3.49 ;
      RECT 57.105 9.55 67.8 9.72 ;
      RECT 67.64 3.69 67.8 9.72 ;
      RECT 57.105 8.83 57.275 9.72 ;
      RECT 68.755 8.94 69.08 9.265 ;
      RECT 53.925 8.94 54.25 9.265 ;
      RECT 67.64 9.03 69.08 9.2 ;
      RECT 57.055 8.83 57.335 9.17 ;
      RECT 53.925 8.97 57.335 9.14 ;
      RECT 67.955 3.66 68.275 3.98 ;
      RECT 67.64 3.69 68.275 3.86 ;
      RECT 64.41 7.775 64.67 8.095 ;
      RECT 64.47 4.035 64.61 8.095 ;
      RECT 64.41 4.035 64.67 4.355 ;
      RECT 63.73 6.075 63.99 6.395 ;
      RECT 63.79 5.055 63.93 6.395 ;
      RECT 63.73 5.055 63.99 5.375 ;
      RECT 62.71 7.775 62.97 8.095 ;
      RECT 62.77 6.505 62.91 8.095 ;
      RECT 62.09 6.505 62.91 6.645 ;
      RECT 62.09 4.035 62.23 6.645 ;
      RECT 62.02 5.43 62.3 5.8 ;
      RECT 62.03 4.035 62.29 4.355 ;
      RECT 59.98 5.43 60.26 5.8 ;
      RECT 60.05 3.695 60.19 5.8 ;
      RECT 59.99 3.695 60.25 4.015 ;
      RECT 59.31 6.075 59.57 6.395 ;
      RECT 59.37 4.035 59.51 6.395 ;
      RECT 59.31 4.035 59.57 4.355 ;
      RECT 50.735 8.565 51.055 8.89 ;
      RECT 50.765 7.98 50.935 8.89 ;
      RECT 50.765 7.98 50.94 8.33 ;
      RECT 50.765 7.98 51.74 8.155 ;
      RECT 51.565 3.26 51.74 8.155 ;
      RECT 44.12 3.5 44.4 3.87 ;
      RECT 44.12 3.64 48.77 3.815 ;
      RECT 48.595 3.32 48.77 3.815 ;
      RECT 49.065 3.29 49.39 3.615 ;
      RECT 51.51 3.26 51.86 3.61 ;
      RECT 48.595 3.32 51.86 3.49 ;
      RECT 39.885 9.55 50.58 9.72 ;
      RECT 50.42 3.69 50.58 9.72 ;
      RECT 39.885 8.83 40.055 9.72 ;
      RECT 51.535 8.94 51.86 9.265 ;
      RECT 36.705 8.94 37.03 9.265 ;
      RECT 50.42 9.03 51.86 9.2 ;
      RECT 39.835 8.83 40.115 9.17 ;
      RECT 36.705 8.97 40.125 9.14 ;
      RECT 50.735 3.66 51.055 3.98 ;
      RECT 50.42 3.69 51.055 3.86 ;
      RECT 47.19 7.775 47.45 8.095 ;
      RECT 47.25 4.035 47.39 8.095 ;
      RECT 47.19 4.035 47.45 4.355 ;
      RECT 46.51 6.075 46.77 6.395 ;
      RECT 46.57 5.055 46.71 6.395 ;
      RECT 46.51 5.055 46.77 5.375 ;
      RECT 45.49 7.775 45.75 8.095 ;
      RECT 45.55 6.505 45.69 8.095 ;
      RECT 44.87 6.505 45.69 6.645 ;
      RECT 44.87 4.035 45.01 6.645 ;
      RECT 44.8 5.43 45.08 5.8 ;
      RECT 44.81 4.035 45.07 4.355 ;
      RECT 42.76 5.43 43.04 5.8 ;
      RECT 42.83 3.695 42.97 5.8 ;
      RECT 42.77 3.695 43.03 4.015 ;
      RECT 42.09 6.075 42.35 6.395 ;
      RECT 42.15 4.035 42.29 6.395 ;
      RECT 42.09 4.035 42.35 4.355 ;
      RECT 33.515 8.565 33.835 8.89 ;
      RECT 33.545 7.98 33.715 8.89 ;
      RECT 33.545 7.98 33.72 8.33 ;
      RECT 33.545 7.98 34.52 8.155 ;
      RECT 34.345 3.26 34.52 8.155 ;
      RECT 26.9 3.5 27.18 3.87 ;
      RECT 26.9 3.64 31.55 3.815 ;
      RECT 31.375 3.32 31.55 3.815 ;
      RECT 31.845 3.29 32.17 3.615 ;
      RECT 34.29 3.26 34.64 3.61 ;
      RECT 31.375 3.32 34.64 3.49 ;
      RECT 22.665 9.55 33.36 9.72 ;
      RECT 33.2 3.69 33.36 9.72 ;
      RECT 22.665 8.83 22.835 9.72 ;
      RECT 34.315 8.94 34.64 9.265 ;
      RECT 19.485 8.94 19.81 9.265 ;
      RECT 33.2 9.03 34.64 9.2 ;
      RECT 22.615 8.83 22.895 9.17 ;
      RECT 19.485 8.97 22.895 9.14 ;
      RECT 33.515 3.66 33.835 3.98 ;
      RECT 33.2 3.69 33.835 3.86 ;
      RECT 29.97 7.775 30.23 8.095 ;
      RECT 30.03 4.035 30.17 8.095 ;
      RECT 29.97 4.035 30.23 4.355 ;
      RECT 29.29 6.075 29.55 6.395 ;
      RECT 29.35 5.055 29.49 6.395 ;
      RECT 29.29 5.055 29.55 5.375 ;
      RECT 28.27 7.775 28.53 8.095 ;
      RECT 28.33 6.505 28.47 8.095 ;
      RECT 27.65 6.505 28.47 6.645 ;
      RECT 27.65 4.035 27.79 6.645 ;
      RECT 27.58 5.43 27.86 5.8 ;
      RECT 27.59 4.035 27.85 4.355 ;
      RECT 25.54 5.43 25.82 5.8 ;
      RECT 25.61 3.695 25.75 5.8 ;
      RECT 25.55 3.695 25.81 4.015 ;
      RECT 24.87 6.075 25.13 6.395 ;
      RECT 24.93 4.035 25.07 6.395 ;
      RECT 24.87 4.035 25.13 4.355 ;
      RECT 16.295 8.565 16.615 8.89 ;
      RECT 16.325 7.98 16.495 8.89 ;
      RECT 16.325 7.98 16.5 8.33 ;
      RECT 16.325 7.98 17.3 8.155 ;
      RECT 17.125 3.26 17.3 8.155 ;
      RECT 9.68 3.5 9.96 3.87 ;
      RECT 9.68 3.64 14.33 3.815 ;
      RECT 14.155 3.32 14.33 3.815 ;
      RECT 14.625 3.29 14.95 3.615 ;
      RECT 17.07 3.26 17.42 3.61 ;
      RECT 14.155 3.32 17.42 3.49 ;
      RECT 5.445 9.55 16.14 9.72 ;
      RECT 15.98 3.69 16.14 9.72 ;
      RECT 1.545 9.28 1.825 9.62 ;
      RECT 5.445 8.83 5.615 9.72 ;
      RECT 1.545 9.345 2.75 9.515 ;
      RECT 2.58 8.97 2.75 9.515 ;
      RECT 17.095 8.94 17.42 9.265 ;
      RECT 15.98 9.03 17.42 9.2 ;
      RECT 5.395 8.83 5.675 9.17 ;
      RECT 2.58 8.97 5.675 9.14 ;
      RECT 16.295 3.66 16.615 3.98 ;
      RECT 15.98 3.69 16.615 3.86 ;
      RECT 12.75 7.775 13.01 8.095 ;
      RECT 12.81 4.035 12.95 8.095 ;
      RECT 12.75 4.035 13.01 4.355 ;
      RECT 12.07 6.075 12.33 6.395 ;
      RECT 12.13 5.055 12.27 6.395 ;
      RECT 12.07 5.055 12.33 5.375 ;
      RECT 11.05 7.775 11.31 8.095 ;
      RECT 11.11 6.505 11.25 8.095 ;
      RECT 10.43 6.505 11.25 6.645 ;
      RECT 10.43 4.035 10.57 6.645 ;
      RECT 10.36 5.43 10.64 5.8 ;
      RECT 10.37 4.035 10.63 4.355 ;
      RECT 8.32 5.43 8.6 5.8 ;
      RECT 8.39 3.695 8.53 5.8 ;
      RECT 8.33 3.695 8.59 4.015 ;
      RECT 7.65 6.075 7.91 6.395 ;
      RECT 7.71 4.035 7.85 6.395 ;
      RECT 7.65 4.035 7.91 4.355 ;
      RECT 80.61 7.065 80.89 7.435 ;
      RECT 80.26 5.03 80.54 5.4 ;
      RECT 79.92 4.35 80.2 4.72 ;
      RECT 79.57 7.065 79.85 7.435 ;
      RECT 78.89 4.69 79.17 5.06 ;
      RECT 78.56 7.755 78.84 8.125 ;
      RECT 73.8 9.285 74.17 9.655 ;
      RECT 63.39 7.065 63.67 7.435 ;
      RECT 63.04 5.03 63.32 5.4 ;
      RECT 62.7 4.35 62.98 4.72 ;
      RECT 62.35 7.065 62.63 7.435 ;
      RECT 61.67 4.69 61.95 5.06 ;
      RECT 61.34 7.755 61.62 8.125 ;
      RECT 56.58 9.285 56.95 9.655 ;
      RECT 46.17 7.065 46.45 7.435 ;
      RECT 45.82 5.03 46.1 5.4 ;
      RECT 45.48 4.35 45.76 4.72 ;
      RECT 45.13 7.065 45.41 7.435 ;
      RECT 44.45 4.69 44.73 5.06 ;
      RECT 44.12 7.755 44.4 8.125 ;
      RECT 39.36 9.285 39.73 9.655 ;
      RECT 28.95 7.065 29.23 7.435 ;
      RECT 28.6 5.03 28.88 5.4 ;
      RECT 28.26 4.35 28.54 4.72 ;
      RECT 27.91 7.065 28.19 7.435 ;
      RECT 27.23 4.69 27.51 5.06 ;
      RECT 26.9 7.755 27.18 8.125 ;
      RECT 22.14 9.285 22.51 9.655 ;
      RECT 11.73 7.065 12.01 7.435 ;
      RECT 11.38 5.03 11.66 5.4 ;
      RECT 11.04 4.35 11.32 4.72 ;
      RECT 10.69 7.065 10.97 7.435 ;
      RECT 10.01 4.69 10.29 5.06 ;
      RECT 9.68 7.755 9.96 8.125 ;
      RECT 4.92 9.285 5.29 9.655 ;
    LAYER via1 ;
      RECT 88.42 9.67 88.57 9.82 ;
      RECT 86.065 9.025 86.215 9.175 ;
      RECT 86.05 3.36 86.2 3.51 ;
      RECT 85.26 3.745 85.41 3.895 ;
      RECT 85.26 8.655 85.41 8.805 ;
      RECT 83.595 3.375 83.745 3.525 ;
      RECT 81.685 4.12 81.835 4.27 ;
      RECT 81.685 7.86 81.835 8.01 ;
      RECT 81.005 5.14 81.155 5.29 ;
      RECT 81.005 6.16 81.155 6.31 ;
      RECT 80.665 7.18 80.815 7.33 ;
      RECT 80.325 5.14 80.475 5.29 ;
      RECT 79.985 4.46 80.135 4.61 ;
      RECT 79.985 7.86 80.135 8.01 ;
      RECT 79.635 7.18 79.785 7.33 ;
      RECT 79.305 4.12 79.455 4.27 ;
      RECT 78.965 4.8 79.115 4.95 ;
      RECT 78.625 3.61 78.775 3.76 ;
      RECT 78.625 7.86 78.775 8.01 ;
      RECT 77.265 3.78 77.415 3.93 ;
      RECT 76.585 4.12 76.735 4.27 ;
      RECT 76.585 6.16 76.735 6.31 ;
      RECT 74.34 8.925 74.49 9.075 ;
      RECT 73.91 9.395 74.06 9.545 ;
      RECT 71.235 9.025 71.385 9.175 ;
      RECT 68.845 9.025 68.995 9.175 ;
      RECT 68.83 3.36 68.98 3.51 ;
      RECT 68.04 3.745 68.19 3.895 ;
      RECT 68.04 8.655 68.19 8.805 ;
      RECT 66.375 3.375 66.525 3.525 ;
      RECT 64.465 4.12 64.615 4.27 ;
      RECT 64.465 7.86 64.615 8.01 ;
      RECT 63.785 5.14 63.935 5.29 ;
      RECT 63.785 6.16 63.935 6.31 ;
      RECT 63.445 7.18 63.595 7.33 ;
      RECT 63.105 5.14 63.255 5.29 ;
      RECT 62.765 4.46 62.915 4.61 ;
      RECT 62.765 7.86 62.915 8.01 ;
      RECT 62.415 7.18 62.565 7.33 ;
      RECT 62.085 4.12 62.235 4.27 ;
      RECT 61.745 4.8 61.895 4.95 ;
      RECT 61.405 3.61 61.555 3.76 ;
      RECT 61.405 7.86 61.555 8.01 ;
      RECT 60.045 3.78 60.195 3.93 ;
      RECT 59.365 4.12 59.515 4.27 ;
      RECT 59.365 6.16 59.515 6.31 ;
      RECT 57.12 8.925 57.27 9.075 ;
      RECT 56.69 9.395 56.84 9.545 ;
      RECT 54.015 9.025 54.165 9.175 ;
      RECT 51.625 9.025 51.775 9.175 ;
      RECT 51.61 3.36 51.76 3.51 ;
      RECT 50.82 3.745 50.97 3.895 ;
      RECT 50.82 8.655 50.97 8.805 ;
      RECT 49.155 3.375 49.305 3.525 ;
      RECT 47.245 4.12 47.395 4.27 ;
      RECT 47.245 7.86 47.395 8.01 ;
      RECT 46.565 5.14 46.715 5.29 ;
      RECT 46.565 6.16 46.715 6.31 ;
      RECT 46.225 7.18 46.375 7.33 ;
      RECT 45.885 5.14 46.035 5.29 ;
      RECT 45.545 4.46 45.695 4.61 ;
      RECT 45.545 7.86 45.695 8.01 ;
      RECT 45.195 7.18 45.345 7.33 ;
      RECT 44.865 4.12 45.015 4.27 ;
      RECT 44.525 4.8 44.675 4.95 ;
      RECT 44.185 3.61 44.335 3.76 ;
      RECT 44.185 7.86 44.335 8.01 ;
      RECT 42.825 3.78 42.975 3.93 ;
      RECT 42.145 4.12 42.295 4.27 ;
      RECT 42.145 6.16 42.295 6.31 ;
      RECT 39.9 8.925 40.05 9.075 ;
      RECT 39.47 9.395 39.62 9.545 ;
      RECT 36.795 9.025 36.945 9.175 ;
      RECT 34.405 9.025 34.555 9.175 ;
      RECT 34.39 3.36 34.54 3.51 ;
      RECT 33.6 3.745 33.75 3.895 ;
      RECT 33.6 8.655 33.75 8.805 ;
      RECT 31.935 3.375 32.085 3.525 ;
      RECT 30.025 4.12 30.175 4.27 ;
      RECT 30.025 7.86 30.175 8.01 ;
      RECT 29.345 5.14 29.495 5.29 ;
      RECT 29.345 6.16 29.495 6.31 ;
      RECT 29.005 7.18 29.155 7.33 ;
      RECT 28.665 5.14 28.815 5.29 ;
      RECT 28.325 4.46 28.475 4.61 ;
      RECT 28.325 7.86 28.475 8.01 ;
      RECT 27.975 7.18 28.125 7.33 ;
      RECT 27.645 4.12 27.795 4.27 ;
      RECT 27.305 4.8 27.455 4.95 ;
      RECT 26.965 3.61 27.115 3.76 ;
      RECT 26.965 7.86 27.115 8.01 ;
      RECT 25.605 3.78 25.755 3.93 ;
      RECT 24.925 4.12 25.075 4.27 ;
      RECT 24.925 6.16 25.075 6.31 ;
      RECT 22.68 8.925 22.83 9.075 ;
      RECT 22.25 9.395 22.4 9.545 ;
      RECT 19.575 9.025 19.725 9.175 ;
      RECT 17.185 9.025 17.335 9.175 ;
      RECT 17.17 3.36 17.32 3.51 ;
      RECT 16.38 3.745 16.53 3.895 ;
      RECT 16.38 8.655 16.53 8.805 ;
      RECT 14.715 3.375 14.865 3.525 ;
      RECT 12.805 4.12 12.955 4.27 ;
      RECT 12.805 7.86 12.955 8.01 ;
      RECT 12.125 5.14 12.275 5.29 ;
      RECT 12.125 6.16 12.275 6.31 ;
      RECT 11.785 7.18 11.935 7.33 ;
      RECT 11.445 5.14 11.595 5.29 ;
      RECT 11.105 4.46 11.255 4.61 ;
      RECT 11.105 7.86 11.255 8.01 ;
      RECT 10.755 7.18 10.905 7.33 ;
      RECT 10.425 4.12 10.575 4.27 ;
      RECT 10.085 4.8 10.235 4.95 ;
      RECT 9.745 3.61 9.895 3.76 ;
      RECT 9.745 7.86 9.895 8.01 ;
      RECT 8.385 3.78 8.535 3.93 ;
      RECT 7.705 4.12 7.855 4.27 ;
      RECT 7.705 6.16 7.855 6.31 ;
      RECT 5.46 8.925 5.61 9.075 ;
      RECT 5.03 9.395 5.18 9.545 ;
      RECT 1.61 9.375 1.76 9.525 ;
      RECT 1.235 8.635 1.385 8.785 ;
    LAYER met1 ;
      RECT 88.3 10.055 88.59 10.285 ;
      RECT 88.36 8.575 88.53 10.285 ;
      RECT 88.33 9.585 88.655 9.91 ;
      RECT 88.3 8.575 88.59 8.805 ;
      RECT 87.895 3.69 88 4.26 ;
      RECT 87.895 4.025 88.22 4.255 ;
      RECT 87.895 4.055 88.39 4.225 ;
      RECT 87.895 3.69 88.085 4.255 ;
      RECT 87.31 3.655 87.6 3.885 ;
      RECT 87.31 3.69 88.085 3.86 ;
      RECT 87.37 2.175 87.54 3.885 ;
      RECT 87.31 2.175 87.6 2.405 ;
      RECT 87.31 10.055 87.6 10.285 ;
      RECT 87.37 8.575 87.54 10.285 ;
      RECT 87.31 8.575 87.6 8.805 ;
      RECT 87.31 8.61 88.165 8.77 ;
      RECT 87.995 8.205 88.165 8.77 ;
      RECT 87.31 8.605 87.705 8.77 ;
      RECT 87.93 8.205 88.22 8.435 ;
      RECT 87.93 8.235 88.39 8.405 ;
      RECT 86.94 4.025 87.23 4.255 ;
      RECT 86.94 4.055 87.4 4.225 ;
      RECT 87.005 2.95 87.17 4.255 ;
      RECT 85.52 2.92 85.81 3.15 ;
      RECT 85.52 2.95 87.17 3.12 ;
      RECT 85.58 2.18 85.75 3.15 ;
      RECT 85.52 2.18 85.81 2.41 ;
      RECT 85.52 10.05 85.81 10.28 ;
      RECT 85.58 9.31 85.75 10.28 ;
      RECT 85.58 9.405 87.17 9.575 ;
      RECT 87 8.205 87.17 9.575 ;
      RECT 85.52 9.31 85.81 9.54 ;
      RECT 86.94 8.205 87.23 8.435 ;
      RECT 86.94 8.235 87.4 8.405 ;
      RECT 85.95 3.26 86.3 3.61 ;
      RECT 85.78 3.32 86.3 3.49 ;
      RECT 85.975 8.94 86.3 9.265 ;
      RECT 85.95 8.94 86.3 9.17 ;
      RECT 85.78 8.97 86.3 9.14 ;
      RECT 85.175 3.66 85.495 3.98 ;
      RECT 85.145 3.66 85.495 3.89 ;
      RECT 84.86 3.69 85.495 3.86 ;
      RECT 85.175 8.565 85.495 8.89 ;
      RECT 85.145 8.57 85.495 8.8 ;
      RECT 84.975 8.6 85.495 8.77 ;
      RECT 80.92 5.085 81.24 5.345 ;
      RECT 81.955 5.1 82.245 5.33 ;
      RECT 80.92 5.145 82.245 5.285 ;
      RECT 80.58 7.125 80.9 7.385 ;
      RECT 81.955 7.14 82.245 7.37 ;
      RECT 82.03 6.845 82.17 7.37 ;
      RECT 80.67 6.845 80.81 7.385 ;
      RECT 80.67 6.845 82.17 6.985 ;
      RECT 81.6 4.065 81.92 4.325 ;
      RECT 81.325 4.125 81.92 4.265 ;
      RECT 78.54 7.805 78.86 8.065 ;
      RECT 77.535 7.82 77.825 8.05 ;
      RECT 77.535 7.865 79.45 8.005 ;
      RECT 79.31 7.525 79.45 8.005 ;
      RECT 79.31 7.525 81.32 7.665 ;
      RECT 81.18 7.14 81.32 7.665 ;
      RECT 81.105 7.14 81.395 7.37 ;
      RECT 80.92 6.105 81.24 6.365 ;
      RECT 78.775 6.12 79.065 6.35 ;
      RECT 78.775 6.165 81.24 6.305 ;
      RECT 80.24 5.085 80.56 5.345 ;
      RECT 77.875 5.1 78.165 5.33 ;
      RECT 77.875 5.145 80.56 5.285 ;
      RECT 79.9 7.805 80.22 8.065 ;
      RECT 79.9 7.865 80.495 8.005 ;
      RECT 79.9 4.405 80.22 4.665 ;
      RECT 79.625 4.465 80.22 4.605 ;
      RECT 79.22 4.065 79.54 4.325 ;
      RECT 78.945 4.125 79.54 4.265 ;
      RECT 78.88 4.745 79.2 5.005 ;
      RECT 76.005 4.76 76.295 4.99 ;
      RECT 76.005 4.805 79.2 4.945 ;
      RECT 78.46 4.085 78.6 4.945 ;
      RECT 78.385 4.085 78.675 4.315 ;
      RECT 78.54 3.555 78.86 3.815 ;
      RECT 78.54 3.57 79.045 3.8 ;
      RECT 78.45 3.615 79.045 3.755 ;
      RECT 77.875 4.085 78.165 4.315 ;
      RECT 77.27 4.13 78.165 4.27 ;
      RECT 77.27 3.725 77.41 4.27 ;
      RECT 77.18 3.725 77.5 3.985 ;
      RECT 76.5 4.065 76.82 4.325 ;
      RECT 76.225 4.125 76.82 4.265 ;
      RECT 76.5 6.105 76.82 6.365 ;
      RECT 76.225 6.165 76.82 6.305 ;
      RECT 74.265 8.86 74.555 9.17 ;
      RECT 74.095 8.97 74.585 9.14 ;
      RECT 74.245 8.86 74.585 9.14 ;
      RECT 73.835 10.05 74.125 10.28 ;
      RECT 73.895 9.28 74.065 10.28 ;
      RECT 73.8 9.28 74.17 9.655 ;
      RECT 71.08 10.055 71.37 10.285 ;
      RECT 71.14 8.575 71.31 10.285 ;
      RECT 71.14 8.94 71.47 9.265 ;
      RECT 71.08 8.575 71.37 8.805 ;
      RECT 70.675 3.69 70.78 4.26 ;
      RECT 70.675 4.025 71 4.255 ;
      RECT 70.675 4.055 71.17 4.225 ;
      RECT 70.675 3.69 70.865 4.255 ;
      RECT 70.09 3.655 70.38 3.885 ;
      RECT 70.09 3.69 70.865 3.86 ;
      RECT 70.15 2.175 70.32 3.885 ;
      RECT 70.09 2.175 70.38 2.405 ;
      RECT 70.09 10.055 70.38 10.285 ;
      RECT 70.15 8.575 70.32 10.285 ;
      RECT 70.09 8.575 70.38 8.805 ;
      RECT 70.09 8.61 70.945 8.77 ;
      RECT 70.775 8.205 70.945 8.77 ;
      RECT 70.09 8.605 70.485 8.77 ;
      RECT 70.71 8.205 71 8.435 ;
      RECT 70.71 8.235 71.17 8.405 ;
      RECT 69.72 4.025 70.01 4.255 ;
      RECT 69.72 4.055 70.18 4.225 ;
      RECT 69.785 2.95 69.95 4.255 ;
      RECT 68.3 2.92 68.59 3.15 ;
      RECT 68.3 2.95 69.95 3.12 ;
      RECT 68.36 2.18 68.53 3.15 ;
      RECT 68.3 2.18 68.59 2.41 ;
      RECT 68.3 10.05 68.59 10.28 ;
      RECT 68.36 9.31 68.53 10.28 ;
      RECT 68.36 9.405 69.95 9.575 ;
      RECT 69.78 8.205 69.95 9.575 ;
      RECT 68.3 9.31 68.59 9.54 ;
      RECT 69.72 8.205 70.01 8.435 ;
      RECT 69.72 8.235 70.18 8.405 ;
      RECT 68.73 3.26 69.08 3.61 ;
      RECT 68.56 3.32 69.08 3.49 ;
      RECT 68.755 8.94 69.08 9.265 ;
      RECT 68.73 8.94 69.08 9.17 ;
      RECT 68.56 8.97 69.08 9.14 ;
      RECT 67.955 3.66 68.275 3.98 ;
      RECT 67.925 3.66 68.275 3.89 ;
      RECT 67.64 3.69 68.275 3.86 ;
      RECT 67.955 8.565 68.275 8.89 ;
      RECT 67.925 8.57 68.275 8.8 ;
      RECT 67.755 8.6 68.275 8.77 ;
      RECT 63.7 5.085 64.02 5.345 ;
      RECT 64.735 5.1 65.025 5.33 ;
      RECT 63.7 5.145 65.025 5.285 ;
      RECT 63.36 7.125 63.68 7.385 ;
      RECT 64.735 7.14 65.025 7.37 ;
      RECT 64.81 6.845 64.95 7.37 ;
      RECT 63.45 6.845 63.59 7.385 ;
      RECT 63.45 6.845 64.95 6.985 ;
      RECT 64.38 4.065 64.7 4.325 ;
      RECT 64.105 4.125 64.7 4.265 ;
      RECT 61.32 7.805 61.64 8.065 ;
      RECT 60.315 7.82 60.605 8.05 ;
      RECT 60.315 7.865 62.23 8.005 ;
      RECT 62.09 7.525 62.23 8.005 ;
      RECT 62.09 7.525 64.1 7.665 ;
      RECT 63.96 7.14 64.1 7.665 ;
      RECT 63.885 7.14 64.175 7.37 ;
      RECT 63.7 6.105 64.02 6.365 ;
      RECT 61.555 6.12 61.845 6.35 ;
      RECT 61.555 6.165 64.02 6.305 ;
      RECT 63.02 5.085 63.34 5.345 ;
      RECT 60.655 5.1 60.945 5.33 ;
      RECT 60.655 5.145 63.34 5.285 ;
      RECT 62.68 7.805 63 8.065 ;
      RECT 62.68 7.865 63.275 8.005 ;
      RECT 62.68 4.405 63 4.665 ;
      RECT 62.405 4.465 63 4.605 ;
      RECT 62 4.065 62.32 4.325 ;
      RECT 61.725 4.125 62.32 4.265 ;
      RECT 61.66 4.745 61.98 5.005 ;
      RECT 58.785 4.76 59.075 4.99 ;
      RECT 58.785 4.805 61.98 4.945 ;
      RECT 61.24 4.085 61.38 4.945 ;
      RECT 61.165 4.085 61.455 4.315 ;
      RECT 61.32 3.555 61.64 3.815 ;
      RECT 61.32 3.57 61.825 3.8 ;
      RECT 61.23 3.615 61.825 3.755 ;
      RECT 60.655 4.085 60.945 4.315 ;
      RECT 60.05 4.13 60.945 4.27 ;
      RECT 60.05 3.725 60.19 4.27 ;
      RECT 59.96 3.725 60.28 3.985 ;
      RECT 59.28 4.065 59.6 4.325 ;
      RECT 59.005 4.125 59.6 4.265 ;
      RECT 59.28 6.105 59.6 6.365 ;
      RECT 59.005 6.165 59.6 6.305 ;
      RECT 57.045 8.86 57.335 9.17 ;
      RECT 56.875 8.97 57.365 9.14 ;
      RECT 57.025 8.86 57.365 9.14 ;
      RECT 56.615 10.05 56.905 10.28 ;
      RECT 56.675 9.28 56.845 10.28 ;
      RECT 56.58 9.28 56.95 9.655 ;
      RECT 53.86 10.055 54.15 10.285 ;
      RECT 53.92 8.575 54.09 10.285 ;
      RECT 53.92 8.94 54.25 9.265 ;
      RECT 53.86 8.575 54.15 8.805 ;
      RECT 53.455 3.69 53.56 4.26 ;
      RECT 53.455 4.025 53.78 4.255 ;
      RECT 53.455 4.055 53.95 4.225 ;
      RECT 53.455 3.69 53.645 4.255 ;
      RECT 52.87 3.655 53.16 3.885 ;
      RECT 52.87 3.69 53.645 3.86 ;
      RECT 52.93 2.175 53.1 3.885 ;
      RECT 52.87 2.175 53.16 2.405 ;
      RECT 52.87 10.055 53.16 10.285 ;
      RECT 52.93 8.575 53.1 10.285 ;
      RECT 52.87 8.575 53.16 8.805 ;
      RECT 52.87 8.61 53.725 8.77 ;
      RECT 53.555 8.205 53.725 8.77 ;
      RECT 52.87 8.605 53.265 8.77 ;
      RECT 53.49 8.205 53.78 8.435 ;
      RECT 53.49 8.235 53.95 8.405 ;
      RECT 52.5 4.025 52.79 4.255 ;
      RECT 52.5 4.055 52.96 4.225 ;
      RECT 52.565 2.95 52.73 4.255 ;
      RECT 51.08 2.92 51.37 3.15 ;
      RECT 51.08 2.95 52.73 3.12 ;
      RECT 51.14 2.18 51.31 3.15 ;
      RECT 51.08 2.18 51.37 2.41 ;
      RECT 51.08 10.05 51.37 10.28 ;
      RECT 51.14 9.31 51.31 10.28 ;
      RECT 51.14 9.405 52.73 9.575 ;
      RECT 52.56 8.205 52.73 9.575 ;
      RECT 51.08 9.31 51.37 9.54 ;
      RECT 52.5 8.205 52.79 8.435 ;
      RECT 52.5 8.235 52.96 8.405 ;
      RECT 51.51 3.26 51.86 3.61 ;
      RECT 51.34 3.32 51.86 3.49 ;
      RECT 51.535 8.94 51.86 9.265 ;
      RECT 51.51 8.94 51.86 9.17 ;
      RECT 51.34 8.97 51.86 9.14 ;
      RECT 50.735 3.66 51.055 3.98 ;
      RECT 50.705 3.66 51.055 3.89 ;
      RECT 50.42 3.69 51.055 3.86 ;
      RECT 50.735 8.565 51.055 8.89 ;
      RECT 50.705 8.57 51.055 8.8 ;
      RECT 50.535 8.6 51.055 8.77 ;
      RECT 46.48 5.085 46.8 5.345 ;
      RECT 47.515 5.1 47.805 5.33 ;
      RECT 46.48 5.145 47.805 5.285 ;
      RECT 46.14 7.125 46.46 7.385 ;
      RECT 47.515 7.14 47.805 7.37 ;
      RECT 47.59 6.845 47.73 7.37 ;
      RECT 46.23 6.845 46.37 7.385 ;
      RECT 46.23 6.845 47.73 6.985 ;
      RECT 47.16 4.065 47.48 4.325 ;
      RECT 46.885 4.125 47.48 4.265 ;
      RECT 44.1 7.805 44.42 8.065 ;
      RECT 43.095 7.82 43.385 8.05 ;
      RECT 43.095 7.865 45.01 8.005 ;
      RECT 44.87 7.525 45.01 8.005 ;
      RECT 44.87 7.525 46.88 7.665 ;
      RECT 46.74 7.14 46.88 7.665 ;
      RECT 46.665 7.14 46.955 7.37 ;
      RECT 46.48 6.105 46.8 6.365 ;
      RECT 44.335 6.12 44.625 6.35 ;
      RECT 44.335 6.165 46.8 6.305 ;
      RECT 45.8 5.085 46.12 5.345 ;
      RECT 43.435 5.1 43.725 5.33 ;
      RECT 43.435 5.145 46.12 5.285 ;
      RECT 45.46 7.805 45.78 8.065 ;
      RECT 45.46 7.865 46.055 8.005 ;
      RECT 45.46 4.405 45.78 4.665 ;
      RECT 45.185 4.465 45.78 4.605 ;
      RECT 44.78 4.065 45.1 4.325 ;
      RECT 44.505 4.125 45.1 4.265 ;
      RECT 44.44 4.745 44.76 5.005 ;
      RECT 41.565 4.76 41.855 4.99 ;
      RECT 41.565 4.805 44.76 4.945 ;
      RECT 44.02 4.085 44.16 4.945 ;
      RECT 43.945 4.085 44.235 4.315 ;
      RECT 44.1 3.555 44.42 3.815 ;
      RECT 44.1 3.57 44.605 3.8 ;
      RECT 44.01 3.615 44.605 3.755 ;
      RECT 43.435 4.085 43.725 4.315 ;
      RECT 42.83 4.13 43.725 4.27 ;
      RECT 42.83 3.725 42.97 4.27 ;
      RECT 42.74 3.725 43.06 3.985 ;
      RECT 42.06 4.065 42.38 4.325 ;
      RECT 41.785 4.125 42.38 4.265 ;
      RECT 42.06 6.105 42.38 6.365 ;
      RECT 41.785 6.165 42.38 6.305 ;
      RECT 39.825 8.86 40.115 9.17 ;
      RECT 39.655 8.97 40.145 9.14 ;
      RECT 39.805 8.86 40.145 9.14 ;
      RECT 39.395 10.05 39.685 10.28 ;
      RECT 39.455 9.28 39.625 10.28 ;
      RECT 39.36 9.28 39.73 9.655 ;
      RECT 36.64 10.055 36.93 10.285 ;
      RECT 36.7 8.575 36.87 10.285 ;
      RECT 36.7 8.94 37.03 9.265 ;
      RECT 36.64 8.575 36.93 8.805 ;
      RECT 36.235 3.69 36.34 4.26 ;
      RECT 36.235 4.025 36.56 4.255 ;
      RECT 36.235 4.055 36.73 4.225 ;
      RECT 36.235 3.69 36.425 4.255 ;
      RECT 35.65 3.655 35.94 3.885 ;
      RECT 35.65 3.69 36.425 3.86 ;
      RECT 35.71 2.175 35.88 3.885 ;
      RECT 35.65 2.175 35.94 2.405 ;
      RECT 35.65 10.055 35.94 10.285 ;
      RECT 35.71 8.575 35.88 10.285 ;
      RECT 35.65 8.575 35.94 8.805 ;
      RECT 35.65 8.61 36.505 8.77 ;
      RECT 36.335 8.205 36.505 8.77 ;
      RECT 35.65 8.605 36.045 8.77 ;
      RECT 36.27 8.205 36.56 8.435 ;
      RECT 36.27 8.235 36.73 8.405 ;
      RECT 35.28 4.025 35.57 4.255 ;
      RECT 35.28 4.055 35.74 4.225 ;
      RECT 35.345 2.95 35.51 4.255 ;
      RECT 33.86 2.92 34.15 3.15 ;
      RECT 33.86 2.95 35.51 3.12 ;
      RECT 33.92 2.18 34.09 3.15 ;
      RECT 33.86 2.18 34.15 2.41 ;
      RECT 33.86 10.05 34.15 10.28 ;
      RECT 33.92 9.31 34.09 10.28 ;
      RECT 33.92 9.405 35.51 9.575 ;
      RECT 35.34 8.205 35.51 9.575 ;
      RECT 33.86 9.31 34.15 9.54 ;
      RECT 35.28 8.205 35.57 8.435 ;
      RECT 35.28 8.235 35.74 8.405 ;
      RECT 34.29 3.26 34.64 3.61 ;
      RECT 34.12 3.32 34.64 3.49 ;
      RECT 34.315 8.94 34.64 9.265 ;
      RECT 34.29 8.94 34.64 9.17 ;
      RECT 34.12 8.97 34.64 9.14 ;
      RECT 33.515 3.66 33.835 3.98 ;
      RECT 33.485 3.66 33.835 3.89 ;
      RECT 33.2 3.69 33.835 3.86 ;
      RECT 33.515 8.565 33.835 8.89 ;
      RECT 33.485 8.57 33.835 8.8 ;
      RECT 33.315 8.6 33.835 8.77 ;
      RECT 29.26 5.085 29.58 5.345 ;
      RECT 30.295 5.1 30.585 5.33 ;
      RECT 29.26 5.145 30.585 5.285 ;
      RECT 28.92 7.125 29.24 7.385 ;
      RECT 30.295 7.14 30.585 7.37 ;
      RECT 30.37 6.845 30.51 7.37 ;
      RECT 29.01 6.845 29.15 7.385 ;
      RECT 29.01 6.845 30.51 6.985 ;
      RECT 29.94 4.065 30.26 4.325 ;
      RECT 29.665 4.125 30.26 4.265 ;
      RECT 26.88 7.805 27.2 8.065 ;
      RECT 25.875 7.82 26.165 8.05 ;
      RECT 25.875 7.865 27.79 8.005 ;
      RECT 27.65 7.525 27.79 8.005 ;
      RECT 27.65 7.525 29.66 7.665 ;
      RECT 29.52 7.14 29.66 7.665 ;
      RECT 29.445 7.14 29.735 7.37 ;
      RECT 29.26 6.105 29.58 6.365 ;
      RECT 27.115 6.12 27.405 6.35 ;
      RECT 27.115 6.165 29.58 6.305 ;
      RECT 28.58 5.085 28.9 5.345 ;
      RECT 26.215 5.1 26.505 5.33 ;
      RECT 26.215 5.145 28.9 5.285 ;
      RECT 28.24 7.805 28.56 8.065 ;
      RECT 28.24 7.865 28.835 8.005 ;
      RECT 28.24 4.405 28.56 4.665 ;
      RECT 27.965 4.465 28.56 4.605 ;
      RECT 27.56 4.065 27.88 4.325 ;
      RECT 27.285 4.125 27.88 4.265 ;
      RECT 27.22 4.745 27.54 5.005 ;
      RECT 24.345 4.76 24.635 4.99 ;
      RECT 24.345 4.805 27.54 4.945 ;
      RECT 26.8 4.085 26.94 4.945 ;
      RECT 26.725 4.085 27.015 4.315 ;
      RECT 26.88 3.555 27.2 3.815 ;
      RECT 26.88 3.57 27.385 3.8 ;
      RECT 26.79 3.615 27.385 3.755 ;
      RECT 26.215 4.085 26.505 4.315 ;
      RECT 25.61 4.13 26.505 4.27 ;
      RECT 25.61 3.725 25.75 4.27 ;
      RECT 25.52 3.725 25.84 3.985 ;
      RECT 24.84 4.065 25.16 4.325 ;
      RECT 24.565 4.125 25.16 4.265 ;
      RECT 24.84 6.105 25.16 6.365 ;
      RECT 24.565 6.165 25.16 6.305 ;
      RECT 22.605 8.86 22.895 9.17 ;
      RECT 22.435 8.97 22.925 9.14 ;
      RECT 22.585 8.86 22.925 9.14 ;
      RECT 22.175 10.05 22.465 10.28 ;
      RECT 22.235 9.28 22.405 10.28 ;
      RECT 22.14 9.28 22.51 9.655 ;
      RECT 19.42 10.055 19.71 10.285 ;
      RECT 19.48 8.575 19.65 10.285 ;
      RECT 19.48 8.94 19.81 9.265 ;
      RECT 19.42 8.575 19.71 8.805 ;
      RECT 19.015 3.69 19.12 4.26 ;
      RECT 19.015 4.025 19.34 4.255 ;
      RECT 19.015 4.055 19.51 4.225 ;
      RECT 19.015 3.69 19.205 4.255 ;
      RECT 18.43 3.655 18.72 3.885 ;
      RECT 18.43 3.69 19.205 3.86 ;
      RECT 18.49 2.175 18.66 3.885 ;
      RECT 18.43 2.175 18.72 2.405 ;
      RECT 18.43 10.055 18.72 10.285 ;
      RECT 18.49 8.575 18.66 10.285 ;
      RECT 18.43 8.575 18.72 8.805 ;
      RECT 18.43 8.61 19.285 8.77 ;
      RECT 19.115 8.205 19.285 8.77 ;
      RECT 18.43 8.605 18.825 8.77 ;
      RECT 19.05 8.205 19.34 8.435 ;
      RECT 19.05 8.235 19.51 8.405 ;
      RECT 18.06 4.025 18.35 4.255 ;
      RECT 18.06 4.055 18.52 4.225 ;
      RECT 18.125 2.95 18.29 4.255 ;
      RECT 16.64 2.92 16.93 3.15 ;
      RECT 16.64 2.95 18.29 3.12 ;
      RECT 16.7 2.18 16.87 3.15 ;
      RECT 16.64 2.18 16.93 2.41 ;
      RECT 16.64 10.05 16.93 10.28 ;
      RECT 16.7 9.31 16.87 10.28 ;
      RECT 16.7 9.405 18.29 9.575 ;
      RECT 18.12 8.205 18.29 9.575 ;
      RECT 16.64 9.31 16.93 9.54 ;
      RECT 18.06 8.205 18.35 8.435 ;
      RECT 18.06 8.235 18.52 8.405 ;
      RECT 17.07 3.26 17.42 3.61 ;
      RECT 16.9 3.32 17.42 3.49 ;
      RECT 17.095 8.94 17.42 9.265 ;
      RECT 17.07 8.94 17.42 9.17 ;
      RECT 16.9 8.97 17.42 9.14 ;
      RECT 16.295 3.66 16.615 3.98 ;
      RECT 16.265 3.66 16.615 3.89 ;
      RECT 15.98 3.69 16.615 3.86 ;
      RECT 16.295 8.565 16.615 8.89 ;
      RECT 16.265 8.57 16.615 8.8 ;
      RECT 16.095 8.6 16.615 8.77 ;
      RECT 12.04 5.085 12.36 5.345 ;
      RECT 13.075 5.1 13.365 5.33 ;
      RECT 12.04 5.145 13.365 5.285 ;
      RECT 11.7 7.125 12.02 7.385 ;
      RECT 13.075 7.14 13.365 7.37 ;
      RECT 13.15 6.845 13.29 7.37 ;
      RECT 11.79 6.845 11.93 7.385 ;
      RECT 11.79 6.845 13.29 6.985 ;
      RECT 12.72 4.065 13.04 4.325 ;
      RECT 12.445 4.125 13.04 4.265 ;
      RECT 9.66 7.805 9.98 8.065 ;
      RECT 8.655 7.82 8.945 8.05 ;
      RECT 8.655 7.865 10.57 8.005 ;
      RECT 10.43 7.525 10.57 8.005 ;
      RECT 10.43 7.525 12.44 7.665 ;
      RECT 12.3 7.14 12.44 7.665 ;
      RECT 12.225 7.14 12.515 7.37 ;
      RECT 12.04 6.105 12.36 6.365 ;
      RECT 9.895 6.12 10.185 6.35 ;
      RECT 9.895 6.165 12.36 6.305 ;
      RECT 11.36 5.085 11.68 5.345 ;
      RECT 8.995 5.1 9.285 5.33 ;
      RECT 8.995 5.145 11.68 5.285 ;
      RECT 11.02 7.805 11.34 8.065 ;
      RECT 11.02 7.865 11.615 8.005 ;
      RECT 11.02 4.405 11.34 4.665 ;
      RECT 10.745 4.465 11.34 4.605 ;
      RECT 10.34 4.065 10.66 4.325 ;
      RECT 10.065 4.125 10.66 4.265 ;
      RECT 10 4.745 10.32 5.005 ;
      RECT 7.125 4.76 7.415 4.99 ;
      RECT 7.125 4.805 10.32 4.945 ;
      RECT 9.58 4.085 9.72 4.945 ;
      RECT 9.505 4.085 9.795 4.315 ;
      RECT 9.66 3.555 9.98 3.815 ;
      RECT 9.66 3.57 10.165 3.8 ;
      RECT 9.57 3.615 10.165 3.755 ;
      RECT 8.995 4.085 9.285 4.315 ;
      RECT 8.39 4.13 9.285 4.27 ;
      RECT 8.39 3.725 8.53 4.27 ;
      RECT 8.3 3.725 8.62 3.985 ;
      RECT 7.62 4.065 7.94 4.325 ;
      RECT 7.345 4.125 7.94 4.265 ;
      RECT 7.62 6.105 7.94 6.365 ;
      RECT 7.345 6.165 7.94 6.305 ;
      RECT 5.385 8.86 5.675 9.17 ;
      RECT 5.215 8.97 5.705 9.14 ;
      RECT 5.365 8.86 5.705 9.14 ;
      RECT 4.955 10.05 5.245 10.28 ;
      RECT 5.015 9.28 5.185 10.28 ;
      RECT 4.92 9.28 5.29 9.655 ;
      RECT 1.545 10.05 1.835 10.28 ;
      RECT 1.605 9.31 1.775 10.28 ;
      RECT 1.515 9.31 1.855 9.59 ;
      RECT 1.14 8.57 1.48 8.85 ;
      RECT 1 8.6 1.48 8.77 ;
      RECT 83.505 3.29 83.83 3.615 ;
      RECT 81.275 7.805 81.92 8.065 ;
      RECT 79.225 7.125 79.87 7.385 ;
      RECT 66.285 3.29 66.61 3.615 ;
      RECT 64.055 7.805 64.7 8.065 ;
      RECT 62.005 7.125 62.65 7.385 ;
      RECT 49.065 3.29 49.39 3.615 ;
      RECT 46.835 7.805 47.48 8.065 ;
      RECT 44.785 7.125 45.43 7.385 ;
      RECT 31.845 3.29 32.17 3.615 ;
      RECT 29.615 7.805 30.26 8.065 ;
      RECT 27.565 7.125 28.21 7.385 ;
      RECT 14.625 3.29 14.95 3.615 ;
      RECT 12.395 7.805 13.04 8.065 ;
      RECT 10.345 7.125 10.99 7.385 ;
    LAYER mcon ;
      RECT 88.36 8.605 88.53 8.775 ;
      RECT 88.36 10.085 88.53 10.255 ;
      RECT 87.99 4.055 88.16 4.225 ;
      RECT 87.99 8.235 88.16 8.405 ;
      RECT 87.37 2.205 87.54 2.375 ;
      RECT 87.37 3.685 87.54 3.855 ;
      RECT 87.37 8.605 87.54 8.775 ;
      RECT 87.37 10.085 87.54 10.255 ;
      RECT 87 4.055 87.17 4.225 ;
      RECT 87 8.235 87.17 8.405 ;
      RECT 86.01 3.32 86.18 3.49 ;
      RECT 86.01 8.97 86.18 9.14 ;
      RECT 85.58 2.21 85.75 2.38 ;
      RECT 85.58 2.95 85.75 3.12 ;
      RECT 85.58 9.34 85.75 9.51 ;
      RECT 85.58 10.08 85.75 10.25 ;
      RECT 85.205 3.69 85.375 3.86 ;
      RECT 85.205 8.6 85.375 8.77 ;
      RECT 82.015 5.13 82.185 5.3 ;
      RECT 82.015 7.17 82.185 7.34 ;
      RECT 81.675 4.11 81.845 4.28 ;
      RECT 81.335 7.85 81.505 8.02 ;
      RECT 81.165 7.17 81.335 7.34 ;
      RECT 80.655 7.17 80.825 7.34 ;
      RECT 79.975 4.45 80.145 4.62 ;
      RECT 79.975 7.85 80.145 8.02 ;
      RECT 79.295 4.11 79.465 4.28 ;
      RECT 79.285 7.17 79.455 7.34 ;
      RECT 78.835 6.15 79.005 6.32 ;
      RECT 78.815 3.6 78.985 3.77 ;
      RECT 78.445 4.115 78.615 4.285 ;
      RECT 77.935 4.115 78.105 4.285 ;
      RECT 77.935 5.13 78.105 5.3 ;
      RECT 77.595 7.85 77.765 8.02 ;
      RECT 76.575 4.11 76.745 4.28 ;
      RECT 76.575 6.15 76.745 6.32 ;
      RECT 76.065 4.79 76.235 4.96 ;
      RECT 74.325 8.97 74.495 9.14 ;
      RECT 73.895 9.34 74.065 9.51 ;
      RECT 73.895 10.08 74.065 10.25 ;
      RECT 71.14 8.605 71.31 8.775 ;
      RECT 71.14 10.085 71.31 10.255 ;
      RECT 70.77 4.055 70.94 4.225 ;
      RECT 70.77 8.235 70.94 8.405 ;
      RECT 70.15 2.205 70.32 2.375 ;
      RECT 70.15 3.685 70.32 3.855 ;
      RECT 70.15 8.605 70.32 8.775 ;
      RECT 70.15 10.085 70.32 10.255 ;
      RECT 69.78 4.055 69.95 4.225 ;
      RECT 69.78 8.235 69.95 8.405 ;
      RECT 68.79 3.32 68.96 3.49 ;
      RECT 68.79 8.97 68.96 9.14 ;
      RECT 68.36 2.21 68.53 2.38 ;
      RECT 68.36 2.95 68.53 3.12 ;
      RECT 68.36 9.34 68.53 9.51 ;
      RECT 68.36 10.08 68.53 10.25 ;
      RECT 67.985 3.69 68.155 3.86 ;
      RECT 67.985 8.6 68.155 8.77 ;
      RECT 64.795 5.13 64.965 5.3 ;
      RECT 64.795 7.17 64.965 7.34 ;
      RECT 64.455 4.11 64.625 4.28 ;
      RECT 64.115 7.85 64.285 8.02 ;
      RECT 63.945 7.17 64.115 7.34 ;
      RECT 63.435 7.17 63.605 7.34 ;
      RECT 62.755 4.45 62.925 4.62 ;
      RECT 62.755 7.85 62.925 8.02 ;
      RECT 62.075 4.11 62.245 4.28 ;
      RECT 62.065 7.17 62.235 7.34 ;
      RECT 61.615 6.15 61.785 6.32 ;
      RECT 61.595 3.6 61.765 3.77 ;
      RECT 61.225 4.115 61.395 4.285 ;
      RECT 60.715 4.115 60.885 4.285 ;
      RECT 60.715 5.13 60.885 5.3 ;
      RECT 60.375 7.85 60.545 8.02 ;
      RECT 59.355 4.11 59.525 4.28 ;
      RECT 59.355 6.15 59.525 6.32 ;
      RECT 58.845 4.79 59.015 4.96 ;
      RECT 57.105 8.97 57.275 9.14 ;
      RECT 56.675 9.34 56.845 9.51 ;
      RECT 56.675 10.08 56.845 10.25 ;
      RECT 53.92 8.605 54.09 8.775 ;
      RECT 53.92 10.085 54.09 10.255 ;
      RECT 53.55 4.055 53.72 4.225 ;
      RECT 53.55 8.235 53.72 8.405 ;
      RECT 52.93 2.205 53.1 2.375 ;
      RECT 52.93 3.685 53.1 3.855 ;
      RECT 52.93 8.605 53.1 8.775 ;
      RECT 52.93 10.085 53.1 10.255 ;
      RECT 52.56 4.055 52.73 4.225 ;
      RECT 52.56 8.235 52.73 8.405 ;
      RECT 51.57 3.32 51.74 3.49 ;
      RECT 51.57 8.97 51.74 9.14 ;
      RECT 51.14 2.21 51.31 2.38 ;
      RECT 51.14 2.95 51.31 3.12 ;
      RECT 51.14 9.34 51.31 9.51 ;
      RECT 51.14 10.08 51.31 10.25 ;
      RECT 50.765 3.69 50.935 3.86 ;
      RECT 50.765 8.6 50.935 8.77 ;
      RECT 47.575 5.13 47.745 5.3 ;
      RECT 47.575 7.17 47.745 7.34 ;
      RECT 47.235 4.11 47.405 4.28 ;
      RECT 46.895 7.85 47.065 8.02 ;
      RECT 46.725 7.17 46.895 7.34 ;
      RECT 46.215 7.17 46.385 7.34 ;
      RECT 45.535 4.45 45.705 4.62 ;
      RECT 45.535 7.85 45.705 8.02 ;
      RECT 44.855 4.11 45.025 4.28 ;
      RECT 44.845 7.17 45.015 7.34 ;
      RECT 44.395 6.15 44.565 6.32 ;
      RECT 44.375 3.6 44.545 3.77 ;
      RECT 44.005 4.115 44.175 4.285 ;
      RECT 43.495 4.115 43.665 4.285 ;
      RECT 43.495 5.13 43.665 5.3 ;
      RECT 43.155 7.85 43.325 8.02 ;
      RECT 42.135 4.11 42.305 4.28 ;
      RECT 42.135 6.15 42.305 6.32 ;
      RECT 41.625 4.79 41.795 4.96 ;
      RECT 39.885 8.97 40.055 9.14 ;
      RECT 39.455 9.34 39.625 9.51 ;
      RECT 39.455 10.08 39.625 10.25 ;
      RECT 36.7 8.605 36.87 8.775 ;
      RECT 36.7 10.085 36.87 10.255 ;
      RECT 36.33 4.055 36.5 4.225 ;
      RECT 36.33 8.235 36.5 8.405 ;
      RECT 35.71 2.205 35.88 2.375 ;
      RECT 35.71 3.685 35.88 3.855 ;
      RECT 35.71 8.605 35.88 8.775 ;
      RECT 35.71 10.085 35.88 10.255 ;
      RECT 35.34 4.055 35.51 4.225 ;
      RECT 35.34 8.235 35.51 8.405 ;
      RECT 34.35 3.32 34.52 3.49 ;
      RECT 34.35 8.97 34.52 9.14 ;
      RECT 33.92 2.21 34.09 2.38 ;
      RECT 33.92 2.95 34.09 3.12 ;
      RECT 33.92 9.34 34.09 9.51 ;
      RECT 33.92 10.08 34.09 10.25 ;
      RECT 33.545 3.69 33.715 3.86 ;
      RECT 33.545 8.6 33.715 8.77 ;
      RECT 30.355 5.13 30.525 5.3 ;
      RECT 30.355 7.17 30.525 7.34 ;
      RECT 30.015 4.11 30.185 4.28 ;
      RECT 29.675 7.85 29.845 8.02 ;
      RECT 29.505 7.17 29.675 7.34 ;
      RECT 28.995 7.17 29.165 7.34 ;
      RECT 28.315 4.45 28.485 4.62 ;
      RECT 28.315 7.85 28.485 8.02 ;
      RECT 27.635 4.11 27.805 4.28 ;
      RECT 27.625 7.17 27.795 7.34 ;
      RECT 27.175 6.15 27.345 6.32 ;
      RECT 27.155 3.6 27.325 3.77 ;
      RECT 26.785 4.115 26.955 4.285 ;
      RECT 26.275 4.115 26.445 4.285 ;
      RECT 26.275 5.13 26.445 5.3 ;
      RECT 25.935 7.85 26.105 8.02 ;
      RECT 24.915 4.11 25.085 4.28 ;
      RECT 24.915 6.15 25.085 6.32 ;
      RECT 24.405 4.79 24.575 4.96 ;
      RECT 22.665 8.97 22.835 9.14 ;
      RECT 22.235 9.34 22.405 9.51 ;
      RECT 22.235 10.08 22.405 10.25 ;
      RECT 19.48 8.605 19.65 8.775 ;
      RECT 19.48 10.085 19.65 10.255 ;
      RECT 19.11 4.055 19.28 4.225 ;
      RECT 19.11 8.235 19.28 8.405 ;
      RECT 18.49 2.205 18.66 2.375 ;
      RECT 18.49 3.685 18.66 3.855 ;
      RECT 18.49 8.605 18.66 8.775 ;
      RECT 18.49 10.085 18.66 10.255 ;
      RECT 18.12 4.055 18.29 4.225 ;
      RECT 18.12 8.235 18.29 8.405 ;
      RECT 17.13 3.32 17.3 3.49 ;
      RECT 17.13 8.97 17.3 9.14 ;
      RECT 16.7 2.21 16.87 2.38 ;
      RECT 16.7 2.95 16.87 3.12 ;
      RECT 16.7 9.34 16.87 9.51 ;
      RECT 16.7 10.08 16.87 10.25 ;
      RECT 16.325 3.69 16.495 3.86 ;
      RECT 16.325 8.6 16.495 8.77 ;
      RECT 13.135 5.13 13.305 5.3 ;
      RECT 13.135 7.17 13.305 7.34 ;
      RECT 12.795 4.11 12.965 4.28 ;
      RECT 12.455 7.85 12.625 8.02 ;
      RECT 12.285 7.17 12.455 7.34 ;
      RECT 11.775 7.17 11.945 7.34 ;
      RECT 11.095 4.45 11.265 4.62 ;
      RECT 11.095 7.85 11.265 8.02 ;
      RECT 10.415 4.11 10.585 4.28 ;
      RECT 10.405 7.17 10.575 7.34 ;
      RECT 9.955 6.15 10.125 6.32 ;
      RECT 9.935 3.6 10.105 3.77 ;
      RECT 9.565 4.115 9.735 4.285 ;
      RECT 9.055 4.115 9.225 4.285 ;
      RECT 9.055 5.13 9.225 5.3 ;
      RECT 8.715 7.85 8.885 8.02 ;
      RECT 7.695 4.11 7.865 4.28 ;
      RECT 7.695 6.15 7.865 6.32 ;
      RECT 7.185 4.79 7.355 4.96 ;
      RECT 5.445 8.97 5.615 9.14 ;
      RECT 5.015 9.34 5.185 9.51 ;
      RECT 5.015 10.08 5.185 10.25 ;
      RECT 1.605 9.34 1.775 9.51 ;
      RECT 1.605 10.08 1.775 10.25 ;
      RECT 1.23 8.6 1.4 8.77 ;
    LAYER li1 ;
      RECT 87.99 3.035 88.16 4.225 ;
      RECT 87.99 3.035 88.46 3.205 ;
      RECT 87.99 9.255 88.46 9.425 ;
      RECT 87.99 8.235 88.16 9.425 ;
      RECT 87 3.035 87.17 4.225 ;
      RECT 87 3.035 87.47 3.205 ;
      RECT 87 9.255 87.47 9.425 ;
      RECT 87 8.235 87.17 9.425 ;
      RECT 85.15 3.93 85.32 5.16 ;
      RECT 85.205 2.15 85.375 4.1 ;
      RECT 85.15 1.87 85.32 2.32 ;
      RECT 85.15 10.14 85.32 10.59 ;
      RECT 85.205 8.36 85.375 10.31 ;
      RECT 85.15 7.3 85.32 8.53 ;
      RECT 84.63 1.87 84.8 5.16 ;
      RECT 84.63 3.37 85.035 3.7 ;
      RECT 84.63 2.53 85.035 2.86 ;
      RECT 84.63 7.3 84.8 10.59 ;
      RECT 84.63 9.6 85.035 9.93 ;
      RECT 84.63 8.76 85.035 9.09 ;
      RECT 82.365 4.79 82.745 5.47 ;
      RECT 82.575 3.66 82.745 5.47 ;
      RECT 80.495 3.66 80.725 4.33 ;
      RECT 80.495 3.66 82.745 3.83 ;
      RECT 82.025 3.34 82.195 3.83 ;
      RECT 82.015 4.45 82.185 5.3 ;
      RECT 81.1 4.45 82.405 4.62 ;
      RECT 82.16 4 82.405 4.62 ;
      RECT 81.1 4.08 81.27 4.62 ;
      RECT 80.895 4.08 81.27 4.25 ;
      RECT 81.075 7.56 81.77 8.19 ;
      RECT 81.6 5.98 81.77 8.19 ;
      RECT 81.505 5.98 81.835 6.96 ;
      RECT 81.105 4.79 81.435 5.47 ;
      RECT 80.195 4.79 80.595 5.47 ;
      RECT 80.195 4.79 81.435 4.96 ;
      RECT 79.695 4.37 80.015 5.47 ;
      RECT 79.695 4.37 80.145 4.62 ;
      RECT 79.695 4.37 80.325 4.54 ;
      RECT 80.155 3.32 80.325 4.54 ;
      RECT 80.155 3.32 81.11 3.49 ;
      RECT 79.695 7.56 80.39 8.19 ;
      RECT 80.22 5.98 80.39 8.19 ;
      RECT 80.125 5.98 80.455 6.96 ;
      RECT 79.715 7.12 80.05 7.37 ;
      RECT 79.17 7.12 79.505 7.37 ;
      RECT 79.17 7.17 80.05 7.34 ;
      RECT 78.83 7.56 79.525 8.19 ;
      RECT 78.83 5.98 79 8.19 ;
      RECT 78.765 5.98 79.095 6.96 ;
      RECT 78.325 4.5 78.655 5.455 ;
      RECT 78.325 4.5 79.005 4.67 ;
      RECT 78.835 3.26 79.005 4.67 ;
      RECT 78.745 3.26 79.075 3.9 ;
      RECT 77.805 4.5 78.135 5.455 ;
      RECT 77.455 4.5 78.135 4.67 ;
      RECT 77.455 3.26 77.625 4.67 ;
      RECT 77.385 3.26 77.715 3.9 ;
      RECT 77.595 7.17 77.765 8.02 ;
      RECT 76.87 7.12 77.205 7.37 ;
      RECT 76.87 7.17 77.765 7.34 ;
      RECT 76.935 4.08 77.285 4.33 ;
      RECT 76.415 4.08 76.745 4.33 ;
      RECT 76.415 4.11 77.285 4.28 ;
      RECT 76.53 7.56 77.225 8.19 ;
      RECT 76.53 5.98 76.7 8.19 ;
      RECT 76.465 5.98 76.795 6.96 ;
      RECT 75.995 4.49 76.325 5.47 ;
      RECT 75.995 3.26 76.245 5.47 ;
      RECT 75.995 3.26 76.325 3.89 ;
      RECT 72.945 7.3 73.115 10.59 ;
      RECT 72.945 9.6 73.35 9.93 ;
      RECT 72.945 8.76 73.35 9.09 ;
      RECT 70.77 3.035 70.94 4.225 ;
      RECT 70.77 3.035 71.24 3.205 ;
      RECT 70.77 9.255 71.24 9.425 ;
      RECT 70.77 8.235 70.94 9.425 ;
      RECT 69.78 3.035 69.95 4.225 ;
      RECT 69.78 3.035 70.25 3.205 ;
      RECT 69.78 9.255 70.25 9.425 ;
      RECT 69.78 8.235 69.95 9.425 ;
      RECT 67.93 3.93 68.1 5.16 ;
      RECT 67.985 2.15 68.155 4.1 ;
      RECT 67.93 1.87 68.1 2.32 ;
      RECT 67.93 10.14 68.1 10.59 ;
      RECT 67.985 8.36 68.155 10.31 ;
      RECT 67.93 7.3 68.1 8.53 ;
      RECT 67.41 1.87 67.58 5.16 ;
      RECT 67.41 3.37 67.815 3.7 ;
      RECT 67.41 2.53 67.815 2.86 ;
      RECT 67.41 7.3 67.58 10.59 ;
      RECT 67.41 9.6 67.815 9.93 ;
      RECT 67.41 8.76 67.815 9.09 ;
      RECT 65.145 4.79 65.525 5.47 ;
      RECT 65.355 3.66 65.525 5.47 ;
      RECT 63.275 3.66 63.505 4.33 ;
      RECT 63.275 3.66 65.525 3.83 ;
      RECT 64.805 3.34 64.975 3.83 ;
      RECT 64.795 4.45 64.965 5.3 ;
      RECT 63.88 4.45 65.185 4.62 ;
      RECT 64.94 4 65.185 4.62 ;
      RECT 63.88 4.08 64.05 4.62 ;
      RECT 63.675 4.08 64.05 4.25 ;
      RECT 63.855 7.56 64.55 8.19 ;
      RECT 64.38 5.98 64.55 8.19 ;
      RECT 64.285 5.98 64.615 6.96 ;
      RECT 63.885 4.79 64.215 5.47 ;
      RECT 62.975 4.79 63.375 5.47 ;
      RECT 62.975 4.79 64.215 4.96 ;
      RECT 62.475 4.37 62.795 5.47 ;
      RECT 62.475 4.37 62.925 4.62 ;
      RECT 62.475 4.37 63.105 4.54 ;
      RECT 62.935 3.32 63.105 4.54 ;
      RECT 62.935 3.32 63.89 3.49 ;
      RECT 62.475 7.56 63.17 8.19 ;
      RECT 63 5.98 63.17 8.19 ;
      RECT 62.905 5.98 63.235 6.96 ;
      RECT 62.495 7.12 62.83 7.37 ;
      RECT 61.95 7.12 62.285 7.37 ;
      RECT 61.95 7.17 62.83 7.34 ;
      RECT 61.61 7.56 62.305 8.19 ;
      RECT 61.61 5.98 61.78 8.19 ;
      RECT 61.545 5.98 61.875 6.96 ;
      RECT 61.105 4.5 61.435 5.455 ;
      RECT 61.105 4.5 61.785 4.67 ;
      RECT 61.615 3.26 61.785 4.67 ;
      RECT 61.525 3.26 61.855 3.9 ;
      RECT 60.585 4.5 60.915 5.455 ;
      RECT 60.235 4.5 60.915 4.67 ;
      RECT 60.235 3.26 60.405 4.67 ;
      RECT 60.165 3.26 60.495 3.9 ;
      RECT 60.375 7.17 60.545 8.02 ;
      RECT 59.65 7.12 59.985 7.37 ;
      RECT 59.65 7.17 60.545 7.34 ;
      RECT 59.715 4.08 60.065 4.33 ;
      RECT 59.195 4.08 59.525 4.33 ;
      RECT 59.195 4.11 60.065 4.28 ;
      RECT 59.31 7.56 60.005 8.19 ;
      RECT 59.31 5.98 59.48 8.19 ;
      RECT 59.245 5.98 59.575 6.96 ;
      RECT 58.775 4.49 59.105 5.47 ;
      RECT 58.775 3.26 59.025 5.47 ;
      RECT 58.775 3.26 59.105 3.89 ;
      RECT 55.725 7.3 55.895 10.59 ;
      RECT 55.725 9.6 56.13 9.93 ;
      RECT 55.725 8.76 56.13 9.09 ;
      RECT 53.55 3.035 53.72 4.225 ;
      RECT 53.55 3.035 54.02 3.205 ;
      RECT 53.55 9.255 54.02 9.425 ;
      RECT 53.55 8.235 53.72 9.425 ;
      RECT 52.56 3.035 52.73 4.225 ;
      RECT 52.56 3.035 53.03 3.205 ;
      RECT 52.56 9.255 53.03 9.425 ;
      RECT 52.56 8.235 52.73 9.425 ;
      RECT 50.71 3.93 50.88 5.16 ;
      RECT 50.765 2.15 50.935 4.1 ;
      RECT 50.71 1.87 50.88 2.32 ;
      RECT 50.71 10.14 50.88 10.59 ;
      RECT 50.765 8.36 50.935 10.31 ;
      RECT 50.71 7.3 50.88 8.53 ;
      RECT 50.19 1.87 50.36 5.16 ;
      RECT 50.19 3.37 50.595 3.7 ;
      RECT 50.19 2.53 50.595 2.86 ;
      RECT 50.19 7.3 50.36 10.59 ;
      RECT 50.19 9.6 50.595 9.93 ;
      RECT 50.19 8.76 50.595 9.09 ;
      RECT 47.925 4.79 48.305 5.47 ;
      RECT 48.135 3.66 48.305 5.47 ;
      RECT 46.055 3.66 46.285 4.33 ;
      RECT 46.055 3.66 48.305 3.83 ;
      RECT 47.585 3.34 47.755 3.83 ;
      RECT 47.575 4.45 47.745 5.3 ;
      RECT 46.66 4.45 47.965 4.62 ;
      RECT 47.72 4 47.965 4.62 ;
      RECT 46.66 4.08 46.83 4.62 ;
      RECT 46.455 4.08 46.83 4.25 ;
      RECT 46.635 7.56 47.33 8.19 ;
      RECT 47.16 5.98 47.33 8.19 ;
      RECT 47.065 5.98 47.395 6.96 ;
      RECT 46.665 4.79 46.995 5.47 ;
      RECT 45.755 4.79 46.155 5.47 ;
      RECT 45.755 4.79 46.995 4.96 ;
      RECT 45.255 4.37 45.575 5.47 ;
      RECT 45.255 4.37 45.705 4.62 ;
      RECT 45.255 4.37 45.885 4.54 ;
      RECT 45.715 3.32 45.885 4.54 ;
      RECT 45.715 3.32 46.67 3.49 ;
      RECT 45.255 7.56 45.95 8.19 ;
      RECT 45.78 5.98 45.95 8.19 ;
      RECT 45.685 5.98 46.015 6.96 ;
      RECT 45.275 7.12 45.61 7.37 ;
      RECT 44.73 7.12 45.065 7.37 ;
      RECT 44.73 7.17 45.61 7.34 ;
      RECT 44.39 7.56 45.085 8.19 ;
      RECT 44.39 5.98 44.56 8.19 ;
      RECT 44.325 5.98 44.655 6.96 ;
      RECT 43.885 4.5 44.215 5.455 ;
      RECT 43.885 4.5 44.565 4.67 ;
      RECT 44.395 3.26 44.565 4.67 ;
      RECT 44.305 3.26 44.635 3.9 ;
      RECT 43.365 4.5 43.695 5.455 ;
      RECT 43.015 4.5 43.695 4.67 ;
      RECT 43.015 3.26 43.185 4.67 ;
      RECT 42.945 3.26 43.275 3.9 ;
      RECT 43.155 7.17 43.325 8.02 ;
      RECT 42.43 7.12 42.765 7.37 ;
      RECT 42.43 7.17 43.325 7.34 ;
      RECT 42.495 4.08 42.845 4.33 ;
      RECT 41.975 4.08 42.305 4.33 ;
      RECT 41.975 4.11 42.845 4.28 ;
      RECT 42.09 7.56 42.785 8.19 ;
      RECT 42.09 5.98 42.26 8.19 ;
      RECT 42.025 5.98 42.355 6.96 ;
      RECT 41.555 4.49 41.885 5.47 ;
      RECT 41.555 3.26 41.805 5.47 ;
      RECT 41.555 3.26 41.885 3.89 ;
      RECT 38.505 7.3 38.675 10.59 ;
      RECT 38.505 9.6 38.91 9.93 ;
      RECT 38.505 8.76 38.91 9.09 ;
      RECT 36.33 3.035 36.5 4.225 ;
      RECT 36.33 3.035 36.8 3.205 ;
      RECT 36.33 9.255 36.8 9.425 ;
      RECT 36.33 8.235 36.5 9.425 ;
      RECT 35.34 3.035 35.51 4.225 ;
      RECT 35.34 3.035 35.81 3.205 ;
      RECT 35.34 9.255 35.81 9.425 ;
      RECT 35.34 8.235 35.51 9.425 ;
      RECT 33.49 3.93 33.66 5.16 ;
      RECT 33.545 2.15 33.715 4.1 ;
      RECT 33.49 1.87 33.66 2.32 ;
      RECT 33.49 10.14 33.66 10.59 ;
      RECT 33.545 8.36 33.715 10.31 ;
      RECT 33.49 7.3 33.66 8.53 ;
      RECT 32.97 1.87 33.14 5.16 ;
      RECT 32.97 3.37 33.375 3.7 ;
      RECT 32.97 2.53 33.375 2.86 ;
      RECT 32.97 7.3 33.14 10.59 ;
      RECT 32.97 9.6 33.375 9.93 ;
      RECT 32.97 8.76 33.375 9.09 ;
      RECT 30.705 4.79 31.085 5.47 ;
      RECT 30.915 3.66 31.085 5.47 ;
      RECT 28.835 3.66 29.065 4.33 ;
      RECT 28.835 3.66 31.085 3.83 ;
      RECT 30.365 3.34 30.535 3.83 ;
      RECT 30.355 4.45 30.525 5.3 ;
      RECT 29.44 4.45 30.745 4.62 ;
      RECT 30.5 4 30.745 4.62 ;
      RECT 29.44 4.08 29.61 4.62 ;
      RECT 29.235 4.08 29.61 4.25 ;
      RECT 29.415 7.56 30.11 8.19 ;
      RECT 29.94 5.98 30.11 8.19 ;
      RECT 29.845 5.98 30.175 6.96 ;
      RECT 29.445 4.79 29.775 5.47 ;
      RECT 28.535 4.79 28.935 5.47 ;
      RECT 28.535 4.79 29.775 4.96 ;
      RECT 28.035 4.37 28.355 5.47 ;
      RECT 28.035 4.37 28.485 4.62 ;
      RECT 28.035 4.37 28.665 4.54 ;
      RECT 28.495 3.32 28.665 4.54 ;
      RECT 28.495 3.32 29.45 3.49 ;
      RECT 28.035 7.56 28.73 8.19 ;
      RECT 28.56 5.98 28.73 8.19 ;
      RECT 28.465 5.98 28.795 6.96 ;
      RECT 28.055 7.12 28.39 7.37 ;
      RECT 27.51 7.12 27.845 7.37 ;
      RECT 27.51 7.17 28.39 7.34 ;
      RECT 27.17 7.56 27.865 8.19 ;
      RECT 27.17 5.98 27.34 8.19 ;
      RECT 27.105 5.98 27.435 6.96 ;
      RECT 26.665 4.5 26.995 5.455 ;
      RECT 26.665 4.5 27.345 4.67 ;
      RECT 27.175 3.26 27.345 4.67 ;
      RECT 27.085 3.26 27.415 3.9 ;
      RECT 26.145 4.5 26.475 5.455 ;
      RECT 25.795 4.5 26.475 4.67 ;
      RECT 25.795 3.26 25.965 4.67 ;
      RECT 25.725 3.26 26.055 3.9 ;
      RECT 25.935 7.17 26.105 8.02 ;
      RECT 25.21 7.12 25.545 7.37 ;
      RECT 25.21 7.17 26.105 7.34 ;
      RECT 25.275 4.08 25.625 4.33 ;
      RECT 24.755 4.08 25.085 4.33 ;
      RECT 24.755 4.11 25.625 4.28 ;
      RECT 24.87 7.56 25.565 8.19 ;
      RECT 24.87 5.98 25.04 8.19 ;
      RECT 24.805 5.98 25.135 6.96 ;
      RECT 24.335 4.49 24.665 5.47 ;
      RECT 24.335 3.26 24.585 5.47 ;
      RECT 24.335 3.26 24.665 3.89 ;
      RECT 21.285 7.3 21.455 10.59 ;
      RECT 21.285 9.6 21.69 9.93 ;
      RECT 21.285 8.76 21.69 9.09 ;
      RECT 19.11 3.035 19.28 4.225 ;
      RECT 19.11 3.035 19.58 3.205 ;
      RECT 19.11 9.255 19.58 9.425 ;
      RECT 19.11 8.235 19.28 9.425 ;
      RECT 18.12 3.035 18.29 4.225 ;
      RECT 18.12 3.035 18.59 3.205 ;
      RECT 18.12 9.255 18.59 9.425 ;
      RECT 18.12 8.235 18.29 9.425 ;
      RECT 16.27 3.93 16.44 5.16 ;
      RECT 16.325 2.15 16.495 4.1 ;
      RECT 16.27 1.87 16.44 2.32 ;
      RECT 16.27 10.14 16.44 10.59 ;
      RECT 16.325 8.36 16.495 10.31 ;
      RECT 16.27 7.3 16.44 8.53 ;
      RECT 15.75 1.87 15.92 5.16 ;
      RECT 15.75 3.37 16.155 3.7 ;
      RECT 15.75 2.53 16.155 2.86 ;
      RECT 15.75 7.3 15.92 10.59 ;
      RECT 15.75 9.6 16.155 9.93 ;
      RECT 15.75 8.76 16.155 9.09 ;
      RECT 13.485 4.79 13.865 5.47 ;
      RECT 13.695 3.66 13.865 5.47 ;
      RECT 11.615 3.66 11.845 4.33 ;
      RECT 11.615 3.66 13.865 3.83 ;
      RECT 13.145 3.34 13.315 3.83 ;
      RECT 13.135 4.45 13.305 5.3 ;
      RECT 12.22 4.45 13.525 4.62 ;
      RECT 13.28 4 13.525 4.62 ;
      RECT 12.22 4.08 12.39 4.62 ;
      RECT 12.015 4.08 12.39 4.25 ;
      RECT 12.195 7.56 12.89 8.19 ;
      RECT 12.72 5.98 12.89 8.19 ;
      RECT 12.625 5.98 12.955 6.96 ;
      RECT 12.225 4.79 12.555 5.47 ;
      RECT 11.315 4.79 11.715 5.47 ;
      RECT 11.315 4.79 12.555 4.96 ;
      RECT 10.815 4.37 11.135 5.47 ;
      RECT 10.815 4.37 11.265 4.62 ;
      RECT 10.815 4.37 11.445 4.54 ;
      RECT 11.275 3.32 11.445 4.54 ;
      RECT 11.275 3.32 12.23 3.49 ;
      RECT 10.815 7.56 11.51 8.19 ;
      RECT 11.34 5.98 11.51 8.19 ;
      RECT 11.245 5.98 11.575 6.96 ;
      RECT 10.835 7.12 11.17 7.37 ;
      RECT 10.29 7.12 10.625 7.37 ;
      RECT 10.29 7.17 11.17 7.34 ;
      RECT 9.95 7.56 10.645 8.19 ;
      RECT 9.95 5.98 10.12 8.19 ;
      RECT 9.885 5.98 10.215 6.96 ;
      RECT 9.445 4.5 9.775 5.455 ;
      RECT 9.445 4.5 10.125 4.67 ;
      RECT 9.955 3.26 10.125 4.67 ;
      RECT 9.865 3.26 10.195 3.9 ;
      RECT 8.925 4.5 9.255 5.455 ;
      RECT 8.575 4.5 9.255 4.67 ;
      RECT 8.575 3.26 8.745 4.67 ;
      RECT 8.505 3.26 8.835 3.9 ;
      RECT 8.715 7.17 8.885 8.02 ;
      RECT 7.99 7.12 8.325 7.37 ;
      RECT 7.99 7.17 8.885 7.34 ;
      RECT 8.055 4.08 8.405 4.33 ;
      RECT 7.535 4.08 7.865 4.33 ;
      RECT 7.535 4.11 8.405 4.28 ;
      RECT 7.65 7.56 8.345 8.19 ;
      RECT 7.65 5.98 7.82 8.19 ;
      RECT 7.585 5.98 7.915 6.96 ;
      RECT 7.115 4.49 7.445 5.47 ;
      RECT 7.115 3.26 7.365 5.47 ;
      RECT 7.115 3.26 7.445 3.89 ;
      RECT 4.065 7.3 4.235 10.59 ;
      RECT 4.065 9.6 4.47 9.93 ;
      RECT 4.065 8.76 4.47 9.09 ;
      RECT 1.175 10.14 1.345 10.59 ;
      RECT 1.23 8.36 1.4 10.31 ;
      RECT 1.175 7.3 1.345 8.53 ;
      RECT 0.655 7.3 0.825 10.59 ;
      RECT 0.655 9.6 1.06 9.93 ;
      RECT 0.655 8.76 1.06 9.09 ;
      RECT 88.36 7.305 88.53 8.775 ;
      RECT 88.36 10.085 88.53 10.595 ;
      RECT 87.37 1.865 87.54 2.375 ;
      RECT 87.37 3.685 87.54 5.155 ;
      RECT 87.37 7.305 87.54 8.775 ;
      RECT 87.37 10.085 87.54 10.595 ;
      RECT 86.01 1.87 86.18 5.16 ;
      RECT 86.01 7.3 86.18 10.59 ;
      RECT 85.58 1.87 85.75 2.38 ;
      RECT 85.58 2.95 85.75 5.16 ;
      RECT 85.58 7.3 85.75 9.51 ;
      RECT 85.58 10.08 85.75 10.59 ;
      RECT 81.94 7.12 82.275 7.39 ;
      RECT 81.44 4.08 81.99 4.28 ;
      RECT 81.095 7.12 81.43 7.37 ;
      RECT 80.56 7.12 80.895 7.39 ;
      RECT 79.175 4.08 79.525 4.33 ;
      RECT 78.315 4.08 78.665 4.33 ;
      RECT 77.795 4.08 78.145 4.33 ;
      RECT 74.325 7.3 74.495 10.59 ;
      RECT 73.895 7.3 74.065 9.51 ;
      RECT 73.895 10.08 74.065 10.59 ;
      RECT 71.14 7.305 71.31 8.775 ;
      RECT 71.14 10.085 71.31 10.595 ;
      RECT 70.15 1.865 70.32 2.375 ;
      RECT 70.15 3.685 70.32 5.155 ;
      RECT 70.15 7.305 70.32 8.775 ;
      RECT 70.15 10.085 70.32 10.595 ;
      RECT 68.79 1.87 68.96 5.16 ;
      RECT 68.79 7.3 68.96 10.59 ;
      RECT 68.36 1.87 68.53 2.38 ;
      RECT 68.36 2.95 68.53 5.16 ;
      RECT 68.36 7.3 68.53 9.51 ;
      RECT 68.36 10.08 68.53 10.59 ;
      RECT 64.72 7.12 65.055 7.39 ;
      RECT 64.22 4.08 64.77 4.28 ;
      RECT 63.875 7.12 64.21 7.37 ;
      RECT 63.34 7.12 63.675 7.39 ;
      RECT 61.955 4.08 62.305 4.33 ;
      RECT 61.095 4.08 61.445 4.33 ;
      RECT 60.575 4.08 60.925 4.33 ;
      RECT 57.105 7.3 57.275 10.59 ;
      RECT 56.675 7.3 56.845 9.51 ;
      RECT 56.675 10.08 56.845 10.59 ;
      RECT 53.92 7.305 54.09 8.775 ;
      RECT 53.92 10.085 54.09 10.595 ;
      RECT 52.93 1.865 53.1 2.375 ;
      RECT 52.93 3.685 53.1 5.155 ;
      RECT 52.93 7.305 53.1 8.775 ;
      RECT 52.93 10.085 53.1 10.595 ;
      RECT 51.57 1.87 51.74 5.16 ;
      RECT 51.57 7.3 51.74 10.59 ;
      RECT 51.14 1.87 51.31 2.38 ;
      RECT 51.14 2.95 51.31 5.16 ;
      RECT 51.14 7.3 51.31 9.51 ;
      RECT 51.14 10.08 51.31 10.59 ;
      RECT 47.5 7.12 47.835 7.39 ;
      RECT 47 4.08 47.55 4.28 ;
      RECT 46.655 7.12 46.99 7.37 ;
      RECT 46.12 7.12 46.455 7.39 ;
      RECT 44.735 4.08 45.085 4.33 ;
      RECT 43.875 4.08 44.225 4.33 ;
      RECT 43.355 4.08 43.705 4.33 ;
      RECT 39.885 7.3 40.055 10.59 ;
      RECT 39.455 7.3 39.625 9.51 ;
      RECT 39.455 10.08 39.625 10.59 ;
      RECT 36.7 7.305 36.87 8.775 ;
      RECT 36.7 10.085 36.87 10.595 ;
      RECT 35.71 1.865 35.88 2.375 ;
      RECT 35.71 3.685 35.88 5.155 ;
      RECT 35.71 7.305 35.88 8.775 ;
      RECT 35.71 10.085 35.88 10.595 ;
      RECT 34.35 1.87 34.52 5.16 ;
      RECT 34.35 7.3 34.52 10.59 ;
      RECT 33.92 1.87 34.09 2.38 ;
      RECT 33.92 2.95 34.09 5.16 ;
      RECT 33.92 7.3 34.09 9.51 ;
      RECT 33.92 10.08 34.09 10.59 ;
      RECT 30.28 7.12 30.615 7.39 ;
      RECT 29.78 4.08 30.33 4.28 ;
      RECT 29.435 7.12 29.77 7.37 ;
      RECT 28.9 7.12 29.235 7.39 ;
      RECT 27.515 4.08 27.865 4.33 ;
      RECT 26.655 4.08 27.005 4.33 ;
      RECT 26.135 4.08 26.485 4.33 ;
      RECT 22.665 7.3 22.835 10.59 ;
      RECT 22.235 7.3 22.405 9.51 ;
      RECT 22.235 10.08 22.405 10.59 ;
      RECT 19.48 7.305 19.65 8.775 ;
      RECT 19.48 10.085 19.65 10.595 ;
      RECT 18.49 1.865 18.66 2.375 ;
      RECT 18.49 3.685 18.66 5.155 ;
      RECT 18.49 7.305 18.66 8.775 ;
      RECT 18.49 10.085 18.66 10.595 ;
      RECT 17.13 1.87 17.3 5.16 ;
      RECT 17.13 7.3 17.3 10.59 ;
      RECT 16.7 1.87 16.87 2.38 ;
      RECT 16.7 2.95 16.87 5.16 ;
      RECT 16.7 7.3 16.87 9.51 ;
      RECT 16.7 10.08 16.87 10.59 ;
      RECT 13.06 7.12 13.395 7.39 ;
      RECT 12.56 4.08 13.11 4.28 ;
      RECT 12.215 7.12 12.55 7.37 ;
      RECT 11.68 7.12 12.015 7.39 ;
      RECT 10.295 4.08 10.645 4.33 ;
      RECT 9.435 4.08 9.785 4.33 ;
      RECT 8.915 4.08 9.265 4.33 ;
      RECT 5.445 7.3 5.615 10.59 ;
      RECT 5.015 7.3 5.185 9.51 ;
      RECT 5.015 10.08 5.185 10.59 ;
      RECT 1.605 7.3 1.775 9.51 ;
      RECT 1.605 10.08 1.775 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  ORIGIN -9.9 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r1 ;
  SIZE 84.43 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 28.485 2.21 28.655 2.38 ;
        RECT 28.48 2.205 28.65 2.375 ;
        RECT 28.48 3.685 28.65 3.855 ;
      LAYER li1 ;
        RECT 28.485 2.21 28.655 2.38 ;
        RECT 28.48 1.865 28.65 2.375 ;
        RECT 28.48 3.685 28.65 5.155 ;
      LAYER met1 ;
        RECT 28.42 3.655 28.71 3.885 ;
        RECT 28.42 2.175 28.71 2.405 ;
        RECT 28.48 2.175 28.65 3.885 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 44.81 2.21 44.98 2.38 ;
        RECT 44.805 2.205 44.975 2.375 ;
        RECT 44.805 3.685 44.975 3.855 ;
      LAYER li1 ;
        RECT 44.81 2.21 44.98 2.38 ;
        RECT 44.805 1.865 44.975 2.375 ;
        RECT 44.805 3.685 44.975 5.155 ;
      LAYER met1 ;
        RECT 44.745 3.655 45.035 3.885 ;
        RECT 44.745 2.175 45.035 2.405 ;
        RECT 44.805 2.175 44.975 3.885 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 61.135 2.21 61.305 2.38 ;
        RECT 61.13 2.205 61.3 2.375 ;
        RECT 61.13 3.685 61.3 3.855 ;
      LAYER li1 ;
        RECT 61.135 2.21 61.305 2.38 ;
        RECT 61.13 1.865 61.3 2.375 ;
        RECT 61.13 3.685 61.3 5.155 ;
      LAYER met1 ;
        RECT 61.07 3.655 61.36 3.885 ;
        RECT 61.07 2.175 61.36 2.405 ;
        RECT 61.13 2.175 61.3 3.885 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 77.46 2.21 77.63 2.38 ;
        RECT 77.455 2.205 77.625 2.375 ;
        RECT 77.455 3.685 77.625 3.855 ;
      LAYER li1 ;
        RECT 77.46 2.21 77.63 2.38 ;
        RECT 77.455 1.865 77.625 2.375 ;
        RECT 77.455 3.685 77.625 5.155 ;
      LAYER met1 ;
        RECT 77.395 3.655 77.685 3.885 ;
        RECT 77.395 2.175 77.685 2.405 ;
        RECT 77.455 2.175 77.625 3.885 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 93.785 2.21 93.955 2.38 ;
        RECT 93.78 2.205 93.95 2.375 ;
        RECT 93.78 3.685 93.95 3.855 ;
      LAYER li1 ;
        RECT 93.785 2.21 93.955 2.38 ;
        RECT 93.78 1.865 93.95 2.375 ;
        RECT 93.78 3.685 93.95 5.155 ;
      LAYER met1 ;
        RECT 93.72 3.655 94.01 3.885 ;
        RECT 93.72 2.175 94.01 2.405 ;
        RECT 93.78 2.175 93.95 3.885 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 24.33 2.955 24.5 4.23 ;
        RECT 24.33 8.23 24.5 9.505 ;
        RECT 18.715 8.23 18.885 9.505 ;
      LAYER met2 ;
        RECT 24.255 4 24.595 4.35 ;
        RECT 24.245 8.125 24.585 8.475 ;
        RECT 24.33 4 24.5 8.475 ;
      LAYER met1 ;
        RECT 24.255 4.06 24.73 4.23 ;
        RECT 24.255 4 24.595 4.35 ;
        RECT 18.655 8.23 24.73 8.4 ;
        RECT 24.245 8.125 24.585 8.475 ;
        RECT 18.655 8.2 18.945 8.43 ;
      LAYER via1 ;
        RECT 24.345 8.225 24.495 8.375 ;
        RECT 24.355 4.1 24.505 4.25 ;
      LAYER mcon ;
        RECT 18.715 8.23 18.885 8.4 ;
        RECT 24.33 8.23 24.5 8.4 ;
        RECT 24.33 4.06 24.5 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 40.655 2.955 40.825 4.23 ;
        RECT 40.655 8.23 40.825 9.505 ;
        RECT 35.04 8.23 35.21 9.505 ;
      LAYER met2 ;
        RECT 40.58 4 40.92 4.35 ;
        RECT 40.57 8.125 40.91 8.475 ;
        RECT 40.655 4 40.825 8.475 ;
      LAYER met1 ;
        RECT 40.58 4.06 41.055 4.23 ;
        RECT 40.58 4 40.92 4.35 ;
        RECT 34.98 8.23 41.055 8.4 ;
        RECT 40.57 8.125 40.91 8.475 ;
        RECT 34.98 8.2 35.27 8.43 ;
      LAYER via1 ;
        RECT 40.67 8.225 40.82 8.375 ;
        RECT 40.68 4.1 40.83 4.25 ;
      LAYER mcon ;
        RECT 35.04 8.23 35.21 8.4 ;
        RECT 40.655 8.23 40.825 8.4 ;
        RECT 40.655 4.06 40.825 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 56.98 2.955 57.15 4.23 ;
        RECT 56.98 8.23 57.15 9.505 ;
        RECT 51.365 8.23 51.535 9.505 ;
      LAYER met2 ;
        RECT 56.905 4 57.245 4.35 ;
        RECT 56.895 8.125 57.235 8.475 ;
        RECT 56.98 4 57.15 8.475 ;
      LAYER met1 ;
        RECT 56.905 4.06 57.38 4.23 ;
        RECT 56.905 4 57.245 4.35 ;
        RECT 51.305 8.23 57.38 8.4 ;
        RECT 56.895 8.125 57.235 8.475 ;
        RECT 51.305 8.2 51.595 8.43 ;
      LAYER via1 ;
        RECT 56.995 8.225 57.145 8.375 ;
        RECT 57.005 4.1 57.155 4.25 ;
      LAYER mcon ;
        RECT 51.365 8.23 51.535 8.4 ;
        RECT 56.98 8.23 57.15 8.4 ;
        RECT 56.98 4.06 57.15 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 73.305 2.955 73.475 4.23 ;
        RECT 73.305 8.23 73.475 9.505 ;
        RECT 67.69 8.23 67.86 9.505 ;
      LAYER met2 ;
        RECT 73.23 4 73.57 4.35 ;
        RECT 73.22 8.125 73.56 8.475 ;
        RECT 73.305 4 73.475 8.475 ;
      LAYER met1 ;
        RECT 73.23 4.06 73.705 4.23 ;
        RECT 73.23 4 73.57 4.35 ;
        RECT 67.63 8.23 73.705 8.4 ;
        RECT 73.22 8.125 73.56 8.475 ;
        RECT 67.63 8.2 67.92 8.43 ;
      LAYER via1 ;
        RECT 73.32 8.225 73.47 8.375 ;
        RECT 73.33 4.1 73.48 4.25 ;
      LAYER mcon ;
        RECT 67.69 8.23 67.86 8.4 ;
        RECT 73.305 8.23 73.475 8.4 ;
        RECT 73.305 4.06 73.475 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 89.63 2.955 89.8 4.23 ;
        RECT 89.63 8.23 89.8 9.505 ;
        RECT 84.015 8.23 84.185 9.505 ;
      LAYER met2 ;
        RECT 89.555 4 89.895 4.35 ;
        RECT 89.545 8.125 89.885 8.475 ;
        RECT 89.63 4 89.8 8.475 ;
      LAYER met1 ;
        RECT 89.555 4.06 90.03 4.23 ;
        RECT 89.555 4 89.895 4.35 ;
        RECT 83.955 8.23 90.03 8.4 ;
        RECT 89.545 8.125 89.885 8.475 ;
        RECT 83.955 8.2 84.245 8.43 ;
      LAYER via1 ;
        RECT 89.645 8.225 89.795 8.375 ;
        RECT 89.655 4.1 89.805 4.25 ;
      LAYER mcon ;
        RECT 84.015 8.23 84.185 8.4 ;
        RECT 89.63 8.23 89.8 8.4 ;
        RECT 89.63 4.06 89.8 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 10.135 8.23 10.305 9.505 ;
      LAYER met1 ;
        RECT 10.075 8.23 10.535 8.4 ;
        RECT 10.075 8.2 10.365 8.43 ;
      LAYER mcon ;
        RECT 10.135 8.23 10.305 8.4 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 9.905 5.43 94.325 7.03 ;
        RECT 92.19 5.425 94.17 7.035 ;
        RECT 93.35 4.695 93.52 7.765 ;
        RECT 92.36 4.695 92.53 7.765 ;
        RECT 89.62 4.7 89.79 7.76 ;
        RECT 87.83 4.93 88 7.03 ;
        RECT 86.87 4.93 87.04 7.03 ;
        RECT 84.43 4.93 84.6 7.03 ;
        RECT 84.005 5.43 84.175 7.76 ;
        RECT 83.43 4.93 83.6 7.03 ;
        RECT 82.47 4.93 82.64 7.03 ;
        RECT 80.03 4.93 80.2 7.03 ;
        RECT 75.865 5.425 77.845 7.035 ;
        RECT 77.025 4.695 77.195 7.765 ;
        RECT 76.035 4.695 76.205 7.765 ;
        RECT 73.295 4.7 73.465 7.76 ;
        RECT 71.505 4.93 71.675 7.03 ;
        RECT 70.545 4.93 70.715 7.03 ;
        RECT 68.105 4.93 68.275 7.03 ;
        RECT 67.68 5.43 67.85 7.76 ;
        RECT 67.105 4.93 67.275 7.03 ;
        RECT 66.145 4.93 66.315 7.03 ;
        RECT 63.705 4.93 63.875 7.03 ;
        RECT 59.54 5.425 61.52 7.035 ;
        RECT 60.7 4.695 60.87 7.765 ;
        RECT 59.71 4.695 59.88 7.765 ;
        RECT 56.97 4.7 57.14 7.76 ;
        RECT 55.18 4.93 55.35 7.03 ;
        RECT 54.22 4.93 54.39 7.03 ;
        RECT 51.78 4.93 51.95 7.03 ;
        RECT 51.355 5.43 51.525 7.76 ;
        RECT 50.78 4.93 50.95 7.03 ;
        RECT 49.82 4.93 49.99 7.03 ;
        RECT 47.38 4.93 47.55 7.03 ;
        RECT 43.215 5.425 45.195 7.035 ;
        RECT 44.375 4.695 44.545 7.765 ;
        RECT 43.385 4.695 43.555 7.765 ;
        RECT 40.645 4.7 40.815 7.76 ;
        RECT 38.855 4.93 39.025 7.03 ;
        RECT 37.895 4.93 38.065 7.03 ;
        RECT 35.455 4.93 35.625 7.03 ;
        RECT 35.03 5.43 35.2 7.76 ;
        RECT 34.455 4.93 34.625 7.03 ;
        RECT 33.495 4.93 33.665 7.03 ;
        RECT 31.055 4.93 31.225 7.03 ;
        RECT 26.89 5.425 28.87 7.035 ;
        RECT 28.05 4.695 28.22 7.765 ;
        RECT 27.06 4.695 27.23 7.765 ;
        RECT 24.32 4.7 24.49 7.76 ;
        RECT 22.53 4.93 22.7 7.03 ;
        RECT 21.57 4.93 21.74 7.03 ;
        RECT 19.13 4.93 19.3 7.03 ;
        RECT 18.705 5.43 18.875 7.76 ;
        RECT 18.13 4.93 18.3 7.03 ;
        RECT 17.17 4.93 17.34 7.03 ;
        RECT 14.73 4.93 14.9 7.03 ;
        RECT 11.935 5.43 12.105 10.59 ;
        RECT 10.125 5.43 10.295 7.76 ;
      LAYER met1 ;
        RECT 9.905 5.43 94.325 7.03 ;
        RECT 92.19 5.425 94.17 7.035 ;
        RECT 78.74 5.275 88.4 7.03 ;
        RECT 75.865 5.425 77.845 7.035 ;
        RECT 62.415 5.275 72.075 7.03 ;
        RECT 59.54 5.425 61.52 7.035 ;
        RECT 46.09 5.275 55.75 7.03 ;
        RECT 43.215 5.425 45.195 7.035 ;
        RECT 29.765 5.275 39.425 7.03 ;
        RECT 26.89 5.425 28.87 7.035 ;
        RECT 13.44 5.275 23.1 7.03 ;
        RECT 11.875 8.94 12.165 9.17 ;
        RECT 11.705 8.97 12.165 9.14 ;
      LAYER mcon ;
        RECT 11.935 8.97 12.105 9.14 ;
        RECT 12.245 6.83 12.415 7 ;
        RECT 13.585 5.43 13.755 5.6 ;
        RECT 14.045 5.43 14.215 5.6 ;
        RECT 14.505 5.43 14.675 5.6 ;
        RECT 14.965 5.43 15.135 5.6 ;
        RECT 15.425 5.43 15.595 5.6 ;
        RECT 15.885 5.43 16.055 5.6 ;
        RECT 16.345 5.43 16.515 5.6 ;
        RECT 16.805 5.43 16.975 5.6 ;
        RECT 17.265 5.43 17.435 5.6 ;
        RECT 17.725 5.43 17.895 5.6 ;
        RECT 18.185 5.43 18.355 5.6 ;
        RECT 18.645 5.43 18.815 5.6 ;
        RECT 19.105 5.43 19.275 5.6 ;
        RECT 19.565 5.43 19.735 5.6 ;
        RECT 20.025 5.43 20.195 5.6 ;
        RECT 20.485 5.43 20.655 5.6 ;
        RECT 20.825 6.83 20.995 7 ;
        RECT 20.945 5.43 21.115 5.6 ;
        RECT 21.405 5.43 21.575 5.6 ;
        RECT 21.865 5.43 22.035 5.6 ;
        RECT 22.325 5.43 22.495 5.6 ;
        RECT 22.785 5.43 22.955 5.6 ;
        RECT 26.44 6.83 26.61 7 ;
        RECT 26.44 5.46 26.61 5.63 ;
        RECT 27.14 6.835 27.31 7.005 ;
        RECT 27.14 5.455 27.31 5.625 ;
        RECT 28.13 6.835 28.3 7.005 ;
        RECT 28.13 5.455 28.3 5.625 ;
        RECT 29.91 5.43 30.08 5.6 ;
        RECT 30.37 5.43 30.54 5.6 ;
        RECT 30.83 5.43 31 5.6 ;
        RECT 31.29 5.43 31.46 5.6 ;
        RECT 31.75 5.43 31.92 5.6 ;
        RECT 32.21 5.43 32.38 5.6 ;
        RECT 32.67 5.43 32.84 5.6 ;
        RECT 33.13 5.43 33.3 5.6 ;
        RECT 33.59 5.43 33.76 5.6 ;
        RECT 34.05 5.43 34.22 5.6 ;
        RECT 34.51 5.43 34.68 5.6 ;
        RECT 34.97 5.43 35.14 5.6 ;
        RECT 35.43 5.43 35.6 5.6 ;
        RECT 35.89 5.43 36.06 5.6 ;
        RECT 36.35 5.43 36.52 5.6 ;
        RECT 36.81 5.43 36.98 5.6 ;
        RECT 37.15 6.83 37.32 7 ;
        RECT 37.27 5.43 37.44 5.6 ;
        RECT 37.73 5.43 37.9 5.6 ;
        RECT 38.19 5.43 38.36 5.6 ;
        RECT 38.65 5.43 38.82 5.6 ;
        RECT 39.11 5.43 39.28 5.6 ;
        RECT 42.765 6.83 42.935 7 ;
        RECT 42.765 5.46 42.935 5.63 ;
        RECT 43.465 6.835 43.635 7.005 ;
        RECT 43.465 5.455 43.635 5.625 ;
        RECT 44.455 6.835 44.625 7.005 ;
        RECT 44.455 5.455 44.625 5.625 ;
        RECT 46.235 5.43 46.405 5.6 ;
        RECT 46.695 5.43 46.865 5.6 ;
        RECT 47.155 5.43 47.325 5.6 ;
        RECT 47.615 5.43 47.785 5.6 ;
        RECT 48.075 5.43 48.245 5.6 ;
        RECT 48.535 5.43 48.705 5.6 ;
        RECT 48.995 5.43 49.165 5.6 ;
        RECT 49.455 5.43 49.625 5.6 ;
        RECT 49.915 5.43 50.085 5.6 ;
        RECT 50.375 5.43 50.545 5.6 ;
        RECT 50.835 5.43 51.005 5.6 ;
        RECT 51.295 5.43 51.465 5.6 ;
        RECT 51.755 5.43 51.925 5.6 ;
        RECT 52.215 5.43 52.385 5.6 ;
        RECT 52.675 5.43 52.845 5.6 ;
        RECT 53.135 5.43 53.305 5.6 ;
        RECT 53.475 6.83 53.645 7 ;
        RECT 53.595 5.43 53.765 5.6 ;
        RECT 54.055 5.43 54.225 5.6 ;
        RECT 54.515 5.43 54.685 5.6 ;
        RECT 54.975 5.43 55.145 5.6 ;
        RECT 55.435 5.43 55.605 5.6 ;
        RECT 59.09 6.83 59.26 7 ;
        RECT 59.09 5.46 59.26 5.63 ;
        RECT 59.79 6.835 59.96 7.005 ;
        RECT 59.79 5.455 59.96 5.625 ;
        RECT 60.78 6.835 60.95 7.005 ;
        RECT 60.78 5.455 60.95 5.625 ;
        RECT 62.56 5.43 62.73 5.6 ;
        RECT 63.02 5.43 63.19 5.6 ;
        RECT 63.48 5.43 63.65 5.6 ;
        RECT 63.94 5.43 64.11 5.6 ;
        RECT 64.4 5.43 64.57 5.6 ;
        RECT 64.86 5.43 65.03 5.6 ;
        RECT 65.32 5.43 65.49 5.6 ;
        RECT 65.78 5.43 65.95 5.6 ;
        RECT 66.24 5.43 66.41 5.6 ;
        RECT 66.7 5.43 66.87 5.6 ;
        RECT 67.16 5.43 67.33 5.6 ;
        RECT 67.62 5.43 67.79 5.6 ;
        RECT 68.08 5.43 68.25 5.6 ;
        RECT 68.54 5.43 68.71 5.6 ;
        RECT 69 5.43 69.17 5.6 ;
        RECT 69.46 5.43 69.63 5.6 ;
        RECT 69.8 6.83 69.97 7 ;
        RECT 69.92 5.43 70.09 5.6 ;
        RECT 70.38 5.43 70.55 5.6 ;
        RECT 70.84 5.43 71.01 5.6 ;
        RECT 71.3 5.43 71.47 5.6 ;
        RECT 71.76 5.43 71.93 5.6 ;
        RECT 75.415 6.83 75.585 7 ;
        RECT 75.415 5.46 75.585 5.63 ;
        RECT 76.115 6.835 76.285 7.005 ;
        RECT 76.115 5.455 76.285 5.625 ;
        RECT 77.105 6.835 77.275 7.005 ;
        RECT 77.105 5.455 77.275 5.625 ;
        RECT 78.885 5.43 79.055 5.6 ;
        RECT 79.345 5.43 79.515 5.6 ;
        RECT 79.805 5.43 79.975 5.6 ;
        RECT 80.265 5.43 80.435 5.6 ;
        RECT 80.725 5.43 80.895 5.6 ;
        RECT 81.185 5.43 81.355 5.6 ;
        RECT 81.645 5.43 81.815 5.6 ;
        RECT 82.105 5.43 82.275 5.6 ;
        RECT 82.565 5.43 82.735 5.6 ;
        RECT 83.025 5.43 83.195 5.6 ;
        RECT 83.485 5.43 83.655 5.6 ;
        RECT 83.945 5.43 84.115 5.6 ;
        RECT 84.405 5.43 84.575 5.6 ;
        RECT 84.865 5.43 85.035 5.6 ;
        RECT 85.325 5.43 85.495 5.6 ;
        RECT 85.785 5.43 85.955 5.6 ;
        RECT 86.125 6.83 86.295 7 ;
        RECT 86.245 5.43 86.415 5.6 ;
        RECT 86.705 5.43 86.875 5.6 ;
        RECT 87.165 5.43 87.335 5.6 ;
        RECT 87.625 5.43 87.795 5.6 ;
        RECT 88.085 5.43 88.255 5.6 ;
        RECT 91.74 6.83 91.91 7 ;
        RECT 91.74 5.46 91.91 5.63 ;
        RECT 92.44 6.835 92.61 7.005 ;
        RECT 92.44 5.455 92.61 5.625 ;
        RECT 93.43 6.835 93.6 7.005 ;
        RECT 93.43 5.455 93.6 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 87.63 4.27 87.96 5 ;
        RECT 71.305 4.27 71.635 5 ;
        RECT 54.98 4.27 55.31 5 ;
        RECT 38.655 4.27 38.985 5 ;
        RECT 22.33 4.27 22.66 5 ;
      LAYER li1 ;
        RECT 9.95 10.86 94.33 12.46 ;
        RECT 93.35 10.235 93.52 12.46 ;
        RECT 92.36 10.235 92.53 12.46 ;
        RECT 89.62 10.23 89.79 12.46 ;
        RECT 84.005 10.23 84.175 12.46 ;
        RECT 77.025 10.235 77.195 12.46 ;
        RECT 76.035 10.235 76.205 12.46 ;
        RECT 73.295 10.23 73.465 12.46 ;
        RECT 67.68 10.23 67.85 12.46 ;
        RECT 60.7 10.235 60.87 12.46 ;
        RECT 59.71 10.235 59.88 12.46 ;
        RECT 56.97 10.23 57.14 12.46 ;
        RECT 51.355 10.23 51.525 12.46 ;
        RECT 44.375 10.235 44.545 12.46 ;
        RECT 43.385 10.235 43.555 12.46 ;
        RECT 40.645 10.23 40.815 12.46 ;
        RECT 35.03 10.23 35.2 12.46 ;
        RECT 28.05 10.235 28.22 12.46 ;
        RECT 27.06 10.235 27.23 12.46 ;
        RECT 24.32 10.23 24.49 12.46 ;
        RECT 18.705 10.23 18.875 12.46 ;
        RECT 10.125 10.23 10.295 12.46 ;
        RECT 9.9 0 94.325 1.6 ;
        RECT 93.35 0 93.52 2.225 ;
        RECT 92.36 0 92.53 2.225 ;
        RECT 89.62 0 89.79 2.23 ;
        RECT 78.74 0 88.555 2.88 ;
        RECT 86.87 0 87.04 3.38 ;
        RECT 84.91 0 85.08 3.38 ;
        RECT 84.84 0 85.08 2.89 ;
        RECT 83.29 0 83.485 2.89 ;
        RECT 82.47 0 82.64 3.38 ;
        RECT 81.51 0 81.68 3.38 ;
        RECT 81.165 0 81.36 2.89 ;
        RECT 80.99 0 81.16 3.38 ;
        RECT 80.03 0 80.2 3.38 ;
        RECT 79.07 0 79.24 3.38 ;
        RECT 78.865 0 79.06 2.89 ;
        RECT 77.025 0 77.195 2.225 ;
        RECT 76.035 0 76.205 2.225 ;
        RECT 73.295 0 73.465 2.23 ;
        RECT 62.415 0 72.23 2.88 ;
        RECT 70.545 0 70.715 3.38 ;
        RECT 68.585 0 68.755 3.38 ;
        RECT 68.515 0 68.755 2.89 ;
        RECT 66.965 0 67.16 2.89 ;
        RECT 66.145 0 66.315 3.38 ;
        RECT 65.185 0 65.355 3.38 ;
        RECT 64.84 0 65.035 2.89 ;
        RECT 64.665 0 64.835 3.38 ;
        RECT 63.705 0 63.875 3.38 ;
        RECT 62.745 0 62.915 3.38 ;
        RECT 62.54 0 62.735 2.89 ;
        RECT 60.7 0 60.87 2.225 ;
        RECT 59.71 0 59.88 2.225 ;
        RECT 56.97 0 57.14 2.23 ;
        RECT 46.09 0 55.905 2.88 ;
        RECT 54.22 0 54.39 3.38 ;
        RECT 52.26 0 52.43 3.38 ;
        RECT 52.19 0 52.43 2.89 ;
        RECT 50.64 0 50.835 2.89 ;
        RECT 49.82 0 49.99 3.38 ;
        RECT 48.86 0 49.03 3.38 ;
        RECT 48.515 0 48.71 2.89 ;
        RECT 48.34 0 48.51 3.38 ;
        RECT 47.38 0 47.55 3.38 ;
        RECT 46.42 0 46.59 3.38 ;
        RECT 46.215 0 46.41 2.89 ;
        RECT 44.375 0 44.545 2.225 ;
        RECT 43.385 0 43.555 2.225 ;
        RECT 40.645 0 40.815 2.23 ;
        RECT 29.765 0 39.58 2.88 ;
        RECT 37.895 0 38.065 3.38 ;
        RECT 35.935 0 36.105 3.38 ;
        RECT 35.865 0 36.105 2.89 ;
        RECT 34.315 0 34.51 2.89 ;
        RECT 33.495 0 33.665 3.38 ;
        RECT 32.535 0 32.705 3.38 ;
        RECT 32.19 0 32.385 2.89 ;
        RECT 32.015 0 32.185 3.38 ;
        RECT 31.055 0 31.225 3.38 ;
        RECT 30.095 0 30.265 3.38 ;
        RECT 29.89 0 30.085 2.89 ;
        RECT 28.05 0 28.22 2.225 ;
        RECT 27.06 0 27.23 2.225 ;
        RECT 24.32 0 24.49 2.23 ;
        RECT 13.44 0 23.255 2.88 ;
        RECT 21.57 0 21.74 3.38 ;
        RECT 19.61 0 19.78 3.38 ;
        RECT 19.54 0 19.78 2.89 ;
        RECT 17.99 0 18.185 2.89 ;
        RECT 17.17 0 17.34 3.38 ;
        RECT 16.21 0 16.38 3.38 ;
        RECT 15.865 0 16.06 2.89 ;
        RECT 15.69 0 15.86 3.38 ;
        RECT 14.73 0 14.9 3.38 ;
        RECT 13.77 0 13.94 3.38 ;
        RECT 13.565 0 13.76 2.89 ;
        RECT 87.83 3.87 88 4.24 ;
        RECT 87.51 3.87 88 4.04 ;
        RECT 85.87 3.87 86.04 4.24 ;
        RECT 85.55 3.87 86.04 4.04 ;
        RECT 85.01 8.36 85.18 10.31 ;
        RECT 84.955 10.14 85.125 10.59 ;
        RECT 84.955 7.3 85.125 8.53 ;
        RECT 71.505 3.87 71.675 4.24 ;
        RECT 71.185 3.87 71.675 4.04 ;
        RECT 69.545 3.87 69.715 4.24 ;
        RECT 69.225 3.87 69.715 4.04 ;
        RECT 68.685 8.36 68.855 10.31 ;
        RECT 68.63 10.14 68.8 10.59 ;
        RECT 68.63 7.3 68.8 8.53 ;
        RECT 55.18 3.87 55.35 4.24 ;
        RECT 54.86 3.87 55.35 4.04 ;
        RECT 53.22 3.87 53.39 4.24 ;
        RECT 52.9 3.87 53.39 4.04 ;
        RECT 52.36 8.36 52.53 10.31 ;
        RECT 52.305 10.14 52.475 10.59 ;
        RECT 52.305 7.3 52.475 8.53 ;
        RECT 38.855 3.87 39.025 4.24 ;
        RECT 38.535 3.87 39.025 4.04 ;
        RECT 36.895 3.87 37.065 4.24 ;
        RECT 36.575 3.87 37.065 4.04 ;
        RECT 36.035 8.36 36.205 10.31 ;
        RECT 35.98 10.14 36.15 10.59 ;
        RECT 35.98 7.3 36.15 8.53 ;
        RECT 22.53 3.87 22.7 4.24 ;
        RECT 22.21 3.87 22.7 4.04 ;
        RECT 20.57 3.87 20.74 4.24 ;
        RECT 20.25 3.87 20.74 4.04 ;
        RECT 19.71 8.36 19.88 10.31 ;
        RECT 19.655 10.14 19.825 10.59 ;
        RECT 19.655 7.3 19.825 8.53 ;
      LAYER met2 ;
        RECT 87.655 4.25 87.935 4.62 ;
        RECT 87.665 3.995 87.925 4.62 ;
        RECT 71.33 4.25 71.61 4.62 ;
        RECT 71.34 3.995 71.6 4.62 ;
        RECT 55.005 4.25 55.285 4.62 ;
        RECT 55.015 3.995 55.275 4.62 ;
        RECT 38.68 4.25 38.96 4.62 ;
        RECT 38.69 3.995 38.95 4.62 ;
        RECT 22.355 4.25 22.635 4.62 ;
        RECT 22.365 3.995 22.625 4.62 ;
      LAYER met1 ;
        RECT 9.95 10.86 94.33 12.46 ;
        RECT 84.95 8.57 85.24 8.8 ;
        RECT 84.575 8.6 85.24 8.77 ;
        RECT 84.575 8.6 84.75 12.46 ;
        RECT 68.625 8.57 68.915 8.8 ;
        RECT 68.25 8.6 68.915 8.77 ;
        RECT 68.25 8.6 68.425 12.46 ;
        RECT 52.3 8.57 52.59 8.8 ;
        RECT 51.925 8.6 52.59 8.77 ;
        RECT 51.925 8.6 52.1 12.46 ;
        RECT 35.975 8.57 36.265 8.8 ;
        RECT 35.6 8.6 36.265 8.77 ;
        RECT 35.6 8.6 35.775 12.46 ;
        RECT 19.65 8.57 19.94 8.8 ;
        RECT 19.275 8.6 19.94 8.77 ;
        RECT 19.275 8.6 19.45 12.46 ;
        RECT 9.9 0 94.325 1.6 ;
        RECT 88.37 0 88.555 4.24 ;
        RECT 87.605 4.085 88.555 4.24 ;
        RECT 87.635 4.055 88.555 4.24 ;
        RECT 78.74 0 88.555 3.035 ;
        RECT 87.635 4.04 88.06 4.27 ;
        RECT 87.635 4.025 87.955 4.285 ;
        RECT 86.145 4.225 87.91 4.35 ;
        RECT 86.145 4.225 87.745 4.365 ;
        RECT 85.81 4.085 86.285 4.27 ;
        RECT 85.81 4.04 86.1 4.27 ;
        RECT 72.045 0 72.23 4.24 ;
        RECT 71.28 4.085 72.23 4.24 ;
        RECT 71.31 4.055 72.23 4.24 ;
        RECT 62.415 0 72.23 3.035 ;
        RECT 71.31 4.04 71.735 4.27 ;
        RECT 71.31 4.025 71.63 4.285 ;
        RECT 69.82 4.225 71.585 4.35 ;
        RECT 69.82 4.225 71.42 4.365 ;
        RECT 69.485 4.085 69.96 4.27 ;
        RECT 69.485 4.04 69.775 4.27 ;
        RECT 55.72 0 55.905 4.24 ;
        RECT 54.955 4.085 55.905 4.24 ;
        RECT 54.985 4.055 55.905 4.24 ;
        RECT 46.09 0 55.905 3.035 ;
        RECT 54.985 4.04 55.41 4.27 ;
        RECT 54.985 4.025 55.305 4.285 ;
        RECT 53.495 4.225 55.26 4.35 ;
        RECT 53.495 4.225 55.095 4.365 ;
        RECT 53.16 4.085 53.635 4.27 ;
        RECT 53.16 4.04 53.45 4.27 ;
        RECT 39.395 0 39.58 4.24 ;
        RECT 38.63 4.085 39.58 4.24 ;
        RECT 38.66 4.055 39.58 4.24 ;
        RECT 29.765 0 39.58 3.035 ;
        RECT 38.66 4.04 39.085 4.27 ;
        RECT 38.66 4.025 38.98 4.285 ;
        RECT 37.17 4.225 38.935 4.35 ;
        RECT 37.17 4.225 38.77 4.365 ;
        RECT 36.835 4.085 37.31 4.27 ;
        RECT 36.835 4.04 37.125 4.27 ;
        RECT 23.07 0 23.255 4.24 ;
        RECT 22.305 4.085 23.255 4.24 ;
        RECT 22.335 4.055 23.255 4.24 ;
        RECT 13.44 0 23.255 3.035 ;
        RECT 22.335 4.04 22.76 4.27 ;
        RECT 22.335 4.025 22.655 4.285 ;
        RECT 20.845 4.225 22.61 4.35 ;
        RECT 20.845 4.225 22.445 4.365 ;
        RECT 20.51 4.085 20.985 4.27 ;
        RECT 20.51 4.04 20.8 4.27 ;
      LAYER via2 ;
        RECT 22.395 4.335 22.595 4.535 ;
        RECT 38.72 4.335 38.92 4.535 ;
        RECT 55.045 4.335 55.245 4.535 ;
        RECT 71.37 4.335 71.57 4.535 ;
        RECT 87.695 4.335 87.895 4.535 ;
      LAYER via1 ;
        RECT 22.42 4.08 22.57 4.23 ;
        RECT 38.745 4.08 38.895 4.23 ;
        RECT 55.07 4.08 55.22 4.23 ;
        RECT 71.395 4.08 71.545 4.23 ;
        RECT 87.72 4.08 87.87 4.23 ;
      LAYER mcon ;
        RECT 10.205 10.89 10.375 11.06 ;
        RECT 10.885 10.89 11.055 11.06 ;
        RECT 11.565 10.89 11.735 11.06 ;
        RECT 12.245 10.89 12.415 11.06 ;
        RECT 13.585 2.71 13.755 2.88 ;
        RECT 14.045 2.71 14.215 2.88 ;
        RECT 14.505 2.71 14.675 2.88 ;
        RECT 14.965 2.71 15.135 2.88 ;
        RECT 15.425 2.71 15.595 2.88 ;
        RECT 15.885 2.71 16.055 2.88 ;
        RECT 16.345 2.71 16.515 2.88 ;
        RECT 16.805 2.71 16.975 2.88 ;
        RECT 17.265 2.71 17.435 2.88 ;
        RECT 17.725 2.71 17.895 2.88 ;
        RECT 18.185 2.71 18.355 2.88 ;
        RECT 18.645 2.71 18.815 2.88 ;
        RECT 18.785 10.89 18.955 11.06 ;
        RECT 19.105 2.71 19.275 2.88 ;
        RECT 19.465 10.89 19.635 11.06 ;
        RECT 19.565 2.71 19.735 2.88 ;
        RECT 19.71 8.6 19.88 8.77 ;
        RECT 20.025 2.71 20.195 2.88 ;
        RECT 20.145 10.89 20.315 11.06 ;
        RECT 20.485 2.71 20.655 2.88 ;
        RECT 20.57 4.07 20.74 4.24 ;
        RECT 20.825 10.89 20.995 11.06 ;
        RECT 20.945 2.71 21.115 2.88 ;
        RECT 21.405 2.71 21.575 2.88 ;
        RECT 21.865 2.71 22.035 2.88 ;
        RECT 22.325 2.71 22.495 2.88 ;
        RECT 22.53 4.07 22.7 4.24 ;
        RECT 22.785 2.71 22.955 2.88 ;
        RECT 24.4 10.89 24.57 11.06 ;
        RECT 24.4 1.4 24.57 1.57 ;
        RECT 25.08 10.89 25.25 11.06 ;
        RECT 25.08 1.4 25.25 1.57 ;
        RECT 25.76 10.89 25.93 11.06 ;
        RECT 25.76 1.4 25.93 1.57 ;
        RECT 26.44 10.89 26.61 11.06 ;
        RECT 26.44 1.4 26.61 1.57 ;
        RECT 27.14 10.895 27.31 11.065 ;
        RECT 27.14 1.395 27.31 1.565 ;
        RECT 28.13 10.895 28.3 11.065 ;
        RECT 28.13 1.395 28.3 1.565 ;
        RECT 29.91 2.71 30.08 2.88 ;
        RECT 30.37 2.71 30.54 2.88 ;
        RECT 30.83 2.71 31 2.88 ;
        RECT 31.29 2.71 31.46 2.88 ;
        RECT 31.75 2.71 31.92 2.88 ;
        RECT 32.21 2.71 32.38 2.88 ;
        RECT 32.67 2.71 32.84 2.88 ;
        RECT 33.13 2.71 33.3 2.88 ;
        RECT 33.59 2.71 33.76 2.88 ;
        RECT 34.05 2.71 34.22 2.88 ;
        RECT 34.51 2.71 34.68 2.88 ;
        RECT 34.97 2.71 35.14 2.88 ;
        RECT 35.11 10.89 35.28 11.06 ;
        RECT 35.43 2.71 35.6 2.88 ;
        RECT 35.79 10.89 35.96 11.06 ;
        RECT 35.89 2.71 36.06 2.88 ;
        RECT 36.035 8.6 36.205 8.77 ;
        RECT 36.35 2.71 36.52 2.88 ;
        RECT 36.47 10.89 36.64 11.06 ;
        RECT 36.81 2.71 36.98 2.88 ;
        RECT 36.895 4.07 37.065 4.24 ;
        RECT 37.15 10.89 37.32 11.06 ;
        RECT 37.27 2.71 37.44 2.88 ;
        RECT 37.73 2.71 37.9 2.88 ;
        RECT 38.19 2.71 38.36 2.88 ;
        RECT 38.65 2.71 38.82 2.88 ;
        RECT 38.855 4.07 39.025 4.24 ;
        RECT 39.11 2.71 39.28 2.88 ;
        RECT 40.725 10.89 40.895 11.06 ;
        RECT 40.725 1.4 40.895 1.57 ;
        RECT 41.405 10.89 41.575 11.06 ;
        RECT 41.405 1.4 41.575 1.57 ;
        RECT 42.085 10.89 42.255 11.06 ;
        RECT 42.085 1.4 42.255 1.57 ;
        RECT 42.765 10.89 42.935 11.06 ;
        RECT 42.765 1.4 42.935 1.57 ;
        RECT 43.465 10.895 43.635 11.065 ;
        RECT 43.465 1.395 43.635 1.565 ;
        RECT 44.455 10.895 44.625 11.065 ;
        RECT 44.455 1.395 44.625 1.565 ;
        RECT 46.235 2.71 46.405 2.88 ;
        RECT 46.695 2.71 46.865 2.88 ;
        RECT 47.155 2.71 47.325 2.88 ;
        RECT 47.615 2.71 47.785 2.88 ;
        RECT 48.075 2.71 48.245 2.88 ;
        RECT 48.535 2.71 48.705 2.88 ;
        RECT 48.995 2.71 49.165 2.88 ;
        RECT 49.455 2.71 49.625 2.88 ;
        RECT 49.915 2.71 50.085 2.88 ;
        RECT 50.375 2.71 50.545 2.88 ;
        RECT 50.835 2.71 51.005 2.88 ;
        RECT 51.295 2.71 51.465 2.88 ;
        RECT 51.435 10.89 51.605 11.06 ;
        RECT 51.755 2.71 51.925 2.88 ;
        RECT 52.115 10.89 52.285 11.06 ;
        RECT 52.215 2.71 52.385 2.88 ;
        RECT 52.36 8.6 52.53 8.77 ;
        RECT 52.675 2.71 52.845 2.88 ;
        RECT 52.795 10.89 52.965 11.06 ;
        RECT 53.135 2.71 53.305 2.88 ;
        RECT 53.22 4.07 53.39 4.24 ;
        RECT 53.475 10.89 53.645 11.06 ;
        RECT 53.595 2.71 53.765 2.88 ;
        RECT 54.055 2.71 54.225 2.88 ;
        RECT 54.515 2.71 54.685 2.88 ;
        RECT 54.975 2.71 55.145 2.88 ;
        RECT 55.18 4.07 55.35 4.24 ;
        RECT 55.435 2.71 55.605 2.88 ;
        RECT 57.05 10.89 57.22 11.06 ;
        RECT 57.05 1.4 57.22 1.57 ;
        RECT 57.73 10.89 57.9 11.06 ;
        RECT 57.73 1.4 57.9 1.57 ;
        RECT 58.41 10.89 58.58 11.06 ;
        RECT 58.41 1.4 58.58 1.57 ;
        RECT 59.09 10.89 59.26 11.06 ;
        RECT 59.09 1.4 59.26 1.57 ;
        RECT 59.79 10.895 59.96 11.065 ;
        RECT 59.79 1.395 59.96 1.565 ;
        RECT 60.78 10.895 60.95 11.065 ;
        RECT 60.78 1.395 60.95 1.565 ;
        RECT 62.56 2.71 62.73 2.88 ;
        RECT 63.02 2.71 63.19 2.88 ;
        RECT 63.48 2.71 63.65 2.88 ;
        RECT 63.94 2.71 64.11 2.88 ;
        RECT 64.4 2.71 64.57 2.88 ;
        RECT 64.86 2.71 65.03 2.88 ;
        RECT 65.32 2.71 65.49 2.88 ;
        RECT 65.78 2.71 65.95 2.88 ;
        RECT 66.24 2.71 66.41 2.88 ;
        RECT 66.7 2.71 66.87 2.88 ;
        RECT 67.16 2.71 67.33 2.88 ;
        RECT 67.62 2.71 67.79 2.88 ;
        RECT 67.76 10.89 67.93 11.06 ;
        RECT 68.08 2.71 68.25 2.88 ;
        RECT 68.44 10.89 68.61 11.06 ;
        RECT 68.54 2.71 68.71 2.88 ;
        RECT 68.685 8.6 68.855 8.77 ;
        RECT 69 2.71 69.17 2.88 ;
        RECT 69.12 10.89 69.29 11.06 ;
        RECT 69.46 2.71 69.63 2.88 ;
        RECT 69.545 4.07 69.715 4.24 ;
        RECT 69.8 10.89 69.97 11.06 ;
        RECT 69.92 2.71 70.09 2.88 ;
        RECT 70.38 2.71 70.55 2.88 ;
        RECT 70.84 2.71 71.01 2.88 ;
        RECT 71.3 2.71 71.47 2.88 ;
        RECT 71.505 4.07 71.675 4.24 ;
        RECT 71.76 2.71 71.93 2.88 ;
        RECT 73.375 10.89 73.545 11.06 ;
        RECT 73.375 1.4 73.545 1.57 ;
        RECT 74.055 10.89 74.225 11.06 ;
        RECT 74.055 1.4 74.225 1.57 ;
        RECT 74.735 10.89 74.905 11.06 ;
        RECT 74.735 1.4 74.905 1.57 ;
        RECT 75.415 10.89 75.585 11.06 ;
        RECT 75.415 1.4 75.585 1.57 ;
        RECT 76.115 10.895 76.285 11.065 ;
        RECT 76.115 1.395 76.285 1.565 ;
        RECT 77.105 10.895 77.275 11.065 ;
        RECT 77.105 1.395 77.275 1.565 ;
        RECT 78.885 2.71 79.055 2.88 ;
        RECT 79.345 2.71 79.515 2.88 ;
        RECT 79.805 2.71 79.975 2.88 ;
        RECT 80.265 2.71 80.435 2.88 ;
        RECT 80.725 2.71 80.895 2.88 ;
        RECT 81.185 2.71 81.355 2.88 ;
        RECT 81.645 2.71 81.815 2.88 ;
        RECT 82.105 2.71 82.275 2.88 ;
        RECT 82.565 2.71 82.735 2.88 ;
        RECT 83.025 2.71 83.195 2.88 ;
        RECT 83.485 2.71 83.655 2.88 ;
        RECT 83.945 2.71 84.115 2.88 ;
        RECT 84.085 10.89 84.255 11.06 ;
        RECT 84.405 2.71 84.575 2.88 ;
        RECT 84.765 10.89 84.935 11.06 ;
        RECT 84.865 2.71 85.035 2.88 ;
        RECT 85.01 8.6 85.18 8.77 ;
        RECT 85.325 2.71 85.495 2.88 ;
        RECT 85.445 10.89 85.615 11.06 ;
        RECT 85.785 2.71 85.955 2.88 ;
        RECT 85.87 4.07 86.04 4.24 ;
        RECT 86.125 10.89 86.295 11.06 ;
        RECT 86.245 2.71 86.415 2.88 ;
        RECT 86.705 2.71 86.875 2.88 ;
        RECT 87.165 2.71 87.335 2.88 ;
        RECT 87.625 2.71 87.795 2.88 ;
        RECT 87.83 4.07 88 4.24 ;
        RECT 88.085 2.71 88.255 2.88 ;
        RECT 89.7 10.89 89.87 11.06 ;
        RECT 89.7 1.4 89.87 1.57 ;
        RECT 90.38 10.89 90.55 11.06 ;
        RECT 90.38 1.4 90.55 1.57 ;
        RECT 91.06 10.89 91.23 11.06 ;
        RECT 91.06 1.4 91.23 1.57 ;
        RECT 91.74 10.89 91.91 11.06 ;
        RECT 91.74 1.4 91.91 1.57 ;
        RECT 92.44 10.895 92.61 11.065 ;
        RECT 92.44 1.395 92.61 1.565 ;
        RECT 93.43 10.895 93.6 11.065 ;
        RECT 93.43 1.395 93.6 1.565 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 85.305 9.34 85.675 9.71 ;
      RECT 85.305 9.375 87.29 9.675 ;
      RECT 86.99 3.575 87.29 9.675 ;
      RECT 83.99 3.31 84.32 4.04 ;
      RECT 83.11 3.31 83.44 4.04 ;
      RECT 86.19 3.575 87.48 3.875 ;
      RECT 87.15 3.145 87.48 3.875 ;
      RECT 83.11 3.575 85.25 3.875 ;
      RECT 84.95 3.26 85.25 3.875 ;
      RECT 86.19 3.275 86.495 3.875 ;
      RECT 84.95 3.26 86.31 3.57 ;
      RECT 83.61 4.83 83.94 5.16 ;
      RECT 82.405 4.845 83.94 5.145 ;
      RECT 82.405 3.725 82.705 5.145 ;
      RECT 82.15 3.71 82.48 4.04 ;
      RECT 68.98 9.34 69.35 9.71 ;
      RECT 68.98 9.375 70.965 9.675 ;
      RECT 70.665 3.575 70.965 9.675 ;
      RECT 67.665 3.31 67.995 4.04 ;
      RECT 66.785 3.31 67.115 4.04 ;
      RECT 69.865 3.575 71.155 3.875 ;
      RECT 70.825 3.145 71.155 3.875 ;
      RECT 66.785 3.575 68.925 3.875 ;
      RECT 68.625 3.26 68.925 3.875 ;
      RECT 69.865 3.275 70.17 3.875 ;
      RECT 68.625 3.26 69.985 3.57 ;
      RECT 67.285 4.83 67.615 5.16 ;
      RECT 66.08 4.845 67.615 5.145 ;
      RECT 66.08 3.725 66.38 5.145 ;
      RECT 65.825 3.71 66.155 4.04 ;
      RECT 52.655 9.34 53.025 9.71 ;
      RECT 52.655 9.375 54.64 9.675 ;
      RECT 54.34 3.575 54.64 9.675 ;
      RECT 51.34 3.31 51.67 4.04 ;
      RECT 50.46 3.31 50.79 4.04 ;
      RECT 53.54 3.575 54.83 3.875 ;
      RECT 54.5 3.145 54.83 3.875 ;
      RECT 50.46 3.575 52.6 3.875 ;
      RECT 52.3 3.26 52.6 3.875 ;
      RECT 53.54 3.275 53.845 3.875 ;
      RECT 52.3 3.26 53.66 3.57 ;
      RECT 50.96 4.83 51.29 5.16 ;
      RECT 49.755 4.845 51.29 5.145 ;
      RECT 49.755 3.725 50.055 5.145 ;
      RECT 49.5 3.71 49.83 4.04 ;
      RECT 36.33 9.34 36.7 9.71 ;
      RECT 36.33 9.375 38.315 9.675 ;
      RECT 38.015 3.575 38.315 9.675 ;
      RECT 35.015 3.31 35.345 4.04 ;
      RECT 34.135 3.31 34.465 4.04 ;
      RECT 37.215 3.575 38.505 3.875 ;
      RECT 38.175 3.145 38.505 3.875 ;
      RECT 34.135 3.575 36.275 3.875 ;
      RECT 35.975 3.26 36.275 3.875 ;
      RECT 37.215 3.275 37.52 3.875 ;
      RECT 35.975 3.26 37.335 3.57 ;
      RECT 34.635 4.83 34.965 5.16 ;
      RECT 33.43 4.845 34.965 5.145 ;
      RECT 33.43 3.725 33.73 5.145 ;
      RECT 33.175 3.71 33.505 4.04 ;
      RECT 20.005 9.34 20.375 9.71 ;
      RECT 20.005 9.375 21.99 9.675 ;
      RECT 21.69 3.575 21.99 9.675 ;
      RECT 18.69 3.31 19.02 4.04 ;
      RECT 17.81 3.31 18.14 4.04 ;
      RECT 20.89 3.575 22.18 3.875 ;
      RECT 21.85 3.145 22.18 3.875 ;
      RECT 17.81 3.575 19.95 3.875 ;
      RECT 19.65 3.26 19.95 3.875 ;
      RECT 20.89 3.275 21.195 3.875 ;
      RECT 19.65 3.26 21.01 3.57 ;
      RECT 18.31 4.83 18.64 5.16 ;
      RECT 17.105 4.845 18.64 5.145 ;
      RECT 17.105 3.725 17.405 5.145 ;
      RECT 16.85 3.71 17.18 4.04 ;
      RECT 85.55 3.87 85.88 4.6 ;
      RECT 81.43 3.71 81.76 4.44 ;
      RECT 80.43 3.15 80.76 3.88 ;
      RECT 78.99 3.87 79.32 4.6 ;
      RECT 69.225 3.87 69.555 4.6 ;
      RECT 65.105 3.71 65.435 4.44 ;
      RECT 64.105 3.15 64.435 3.88 ;
      RECT 62.665 3.87 62.995 4.6 ;
      RECT 52.9 3.87 53.23 4.6 ;
      RECT 48.78 3.71 49.11 4.44 ;
      RECT 47.78 3.15 48.11 3.88 ;
      RECT 46.34 3.87 46.67 4.6 ;
      RECT 36.575 3.87 36.905 4.6 ;
      RECT 32.455 3.71 32.785 4.44 ;
      RECT 31.455 3.15 31.785 3.88 ;
      RECT 30.015 3.87 30.345 4.6 ;
      RECT 20.25 3.87 20.58 4.6 ;
      RECT 16.13 3.71 16.46 4.44 ;
      RECT 15.13 3.15 15.46 3.88 ;
      RECT 13.69 3.87 14.02 4.6 ;
    LAYER via2 ;
      RECT 87.215 3.61 87.415 3.81 ;
      RECT 85.615 4.335 85.815 4.535 ;
      RECT 85.39 9.425 85.59 9.625 ;
      RECT 84.055 3.775 84.255 3.975 ;
      RECT 83.675 4.895 83.875 5.095 ;
      RECT 83.175 3.775 83.375 3.975 ;
      RECT 82.215 3.775 82.415 3.975 ;
      RECT 81.495 3.775 81.695 3.975 ;
      RECT 80.495 3.215 80.695 3.415 ;
      RECT 79.055 4.335 79.255 4.535 ;
      RECT 70.89 3.61 71.09 3.81 ;
      RECT 69.29 4.335 69.49 4.535 ;
      RECT 69.065 9.425 69.265 9.625 ;
      RECT 67.73 3.775 67.93 3.975 ;
      RECT 67.35 4.895 67.55 5.095 ;
      RECT 66.85 3.775 67.05 3.975 ;
      RECT 65.89 3.775 66.09 3.975 ;
      RECT 65.17 3.775 65.37 3.975 ;
      RECT 64.17 3.215 64.37 3.415 ;
      RECT 62.73 4.335 62.93 4.535 ;
      RECT 54.565 3.61 54.765 3.81 ;
      RECT 52.965 4.335 53.165 4.535 ;
      RECT 52.74 9.425 52.94 9.625 ;
      RECT 51.405 3.775 51.605 3.975 ;
      RECT 51.025 4.895 51.225 5.095 ;
      RECT 50.525 3.775 50.725 3.975 ;
      RECT 49.565 3.775 49.765 3.975 ;
      RECT 48.845 3.775 49.045 3.975 ;
      RECT 47.845 3.215 48.045 3.415 ;
      RECT 46.405 4.335 46.605 4.535 ;
      RECT 38.24 3.61 38.44 3.81 ;
      RECT 36.64 4.335 36.84 4.535 ;
      RECT 36.415 9.425 36.615 9.625 ;
      RECT 35.08 3.775 35.28 3.975 ;
      RECT 34.7 4.895 34.9 5.095 ;
      RECT 34.2 3.775 34.4 3.975 ;
      RECT 33.24 3.775 33.44 3.975 ;
      RECT 32.52 3.775 32.72 3.975 ;
      RECT 31.52 3.215 31.72 3.415 ;
      RECT 30.08 4.335 30.28 4.535 ;
      RECT 21.915 3.61 22.115 3.81 ;
      RECT 20.315 4.335 20.515 4.535 ;
      RECT 20.09 9.425 20.29 9.625 ;
      RECT 18.755 3.775 18.955 3.975 ;
      RECT 18.375 4.895 18.575 5.095 ;
      RECT 17.875 3.775 18.075 3.975 ;
      RECT 16.915 3.775 17.115 3.975 ;
      RECT 16.195 3.775 16.395 3.975 ;
      RECT 15.195 3.215 15.395 3.415 ;
      RECT 13.755 4.335 13.955 4.535 ;
    LAYER met2 ;
      RECT 11.13 10.685 93.955 10.855 ;
      RECT 93.785 9.56 93.955 10.855 ;
      RECT 11.13 8.54 11.3 10.855 ;
      RECT 93.755 9.56 94.105 9.91 ;
      RECT 11.07 8.54 11.36 8.89 ;
      RECT 90.595 8.505 90.915 8.83 ;
      RECT 90.625 7.98 90.795 8.83 ;
      RECT 90.625 7.98 90.8 8.33 ;
      RECT 90.625 7.98 91.6 8.155 ;
      RECT 91.425 3.26 91.6 8.155 ;
      RECT 91.37 3.26 91.72 3.61 ;
      RECT 91.395 8.94 91.72 9.265 ;
      RECT 90.28 9.03 91.72 9.2 ;
      RECT 90.28 3.69 90.44 9.2 ;
      RECT 90.595 3.66 90.915 3.98 ;
      RECT 90.28 3.69 90.915 3.86 ;
      RECT 80.455 3.13 80.735 3.5 ;
      RECT 80.49 2.585 80.66 3.5 ;
      RECT 89.065 2.585 89.235 3.11 ;
      RECT 88.975 2.755 89.315 3.105 ;
      RECT 80.49 2.585 89.235 2.755 ;
      RECT 85.695 3.69 85.975 4.06 ;
      RECT 84.625 3.715 84.885 4.035 ;
      RECT 87.175 3.525 87.455 3.895 ;
      RECT 87.785 3.435 88.045 3.755 ;
      RECT 84.685 2.875 84.825 4.035 ;
      RECT 85.765 2.875 85.905 4.06 ;
      RECT 86.885 3.525 88.045 3.665 ;
      RECT 86.885 2.875 87.025 3.665 ;
      RECT 84.685 2.875 87.025 3.015 ;
      RECT 84.715 5.015 86.89 5.18 ;
      RECT 86.745 3.895 86.89 5.18 ;
      RECT 83.635 4.81 83.915 5.18 ;
      RECT 83.635 4.925 84.855 5.065 ;
      RECT 86.465 3.895 86.89 4.035 ;
      RECT 86.465 3.715 86.725 4.035 ;
      RECT 79.805 5.295 83.465 5.435 ;
      RECT 83.325 4.48 83.465 5.435 ;
      RECT 79.805 4.365 79.945 5.435 ;
      RECT 86.345 4.555 86.605 4.875 ;
      RECT 83.325 4.48 85.855 4.62 ;
      RECT 85.575 4.25 85.855 4.62 ;
      RECT 79.805 4.365 80.255 4.62 ;
      RECT 79.975 4.25 80.255 4.62 ;
      RECT 86.345 4.365 86.545 4.875 ;
      RECT 85.575 4.365 86.545 4.505 ;
      RECT 86.145 3.155 86.285 4.505 ;
      RECT 86.085 3.155 86.345 3.475 ;
      RECT 77.405 8.94 77.755 9.29 ;
      RECT 85.96 8.895 86.31 9.245 ;
      RECT 77.405 8.97 86.31 9.17 ;
      RECT 79.985 3.715 80.245 4.035 ;
      RECT 79.985 3.805 81.025 3.945 ;
      RECT 80.885 3.015 81.025 3.945 ;
      RECT 83.645 3.155 83.905 3.475 ;
      RECT 80.885 3.015 83.845 3.155 ;
      RECT 83.025 3.995 83.285 4.315 ;
      RECT 83.025 3.995 83.345 4.225 ;
      RECT 83.135 3.69 83.415 4.06 ;
      RECT 82.725 4.555 83.045 4.875 ;
      RECT 82.725 3.435 82.865 4.875 ;
      RECT 82.665 3.435 82.925 3.755 ;
      RECT 80.225 4.835 80.485 5.155 ;
      RECT 80.225 4.925 81.905 5.065 ;
      RECT 81.765 4.645 81.905 5.065 ;
      RECT 81.765 4.645 82.205 4.875 ;
      RECT 81.945 4.555 82.205 4.875 ;
      RECT 81.265 3.715 81.665 4.225 ;
      RECT 81.455 3.69 81.735 4.06 ;
      RECT 81.205 3.715 81.735 4.035 ;
      RECT 74.27 8.505 74.59 8.83 ;
      RECT 74.3 7.98 74.47 8.83 ;
      RECT 74.3 7.98 74.475 8.33 ;
      RECT 74.3 7.98 75.275 8.155 ;
      RECT 75.1 3.26 75.275 8.155 ;
      RECT 75.045 3.26 75.395 3.61 ;
      RECT 75.07 8.94 75.395 9.265 ;
      RECT 73.955 9.03 75.395 9.2 ;
      RECT 73.955 3.69 74.115 9.2 ;
      RECT 74.27 3.66 74.59 3.98 ;
      RECT 73.955 3.69 74.59 3.86 ;
      RECT 64.13 3.13 64.41 3.5 ;
      RECT 64.165 2.585 64.335 3.5 ;
      RECT 72.74 2.585 72.91 3.11 ;
      RECT 72.65 2.755 72.99 3.105 ;
      RECT 64.165 2.585 72.91 2.755 ;
      RECT 69.37 3.69 69.65 4.06 ;
      RECT 68.3 3.715 68.56 4.035 ;
      RECT 70.85 3.525 71.13 3.895 ;
      RECT 71.46 3.435 71.72 3.755 ;
      RECT 68.36 2.875 68.5 4.035 ;
      RECT 69.44 2.875 69.58 4.06 ;
      RECT 70.56 3.525 71.72 3.665 ;
      RECT 70.56 2.875 70.7 3.665 ;
      RECT 68.36 2.875 70.7 3.015 ;
      RECT 68.39 5.015 70.565 5.18 ;
      RECT 70.42 3.895 70.565 5.18 ;
      RECT 67.31 4.81 67.59 5.18 ;
      RECT 67.31 4.925 68.53 5.065 ;
      RECT 70.14 3.895 70.565 4.035 ;
      RECT 70.14 3.715 70.4 4.035 ;
      RECT 63.48 5.295 67.14 5.435 ;
      RECT 67 4.48 67.14 5.435 ;
      RECT 63.48 4.365 63.62 5.435 ;
      RECT 70.02 4.555 70.28 4.875 ;
      RECT 67 4.48 69.53 4.62 ;
      RECT 69.25 4.25 69.53 4.62 ;
      RECT 63.48 4.365 63.93 4.62 ;
      RECT 63.65 4.25 63.93 4.62 ;
      RECT 70.02 4.365 70.22 4.875 ;
      RECT 69.25 4.365 70.22 4.505 ;
      RECT 69.82 3.155 69.96 4.505 ;
      RECT 69.76 3.155 70.02 3.475 ;
      RECT 61.08 8.94 61.43 9.29 ;
      RECT 69.63 8.895 69.98 9.245 ;
      RECT 61.08 8.97 69.98 9.17 ;
      RECT 63.66 3.715 63.92 4.035 ;
      RECT 63.66 3.805 64.7 3.945 ;
      RECT 64.56 3.015 64.7 3.945 ;
      RECT 67.32 3.155 67.58 3.475 ;
      RECT 64.56 3.015 67.52 3.155 ;
      RECT 66.7 3.995 66.96 4.315 ;
      RECT 66.7 3.995 67.02 4.225 ;
      RECT 66.81 3.69 67.09 4.06 ;
      RECT 66.4 4.555 66.72 4.875 ;
      RECT 66.4 3.435 66.54 4.875 ;
      RECT 66.34 3.435 66.6 3.755 ;
      RECT 63.9 4.835 64.16 5.155 ;
      RECT 63.9 4.925 65.58 5.065 ;
      RECT 65.44 4.645 65.58 5.065 ;
      RECT 65.44 4.645 65.88 4.875 ;
      RECT 65.62 4.555 65.88 4.875 ;
      RECT 64.94 3.715 65.34 4.225 ;
      RECT 65.13 3.69 65.41 4.06 ;
      RECT 64.88 3.715 65.41 4.035 ;
      RECT 57.945 8.505 58.265 8.83 ;
      RECT 57.975 7.98 58.145 8.83 ;
      RECT 57.975 7.98 58.15 8.33 ;
      RECT 57.975 7.98 58.95 8.155 ;
      RECT 58.775 3.26 58.95 8.155 ;
      RECT 58.72 3.26 59.07 3.61 ;
      RECT 58.745 8.94 59.07 9.265 ;
      RECT 57.63 9.03 59.07 9.2 ;
      RECT 57.63 3.69 57.79 9.2 ;
      RECT 57.945 3.66 58.265 3.98 ;
      RECT 57.63 3.69 58.265 3.86 ;
      RECT 47.805 3.13 48.085 3.5 ;
      RECT 47.84 2.585 48.01 3.5 ;
      RECT 56.415 2.585 56.585 3.11 ;
      RECT 56.325 2.755 56.665 3.105 ;
      RECT 47.84 2.585 56.585 2.755 ;
      RECT 53.045 3.69 53.325 4.06 ;
      RECT 51.975 3.715 52.235 4.035 ;
      RECT 54.525 3.525 54.805 3.895 ;
      RECT 55.135 3.435 55.395 3.755 ;
      RECT 52.035 2.875 52.175 4.035 ;
      RECT 53.115 2.875 53.255 4.06 ;
      RECT 54.235 3.525 55.395 3.665 ;
      RECT 54.235 2.875 54.375 3.665 ;
      RECT 52.035 2.875 54.375 3.015 ;
      RECT 52.065 5.015 54.24 5.18 ;
      RECT 54.095 3.895 54.24 5.18 ;
      RECT 50.985 4.81 51.265 5.18 ;
      RECT 50.985 4.925 52.205 5.065 ;
      RECT 53.815 3.895 54.24 4.035 ;
      RECT 53.815 3.715 54.075 4.035 ;
      RECT 47.155 5.295 50.815 5.435 ;
      RECT 50.675 4.48 50.815 5.435 ;
      RECT 47.155 4.365 47.295 5.435 ;
      RECT 53.695 4.555 53.955 4.875 ;
      RECT 50.675 4.48 53.205 4.62 ;
      RECT 52.925 4.25 53.205 4.62 ;
      RECT 47.155 4.365 47.605 4.62 ;
      RECT 47.325 4.25 47.605 4.62 ;
      RECT 53.695 4.365 53.895 4.875 ;
      RECT 52.925 4.365 53.895 4.505 ;
      RECT 53.495 3.155 53.635 4.505 ;
      RECT 53.435 3.155 53.695 3.475 ;
      RECT 44.8 8.945 45.15 9.295 ;
      RECT 53.305 8.9 53.655 9.25 ;
      RECT 44.8 8.975 53.655 9.175 ;
      RECT 47.335 3.715 47.595 4.035 ;
      RECT 47.335 3.805 48.375 3.945 ;
      RECT 48.235 3.015 48.375 3.945 ;
      RECT 50.995 3.155 51.255 3.475 ;
      RECT 48.235 3.015 51.195 3.155 ;
      RECT 50.375 3.995 50.635 4.315 ;
      RECT 50.375 3.995 50.695 4.225 ;
      RECT 50.485 3.69 50.765 4.06 ;
      RECT 50.075 4.555 50.395 4.875 ;
      RECT 50.075 3.435 50.215 4.875 ;
      RECT 50.015 3.435 50.275 3.755 ;
      RECT 47.575 4.835 47.835 5.155 ;
      RECT 47.575 4.925 49.255 5.065 ;
      RECT 49.115 4.645 49.255 5.065 ;
      RECT 49.115 4.645 49.555 4.875 ;
      RECT 49.295 4.555 49.555 4.875 ;
      RECT 48.615 3.715 49.015 4.225 ;
      RECT 48.805 3.69 49.085 4.06 ;
      RECT 48.555 3.715 49.085 4.035 ;
      RECT 41.62 8.505 41.94 8.83 ;
      RECT 41.65 7.98 41.82 8.83 ;
      RECT 41.65 7.98 41.825 8.33 ;
      RECT 41.65 7.98 42.625 8.155 ;
      RECT 42.45 3.26 42.625 8.155 ;
      RECT 42.395 3.26 42.745 3.61 ;
      RECT 42.42 8.94 42.745 9.265 ;
      RECT 41.305 9.03 42.745 9.2 ;
      RECT 41.305 3.69 41.465 9.2 ;
      RECT 41.62 3.66 41.94 3.98 ;
      RECT 41.305 3.69 41.94 3.86 ;
      RECT 31.48 3.13 31.76 3.5 ;
      RECT 31.515 2.585 31.685 3.5 ;
      RECT 40.09 2.585 40.26 3.11 ;
      RECT 40 2.755 40.34 3.105 ;
      RECT 31.515 2.585 40.26 2.755 ;
      RECT 36.72 3.69 37 4.06 ;
      RECT 35.65 3.715 35.91 4.035 ;
      RECT 38.2 3.525 38.48 3.895 ;
      RECT 38.81 3.435 39.07 3.755 ;
      RECT 35.71 2.875 35.85 4.035 ;
      RECT 36.79 2.875 36.93 4.06 ;
      RECT 37.91 3.525 39.07 3.665 ;
      RECT 37.91 2.875 38.05 3.665 ;
      RECT 35.71 2.875 38.05 3.015 ;
      RECT 35.74 5.015 37.915 5.18 ;
      RECT 37.77 3.895 37.915 5.18 ;
      RECT 34.66 4.81 34.94 5.18 ;
      RECT 34.66 4.925 35.88 5.065 ;
      RECT 37.49 3.895 37.915 4.035 ;
      RECT 37.49 3.715 37.75 4.035 ;
      RECT 30.83 5.295 34.49 5.435 ;
      RECT 34.35 4.48 34.49 5.435 ;
      RECT 30.83 4.365 30.97 5.435 ;
      RECT 37.37 4.555 37.63 4.875 ;
      RECT 34.35 4.48 36.88 4.62 ;
      RECT 36.6 4.25 36.88 4.62 ;
      RECT 30.83 4.365 31.28 4.62 ;
      RECT 31 4.25 31.28 4.62 ;
      RECT 37.37 4.365 37.57 4.875 ;
      RECT 36.6 4.365 37.57 4.505 ;
      RECT 37.17 3.155 37.31 4.505 ;
      RECT 37.11 3.155 37.37 3.475 ;
      RECT 28.475 8.94 28.825 9.29 ;
      RECT 36.98 8.895 37.33 9.245 ;
      RECT 28.475 8.97 37.33 9.17 ;
      RECT 31.01 3.715 31.27 4.035 ;
      RECT 31.01 3.805 32.05 3.945 ;
      RECT 31.91 3.015 32.05 3.945 ;
      RECT 34.67 3.155 34.93 3.475 ;
      RECT 31.91 3.015 34.87 3.155 ;
      RECT 34.05 3.995 34.31 4.315 ;
      RECT 34.05 3.995 34.37 4.225 ;
      RECT 34.16 3.69 34.44 4.06 ;
      RECT 33.75 4.555 34.07 4.875 ;
      RECT 33.75 3.435 33.89 4.875 ;
      RECT 33.69 3.435 33.95 3.755 ;
      RECT 31.25 4.835 31.51 5.155 ;
      RECT 31.25 4.925 32.93 5.065 ;
      RECT 32.79 4.645 32.93 5.065 ;
      RECT 32.79 4.645 33.23 4.875 ;
      RECT 32.97 4.555 33.23 4.875 ;
      RECT 32.29 3.715 32.69 4.225 ;
      RECT 32.48 3.69 32.76 4.06 ;
      RECT 32.23 3.715 32.76 4.035 ;
      RECT 25.295 8.505 25.615 8.83 ;
      RECT 25.325 7.98 25.495 8.83 ;
      RECT 25.325 7.98 25.5 8.33 ;
      RECT 25.325 7.98 26.3 8.155 ;
      RECT 26.125 3.26 26.3 8.155 ;
      RECT 26.07 3.26 26.42 3.61 ;
      RECT 26.095 8.94 26.42 9.265 ;
      RECT 24.98 9.03 26.42 9.2 ;
      RECT 24.98 3.69 25.14 9.2 ;
      RECT 25.295 3.66 25.615 3.98 ;
      RECT 24.98 3.69 25.615 3.86 ;
      RECT 15.155 3.13 15.435 3.5 ;
      RECT 15.19 2.585 15.36 3.5 ;
      RECT 23.765 2.585 23.935 3.11 ;
      RECT 23.675 2.755 24.015 3.105 ;
      RECT 15.19 2.585 23.935 2.755 ;
      RECT 20.395 3.69 20.675 4.06 ;
      RECT 19.325 3.715 19.585 4.035 ;
      RECT 21.875 3.525 22.155 3.895 ;
      RECT 22.485 3.435 22.745 3.755 ;
      RECT 19.385 2.875 19.525 4.035 ;
      RECT 20.465 2.875 20.605 4.06 ;
      RECT 21.585 3.525 22.745 3.665 ;
      RECT 21.585 2.875 21.725 3.665 ;
      RECT 19.385 2.875 21.725 3.015 ;
      RECT 11.445 9.28 11.735 9.63 ;
      RECT 11.445 9.335 12.73 9.51 ;
      RECT 12.555 8.97 12.73 9.51 ;
      RECT 21.49 8.89 21.84 9.24 ;
      RECT 12.555 8.97 21.84 9.145 ;
      RECT 19.415 5.015 21.59 5.18 ;
      RECT 21.445 3.895 21.59 5.18 ;
      RECT 18.335 4.81 18.615 5.18 ;
      RECT 18.335 4.925 19.555 5.065 ;
      RECT 21.165 3.895 21.59 4.035 ;
      RECT 21.165 3.715 21.425 4.035 ;
      RECT 14.505 5.295 18.165 5.435 ;
      RECT 18.025 4.48 18.165 5.435 ;
      RECT 14.505 4.365 14.645 5.435 ;
      RECT 21.045 4.555 21.305 4.875 ;
      RECT 18.025 4.48 20.555 4.62 ;
      RECT 20.275 4.25 20.555 4.62 ;
      RECT 14.505 4.365 14.955 4.62 ;
      RECT 14.675 4.25 14.955 4.62 ;
      RECT 21.045 4.365 21.245 4.875 ;
      RECT 20.275 4.365 21.245 4.505 ;
      RECT 20.845 3.155 20.985 4.505 ;
      RECT 20.785 3.155 21.045 3.475 ;
      RECT 14.685 3.715 14.945 4.035 ;
      RECT 14.685 3.805 15.725 3.945 ;
      RECT 15.585 3.015 15.725 3.945 ;
      RECT 18.345 3.155 18.605 3.475 ;
      RECT 15.585 3.015 18.545 3.155 ;
      RECT 17.725 3.995 17.985 4.315 ;
      RECT 17.725 3.995 18.045 4.225 ;
      RECT 17.835 3.69 18.115 4.06 ;
      RECT 17.425 4.555 17.745 4.875 ;
      RECT 17.425 3.435 17.565 4.875 ;
      RECT 17.365 3.435 17.625 3.755 ;
      RECT 14.925 4.835 15.185 5.155 ;
      RECT 14.925 4.925 16.605 5.065 ;
      RECT 16.465 4.645 16.605 5.065 ;
      RECT 16.465 4.645 16.905 4.875 ;
      RECT 16.645 4.555 16.905 4.875 ;
      RECT 15.965 3.715 16.365 4.225 ;
      RECT 16.155 3.69 16.435 4.06 ;
      RECT 15.905 3.715 16.435 4.035 ;
      RECT 85.305 9.34 85.675 9.71 ;
      RECT 84.015 3.69 84.295 4.06 ;
      RECT 82.175 3.69 82.455 4.06 ;
      RECT 79.015 4.25 79.295 4.62 ;
      RECT 68.98 9.34 69.35 9.71 ;
      RECT 67.69 3.69 67.97 4.06 ;
      RECT 65.85 3.69 66.13 4.06 ;
      RECT 62.69 4.25 62.97 4.62 ;
      RECT 52.655 9.34 53.025 9.71 ;
      RECT 51.365 3.69 51.645 4.06 ;
      RECT 49.525 3.69 49.805 4.06 ;
      RECT 46.365 4.25 46.645 4.62 ;
      RECT 36.33 9.34 36.7 9.71 ;
      RECT 35.04 3.69 35.32 4.06 ;
      RECT 33.2 3.69 33.48 4.06 ;
      RECT 30.04 4.25 30.32 4.62 ;
      RECT 20.005 9.34 20.375 9.71 ;
      RECT 18.715 3.69 18.995 4.06 ;
      RECT 16.875 3.69 17.155 4.06 ;
      RECT 13.715 4.25 13.995 4.62 ;
    LAYER via1 ;
      RECT 93.855 9.66 94.005 9.81 ;
      RECT 91.485 9.025 91.635 9.175 ;
      RECT 91.47 3.36 91.62 3.51 ;
      RECT 90.68 3.745 90.83 3.895 ;
      RECT 90.68 8.61 90.83 8.76 ;
      RECT 89.075 2.855 89.225 3.005 ;
      RECT 87.84 3.52 87.99 3.67 ;
      RECT 86.52 3.8 86.67 3.95 ;
      RECT 86.4 4.64 86.55 4.79 ;
      RECT 86.14 3.24 86.29 3.39 ;
      RECT 86.06 8.995 86.21 9.145 ;
      RECT 85.415 9.45 85.565 9.6 ;
      RECT 84.68 3.8 84.83 3.95 ;
      RECT 84.08 3.8 84.23 3.95 ;
      RECT 83.7 3.24 83.85 3.39 ;
      RECT 83.08 4.08 83.23 4.23 ;
      RECT 82.84 4.64 82.99 4.79 ;
      RECT 82.72 3.52 82.87 3.67 ;
      RECT 82.24 3.8 82.39 3.95 ;
      RECT 82 4.64 82.15 4.79 ;
      RECT 81.26 3.8 81.41 3.95 ;
      RECT 80.52 3.24 80.67 3.39 ;
      RECT 80.28 4.92 80.43 5.07 ;
      RECT 80.04 3.8 80.19 3.95 ;
      RECT 80.04 4.36 80.19 4.51 ;
      RECT 79.08 4.36 79.23 4.51 ;
      RECT 77.505 9.04 77.655 9.19 ;
      RECT 75.16 9.025 75.31 9.175 ;
      RECT 75.145 3.36 75.295 3.51 ;
      RECT 74.355 3.745 74.505 3.895 ;
      RECT 74.355 8.61 74.505 8.76 ;
      RECT 72.75 2.855 72.9 3.005 ;
      RECT 71.515 3.52 71.665 3.67 ;
      RECT 70.195 3.8 70.345 3.95 ;
      RECT 70.075 4.64 70.225 4.79 ;
      RECT 69.815 3.24 69.965 3.39 ;
      RECT 69.73 8.995 69.88 9.145 ;
      RECT 69.09 9.45 69.24 9.6 ;
      RECT 68.355 3.8 68.505 3.95 ;
      RECT 67.755 3.8 67.905 3.95 ;
      RECT 67.375 3.24 67.525 3.39 ;
      RECT 66.755 4.08 66.905 4.23 ;
      RECT 66.515 4.64 66.665 4.79 ;
      RECT 66.395 3.52 66.545 3.67 ;
      RECT 65.915 3.8 66.065 3.95 ;
      RECT 65.675 4.64 65.825 4.79 ;
      RECT 64.935 3.8 65.085 3.95 ;
      RECT 64.195 3.24 64.345 3.39 ;
      RECT 63.955 4.92 64.105 5.07 ;
      RECT 63.715 3.8 63.865 3.95 ;
      RECT 63.715 4.36 63.865 4.51 ;
      RECT 62.755 4.36 62.905 4.51 ;
      RECT 61.18 9.04 61.33 9.19 ;
      RECT 58.835 9.025 58.985 9.175 ;
      RECT 58.82 3.36 58.97 3.51 ;
      RECT 58.03 3.745 58.18 3.895 ;
      RECT 58.03 8.61 58.18 8.76 ;
      RECT 56.425 2.855 56.575 3.005 ;
      RECT 55.19 3.52 55.34 3.67 ;
      RECT 53.87 3.8 54.02 3.95 ;
      RECT 53.75 4.64 53.9 4.79 ;
      RECT 53.49 3.24 53.64 3.39 ;
      RECT 53.405 9 53.555 9.15 ;
      RECT 52.765 9.45 52.915 9.6 ;
      RECT 52.03 3.8 52.18 3.95 ;
      RECT 51.43 3.8 51.58 3.95 ;
      RECT 51.05 3.24 51.2 3.39 ;
      RECT 50.43 4.08 50.58 4.23 ;
      RECT 50.19 4.64 50.34 4.79 ;
      RECT 50.07 3.52 50.22 3.67 ;
      RECT 49.59 3.8 49.74 3.95 ;
      RECT 49.35 4.64 49.5 4.79 ;
      RECT 48.61 3.8 48.76 3.95 ;
      RECT 47.87 3.24 48.02 3.39 ;
      RECT 47.63 4.92 47.78 5.07 ;
      RECT 47.39 3.8 47.54 3.95 ;
      RECT 47.39 4.36 47.54 4.51 ;
      RECT 46.43 4.36 46.58 4.51 ;
      RECT 44.9 9.045 45.05 9.195 ;
      RECT 42.51 9.025 42.66 9.175 ;
      RECT 42.495 3.36 42.645 3.51 ;
      RECT 41.705 3.745 41.855 3.895 ;
      RECT 41.705 8.61 41.855 8.76 ;
      RECT 40.1 2.855 40.25 3.005 ;
      RECT 38.865 3.52 39.015 3.67 ;
      RECT 37.545 3.8 37.695 3.95 ;
      RECT 37.425 4.64 37.575 4.79 ;
      RECT 37.165 3.24 37.315 3.39 ;
      RECT 37.08 8.995 37.23 9.145 ;
      RECT 36.44 9.45 36.59 9.6 ;
      RECT 35.705 3.8 35.855 3.95 ;
      RECT 35.105 3.8 35.255 3.95 ;
      RECT 34.725 3.24 34.875 3.39 ;
      RECT 34.105 4.08 34.255 4.23 ;
      RECT 33.865 4.64 34.015 4.79 ;
      RECT 33.745 3.52 33.895 3.67 ;
      RECT 33.265 3.8 33.415 3.95 ;
      RECT 33.025 4.64 33.175 4.79 ;
      RECT 32.285 3.8 32.435 3.95 ;
      RECT 31.545 3.24 31.695 3.39 ;
      RECT 31.305 4.92 31.455 5.07 ;
      RECT 31.065 3.8 31.215 3.95 ;
      RECT 31.065 4.36 31.215 4.51 ;
      RECT 30.105 4.36 30.255 4.51 ;
      RECT 28.575 9.04 28.725 9.19 ;
      RECT 26.185 9.025 26.335 9.175 ;
      RECT 26.17 3.36 26.32 3.51 ;
      RECT 25.38 3.745 25.53 3.895 ;
      RECT 25.38 8.61 25.53 8.76 ;
      RECT 23.775 2.855 23.925 3.005 ;
      RECT 22.54 3.52 22.69 3.67 ;
      RECT 21.59 8.99 21.74 9.14 ;
      RECT 21.22 3.8 21.37 3.95 ;
      RECT 21.1 4.64 21.25 4.79 ;
      RECT 20.84 3.24 20.99 3.39 ;
      RECT 20.115 9.45 20.265 9.6 ;
      RECT 19.38 3.8 19.53 3.95 ;
      RECT 18.78 3.8 18.93 3.95 ;
      RECT 18.4 3.24 18.55 3.39 ;
      RECT 17.78 4.08 17.93 4.23 ;
      RECT 17.54 4.64 17.69 4.79 ;
      RECT 17.42 3.52 17.57 3.67 ;
      RECT 16.94 3.8 17.09 3.95 ;
      RECT 16.7 4.64 16.85 4.79 ;
      RECT 15.96 3.8 16.11 3.95 ;
      RECT 15.22 3.24 15.37 3.39 ;
      RECT 14.98 4.92 15.13 5.07 ;
      RECT 14.74 3.8 14.89 3.95 ;
      RECT 14.74 4.36 14.89 4.51 ;
      RECT 13.78 4.36 13.93 4.51 ;
      RECT 11.515 9.38 11.665 9.53 ;
      RECT 11.14 8.64 11.29 8.79 ;
    LAYER met1 ;
      RECT 93.72 10.055 94.01 10.285 ;
      RECT 93.78 8.575 93.95 10.285 ;
      RECT 93.755 9.56 94.105 9.91 ;
      RECT 93.72 8.575 94.01 8.805 ;
      RECT 93.315 3.69 93.42 4.26 ;
      RECT 93.315 4.025 93.64 4.255 ;
      RECT 93.315 4.055 93.81 4.225 ;
      RECT 93.315 3.69 93.505 4.255 ;
      RECT 92.73 3.655 93.02 3.885 ;
      RECT 92.73 3.69 93.505 3.86 ;
      RECT 92.79 2.175 92.96 3.885 ;
      RECT 92.73 2.175 93.02 2.405 ;
      RECT 92.73 10.055 93.02 10.285 ;
      RECT 92.79 8.575 92.96 10.285 ;
      RECT 92.73 8.575 93.02 8.805 ;
      RECT 92.73 8.61 93.585 8.77 ;
      RECT 93.415 8.205 93.585 8.77 ;
      RECT 92.73 8.605 93.125 8.77 ;
      RECT 93.35 8.205 93.64 8.435 ;
      RECT 93.35 8.235 93.81 8.405 ;
      RECT 92.36 4.025 92.65 4.255 ;
      RECT 92.36 4.055 92.82 4.225 ;
      RECT 92.425 2.95 92.59 4.255 ;
      RECT 90.94 2.92 91.23 3.15 ;
      RECT 90.94 2.95 92.59 3.12 ;
      RECT 91 2.18 91.17 3.15 ;
      RECT 90.94 2.18 91.23 2.41 ;
      RECT 90.94 10.05 91.23 10.28 ;
      RECT 91 9.31 91.17 10.28 ;
      RECT 91 9.405 92.59 9.575 ;
      RECT 92.42 8.205 92.59 9.575 ;
      RECT 90.94 9.31 91.23 9.54 ;
      RECT 92.36 8.205 92.65 8.435 ;
      RECT 92.36 8.235 92.82 8.405 ;
      RECT 91.37 3.26 91.72 3.61 ;
      RECT 89.065 3.32 91.72 3.49 ;
      RECT 89.065 2.755 89.235 3.49 ;
      RECT 88.975 2.755 89.315 3.105 ;
      RECT 91.395 8.94 91.72 9.265 ;
      RECT 85.96 8.895 86.31 9.245 ;
      RECT 91.37 8.94 91.72 9.17 ;
      RECT 85.755 8.94 86.31 9.17 ;
      RECT 85.585 8.97 91.72 9.14 ;
      RECT 90.595 3.66 90.915 3.98 ;
      RECT 90.565 3.66 90.915 3.89 ;
      RECT 90.395 3.69 90.915 3.86 ;
      RECT 90.595 8.54 90.915 8.83 ;
      RECT 90.565 8.57 90.915 8.8 ;
      RECT 90.395 8.6 90.915 8.77 ;
      RECT 87.05 3.76 87.34 3.99 ;
      RECT 87.05 3.76 87.505 3.945 ;
      RECT 87.365 3.665 87.985 3.805 ;
      RECT 87.755 3.465 88.075 3.725 ;
      RECT 86.435 3.745 86.755 4.005 ;
      RECT 86.435 3.745 86.9 3.99 ;
      RECT 86.76 3.365 86.9 3.99 ;
      RECT 86.76 3.365 87.025 3.505 ;
      RECT 87.29 3.2 87.58 3.43 ;
      RECT 86.885 3.245 87.58 3.385 ;
      RECT 86.33 4.585 86.62 5.11 ;
      RECT 86.315 4.585 86.635 4.845 ;
      RECT 86.055 3.185 86.375 3.445 ;
      RECT 86.055 3.2 86.62 3.43 ;
      RECT 85.33 4.88 85.62 5.11 ;
      RECT 85.525 3.525 85.665 5.065 ;
      RECT 85.57 3.48 85.86 3.71 ;
      RECT 85.165 3.525 85.86 3.665 ;
      RECT 85.165 3.365 85.305 3.665 ;
      RECT 83.705 3.365 85.305 3.505 ;
      RECT 83.615 3.185 83.935 3.445 ;
      RECT 83.615 3.2 84.18 3.445 ;
      RECT 85.325 10.05 85.615 10.28 ;
      RECT 85.385 9.31 85.555 10.28 ;
      RECT 85.305 9.36 85.675 9.71 ;
      RECT 85.305 9.34 85.615 9.71 ;
      RECT 85.325 9.31 85.615 9.71 ;
      RECT 82.725 4.225 85.305 4.365 ;
      RECT 85.09 4.04 85.38 4.27 ;
      RECT 82.65 4.04 83.315 4.27 ;
      RECT 82.995 4.025 83.315 4.365 ;
      RECT 83.995 3.745 84.315 4.005 ;
      RECT 83.995 3.76 84.42 3.99 ;
      RECT 82.635 3.465 82.955 3.725 ;
      RECT 83.13 3.48 83.42 3.71 ;
      RECT 82.635 3.525 83.42 3.665 ;
      RECT 82.755 4.585 83.075 4.845 ;
      RECT 81.915 4.585 82.235 4.845 ;
      RECT 82.755 4.6 83.18 4.83 ;
      RECT 81.915 4.645 83.18 4.785 ;
      RECT 81.45 4.32 81.74 4.55 ;
      RECT 81.525 3.245 81.665 4.55 ;
      RECT 81.175 3.745 81.665 4.005 ;
      RECT 80.93 3.76 81.665 3.99 ;
      RECT 81.93 3.2 82.22 3.43 ;
      RECT 81.525 3.245 82.22 3.385 ;
      RECT 80.69 4.6 80.98 4.83 ;
      RECT 80.69 4.6 81.145 4.785 ;
      RECT 81.005 4.225 81.145 4.785 ;
      RECT 80.645 4.225 81.145 4.365 ;
      RECT 80.645 3.245 80.785 4.365 ;
      RECT 80.435 3.185 80.755 3.445 ;
      RECT 80.195 4.865 80.515 5.125 ;
      RECT 79.49 4.88 79.78 5.11 ;
      RECT 79.49 4.925 80.515 5.065 ;
      RECT 79.565 4.875 79.825 5.065 ;
      RECT 79.955 3.745 80.275 4.005 ;
      RECT 79.955 3.76 80.5 3.99 ;
      RECT 79.955 4.305 80.275 4.565 ;
      RECT 79.955 4.32 80.5 4.55 ;
      RECT 78.995 4.305 79.315 4.565 ;
      RECT 79.085 3.245 79.225 4.565 ;
      RECT 79.49 3.2 79.78 3.43 ;
      RECT 79.085 3.245 79.78 3.385 ;
      RECT 77.395 10.055 77.685 10.285 ;
      RECT 77.455 8.575 77.625 10.285 ;
      RECT 77.405 8.94 77.755 9.29 ;
      RECT 77.395 8.575 77.685 8.805 ;
      RECT 76.99 3.69 77.095 4.26 ;
      RECT 76.99 4.025 77.315 4.255 ;
      RECT 76.99 4.055 77.485 4.225 ;
      RECT 76.99 3.69 77.18 4.255 ;
      RECT 76.405 3.655 76.695 3.885 ;
      RECT 76.405 3.69 77.18 3.86 ;
      RECT 76.465 2.175 76.635 3.885 ;
      RECT 76.405 2.175 76.695 2.405 ;
      RECT 76.405 10.055 76.695 10.285 ;
      RECT 76.465 8.575 76.635 10.285 ;
      RECT 76.405 8.575 76.695 8.805 ;
      RECT 76.405 8.61 77.26 8.77 ;
      RECT 77.09 8.205 77.26 8.77 ;
      RECT 76.405 8.605 76.8 8.77 ;
      RECT 77.025 8.205 77.315 8.435 ;
      RECT 77.025 8.235 77.485 8.405 ;
      RECT 76.035 4.025 76.325 4.255 ;
      RECT 76.035 4.055 76.495 4.225 ;
      RECT 76.1 2.95 76.265 4.255 ;
      RECT 74.615 2.92 74.905 3.15 ;
      RECT 74.615 2.95 76.265 3.12 ;
      RECT 74.675 2.18 74.845 3.15 ;
      RECT 74.615 2.18 74.905 2.41 ;
      RECT 74.615 10.05 74.905 10.28 ;
      RECT 74.675 9.31 74.845 10.28 ;
      RECT 74.675 9.405 76.265 9.575 ;
      RECT 76.095 8.205 76.265 9.575 ;
      RECT 74.615 9.31 74.905 9.54 ;
      RECT 76.035 8.205 76.325 8.435 ;
      RECT 76.035 8.235 76.495 8.405 ;
      RECT 75.045 3.26 75.395 3.61 ;
      RECT 72.74 3.32 75.395 3.49 ;
      RECT 72.74 2.755 72.91 3.49 ;
      RECT 72.65 2.755 72.99 3.105 ;
      RECT 75.07 8.94 75.395 9.265 ;
      RECT 69.63 8.895 69.98 9.245 ;
      RECT 75.045 8.94 75.395 9.17 ;
      RECT 69.43 8.94 69.98 9.17 ;
      RECT 69.26 8.97 75.395 9.14 ;
      RECT 74.27 3.66 74.59 3.98 ;
      RECT 74.24 3.66 74.59 3.89 ;
      RECT 74.07 3.69 74.59 3.86 ;
      RECT 74.27 8.54 74.59 8.83 ;
      RECT 74.24 8.57 74.59 8.8 ;
      RECT 74.07 8.6 74.59 8.77 ;
      RECT 70.725 3.76 71.015 3.99 ;
      RECT 70.725 3.76 71.18 3.945 ;
      RECT 71.04 3.665 71.66 3.805 ;
      RECT 71.43 3.465 71.75 3.725 ;
      RECT 70.11 3.745 70.43 4.005 ;
      RECT 70.11 3.745 70.575 3.99 ;
      RECT 70.435 3.365 70.575 3.99 ;
      RECT 70.435 3.365 70.7 3.505 ;
      RECT 70.965 3.2 71.255 3.43 ;
      RECT 70.56 3.245 71.255 3.385 ;
      RECT 70.005 4.585 70.295 5.11 ;
      RECT 69.99 4.585 70.31 4.845 ;
      RECT 69.73 3.185 70.05 3.445 ;
      RECT 69.73 3.2 70.295 3.43 ;
      RECT 69.005 4.88 69.295 5.11 ;
      RECT 69.2 3.525 69.34 5.065 ;
      RECT 69.245 3.48 69.535 3.71 ;
      RECT 68.84 3.525 69.535 3.665 ;
      RECT 68.84 3.365 68.98 3.665 ;
      RECT 67.38 3.365 68.98 3.505 ;
      RECT 67.29 3.185 67.61 3.445 ;
      RECT 67.29 3.2 67.855 3.445 ;
      RECT 69 10.05 69.29 10.28 ;
      RECT 69.06 9.31 69.23 10.28 ;
      RECT 68.98 9.36 69.35 9.71 ;
      RECT 68.98 9.34 69.29 9.71 ;
      RECT 69 9.31 69.29 9.71 ;
      RECT 66.4 4.225 68.98 4.365 ;
      RECT 68.765 4.04 69.055 4.27 ;
      RECT 66.325 4.04 66.99 4.27 ;
      RECT 66.67 4.025 66.99 4.365 ;
      RECT 67.67 3.745 67.99 4.005 ;
      RECT 67.67 3.76 68.095 3.99 ;
      RECT 66.31 3.465 66.63 3.725 ;
      RECT 66.805 3.48 67.095 3.71 ;
      RECT 66.31 3.525 67.095 3.665 ;
      RECT 66.43 4.585 66.75 4.845 ;
      RECT 65.59 4.585 65.91 4.845 ;
      RECT 66.43 4.6 66.855 4.83 ;
      RECT 65.59 4.645 66.855 4.785 ;
      RECT 65.125 4.32 65.415 4.55 ;
      RECT 65.2 3.245 65.34 4.55 ;
      RECT 64.85 3.745 65.34 4.005 ;
      RECT 64.605 3.76 65.34 3.99 ;
      RECT 65.605 3.2 65.895 3.43 ;
      RECT 65.2 3.245 65.895 3.385 ;
      RECT 64.365 4.6 64.655 4.83 ;
      RECT 64.365 4.6 64.82 4.785 ;
      RECT 64.68 4.225 64.82 4.785 ;
      RECT 64.32 4.225 64.82 4.365 ;
      RECT 64.32 3.245 64.46 4.365 ;
      RECT 64.11 3.185 64.43 3.445 ;
      RECT 63.87 4.865 64.19 5.125 ;
      RECT 63.165 4.88 63.455 5.11 ;
      RECT 63.165 4.925 64.19 5.065 ;
      RECT 63.24 4.875 63.5 5.065 ;
      RECT 63.63 3.745 63.95 4.005 ;
      RECT 63.63 3.76 64.175 3.99 ;
      RECT 63.63 4.305 63.95 4.565 ;
      RECT 63.63 4.32 64.175 4.55 ;
      RECT 62.67 4.305 62.99 4.565 ;
      RECT 62.76 3.245 62.9 4.565 ;
      RECT 63.165 3.2 63.455 3.43 ;
      RECT 62.76 3.245 63.455 3.385 ;
      RECT 61.07 10.055 61.36 10.285 ;
      RECT 61.13 8.575 61.3 10.285 ;
      RECT 61.08 8.94 61.43 9.29 ;
      RECT 61.07 8.575 61.36 8.805 ;
      RECT 60.665 3.69 60.77 4.26 ;
      RECT 60.665 4.025 60.99 4.255 ;
      RECT 60.665 4.055 61.16 4.225 ;
      RECT 60.665 3.69 60.855 4.255 ;
      RECT 60.08 3.655 60.37 3.885 ;
      RECT 60.08 3.69 60.855 3.86 ;
      RECT 60.14 2.175 60.31 3.885 ;
      RECT 60.08 2.175 60.37 2.405 ;
      RECT 60.08 10.055 60.37 10.285 ;
      RECT 60.14 8.575 60.31 10.285 ;
      RECT 60.08 8.575 60.37 8.805 ;
      RECT 60.08 8.61 60.935 8.77 ;
      RECT 60.765 8.205 60.935 8.77 ;
      RECT 60.08 8.605 60.475 8.77 ;
      RECT 60.7 8.205 60.99 8.435 ;
      RECT 60.7 8.235 61.16 8.405 ;
      RECT 59.71 4.025 60 4.255 ;
      RECT 59.71 4.055 60.17 4.225 ;
      RECT 59.775 2.95 59.94 4.255 ;
      RECT 58.29 2.92 58.58 3.15 ;
      RECT 58.29 2.95 59.94 3.12 ;
      RECT 58.35 2.18 58.52 3.15 ;
      RECT 58.29 2.18 58.58 2.41 ;
      RECT 58.29 10.05 58.58 10.28 ;
      RECT 58.35 9.31 58.52 10.28 ;
      RECT 58.35 9.405 59.94 9.575 ;
      RECT 59.77 8.205 59.94 9.575 ;
      RECT 58.29 9.31 58.58 9.54 ;
      RECT 59.71 8.205 60 8.435 ;
      RECT 59.71 8.235 60.17 8.405 ;
      RECT 58.72 3.26 59.07 3.61 ;
      RECT 56.415 3.32 59.07 3.49 ;
      RECT 56.415 2.755 56.585 3.49 ;
      RECT 56.325 2.755 56.665 3.105 ;
      RECT 58.745 8.94 59.07 9.265 ;
      RECT 53.305 8.9 53.655 9.25 ;
      RECT 58.72 8.94 59.07 9.17 ;
      RECT 53.105 8.94 53.655 9.17 ;
      RECT 52.935 8.97 59.07 9.14 ;
      RECT 57.945 3.66 58.265 3.98 ;
      RECT 57.915 3.66 58.265 3.89 ;
      RECT 57.745 3.69 58.265 3.86 ;
      RECT 57.945 8.54 58.265 8.83 ;
      RECT 57.915 8.57 58.265 8.8 ;
      RECT 57.745 8.6 58.265 8.77 ;
      RECT 54.4 3.76 54.69 3.99 ;
      RECT 54.4 3.76 54.855 3.945 ;
      RECT 54.715 3.665 55.335 3.805 ;
      RECT 55.105 3.465 55.425 3.725 ;
      RECT 53.785 3.745 54.105 4.005 ;
      RECT 53.785 3.745 54.25 3.99 ;
      RECT 54.11 3.365 54.25 3.99 ;
      RECT 54.11 3.365 54.375 3.505 ;
      RECT 54.64 3.2 54.93 3.43 ;
      RECT 54.235 3.245 54.93 3.385 ;
      RECT 53.68 4.585 53.97 5.11 ;
      RECT 53.665 4.585 53.985 4.845 ;
      RECT 53.405 3.185 53.725 3.445 ;
      RECT 53.405 3.2 53.97 3.43 ;
      RECT 52.68 4.88 52.97 5.11 ;
      RECT 52.875 3.525 53.015 5.065 ;
      RECT 52.92 3.48 53.21 3.71 ;
      RECT 52.515 3.525 53.21 3.665 ;
      RECT 52.515 3.365 52.655 3.665 ;
      RECT 51.055 3.365 52.655 3.505 ;
      RECT 50.965 3.185 51.285 3.445 ;
      RECT 50.965 3.2 51.53 3.445 ;
      RECT 52.675 10.05 52.965 10.28 ;
      RECT 52.735 9.31 52.905 10.28 ;
      RECT 52.655 9.36 53.025 9.71 ;
      RECT 52.655 9.34 52.965 9.71 ;
      RECT 52.675 9.31 52.965 9.71 ;
      RECT 50.075 4.225 52.655 4.365 ;
      RECT 52.44 4.04 52.73 4.27 ;
      RECT 50 4.04 50.665 4.27 ;
      RECT 50.345 4.025 50.665 4.365 ;
      RECT 51.345 3.745 51.665 4.005 ;
      RECT 51.345 3.76 51.77 3.99 ;
      RECT 49.985 3.465 50.305 3.725 ;
      RECT 50.48 3.48 50.77 3.71 ;
      RECT 49.985 3.525 50.77 3.665 ;
      RECT 50.105 4.585 50.425 4.845 ;
      RECT 49.265 4.585 49.585 4.845 ;
      RECT 50.105 4.6 50.53 4.83 ;
      RECT 49.265 4.645 50.53 4.785 ;
      RECT 48.8 4.32 49.09 4.55 ;
      RECT 48.875 3.245 49.015 4.55 ;
      RECT 48.525 3.745 49.015 4.005 ;
      RECT 48.28 3.76 49.015 3.99 ;
      RECT 49.28 3.2 49.57 3.43 ;
      RECT 48.875 3.245 49.57 3.385 ;
      RECT 48.04 4.6 48.33 4.83 ;
      RECT 48.04 4.6 48.495 4.785 ;
      RECT 48.355 4.225 48.495 4.785 ;
      RECT 47.995 4.225 48.495 4.365 ;
      RECT 47.995 3.245 48.135 4.365 ;
      RECT 47.785 3.185 48.105 3.445 ;
      RECT 47.545 4.865 47.865 5.125 ;
      RECT 46.84 4.88 47.13 5.11 ;
      RECT 46.84 4.925 47.865 5.065 ;
      RECT 46.915 4.875 47.175 5.065 ;
      RECT 47.305 3.745 47.625 4.005 ;
      RECT 47.305 3.76 47.85 3.99 ;
      RECT 47.305 4.305 47.625 4.565 ;
      RECT 47.305 4.32 47.85 4.55 ;
      RECT 46.345 4.305 46.665 4.565 ;
      RECT 46.435 3.245 46.575 4.565 ;
      RECT 46.84 3.2 47.13 3.43 ;
      RECT 46.435 3.245 47.13 3.385 ;
      RECT 44.745 10.055 45.035 10.285 ;
      RECT 44.805 8.575 44.975 10.285 ;
      RECT 44.795 8.945 45.15 9.3 ;
      RECT 44.745 8.575 45.035 8.805 ;
      RECT 44.34 3.69 44.445 4.26 ;
      RECT 44.34 4.025 44.665 4.255 ;
      RECT 44.34 4.055 44.835 4.225 ;
      RECT 44.34 3.69 44.53 4.255 ;
      RECT 43.755 3.655 44.045 3.885 ;
      RECT 43.755 3.69 44.53 3.86 ;
      RECT 43.815 2.175 43.985 3.885 ;
      RECT 43.755 2.175 44.045 2.405 ;
      RECT 43.755 10.055 44.045 10.285 ;
      RECT 43.815 8.575 43.985 10.285 ;
      RECT 43.755 8.575 44.045 8.805 ;
      RECT 43.755 8.61 44.61 8.77 ;
      RECT 44.44 8.205 44.61 8.77 ;
      RECT 43.755 8.605 44.15 8.77 ;
      RECT 44.375 8.205 44.665 8.435 ;
      RECT 44.375 8.235 44.835 8.405 ;
      RECT 43.385 4.025 43.675 4.255 ;
      RECT 43.385 4.055 43.845 4.225 ;
      RECT 43.45 2.95 43.615 4.255 ;
      RECT 41.965 2.92 42.255 3.15 ;
      RECT 41.965 2.95 43.615 3.12 ;
      RECT 42.025 2.18 42.195 3.15 ;
      RECT 41.965 2.18 42.255 2.41 ;
      RECT 41.965 10.05 42.255 10.28 ;
      RECT 42.025 9.31 42.195 10.28 ;
      RECT 42.025 9.405 43.615 9.575 ;
      RECT 43.445 8.205 43.615 9.575 ;
      RECT 41.965 9.31 42.255 9.54 ;
      RECT 43.385 8.205 43.675 8.435 ;
      RECT 43.385 8.235 43.845 8.405 ;
      RECT 42.395 3.26 42.745 3.61 ;
      RECT 40.09 3.32 42.745 3.49 ;
      RECT 40.09 2.755 40.26 3.49 ;
      RECT 40 2.755 40.34 3.105 ;
      RECT 42.42 8.94 42.745 9.265 ;
      RECT 36.98 8.895 37.33 9.245 ;
      RECT 42.395 8.94 42.745 9.17 ;
      RECT 36.78 8.94 37.33 9.17 ;
      RECT 36.61 8.97 42.745 9.14 ;
      RECT 41.62 3.66 41.94 3.98 ;
      RECT 41.59 3.66 41.94 3.89 ;
      RECT 41.42 3.69 41.94 3.86 ;
      RECT 41.62 8.54 41.94 8.83 ;
      RECT 41.59 8.57 41.94 8.8 ;
      RECT 41.42 8.6 41.94 8.77 ;
      RECT 38.075 3.76 38.365 3.99 ;
      RECT 38.075 3.76 38.53 3.945 ;
      RECT 38.39 3.665 39.01 3.805 ;
      RECT 38.78 3.465 39.1 3.725 ;
      RECT 37.46 3.745 37.78 4.005 ;
      RECT 37.46 3.745 37.925 3.99 ;
      RECT 37.785 3.365 37.925 3.99 ;
      RECT 37.785 3.365 38.05 3.505 ;
      RECT 38.315 3.2 38.605 3.43 ;
      RECT 37.91 3.245 38.605 3.385 ;
      RECT 37.355 4.585 37.645 5.11 ;
      RECT 37.34 4.585 37.66 4.845 ;
      RECT 37.08 3.185 37.4 3.445 ;
      RECT 37.08 3.2 37.645 3.43 ;
      RECT 36.355 4.88 36.645 5.11 ;
      RECT 36.55 3.525 36.69 5.065 ;
      RECT 36.595 3.48 36.885 3.71 ;
      RECT 36.19 3.525 36.885 3.665 ;
      RECT 36.19 3.365 36.33 3.665 ;
      RECT 34.73 3.365 36.33 3.505 ;
      RECT 34.64 3.185 34.96 3.445 ;
      RECT 34.64 3.2 35.205 3.445 ;
      RECT 36.35 10.05 36.64 10.28 ;
      RECT 36.41 9.31 36.58 10.28 ;
      RECT 36.33 9.36 36.7 9.71 ;
      RECT 36.33 9.34 36.64 9.71 ;
      RECT 36.35 9.31 36.64 9.71 ;
      RECT 33.75 4.225 36.33 4.365 ;
      RECT 36.115 4.04 36.405 4.27 ;
      RECT 33.675 4.04 34.34 4.27 ;
      RECT 34.02 4.025 34.34 4.365 ;
      RECT 35.02 3.745 35.34 4.005 ;
      RECT 35.02 3.76 35.445 3.99 ;
      RECT 33.66 3.465 33.98 3.725 ;
      RECT 34.155 3.48 34.445 3.71 ;
      RECT 33.66 3.525 34.445 3.665 ;
      RECT 33.78 4.585 34.1 4.845 ;
      RECT 32.94 4.585 33.26 4.845 ;
      RECT 33.78 4.6 34.205 4.83 ;
      RECT 32.94 4.645 34.205 4.785 ;
      RECT 32.475 4.32 32.765 4.55 ;
      RECT 32.55 3.245 32.69 4.55 ;
      RECT 32.2 3.745 32.69 4.005 ;
      RECT 31.955 3.76 32.69 3.99 ;
      RECT 32.955 3.2 33.245 3.43 ;
      RECT 32.55 3.245 33.245 3.385 ;
      RECT 31.715 4.6 32.005 4.83 ;
      RECT 31.715 4.6 32.17 4.785 ;
      RECT 32.03 4.225 32.17 4.785 ;
      RECT 31.67 4.225 32.17 4.365 ;
      RECT 31.67 3.245 31.81 4.365 ;
      RECT 31.46 3.185 31.78 3.445 ;
      RECT 31.22 4.865 31.54 5.125 ;
      RECT 30.515 4.88 30.805 5.11 ;
      RECT 30.515 4.925 31.54 5.065 ;
      RECT 30.59 4.875 30.85 5.065 ;
      RECT 30.98 3.745 31.3 4.005 ;
      RECT 30.98 3.76 31.525 3.99 ;
      RECT 30.98 4.305 31.3 4.565 ;
      RECT 30.98 4.32 31.525 4.55 ;
      RECT 30.02 4.305 30.34 4.565 ;
      RECT 30.11 3.245 30.25 4.565 ;
      RECT 30.515 3.2 30.805 3.43 ;
      RECT 30.11 3.245 30.805 3.385 ;
      RECT 28.42 10.055 28.71 10.285 ;
      RECT 28.48 8.575 28.65 10.285 ;
      RECT 28.475 8.94 28.825 9.29 ;
      RECT 28.42 8.575 28.71 8.805 ;
      RECT 28.015 3.69 28.12 4.26 ;
      RECT 28.015 4.025 28.34 4.255 ;
      RECT 28.015 4.055 28.51 4.225 ;
      RECT 28.015 3.69 28.205 4.255 ;
      RECT 27.43 3.655 27.72 3.885 ;
      RECT 27.43 3.69 28.205 3.86 ;
      RECT 27.49 2.175 27.66 3.885 ;
      RECT 27.43 2.175 27.72 2.405 ;
      RECT 27.43 10.055 27.72 10.285 ;
      RECT 27.49 8.575 27.66 10.285 ;
      RECT 27.43 8.575 27.72 8.805 ;
      RECT 27.43 8.61 28.285 8.77 ;
      RECT 28.115 8.205 28.285 8.77 ;
      RECT 27.43 8.605 27.825 8.77 ;
      RECT 28.05 8.205 28.34 8.435 ;
      RECT 28.05 8.235 28.51 8.405 ;
      RECT 27.06 4.025 27.35 4.255 ;
      RECT 27.06 4.055 27.52 4.225 ;
      RECT 27.125 2.95 27.29 4.255 ;
      RECT 25.64 2.92 25.93 3.15 ;
      RECT 25.64 2.95 27.29 3.12 ;
      RECT 25.7 2.18 25.87 3.15 ;
      RECT 25.64 2.18 25.93 2.41 ;
      RECT 25.64 10.05 25.93 10.28 ;
      RECT 25.7 9.31 25.87 10.28 ;
      RECT 25.7 9.405 27.29 9.575 ;
      RECT 27.12 8.205 27.29 9.575 ;
      RECT 25.64 9.31 25.93 9.54 ;
      RECT 27.06 8.205 27.35 8.435 ;
      RECT 27.06 8.235 27.52 8.405 ;
      RECT 26.07 3.26 26.42 3.61 ;
      RECT 23.765 3.32 26.42 3.49 ;
      RECT 23.765 2.755 23.935 3.49 ;
      RECT 23.675 2.755 24.015 3.105 ;
      RECT 26.095 8.94 26.42 9.265 ;
      RECT 21.49 8.89 21.84 9.24 ;
      RECT 26.07 8.94 26.42 9.17 ;
      RECT 20.455 8.94 20.745 9.17 ;
      RECT 20.285 8.97 26.42 9.14 ;
      RECT 25.295 3.66 25.615 3.98 ;
      RECT 25.265 3.66 25.615 3.89 ;
      RECT 25.095 3.69 25.615 3.86 ;
      RECT 25.295 8.54 25.615 8.83 ;
      RECT 25.265 8.57 25.615 8.8 ;
      RECT 25.095 8.6 25.615 8.77 ;
      RECT 21.75 3.76 22.04 3.99 ;
      RECT 21.75 3.76 22.205 3.945 ;
      RECT 22.065 3.665 22.685 3.805 ;
      RECT 22.455 3.465 22.775 3.725 ;
      RECT 21.135 3.745 21.455 4.005 ;
      RECT 21.135 3.745 21.6 3.99 ;
      RECT 21.46 3.365 21.6 3.99 ;
      RECT 21.46 3.365 21.725 3.505 ;
      RECT 21.99 3.2 22.28 3.43 ;
      RECT 21.585 3.245 22.28 3.385 ;
      RECT 21.03 4.585 21.32 5.11 ;
      RECT 21.015 4.585 21.335 4.845 ;
      RECT 20.755 3.185 21.075 3.445 ;
      RECT 20.755 3.2 21.32 3.43 ;
      RECT 20.03 4.88 20.32 5.11 ;
      RECT 20.225 3.525 20.365 5.065 ;
      RECT 20.27 3.48 20.56 3.71 ;
      RECT 19.865 3.525 20.56 3.665 ;
      RECT 19.865 3.365 20.005 3.665 ;
      RECT 18.405 3.365 20.005 3.505 ;
      RECT 18.315 3.185 18.635 3.445 ;
      RECT 18.315 3.2 18.88 3.445 ;
      RECT 20.025 10.05 20.315 10.28 ;
      RECT 20.085 9.31 20.255 10.28 ;
      RECT 20.005 9.36 20.375 9.71 ;
      RECT 20.005 9.34 20.315 9.71 ;
      RECT 20.025 9.31 20.315 9.71 ;
      RECT 17.425 4.225 20.005 4.365 ;
      RECT 19.79 4.04 20.08 4.27 ;
      RECT 17.35 4.04 18.015 4.27 ;
      RECT 17.695 4.025 18.015 4.365 ;
      RECT 18.695 3.745 19.015 4.005 ;
      RECT 18.695 3.76 19.12 3.99 ;
      RECT 17.335 3.465 17.655 3.725 ;
      RECT 17.83 3.48 18.12 3.71 ;
      RECT 17.335 3.525 18.12 3.665 ;
      RECT 17.455 4.585 17.775 4.845 ;
      RECT 16.615 4.585 16.935 4.845 ;
      RECT 17.455 4.6 17.88 4.83 ;
      RECT 16.615 4.645 17.88 4.785 ;
      RECT 16.15 4.32 16.44 4.55 ;
      RECT 16.225 3.245 16.365 4.55 ;
      RECT 15.875 3.745 16.365 4.005 ;
      RECT 15.63 3.76 16.365 3.99 ;
      RECT 16.63 3.2 16.92 3.43 ;
      RECT 16.225 3.245 16.92 3.385 ;
      RECT 15.39 4.6 15.68 4.83 ;
      RECT 15.39 4.6 15.845 4.785 ;
      RECT 15.705 4.225 15.845 4.785 ;
      RECT 15.345 4.225 15.845 4.365 ;
      RECT 15.345 3.245 15.485 4.365 ;
      RECT 15.135 3.185 15.455 3.445 ;
      RECT 14.895 4.865 15.215 5.125 ;
      RECT 14.19 4.88 14.48 5.11 ;
      RECT 14.19 4.925 15.215 5.065 ;
      RECT 14.265 4.875 14.525 5.065 ;
      RECT 14.655 3.745 14.975 4.005 ;
      RECT 14.655 3.76 15.2 3.99 ;
      RECT 14.655 4.305 14.975 4.565 ;
      RECT 14.655 4.32 15.2 4.55 ;
      RECT 13.695 4.305 14.015 4.565 ;
      RECT 13.785 3.245 13.925 4.565 ;
      RECT 14.19 3.2 14.48 3.43 ;
      RECT 13.785 3.245 14.48 3.385 ;
      RECT 11.445 10.05 11.735 10.28 ;
      RECT 11.505 9.31 11.675 10.28 ;
      RECT 11.415 9.31 11.765 9.6 ;
      RECT 11.04 8.57 11.39 8.86 ;
      RECT 10.9 8.6 11.39 8.77 ;
      RECT 84.595 3.745 84.915 4.005 ;
      RECT 82.155 3.745 82.475 4.005 ;
      RECT 68.27 3.745 68.59 4.005 ;
      RECT 65.83 3.745 66.15 4.005 ;
      RECT 51.945 3.745 52.265 4.005 ;
      RECT 49.505 3.745 49.825 4.005 ;
      RECT 35.62 3.745 35.94 4.005 ;
      RECT 33.18 3.745 33.5 4.005 ;
      RECT 19.295 3.745 19.615 4.005 ;
      RECT 16.855 3.745 17.175 4.005 ;
    LAYER mcon ;
      RECT 93.78 8.605 93.95 8.775 ;
      RECT 93.785 8.6 93.955 8.77 ;
      RECT 77.455 8.605 77.625 8.775 ;
      RECT 77.46 8.6 77.63 8.77 ;
      RECT 61.13 8.605 61.3 8.775 ;
      RECT 61.135 8.6 61.305 8.77 ;
      RECT 44.805 8.605 44.975 8.775 ;
      RECT 44.81 8.6 44.98 8.77 ;
      RECT 28.48 8.605 28.65 8.775 ;
      RECT 28.485 8.6 28.655 8.77 ;
      RECT 93.78 10.085 93.95 10.255 ;
      RECT 93.41 4.055 93.58 4.225 ;
      RECT 93.41 8.235 93.58 8.405 ;
      RECT 92.79 2.205 92.96 2.375 ;
      RECT 92.79 3.685 92.96 3.855 ;
      RECT 92.79 8.605 92.96 8.775 ;
      RECT 92.79 10.085 92.96 10.255 ;
      RECT 92.42 4.055 92.59 4.225 ;
      RECT 92.42 8.235 92.59 8.405 ;
      RECT 91.43 3.32 91.6 3.49 ;
      RECT 91.43 8.97 91.6 9.14 ;
      RECT 91 2.21 91.17 2.38 ;
      RECT 91 2.95 91.17 3.12 ;
      RECT 91 9.34 91.17 9.51 ;
      RECT 91 10.08 91.17 10.25 ;
      RECT 90.625 3.69 90.795 3.86 ;
      RECT 90.625 8.6 90.795 8.77 ;
      RECT 87.35 3.23 87.52 3.4 ;
      RECT 87.11 3.79 87.28 3.96 ;
      RECT 86.63 3.79 86.8 3.96 ;
      RECT 86.39 3.23 86.56 3.4 ;
      RECT 86.39 4.91 86.56 5.08 ;
      RECT 85.815 8.97 85.985 9.14 ;
      RECT 85.63 3.51 85.8 3.68 ;
      RECT 85.39 4.91 85.56 5.08 ;
      RECT 85.385 9.34 85.555 9.51 ;
      RECT 85.385 10.08 85.555 10.25 ;
      RECT 85.15 4.07 85.32 4.24 ;
      RECT 84.67 3.79 84.84 3.96 ;
      RECT 84.19 3.79 84.36 3.96 ;
      RECT 83.95 3.23 84.12 3.4 ;
      RECT 83.19 3.51 83.36 3.68 ;
      RECT 82.95 4.63 83.12 4.8 ;
      RECT 82.71 4.07 82.88 4.24 ;
      RECT 82.23 3.79 82.4 3.96 ;
      RECT 81.99 3.23 82.16 3.4 ;
      RECT 81.99 4.63 82.16 4.8 ;
      RECT 81.51 4.35 81.68 4.52 ;
      RECT 80.99 3.79 81.16 3.96 ;
      RECT 80.75 4.63 80.92 4.8 ;
      RECT 80.51 3.23 80.68 3.4 ;
      RECT 80.27 3.79 80.44 3.96 ;
      RECT 80.27 4.35 80.44 4.52 ;
      RECT 79.55 3.23 79.72 3.4 ;
      RECT 79.55 4.91 79.72 5.08 ;
      RECT 79.07 4.35 79.24 4.52 ;
      RECT 77.455 10.085 77.625 10.255 ;
      RECT 77.085 4.055 77.255 4.225 ;
      RECT 77.085 8.235 77.255 8.405 ;
      RECT 76.465 2.205 76.635 2.375 ;
      RECT 76.465 3.685 76.635 3.855 ;
      RECT 76.465 8.605 76.635 8.775 ;
      RECT 76.465 10.085 76.635 10.255 ;
      RECT 76.095 4.055 76.265 4.225 ;
      RECT 76.095 8.235 76.265 8.405 ;
      RECT 75.105 3.32 75.275 3.49 ;
      RECT 75.105 8.97 75.275 9.14 ;
      RECT 74.675 2.21 74.845 2.38 ;
      RECT 74.675 2.95 74.845 3.12 ;
      RECT 74.675 9.34 74.845 9.51 ;
      RECT 74.675 10.08 74.845 10.25 ;
      RECT 74.3 3.69 74.47 3.86 ;
      RECT 74.3 8.6 74.47 8.77 ;
      RECT 71.025 3.23 71.195 3.4 ;
      RECT 70.785 3.79 70.955 3.96 ;
      RECT 70.305 3.79 70.475 3.96 ;
      RECT 70.065 3.23 70.235 3.4 ;
      RECT 70.065 4.91 70.235 5.08 ;
      RECT 69.49 8.97 69.66 9.14 ;
      RECT 69.305 3.51 69.475 3.68 ;
      RECT 69.065 4.91 69.235 5.08 ;
      RECT 69.06 9.34 69.23 9.51 ;
      RECT 69.06 10.08 69.23 10.25 ;
      RECT 68.825 4.07 68.995 4.24 ;
      RECT 68.345 3.79 68.515 3.96 ;
      RECT 67.865 3.79 68.035 3.96 ;
      RECT 67.625 3.23 67.795 3.4 ;
      RECT 66.865 3.51 67.035 3.68 ;
      RECT 66.625 4.63 66.795 4.8 ;
      RECT 66.385 4.07 66.555 4.24 ;
      RECT 65.905 3.79 66.075 3.96 ;
      RECT 65.665 3.23 65.835 3.4 ;
      RECT 65.665 4.63 65.835 4.8 ;
      RECT 65.185 4.35 65.355 4.52 ;
      RECT 64.665 3.79 64.835 3.96 ;
      RECT 64.425 4.63 64.595 4.8 ;
      RECT 64.185 3.23 64.355 3.4 ;
      RECT 63.945 3.79 64.115 3.96 ;
      RECT 63.945 4.35 64.115 4.52 ;
      RECT 63.225 3.23 63.395 3.4 ;
      RECT 63.225 4.91 63.395 5.08 ;
      RECT 62.745 4.35 62.915 4.52 ;
      RECT 61.13 10.085 61.3 10.255 ;
      RECT 60.76 4.055 60.93 4.225 ;
      RECT 60.76 8.235 60.93 8.405 ;
      RECT 60.14 2.205 60.31 2.375 ;
      RECT 60.14 3.685 60.31 3.855 ;
      RECT 60.14 8.605 60.31 8.775 ;
      RECT 60.14 10.085 60.31 10.255 ;
      RECT 59.77 4.055 59.94 4.225 ;
      RECT 59.77 8.235 59.94 8.405 ;
      RECT 58.78 3.32 58.95 3.49 ;
      RECT 58.78 8.97 58.95 9.14 ;
      RECT 58.35 2.21 58.52 2.38 ;
      RECT 58.35 2.95 58.52 3.12 ;
      RECT 58.35 9.34 58.52 9.51 ;
      RECT 58.35 10.08 58.52 10.25 ;
      RECT 57.975 3.69 58.145 3.86 ;
      RECT 57.975 8.6 58.145 8.77 ;
      RECT 54.7 3.23 54.87 3.4 ;
      RECT 54.46 3.79 54.63 3.96 ;
      RECT 53.98 3.79 54.15 3.96 ;
      RECT 53.74 3.23 53.91 3.4 ;
      RECT 53.74 4.91 53.91 5.08 ;
      RECT 53.165 8.97 53.335 9.14 ;
      RECT 52.98 3.51 53.15 3.68 ;
      RECT 52.74 4.91 52.91 5.08 ;
      RECT 52.735 9.34 52.905 9.51 ;
      RECT 52.735 10.08 52.905 10.25 ;
      RECT 52.5 4.07 52.67 4.24 ;
      RECT 52.02 3.79 52.19 3.96 ;
      RECT 51.54 3.79 51.71 3.96 ;
      RECT 51.3 3.23 51.47 3.4 ;
      RECT 50.54 3.51 50.71 3.68 ;
      RECT 50.3 4.63 50.47 4.8 ;
      RECT 50.06 4.07 50.23 4.24 ;
      RECT 49.58 3.79 49.75 3.96 ;
      RECT 49.34 3.23 49.51 3.4 ;
      RECT 49.34 4.63 49.51 4.8 ;
      RECT 48.86 4.35 49.03 4.52 ;
      RECT 48.34 3.79 48.51 3.96 ;
      RECT 48.1 4.63 48.27 4.8 ;
      RECT 47.86 3.23 48.03 3.4 ;
      RECT 47.62 3.79 47.79 3.96 ;
      RECT 47.62 4.35 47.79 4.52 ;
      RECT 46.9 3.23 47.07 3.4 ;
      RECT 46.9 4.91 47.07 5.08 ;
      RECT 46.42 4.35 46.59 4.52 ;
      RECT 44.805 10.085 44.975 10.255 ;
      RECT 44.435 4.055 44.605 4.225 ;
      RECT 44.435 8.235 44.605 8.405 ;
      RECT 43.815 2.205 43.985 2.375 ;
      RECT 43.815 3.685 43.985 3.855 ;
      RECT 43.815 8.605 43.985 8.775 ;
      RECT 43.815 10.085 43.985 10.255 ;
      RECT 43.445 4.055 43.615 4.225 ;
      RECT 43.445 8.235 43.615 8.405 ;
      RECT 42.455 3.32 42.625 3.49 ;
      RECT 42.455 8.97 42.625 9.14 ;
      RECT 42.025 2.21 42.195 2.38 ;
      RECT 42.025 2.95 42.195 3.12 ;
      RECT 42.025 9.34 42.195 9.51 ;
      RECT 42.025 10.08 42.195 10.25 ;
      RECT 41.65 3.69 41.82 3.86 ;
      RECT 41.65 8.6 41.82 8.77 ;
      RECT 38.375 3.23 38.545 3.4 ;
      RECT 38.135 3.79 38.305 3.96 ;
      RECT 37.655 3.79 37.825 3.96 ;
      RECT 37.415 3.23 37.585 3.4 ;
      RECT 37.415 4.91 37.585 5.08 ;
      RECT 36.84 8.97 37.01 9.14 ;
      RECT 36.655 3.51 36.825 3.68 ;
      RECT 36.415 4.91 36.585 5.08 ;
      RECT 36.41 9.34 36.58 9.51 ;
      RECT 36.41 10.08 36.58 10.25 ;
      RECT 36.175 4.07 36.345 4.24 ;
      RECT 35.695 3.79 35.865 3.96 ;
      RECT 35.215 3.79 35.385 3.96 ;
      RECT 34.975 3.23 35.145 3.4 ;
      RECT 34.215 3.51 34.385 3.68 ;
      RECT 33.975 4.63 34.145 4.8 ;
      RECT 33.735 4.07 33.905 4.24 ;
      RECT 33.255 3.79 33.425 3.96 ;
      RECT 33.015 3.23 33.185 3.4 ;
      RECT 33.015 4.63 33.185 4.8 ;
      RECT 32.535 4.35 32.705 4.52 ;
      RECT 32.015 3.79 32.185 3.96 ;
      RECT 31.775 4.63 31.945 4.8 ;
      RECT 31.535 3.23 31.705 3.4 ;
      RECT 31.295 3.79 31.465 3.96 ;
      RECT 31.295 4.35 31.465 4.52 ;
      RECT 30.575 3.23 30.745 3.4 ;
      RECT 30.575 4.91 30.745 5.08 ;
      RECT 30.095 4.35 30.265 4.52 ;
      RECT 28.48 10.085 28.65 10.255 ;
      RECT 28.11 4.055 28.28 4.225 ;
      RECT 28.11 8.235 28.28 8.405 ;
      RECT 27.49 2.205 27.66 2.375 ;
      RECT 27.49 3.685 27.66 3.855 ;
      RECT 27.49 8.605 27.66 8.775 ;
      RECT 27.49 10.085 27.66 10.255 ;
      RECT 27.12 4.055 27.29 4.225 ;
      RECT 27.12 8.235 27.29 8.405 ;
      RECT 26.13 3.32 26.3 3.49 ;
      RECT 26.13 8.97 26.3 9.14 ;
      RECT 25.7 2.21 25.87 2.38 ;
      RECT 25.7 2.95 25.87 3.12 ;
      RECT 25.7 9.34 25.87 9.51 ;
      RECT 25.7 10.08 25.87 10.25 ;
      RECT 25.325 3.69 25.495 3.86 ;
      RECT 25.325 8.6 25.495 8.77 ;
      RECT 22.05 3.23 22.22 3.4 ;
      RECT 21.81 3.79 21.98 3.96 ;
      RECT 21.33 3.79 21.5 3.96 ;
      RECT 21.09 3.23 21.26 3.4 ;
      RECT 21.09 4.91 21.26 5.08 ;
      RECT 20.515 8.97 20.685 9.14 ;
      RECT 20.33 3.51 20.5 3.68 ;
      RECT 20.09 4.91 20.26 5.08 ;
      RECT 20.085 9.34 20.255 9.51 ;
      RECT 20.085 10.08 20.255 10.25 ;
      RECT 19.85 4.07 20.02 4.24 ;
      RECT 19.37 3.79 19.54 3.96 ;
      RECT 18.89 3.79 19.06 3.96 ;
      RECT 18.65 3.23 18.82 3.4 ;
      RECT 17.89 3.51 18.06 3.68 ;
      RECT 17.65 4.63 17.82 4.8 ;
      RECT 17.41 4.07 17.58 4.24 ;
      RECT 16.93 3.79 17.1 3.96 ;
      RECT 16.69 3.23 16.86 3.4 ;
      RECT 16.69 4.63 16.86 4.8 ;
      RECT 16.21 4.35 16.38 4.52 ;
      RECT 15.69 3.79 15.86 3.96 ;
      RECT 15.45 4.63 15.62 4.8 ;
      RECT 15.21 3.23 15.38 3.4 ;
      RECT 14.97 3.79 15.14 3.96 ;
      RECT 14.97 4.35 15.14 4.52 ;
      RECT 14.25 3.23 14.42 3.4 ;
      RECT 14.25 4.91 14.42 5.08 ;
      RECT 13.77 4.35 13.94 4.52 ;
      RECT 11.505 9.34 11.675 9.51 ;
      RECT 11.505 10.08 11.675 10.25 ;
      RECT 11.13 8.6 11.3 8.77 ;
    LAYER li1 ;
      RECT 93.78 7.305 93.95 8.775 ;
      RECT 93.78 8.6 93.955 8.77 ;
      RECT 93.41 3.035 93.58 4.225 ;
      RECT 93.41 3.035 93.88 3.205 ;
      RECT 93.41 9.255 93.88 9.425 ;
      RECT 93.41 8.235 93.58 9.425 ;
      RECT 92.42 3.035 92.59 4.225 ;
      RECT 92.42 3.035 92.89 3.205 ;
      RECT 92.42 9.255 92.89 9.425 ;
      RECT 92.42 8.235 92.59 9.425 ;
      RECT 90.57 3.93 90.74 5.16 ;
      RECT 90.625 2.15 90.795 4.1 ;
      RECT 90.57 1.87 90.74 2.32 ;
      RECT 90.57 10.14 90.74 10.59 ;
      RECT 90.625 8.36 90.795 10.31 ;
      RECT 90.57 7.3 90.74 8.53 ;
      RECT 90.05 1.87 90.22 5.16 ;
      RECT 90.05 3.37 90.455 3.7 ;
      RECT 90.05 2.53 90.455 2.86 ;
      RECT 90.05 7.3 90.22 10.59 ;
      RECT 90.05 9.6 90.455 9.93 ;
      RECT 90.05 8.76 90.455 9.09 ;
      RECT 87.35 3.13 87.52 3.4 ;
      RECT 87.35 3.13 88.08 3.3 ;
      RECT 87.27 4.52 87.6 4.69 ;
      RECT 86.51 4.35 87.52 4.52 ;
      RECT 86.51 3.87 86.68 4.52 ;
      RECT 86.63 3.79 86.8 4.12 ;
      RECT 85.79 4.52 86.12 4.69 ;
      RECT 83.87 4.52 85.16 4.69 ;
      RECT 84.91 4.435 86.04 4.605 ;
      RECT 85.63 3.51 86.04 3.68 ;
      RECT 85.87 3.05 86.04 3.68 ;
      RECT 84.435 7.3 84.605 10.59 ;
      RECT 84.435 9.6 84.84 9.93 ;
      RECT 84.435 8.76 84.84 9.09 ;
      RECT 83.11 3.87 84.44 4.04 ;
      RECT 84.19 3.79 84.36 4.04 ;
      RECT 83.19 3.47 83.36 3.68 ;
      RECT 83.19 3.47 83.68 3.64 ;
      RECT 81.87 4.63 82.16 4.8 ;
      RECT 81.87 3.87 82.04 4.8 ;
      RECT 81.67 3.87 82.04 4.04 ;
      RECT 80.67 3.87 81.16 4.04 ;
      RECT 80.99 3.79 81.16 4.04 ;
      RECT 80.75 4.63 81.16 4.8 ;
      RECT 80.99 4.44 81.16 4.8 ;
      RECT 79.79 4.35 80.44 4.52 ;
      RECT 79.79 3.79 79.96 4.52 ;
      RECT 79.43 4.91 79.72 5.08 ;
      RECT 79.43 3.87 79.6 5.08 ;
      RECT 79.23 3.87 79.6 4.04 ;
      RECT 77.455 7.305 77.625 8.775 ;
      RECT 77.455 8.6 77.63 8.77 ;
      RECT 77.085 3.035 77.255 4.225 ;
      RECT 77.085 3.035 77.555 3.205 ;
      RECT 77.085 9.255 77.555 9.425 ;
      RECT 77.085 8.235 77.255 9.425 ;
      RECT 76.095 3.035 76.265 4.225 ;
      RECT 76.095 3.035 76.565 3.205 ;
      RECT 76.095 9.255 76.565 9.425 ;
      RECT 76.095 8.235 76.265 9.425 ;
      RECT 74.245 3.93 74.415 5.16 ;
      RECT 74.3 2.15 74.47 4.1 ;
      RECT 74.245 1.87 74.415 2.32 ;
      RECT 74.245 10.14 74.415 10.59 ;
      RECT 74.3 8.36 74.47 10.31 ;
      RECT 74.245 7.3 74.415 8.53 ;
      RECT 73.725 1.87 73.895 5.16 ;
      RECT 73.725 3.37 74.13 3.7 ;
      RECT 73.725 2.53 74.13 2.86 ;
      RECT 73.725 7.3 73.895 10.59 ;
      RECT 73.725 9.6 74.13 9.93 ;
      RECT 73.725 8.76 74.13 9.09 ;
      RECT 71.025 3.13 71.195 3.4 ;
      RECT 71.025 3.13 71.755 3.3 ;
      RECT 70.945 4.52 71.275 4.69 ;
      RECT 70.185 4.35 71.195 4.52 ;
      RECT 70.185 3.87 70.355 4.52 ;
      RECT 70.305 3.79 70.475 4.12 ;
      RECT 69.465 4.52 69.795 4.69 ;
      RECT 67.545 4.52 68.835 4.69 ;
      RECT 68.585 4.435 69.715 4.605 ;
      RECT 69.305 3.51 69.715 3.68 ;
      RECT 69.545 3.05 69.715 3.68 ;
      RECT 68.11 7.3 68.28 10.59 ;
      RECT 68.11 9.6 68.515 9.93 ;
      RECT 68.11 8.76 68.515 9.09 ;
      RECT 66.785 3.87 68.115 4.04 ;
      RECT 67.865 3.79 68.035 4.04 ;
      RECT 66.865 3.47 67.035 3.68 ;
      RECT 66.865 3.47 67.355 3.64 ;
      RECT 65.545 4.63 65.835 4.8 ;
      RECT 65.545 3.87 65.715 4.8 ;
      RECT 65.345 3.87 65.715 4.04 ;
      RECT 64.345 3.87 64.835 4.04 ;
      RECT 64.665 3.79 64.835 4.04 ;
      RECT 64.425 4.63 64.835 4.8 ;
      RECT 64.665 4.44 64.835 4.8 ;
      RECT 63.465 4.35 64.115 4.52 ;
      RECT 63.465 3.79 63.635 4.52 ;
      RECT 63.105 4.91 63.395 5.08 ;
      RECT 63.105 3.87 63.275 5.08 ;
      RECT 62.905 3.87 63.275 4.04 ;
      RECT 61.13 7.305 61.3 8.775 ;
      RECT 61.13 8.6 61.305 8.77 ;
      RECT 60.76 3.035 60.93 4.225 ;
      RECT 60.76 3.035 61.23 3.205 ;
      RECT 60.76 9.255 61.23 9.425 ;
      RECT 60.76 8.235 60.93 9.425 ;
      RECT 59.77 3.035 59.94 4.225 ;
      RECT 59.77 3.035 60.24 3.205 ;
      RECT 59.77 9.255 60.24 9.425 ;
      RECT 59.77 8.235 59.94 9.425 ;
      RECT 57.92 3.93 58.09 5.16 ;
      RECT 57.975 2.15 58.145 4.1 ;
      RECT 57.92 1.87 58.09 2.32 ;
      RECT 57.92 10.14 58.09 10.59 ;
      RECT 57.975 8.36 58.145 10.31 ;
      RECT 57.92 7.3 58.09 8.53 ;
      RECT 57.4 1.87 57.57 5.16 ;
      RECT 57.4 3.37 57.805 3.7 ;
      RECT 57.4 2.53 57.805 2.86 ;
      RECT 57.4 7.3 57.57 10.59 ;
      RECT 57.4 9.6 57.805 9.93 ;
      RECT 57.4 8.76 57.805 9.09 ;
      RECT 54.7 3.13 54.87 3.4 ;
      RECT 54.7 3.13 55.43 3.3 ;
      RECT 54.62 4.52 54.95 4.69 ;
      RECT 53.86 4.35 54.87 4.52 ;
      RECT 53.86 3.87 54.03 4.52 ;
      RECT 53.98 3.79 54.15 4.12 ;
      RECT 53.14 4.52 53.47 4.69 ;
      RECT 51.22 4.52 52.51 4.69 ;
      RECT 52.26 4.435 53.39 4.605 ;
      RECT 52.98 3.51 53.39 3.68 ;
      RECT 53.22 3.05 53.39 3.68 ;
      RECT 51.785 7.3 51.955 10.59 ;
      RECT 51.785 9.6 52.19 9.93 ;
      RECT 51.785 8.76 52.19 9.09 ;
      RECT 50.46 3.87 51.79 4.04 ;
      RECT 51.54 3.79 51.71 4.04 ;
      RECT 50.54 3.47 50.71 3.68 ;
      RECT 50.54 3.47 51.03 3.64 ;
      RECT 49.22 4.63 49.51 4.8 ;
      RECT 49.22 3.87 49.39 4.8 ;
      RECT 49.02 3.87 49.39 4.04 ;
      RECT 48.02 3.87 48.51 4.04 ;
      RECT 48.34 3.79 48.51 4.04 ;
      RECT 48.1 4.63 48.51 4.8 ;
      RECT 48.34 4.44 48.51 4.8 ;
      RECT 47.14 4.35 47.79 4.52 ;
      RECT 47.14 3.79 47.31 4.52 ;
      RECT 46.78 4.91 47.07 5.08 ;
      RECT 46.78 3.87 46.95 5.08 ;
      RECT 46.58 3.87 46.95 4.04 ;
      RECT 44.805 7.305 44.975 8.775 ;
      RECT 44.805 8.6 44.98 8.77 ;
      RECT 44.435 3.035 44.605 4.225 ;
      RECT 44.435 3.035 44.905 3.205 ;
      RECT 44.435 9.255 44.905 9.425 ;
      RECT 44.435 8.235 44.605 9.425 ;
      RECT 43.445 3.035 43.615 4.225 ;
      RECT 43.445 3.035 43.915 3.205 ;
      RECT 43.445 9.255 43.915 9.425 ;
      RECT 43.445 8.235 43.615 9.425 ;
      RECT 41.595 3.93 41.765 5.16 ;
      RECT 41.65 2.15 41.82 4.1 ;
      RECT 41.595 1.87 41.765 2.32 ;
      RECT 41.595 10.14 41.765 10.59 ;
      RECT 41.65 8.36 41.82 10.31 ;
      RECT 41.595 7.3 41.765 8.53 ;
      RECT 41.075 1.87 41.245 5.16 ;
      RECT 41.075 3.37 41.48 3.7 ;
      RECT 41.075 2.53 41.48 2.86 ;
      RECT 41.075 7.3 41.245 10.59 ;
      RECT 41.075 9.6 41.48 9.93 ;
      RECT 41.075 8.76 41.48 9.09 ;
      RECT 38.375 3.13 38.545 3.4 ;
      RECT 38.375 3.13 39.105 3.3 ;
      RECT 38.295 4.52 38.625 4.69 ;
      RECT 37.535 4.35 38.545 4.52 ;
      RECT 37.535 3.87 37.705 4.52 ;
      RECT 37.655 3.79 37.825 4.12 ;
      RECT 36.815 4.52 37.145 4.69 ;
      RECT 34.895 4.52 36.185 4.69 ;
      RECT 35.935 4.435 37.065 4.605 ;
      RECT 36.655 3.51 37.065 3.68 ;
      RECT 36.895 3.05 37.065 3.68 ;
      RECT 35.46 7.3 35.63 10.59 ;
      RECT 35.46 9.6 35.865 9.93 ;
      RECT 35.46 8.76 35.865 9.09 ;
      RECT 34.135 3.87 35.465 4.04 ;
      RECT 35.215 3.79 35.385 4.04 ;
      RECT 34.215 3.47 34.385 3.68 ;
      RECT 34.215 3.47 34.705 3.64 ;
      RECT 32.895 4.63 33.185 4.8 ;
      RECT 32.895 3.87 33.065 4.8 ;
      RECT 32.695 3.87 33.065 4.04 ;
      RECT 31.695 3.87 32.185 4.04 ;
      RECT 32.015 3.79 32.185 4.04 ;
      RECT 31.775 4.63 32.185 4.8 ;
      RECT 32.015 4.44 32.185 4.8 ;
      RECT 30.815 4.35 31.465 4.52 ;
      RECT 30.815 3.79 30.985 4.52 ;
      RECT 30.455 4.91 30.745 5.08 ;
      RECT 30.455 3.87 30.625 5.08 ;
      RECT 30.255 3.87 30.625 4.04 ;
      RECT 28.48 7.305 28.65 8.775 ;
      RECT 28.48 8.6 28.655 8.77 ;
      RECT 28.11 3.035 28.28 4.225 ;
      RECT 28.11 3.035 28.58 3.205 ;
      RECT 28.11 9.255 28.58 9.425 ;
      RECT 28.11 8.235 28.28 9.425 ;
      RECT 27.12 3.035 27.29 4.225 ;
      RECT 27.12 3.035 27.59 3.205 ;
      RECT 27.12 9.255 27.59 9.425 ;
      RECT 27.12 8.235 27.29 9.425 ;
      RECT 25.27 3.93 25.44 5.16 ;
      RECT 25.325 2.15 25.495 4.1 ;
      RECT 25.27 1.87 25.44 2.32 ;
      RECT 25.27 10.14 25.44 10.59 ;
      RECT 25.325 8.36 25.495 10.31 ;
      RECT 25.27 7.3 25.44 8.53 ;
      RECT 24.75 1.87 24.92 5.16 ;
      RECT 24.75 3.37 25.155 3.7 ;
      RECT 24.75 2.53 25.155 2.86 ;
      RECT 24.75 7.3 24.92 10.59 ;
      RECT 24.75 9.6 25.155 9.93 ;
      RECT 24.75 8.76 25.155 9.09 ;
      RECT 22.05 3.13 22.22 3.4 ;
      RECT 22.05 3.13 22.78 3.3 ;
      RECT 21.97 4.52 22.3 4.69 ;
      RECT 21.21 4.35 22.22 4.52 ;
      RECT 21.21 3.87 21.38 4.52 ;
      RECT 21.33 3.79 21.5 4.12 ;
      RECT 20.49 4.52 20.82 4.69 ;
      RECT 18.57 4.52 19.86 4.69 ;
      RECT 19.61 4.435 20.74 4.605 ;
      RECT 20.33 3.51 20.74 3.68 ;
      RECT 20.57 3.05 20.74 3.68 ;
      RECT 19.135 7.3 19.305 10.59 ;
      RECT 19.135 9.6 19.54 9.93 ;
      RECT 19.135 8.76 19.54 9.09 ;
      RECT 17.81 3.87 19.14 4.04 ;
      RECT 18.89 3.79 19.06 4.04 ;
      RECT 17.89 3.47 18.06 3.68 ;
      RECT 17.89 3.47 18.38 3.64 ;
      RECT 16.57 4.63 16.86 4.8 ;
      RECT 16.57 3.87 16.74 4.8 ;
      RECT 16.37 3.87 16.74 4.04 ;
      RECT 15.37 3.87 15.86 4.04 ;
      RECT 15.69 3.79 15.86 4.04 ;
      RECT 15.45 4.63 15.86 4.8 ;
      RECT 15.69 4.44 15.86 4.8 ;
      RECT 14.49 4.35 15.14 4.52 ;
      RECT 14.49 3.79 14.66 4.52 ;
      RECT 14.13 4.91 14.42 5.08 ;
      RECT 14.13 3.87 14.3 5.08 ;
      RECT 13.93 3.87 14.3 4.04 ;
      RECT 11.075 10.14 11.245 10.59 ;
      RECT 11.13 8.36 11.3 10.31 ;
      RECT 11.075 7.3 11.245 8.53 ;
      RECT 10.555 7.3 10.725 10.59 ;
      RECT 10.555 9.6 10.96 9.93 ;
      RECT 10.555 8.76 10.96 9.09 ;
      RECT 93.78 10.085 93.95 10.595 ;
      RECT 92.79 1.865 92.96 2.375 ;
      RECT 92.79 3.685 92.96 5.155 ;
      RECT 92.79 7.305 92.96 8.775 ;
      RECT 92.79 10.085 92.96 10.595 ;
      RECT 91.43 1.87 91.6 5.16 ;
      RECT 91.43 7.3 91.6 10.59 ;
      RECT 91 1.87 91.17 2.38 ;
      RECT 91 2.95 91.17 5.16 ;
      RECT 91 7.3 91.17 9.51 ;
      RECT 91 10.08 91.17 10.59 ;
      RECT 87.11 3.79 87.28 4.12 ;
      RECT 86.39 3.05 86.56 3.4 ;
      RECT 86.39 4.78 86.56 5.11 ;
      RECT 85.815 7.3 85.985 10.59 ;
      RECT 85.39 4.78 85.56 5.11 ;
      RECT 85.385 7.3 85.555 9.51 ;
      RECT 85.385 10.08 85.555 10.59 ;
      RECT 85.15 3.79 85.32 4.24 ;
      RECT 84.67 3.79 84.84 4.12 ;
      RECT 83.95 3.05 84.12 3.4 ;
      RECT 82.95 4.44 83.12 4.8 ;
      RECT 82.71 3.79 82.88 4.24 ;
      RECT 82.23 3.79 82.4 4.12 ;
      RECT 81.99 3.05 82.16 3.4 ;
      RECT 81.51 4.35 81.68 4.77 ;
      RECT 80.51 3.05 80.68 3.4 ;
      RECT 80.27 3.79 80.44 4.12 ;
      RECT 79.55 3.05 79.72 3.4 ;
      RECT 79.07 4.35 79.24 4.77 ;
      RECT 77.455 10.085 77.625 10.595 ;
      RECT 76.465 1.865 76.635 2.375 ;
      RECT 76.465 3.685 76.635 5.155 ;
      RECT 76.465 7.305 76.635 8.775 ;
      RECT 76.465 10.085 76.635 10.595 ;
      RECT 75.105 1.87 75.275 5.16 ;
      RECT 75.105 7.3 75.275 10.59 ;
      RECT 74.675 1.87 74.845 2.38 ;
      RECT 74.675 2.95 74.845 5.16 ;
      RECT 74.675 7.3 74.845 9.51 ;
      RECT 74.675 10.08 74.845 10.59 ;
      RECT 70.785 3.79 70.955 4.12 ;
      RECT 70.065 3.05 70.235 3.4 ;
      RECT 70.065 4.78 70.235 5.11 ;
      RECT 69.49 7.3 69.66 10.59 ;
      RECT 69.065 4.78 69.235 5.11 ;
      RECT 69.06 7.3 69.23 9.51 ;
      RECT 69.06 10.08 69.23 10.59 ;
      RECT 68.825 3.79 68.995 4.24 ;
      RECT 68.345 3.79 68.515 4.12 ;
      RECT 67.625 3.05 67.795 3.4 ;
      RECT 66.625 4.44 66.795 4.8 ;
      RECT 66.385 3.79 66.555 4.24 ;
      RECT 65.905 3.79 66.075 4.12 ;
      RECT 65.665 3.05 65.835 3.4 ;
      RECT 65.185 4.35 65.355 4.77 ;
      RECT 64.185 3.05 64.355 3.4 ;
      RECT 63.945 3.79 64.115 4.12 ;
      RECT 63.225 3.05 63.395 3.4 ;
      RECT 62.745 4.35 62.915 4.77 ;
      RECT 61.13 10.085 61.3 10.595 ;
      RECT 60.14 1.865 60.31 2.375 ;
      RECT 60.14 3.685 60.31 5.155 ;
      RECT 60.14 7.305 60.31 8.775 ;
      RECT 60.14 10.085 60.31 10.595 ;
      RECT 58.78 1.87 58.95 5.16 ;
      RECT 58.78 7.3 58.95 10.59 ;
      RECT 58.35 1.87 58.52 2.38 ;
      RECT 58.35 2.95 58.52 5.16 ;
      RECT 58.35 7.3 58.52 9.51 ;
      RECT 58.35 10.08 58.52 10.59 ;
      RECT 54.46 3.79 54.63 4.12 ;
      RECT 53.74 3.05 53.91 3.4 ;
      RECT 53.74 4.78 53.91 5.11 ;
      RECT 53.165 7.3 53.335 10.59 ;
      RECT 52.74 4.78 52.91 5.11 ;
      RECT 52.735 7.3 52.905 9.51 ;
      RECT 52.735 10.08 52.905 10.59 ;
      RECT 52.5 3.79 52.67 4.24 ;
      RECT 52.02 3.79 52.19 4.12 ;
      RECT 51.3 3.05 51.47 3.4 ;
      RECT 50.3 4.44 50.47 4.8 ;
      RECT 50.06 3.79 50.23 4.24 ;
      RECT 49.58 3.79 49.75 4.12 ;
      RECT 49.34 3.05 49.51 3.4 ;
      RECT 48.86 4.35 49.03 4.77 ;
      RECT 47.86 3.05 48.03 3.4 ;
      RECT 47.62 3.79 47.79 4.12 ;
      RECT 46.9 3.05 47.07 3.4 ;
      RECT 46.42 4.35 46.59 4.77 ;
      RECT 44.805 10.085 44.975 10.595 ;
      RECT 43.815 1.865 43.985 2.375 ;
      RECT 43.815 3.685 43.985 5.155 ;
      RECT 43.815 7.305 43.985 8.775 ;
      RECT 43.815 10.085 43.985 10.595 ;
      RECT 42.455 1.87 42.625 5.16 ;
      RECT 42.455 7.3 42.625 10.59 ;
      RECT 42.025 1.87 42.195 2.38 ;
      RECT 42.025 2.95 42.195 5.16 ;
      RECT 42.025 7.3 42.195 9.51 ;
      RECT 42.025 10.08 42.195 10.59 ;
      RECT 38.135 3.79 38.305 4.12 ;
      RECT 37.415 3.05 37.585 3.4 ;
      RECT 37.415 4.78 37.585 5.11 ;
      RECT 36.84 7.3 37.01 10.59 ;
      RECT 36.415 4.78 36.585 5.11 ;
      RECT 36.41 7.3 36.58 9.51 ;
      RECT 36.41 10.08 36.58 10.59 ;
      RECT 36.175 3.79 36.345 4.24 ;
      RECT 35.695 3.79 35.865 4.12 ;
      RECT 34.975 3.05 35.145 3.4 ;
      RECT 33.975 4.44 34.145 4.8 ;
      RECT 33.735 3.79 33.905 4.24 ;
      RECT 33.255 3.79 33.425 4.12 ;
      RECT 33.015 3.05 33.185 3.4 ;
      RECT 32.535 4.35 32.705 4.77 ;
      RECT 31.535 3.05 31.705 3.4 ;
      RECT 31.295 3.79 31.465 4.12 ;
      RECT 30.575 3.05 30.745 3.4 ;
      RECT 30.095 4.35 30.265 4.77 ;
      RECT 28.48 10.085 28.65 10.595 ;
      RECT 27.49 1.865 27.66 2.375 ;
      RECT 27.49 3.685 27.66 5.155 ;
      RECT 27.49 7.305 27.66 8.775 ;
      RECT 27.49 10.085 27.66 10.595 ;
      RECT 26.13 1.87 26.3 5.16 ;
      RECT 26.13 7.3 26.3 10.59 ;
      RECT 25.7 1.87 25.87 2.38 ;
      RECT 25.7 2.95 25.87 5.16 ;
      RECT 25.7 7.3 25.87 9.51 ;
      RECT 25.7 10.08 25.87 10.59 ;
      RECT 21.81 3.79 21.98 4.12 ;
      RECT 21.09 3.05 21.26 3.4 ;
      RECT 21.09 4.78 21.26 5.11 ;
      RECT 20.515 7.3 20.685 10.59 ;
      RECT 20.09 4.78 20.26 5.11 ;
      RECT 20.085 7.3 20.255 9.51 ;
      RECT 20.085 10.08 20.255 10.59 ;
      RECT 19.85 3.79 20.02 4.24 ;
      RECT 19.37 3.79 19.54 4.12 ;
      RECT 18.65 3.05 18.82 3.4 ;
      RECT 17.65 4.44 17.82 4.8 ;
      RECT 17.41 3.79 17.58 4.24 ;
      RECT 16.93 3.79 17.1 4.12 ;
      RECT 16.69 3.05 16.86 3.4 ;
      RECT 16.21 4.35 16.38 4.77 ;
      RECT 15.21 3.05 15.38 3.4 ;
      RECT 14.97 3.79 15.14 4.12 ;
      RECT 14.25 3.05 14.42 3.4 ;
      RECT 13.77 4.35 13.94 4.77 ;
      RECT 11.505 7.3 11.675 9.51 ;
      RECT 11.505 10.08 11.675 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  ORIGIN -9.9 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r2 ;
  SIZE 84.425 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 28.48 2.21 28.65 2.38 ;
        RECT 28.475 2.205 28.645 2.375 ;
        RECT 28.475 3.685 28.645 3.855 ;
      LAYER li1 ;
        RECT 28.48 2.21 28.65 2.38 ;
        RECT 28.475 1.865 28.645 2.375 ;
        RECT 28.475 3.685 28.645 5.155 ;
      LAYER met1 ;
        RECT 28.415 3.655 28.705 3.885 ;
        RECT 28.415 2.175 28.705 2.405 ;
        RECT 28.475 2.175 28.645 3.885 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 44.805 2.21 44.975 2.38 ;
        RECT 44.8 2.205 44.97 2.375 ;
        RECT 44.8 3.685 44.97 3.855 ;
      LAYER li1 ;
        RECT 44.805 2.21 44.975 2.38 ;
        RECT 44.8 1.865 44.97 2.375 ;
        RECT 44.8 3.685 44.97 5.155 ;
      LAYER met1 ;
        RECT 44.74 3.655 45.03 3.885 ;
        RECT 44.74 2.175 45.03 2.405 ;
        RECT 44.8 2.175 44.97 3.885 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 61.13 2.21 61.3 2.38 ;
        RECT 61.125 2.205 61.295 2.375 ;
        RECT 61.125 3.685 61.295 3.855 ;
      LAYER li1 ;
        RECT 61.13 2.21 61.3 2.38 ;
        RECT 61.125 1.865 61.295 2.375 ;
        RECT 61.125 3.685 61.295 5.155 ;
      LAYER met1 ;
        RECT 61.065 3.655 61.355 3.885 ;
        RECT 61.065 2.175 61.355 2.405 ;
        RECT 61.125 2.175 61.295 3.885 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 77.455 2.21 77.625 2.38 ;
        RECT 77.45 2.205 77.62 2.375 ;
        RECT 77.45 3.685 77.62 3.855 ;
      LAYER li1 ;
        RECT 77.455 2.21 77.625 2.38 ;
        RECT 77.45 1.865 77.62 2.375 ;
        RECT 77.45 3.685 77.62 5.155 ;
      LAYER met1 ;
        RECT 77.39 3.655 77.68 3.885 ;
        RECT 77.39 2.175 77.68 2.405 ;
        RECT 77.45 2.175 77.62 3.885 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 93.78 2.21 93.95 2.38 ;
        RECT 93.775 2.205 93.945 2.375 ;
        RECT 93.775 3.685 93.945 3.855 ;
      LAYER li1 ;
        RECT 93.78 2.21 93.95 2.38 ;
        RECT 93.775 1.865 93.945 2.375 ;
        RECT 93.775 3.685 93.945 5.155 ;
      LAYER met1 ;
        RECT 93.715 3.655 94.005 3.885 ;
        RECT 93.715 2.175 94.005 2.405 ;
        RECT 93.775 2.175 93.945 3.885 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 24.325 2.955 24.495 4.23 ;
        RECT 24.325 8.23 24.495 9.505 ;
        RECT 18.71 8.23 18.88 9.505 ;
      LAYER met2 ;
        RECT 24.25 4 24.59 4.35 ;
        RECT 24.24 8.125 24.58 8.475 ;
        RECT 24.325 4 24.495 8.475 ;
      LAYER met1 ;
        RECT 24.25 4.06 24.725 4.23 ;
        RECT 24.25 4 24.59 4.35 ;
        RECT 18.65 8.23 24.725 8.4 ;
        RECT 24.24 8.125 24.58 8.475 ;
        RECT 18.65 8.2 18.94 8.43 ;
      LAYER via1 ;
        RECT 24.34 8.225 24.49 8.375 ;
        RECT 24.35 4.1 24.5 4.25 ;
      LAYER mcon ;
        RECT 18.71 8.23 18.88 8.4 ;
        RECT 24.325 8.23 24.495 8.4 ;
        RECT 24.325 4.06 24.495 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 40.65 2.955 40.82 4.23 ;
        RECT 40.65 8.23 40.82 9.505 ;
        RECT 35.035 8.23 35.205 9.505 ;
      LAYER met2 ;
        RECT 40.575 4 40.915 4.35 ;
        RECT 40.565 8.125 40.905 8.475 ;
        RECT 40.65 4 40.82 8.475 ;
      LAYER met1 ;
        RECT 40.575 4.06 41.05 4.23 ;
        RECT 40.575 4 40.915 4.35 ;
        RECT 34.975 8.23 41.05 8.4 ;
        RECT 40.565 8.125 40.905 8.475 ;
        RECT 34.975 8.2 35.265 8.43 ;
      LAYER via1 ;
        RECT 40.665 8.225 40.815 8.375 ;
        RECT 40.675 4.1 40.825 4.25 ;
      LAYER mcon ;
        RECT 35.035 8.23 35.205 8.4 ;
        RECT 40.65 8.23 40.82 8.4 ;
        RECT 40.65 4.06 40.82 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 56.975 2.955 57.145 4.23 ;
        RECT 56.975 8.23 57.145 9.505 ;
        RECT 51.36 8.23 51.53 9.505 ;
      LAYER met2 ;
        RECT 56.9 4 57.24 4.35 ;
        RECT 56.89 8.125 57.23 8.475 ;
        RECT 56.975 4 57.145 8.475 ;
      LAYER met1 ;
        RECT 56.9 4.06 57.375 4.23 ;
        RECT 56.9 4 57.24 4.35 ;
        RECT 51.3 8.23 57.375 8.4 ;
        RECT 56.89 8.125 57.23 8.475 ;
        RECT 51.3 8.2 51.59 8.43 ;
      LAYER via1 ;
        RECT 56.99 8.225 57.14 8.375 ;
        RECT 57 4.1 57.15 4.25 ;
      LAYER mcon ;
        RECT 51.36 8.23 51.53 8.4 ;
        RECT 56.975 8.23 57.145 8.4 ;
        RECT 56.975 4.06 57.145 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 73.3 2.955 73.47 4.23 ;
        RECT 73.3 8.23 73.47 9.505 ;
        RECT 67.685 8.23 67.855 9.505 ;
      LAYER met2 ;
        RECT 73.225 4 73.565 4.35 ;
        RECT 73.215 8.125 73.555 8.475 ;
        RECT 73.3 4 73.47 8.475 ;
      LAYER met1 ;
        RECT 73.225 4.06 73.7 4.23 ;
        RECT 73.225 4 73.565 4.35 ;
        RECT 67.625 8.23 73.7 8.4 ;
        RECT 73.215 8.125 73.555 8.475 ;
        RECT 67.625 8.2 67.915 8.43 ;
      LAYER via1 ;
        RECT 73.315 8.225 73.465 8.375 ;
        RECT 73.325 4.1 73.475 4.25 ;
      LAYER mcon ;
        RECT 67.685 8.23 67.855 8.4 ;
        RECT 73.3 8.23 73.47 8.4 ;
        RECT 73.3 4.06 73.47 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 89.625 2.955 89.795 4.23 ;
        RECT 89.625 8.23 89.795 9.505 ;
        RECT 84.01 8.23 84.18 9.505 ;
      LAYER met2 ;
        RECT 89.55 4 89.89 4.35 ;
        RECT 89.54 8.125 89.88 8.475 ;
        RECT 89.625 4 89.795 8.475 ;
      LAYER met1 ;
        RECT 89.55 4.06 90.025 4.23 ;
        RECT 89.55 4 89.89 4.35 ;
        RECT 83.95 8.23 90.025 8.4 ;
        RECT 89.54 8.125 89.88 8.475 ;
        RECT 83.95 8.2 84.24 8.43 ;
      LAYER via1 ;
        RECT 89.64 8.225 89.79 8.375 ;
        RECT 89.65 4.1 89.8 4.25 ;
      LAYER mcon ;
        RECT 84.01 8.23 84.18 8.4 ;
        RECT 89.625 8.23 89.795 8.4 ;
        RECT 89.625 4.06 89.795 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 10.13 8.23 10.3 9.505 ;
      LAYER met1 ;
        RECT 10.07 8.23 10.53 8.4 ;
        RECT 10.07 8.2 10.36 8.43 ;
      LAYER mcon ;
        RECT 10.13 8.23 10.3 8.4 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 9.9 5.435 94.32 7.035 ;
        RECT 12.69 5.43 94.32 7.035 ;
        RECT 92.185 5.425 94.165 7.035 ;
        RECT 93.345 4.695 93.515 7.765 ;
        RECT 92.355 4.695 92.525 7.765 ;
        RECT 89.615 4.7 89.785 7.76 ;
        RECT 78.735 5.33 88.395 7.035 ;
        RECT 87.825 4.83 87.995 7.035 ;
        RECT 86.865 4.83 87.035 7.035 ;
        RECT 84.425 4.83 84.595 7.035 ;
        RECT 84 5.33 84.17 7.76 ;
        RECT 83.425 4.83 83.595 7.035 ;
        RECT 82.465 4.83 82.635 7.035 ;
        RECT 80.025 4.83 80.195 7.035 ;
        RECT 75.86 5.425 77.84 7.035 ;
        RECT 77.02 4.695 77.19 7.765 ;
        RECT 76.03 4.695 76.2 7.765 ;
        RECT 73.29 4.7 73.46 7.76 ;
        RECT 62.41 5.33 72.07 7.035 ;
        RECT 71.5 4.83 71.67 7.035 ;
        RECT 70.54 4.83 70.71 7.035 ;
        RECT 68.1 4.83 68.27 7.035 ;
        RECT 67.675 5.33 67.845 7.76 ;
        RECT 67.1 4.83 67.27 7.035 ;
        RECT 66.14 4.83 66.31 7.035 ;
        RECT 63.7 4.83 63.87 7.035 ;
        RECT 59.535 5.425 61.515 7.035 ;
        RECT 60.695 4.695 60.865 7.765 ;
        RECT 59.705 4.695 59.875 7.765 ;
        RECT 56.965 4.7 57.135 7.76 ;
        RECT 46.085 5.33 55.745 7.035 ;
        RECT 55.175 4.83 55.345 7.035 ;
        RECT 54.215 4.83 54.385 7.035 ;
        RECT 51.775 4.83 51.945 7.035 ;
        RECT 51.35 5.33 51.52 7.76 ;
        RECT 50.775 4.83 50.945 7.035 ;
        RECT 49.815 4.83 49.985 7.035 ;
        RECT 47.375 4.83 47.545 7.035 ;
        RECT 43.21 5.425 45.19 7.035 ;
        RECT 44.37 4.695 44.54 7.765 ;
        RECT 43.38 4.695 43.55 7.765 ;
        RECT 40.64 4.7 40.81 7.76 ;
        RECT 29.76 5.33 39.42 7.035 ;
        RECT 38.85 4.83 39.02 7.035 ;
        RECT 37.89 4.83 38.06 7.035 ;
        RECT 35.45 4.83 35.62 7.035 ;
        RECT 35.025 5.33 35.195 7.76 ;
        RECT 34.45 4.83 34.62 7.035 ;
        RECT 33.49 4.83 33.66 7.035 ;
        RECT 31.05 4.83 31.22 7.035 ;
        RECT 26.885 5.425 28.865 7.035 ;
        RECT 28.045 4.695 28.215 7.765 ;
        RECT 27.055 4.695 27.225 7.765 ;
        RECT 24.315 4.7 24.485 7.76 ;
        RECT 13.435 5.33 23.095 7.035 ;
        RECT 22.525 4.83 22.695 7.035 ;
        RECT 21.565 4.83 21.735 7.035 ;
        RECT 19.125 4.83 19.295 7.035 ;
        RECT 18.7 5.33 18.87 7.76 ;
        RECT 18.125 4.83 18.295 7.035 ;
        RECT 17.165 4.83 17.335 7.035 ;
        RECT 14.725 4.83 14.895 7.035 ;
        RECT 11.93 5.435 12.1 10.59 ;
        RECT 10.12 5.435 10.29 7.76 ;
      LAYER met1 ;
        RECT 9.9 5.435 94.32 7.035 ;
        RECT 12.69 5.43 94.32 7.035 ;
        RECT 92.185 5.425 94.165 7.035 ;
        RECT 78.735 5.175 88.395 7.035 ;
        RECT 75.86 5.425 77.84 7.035 ;
        RECT 62.41 5.175 72.07 7.035 ;
        RECT 59.535 5.425 61.515 7.035 ;
        RECT 46.085 5.175 55.745 7.035 ;
        RECT 43.21 5.425 45.19 7.035 ;
        RECT 29.76 5.175 39.42 7.035 ;
        RECT 26.885 5.425 28.865 7.035 ;
        RECT 13.435 5.175 23.095 7.035 ;
        RECT 11.87 8.94 12.16 9.17 ;
        RECT 11.7 8.97 12.16 9.14 ;
      LAYER mcon ;
        RECT 11.93 8.97 12.1 9.14 ;
        RECT 12.24 6.83 12.41 7 ;
        RECT 13.58 5.33 13.75 5.5 ;
        RECT 14.04 5.33 14.21 5.5 ;
        RECT 14.5 5.33 14.67 5.5 ;
        RECT 14.96 5.33 15.13 5.5 ;
        RECT 15.42 5.33 15.59 5.5 ;
        RECT 15.88 5.33 16.05 5.5 ;
        RECT 16.34 5.33 16.51 5.5 ;
        RECT 16.8 5.33 16.97 5.5 ;
        RECT 17.26 5.33 17.43 5.5 ;
        RECT 17.72 5.33 17.89 5.5 ;
        RECT 18.18 5.33 18.35 5.5 ;
        RECT 18.64 5.33 18.81 5.5 ;
        RECT 19.1 5.33 19.27 5.5 ;
        RECT 19.56 5.33 19.73 5.5 ;
        RECT 20.02 5.33 20.19 5.5 ;
        RECT 20.48 5.33 20.65 5.5 ;
        RECT 20.82 6.83 20.99 7 ;
        RECT 20.94 5.33 21.11 5.5 ;
        RECT 21.4 5.33 21.57 5.5 ;
        RECT 21.86 5.33 22.03 5.5 ;
        RECT 22.32 5.33 22.49 5.5 ;
        RECT 22.78 5.33 22.95 5.5 ;
        RECT 26.435 6.83 26.605 7 ;
        RECT 26.435 5.46 26.605 5.63 ;
        RECT 27.135 6.835 27.305 7.005 ;
        RECT 27.135 5.455 27.305 5.625 ;
        RECT 28.125 6.835 28.295 7.005 ;
        RECT 28.125 5.455 28.295 5.625 ;
        RECT 29.905 5.33 30.075 5.5 ;
        RECT 30.365 5.33 30.535 5.5 ;
        RECT 30.825 5.33 30.995 5.5 ;
        RECT 31.285 5.33 31.455 5.5 ;
        RECT 31.745 5.33 31.915 5.5 ;
        RECT 32.205 5.33 32.375 5.5 ;
        RECT 32.665 5.33 32.835 5.5 ;
        RECT 33.125 5.33 33.295 5.5 ;
        RECT 33.585 5.33 33.755 5.5 ;
        RECT 34.045 5.33 34.215 5.5 ;
        RECT 34.505 5.33 34.675 5.5 ;
        RECT 34.965 5.33 35.135 5.5 ;
        RECT 35.425 5.33 35.595 5.5 ;
        RECT 35.885 5.33 36.055 5.5 ;
        RECT 36.345 5.33 36.515 5.5 ;
        RECT 36.805 5.33 36.975 5.5 ;
        RECT 37.145 6.83 37.315 7 ;
        RECT 37.265 5.33 37.435 5.5 ;
        RECT 37.725 5.33 37.895 5.5 ;
        RECT 38.185 5.33 38.355 5.5 ;
        RECT 38.645 5.33 38.815 5.5 ;
        RECT 39.105 5.33 39.275 5.5 ;
        RECT 42.76 6.83 42.93 7 ;
        RECT 42.76 5.46 42.93 5.63 ;
        RECT 43.46 6.835 43.63 7.005 ;
        RECT 43.46 5.455 43.63 5.625 ;
        RECT 44.45 6.835 44.62 7.005 ;
        RECT 44.45 5.455 44.62 5.625 ;
        RECT 46.23 5.33 46.4 5.5 ;
        RECT 46.69 5.33 46.86 5.5 ;
        RECT 47.15 5.33 47.32 5.5 ;
        RECT 47.61 5.33 47.78 5.5 ;
        RECT 48.07 5.33 48.24 5.5 ;
        RECT 48.53 5.33 48.7 5.5 ;
        RECT 48.99 5.33 49.16 5.5 ;
        RECT 49.45 5.33 49.62 5.5 ;
        RECT 49.91 5.33 50.08 5.5 ;
        RECT 50.37 5.33 50.54 5.5 ;
        RECT 50.83 5.33 51 5.5 ;
        RECT 51.29 5.33 51.46 5.5 ;
        RECT 51.75 5.33 51.92 5.5 ;
        RECT 52.21 5.33 52.38 5.5 ;
        RECT 52.67 5.33 52.84 5.5 ;
        RECT 53.13 5.33 53.3 5.5 ;
        RECT 53.47 6.83 53.64 7 ;
        RECT 53.59 5.33 53.76 5.5 ;
        RECT 54.05 5.33 54.22 5.5 ;
        RECT 54.51 5.33 54.68 5.5 ;
        RECT 54.97 5.33 55.14 5.5 ;
        RECT 55.43 5.33 55.6 5.5 ;
        RECT 59.085 6.83 59.255 7 ;
        RECT 59.085 5.46 59.255 5.63 ;
        RECT 59.785 6.835 59.955 7.005 ;
        RECT 59.785 5.455 59.955 5.625 ;
        RECT 60.775 6.835 60.945 7.005 ;
        RECT 60.775 5.455 60.945 5.625 ;
        RECT 62.555 5.33 62.725 5.5 ;
        RECT 63.015 5.33 63.185 5.5 ;
        RECT 63.475 5.33 63.645 5.5 ;
        RECT 63.935 5.33 64.105 5.5 ;
        RECT 64.395 5.33 64.565 5.5 ;
        RECT 64.855 5.33 65.025 5.5 ;
        RECT 65.315 5.33 65.485 5.5 ;
        RECT 65.775 5.33 65.945 5.5 ;
        RECT 66.235 5.33 66.405 5.5 ;
        RECT 66.695 5.33 66.865 5.5 ;
        RECT 67.155 5.33 67.325 5.5 ;
        RECT 67.615 5.33 67.785 5.5 ;
        RECT 68.075 5.33 68.245 5.5 ;
        RECT 68.535 5.33 68.705 5.5 ;
        RECT 68.995 5.33 69.165 5.5 ;
        RECT 69.455 5.33 69.625 5.5 ;
        RECT 69.795 6.83 69.965 7 ;
        RECT 69.915 5.33 70.085 5.5 ;
        RECT 70.375 5.33 70.545 5.5 ;
        RECT 70.835 5.33 71.005 5.5 ;
        RECT 71.295 5.33 71.465 5.5 ;
        RECT 71.755 5.33 71.925 5.5 ;
        RECT 75.41 6.83 75.58 7 ;
        RECT 75.41 5.46 75.58 5.63 ;
        RECT 76.11 6.835 76.28 7.005 ;
        RECT 76.11 5.455 76.28 5.625 ;
        RECT 77.1 6.835 77.27 7.005 ;
        RECT 77.1 5.455 77.27 5.625 ;
        RECT 78.88 5.33 79.05 5.5 ;
        RECT 79.34 5.33 79.51 5.5 ;
        RECT 79.8 5.33 79.97 5.5 ;
        RECT 80.26 5.33 80.43 5.5 ;
        RECT 80.72 5.33 80.89 5.5 ;
        RECT 81.18 5.33 81.35 5.5 ;
        RECT 81.64 5.33 81.81 5.5 ;
        RECT 82.1 5.33 82.27 5.5 ;
        RECT 82.56 5.33 82.73 5.5 ;
        RECT 83.02 5.33 83.19 5.5 ;
        RECT 83.48 5.33 83.65 5.5 ;
        RECT 83.94 5.33 84.11 5.5 ;
        RECT 84.4 5.33 84.57 5.5 ;
        RECT 84.86 5.33 85.03 5.5 ;
        RECT 85.32 5.33 85.49 5.5 ;
        RECT 85.78 5.33 85.95 5.5 ;
        RECT 86.12 6.83 86.29 7 ;
        RECT 86.24 5.33 86.41 5.5 ;
        RECT 86.7 5.33 86.87 5.5 ;
        RECT 87.16 5.33 87.33 5.5 ;
        RECT 87.62 5.33 87.79 5.5 ;
        RECT 88.08 5.33 88.25 5.5 ;
        RECT 91.735 6.83 91.905 7 ;
        RECT 91.735 5.46 91.905 5.63 ;
        RECT 92.435 6.835 92.605 7.005 ;
        RECT 92.435 5.455 92.605 5.625 ;
        RECT 93.425 6.835 93.595 7.005 ;
        RECT 93.425 5.455 93.595 5.625 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 85.3 9.34 85.67 9.71 ;
      RECT 85.3 9.375 87.285 9.675 ;
      RECT 86.985 3.575 87.285 9.675 ;
      RECT 83.985 3.21 84.315 3.94 ;
      RECT 83.105 3.21 83.435 3.94 ;
      RECT 86.185 3.575 87.285 3.875 ;
      RECT 83.105 3.575 85.245 3.875 ;
      RECT 84.945 3.26 85.245 3.875 ;
      RECT 87.145 3.045 87.475 3.775 ;
      RECT 86.185 3.275 86.49 3.875 ;
      RECT 84.945 3.26 86.305 3.57 ;
      RECT 83.605 4.73 83.935 5.06 ;
      RECT 82.4 4.745 83.935 5.045 ;
      RECT 82.4 3.625 82.7 5.045 ;
      RECT 82.145 3.61 82.475 3.94 ;
      RECT 68.975 9.34 69.345 9.71 ;
      RECT 68.975 9.375 70.96 9.675 ;
      RECT 70.66 3.575 70.96 9.675 ;
      RECT 67.66 3.21 67.99 3.94 ;
      RECT 66.78 3.21 67.11 3.94 ;
      RECT 69.86 3.575 70.96 3.875 ;
      RECT 66.78 3.575 68.92 3.875 ;
      RECT 68.62 3.26 68.92 3.875 ;
      RECT 70.82 3.045 71.15 3.775 ;
      RECT 69.86 3.275 70.165 3.875 ;
      RECT 68.62 3.26 69.98 3.57 ;
      RECT 67.28 4.73 67.61 5.06 ;
      RECT 66.075 4.745 67.61 5.045 ;
      RECT 66.075 3.625 66.375 5.045 ;
      RECT 65.82 3.61 66.15 3.94 ;
      RECT 52.65 9.34 53.02 9.71 ;
      RECT 52.65 9.375 54.635 9.675 ;
      RECT 54.335 3.575 54.635 9.675 ;
      RECT 51.335 3.21 51.665 3.94 ;
      RECT 50.455 3.21 50.785 3.94 ;
      RECT 53.535 3.575 54.635 3.875 ;
      RECT 50.455 3.575 52.595 3.875 ;
      RECT 52.295 3.26 52.595 3.875 ;
      RECT 54.495 3.045 54.825 3.775 ;
      RECT 53.535 3.275 53.84 3.875 ;
      RECT 52.295 3.26 53.655 3.57 ;
      RECT 50.955 4.73 51.285 5.06 ;
      RECT 49.75 4.745 51.285 5.045 ;
      RECT 49.75 3.625 50.05 5.045 ;
      RECT 49.495 3.61 49.825 3.94 ;
      RECT 36.325 9.34 36.695 9.71 ;
      RECT 36.325 9.375 38.31 9.675 ;
      RECT 38.01 3.575 38.31 9.675 ;
      RECT 35.01 3.21 35.34 3.94 ;
      RECT 34.13 3.21 34.46 3.94 ;
      RECT 37.21 3.575 38.31 3.875 ;
      RECT 34.13 3.575 36.27 3.875 ;
      RECT 35.97 3.26 36.27 3.875 ;
      RECT 38.17 3.045 38.5 3.775 ;
      RECT 37.21 3.275 37.515 3.875 ;
      RECT 35.97 3.26 37.33 3.57 ;
      RECT 34.63 4.73 34.96 5.06 ;
      RECT 33.425 4.745 34.96 5.045 ;
      RECT 33.425 3.625 33.725 5.045 ;
      RECT 33.17 3.61 33.5 3.94 ;
      RECT 20 9.34 20.37 9.71 ;
      RECT 20 9.375 21.985 9.675 ;
      RECT 21.685 3.575 21.985 9.675 ;
      RECT 18.685 3.21 19.015 3.94 ;
      RECT 17.805 3.21 18.135 3.94 ;
      RECT 20.885 3.575 21.985 3.875 ;
      RECT 17.805 3.575 19.945 3.875 ;
      RECT 19.645 3.26 19.945 3.875 ;
      RECT 21.845 3.045 22.175 3.775 ;
      RECT 20.885 3.275 21.19 3.875 ;
      RECT 19.645 3.26 21.005 3.57 ;
      RECT 18.305 4.73 18.635 5.06 ;
      RECT 17.1 4.745 18.635 5.045 ;
      RECT 17.1 3.625 17.4 5.045 ;
      RECT 16.845 3.61 17.175 3.94 ;
      RECT 87.625 4.17 87.955 4.9 ;
      RECT 85.545 3.77 85.875 4.5 ;
      RECT 81.425 3.61 81.755 4.34 ;
      RECT 80.425 3.05 80.755 3.78 ;
      RECT 78.985 3.77 79.315 4.5 ;
      RECT 71.3 4.17 71.63 4.9 ;
      RECT 69.22 3.77 69.55 4.5 ;
      RECT 65.1 3.61 65.43 4.34 ;
      RECT 64.1 3.05 64.43 3.78 ;
      RECT 62.66 3.77 62.99 4.5 ;
      RECT 54.975 4.17 55.305 4.9 ;
      RECT 52.895 3.77 53.225 4.5 ;
      RECT 48.775 3.61 49.105 4.34 ;
      RECT 47.775 3.05 48.105 3.78 ;
      RECT 46.335 3.77 46.665 4.5 ;
      RECT 38.65 4.17 38.98 4.9 ;
      RECT 36.57 3.77 36.9 4.5 ;
      RECT 32.45 3.61 32.78 4.34 ;
      RECT 31.45 3.05 31.78 3.78 ;
      RECT 30.01 3.77 30.34 4.5 ;
      RECT 22.325 4.17 22.655 4.9 ;
      RECT 20.245 3.77 20.575 4.5 ;
      RECT 16.125 3.61 16.455 4.34 ;
      RECT 15.125 3.05 15.455 3.78 ;
      RECT 13.685 3.77 14.015 4.5 ;
      RECT 9.905 10.785 10.71 11.165 ;
      RECT 9.9 0 10.705 0.38 ;
    LAYER via2 ;
      RECT 87.69 4.235 87.89 4.435 ;
      RECT 87.21 3.51 87.41 3.71 ;
      RECT 85.61 4.235 85.81 4.435 ;
      RECT 85.385 9.425 85.585 9.625 ;
      RECT 84.05 3.675 84.25 3.875 ;
      RECT 83.67 4.795 83.87 4.995 ;
      RECT 83.17 3.675 83.37 3.875 ;
      RECT 82.21 3.675 82.41 3.875 ;
      RECT 81.49 3.675 81.69 3.875 ;
      RECT 80.49 3.115 80.69 3.315 ;
      RECT 79.05 4.235 79.25 4.435 ;
      RECT 71.365 4.235 71.565 4.435 ;
      RECT 70.885 3.51 71.085 3.71 ;
      RECT 69.285 4.235 69.485 4.435 ;
      RECT 69.06 9.425 69.26 9.625 ;
      RECT 67.725 3.675 67.925 3.875 ;
      RECT 67.345 4.795 67.545 4.995 ;
      RECT 66.845 3.675 67.045 3.875 ;
      RECT 65.885 3.675 66.085 3.875 ;
      RECT 65.165 3.675 65.365 3.875 ;
      RECT 64.165 3.115 64.365 3.315 ;
      RECT 62.725 4.235 62.925 4.435 ;
      RECT 55.04 4.235 55.24 4.435 ;
      RECT 54.56 3.51 54.76 3.71 ;
      RECT 52.96 4.235 53.16 4.435 ;
      RECT 52.735 9.425 52.935 9.625 ;
      RECT 51.4 3.675 51.6 3.875 ;
      RECT 51.02 4.795 51.22 4.995 ;
      RECT 50.52 3.675 50.72 3.875 ;
      RECT 49.56 3.675 49.76 3.875 ;
      RECT 48.84 3.675 49.04 3.875 ;
      RECT 47.84 3.115 48.04 3.315 ;
      RECT 46.4 4.235 46.6 4.435 ;
      RECT 38.715 4.235 38.915 4.435 ;
      RECT 38.235 3.51 38.435 3.71 ;
      RECT 36.635 4.235 36.835 4.435 ;
      RECT 36.41 9.425 36.61 9.625 ;
      RECT 35.075 3.675 35.275 3.875 ;
      RECT 34.695 4.795 34.895 4.995 ;
      RECT 34.195 3.675 34.395 3.875 ;
      RECT 33.235 3.675 33.435 3.875 ;
      RECT 32.515 3.675 32.715 3.875 ;
      RECT 31.515 3.115 31.715 3.315 ;
      RECT 30.075 4.235 30.275 4.435 ;
      RECT 22.39 4.235 22.59 4.435 ;
      RECT 21.91 3.51 22.11 3.71 ;
      RECT 20.31 4.235 20.51 4.435 ;
      RECT 20.085 9.425 20.285 9.625 ;
      RECT 18.75 3.675 18.95 3.875 ;
      RECT 18.37 4.795 18.57 4.995 ;
      RECT 17.87 3.675 18.07 3.875 ;
      RECT 16.91 3.675 17.11 3.875 ;
      RECT 16.19 3.675 16.39 3.875 ;
      RECT 15.19 3.115 15.39 3.315 ;
      RECT 13.75 4.235 13.95 4.435 ;
      RECT 10.185 10.875 10.385 11.075 ;
      RECT 10.18 0.09 10.38 0.29 ;
    LAYER met2 ;
      RECT 11.125 10.685 93.95 10.855 ;
      RECT 93.78 9.56 93.95 10.855 ;
      RECT 11.125 8.54 11.295 10.855 ;
      RECT 93.75 9.56 94.1 9.91 ;
      RECT 11.065 8.54 11.355 8.89 ;
      RECT 90.59 8.505 90.91 8.83 ;
      RECT 90.62 7.98 90.79 8.83 ;
      RECT 90.62 7.98 90.795 8.33 ;
      RECT 90.62 7.98 91.595 8.155 ;
      RECT 91.42 3.26 91.595 8.155 ;
      RECT 91.365 3.26 91.715 3.61 ;
      RECT 91.39 8.94 91.715 9.265 ;
      RECT 90.275 9.03 91.715 9.2 ;
      RECT 90.275 3.69 90.435 9.2 ;
      RECT 90.59 3.66 90.91 3.98 ;
      RECT 90.275 3.69 90.91 3.86 ;
      RECT 79.01 4.15 79.29 4.52 ;
      RECT 79.065 2.585 79.235 4.52 ;
      RECT 89.06 2.585 89.23 3.11 ;
      RECT 88.97 2.755 89.31 3.105 ;
      RECT 79.065 2.585 89.23 2.755 ;
      RECT 85.69 3.59 85.97 3.96 ;
      RECT 84.62 3.615 84.88 3.935 ;
      RECT 87.17 3.425 87.45 3.795 ;
      RECT 87.78 3.335 88.04 3.655 ;
      RECT 84.68 2.775 84.82 3.935 ;
      RECT 85.76 2.775 85.9 3.96 ;
      RECT 86.88 3.425 88.04 3.565 ;
      RECT 86.88 2.775 87.02 3.565 ;
      RECT 84.68 2.775 87.02 2.915 ;
      RECT 87.65 4.15 87.93 4.52 ;
      RECT 87.66 3.895 87.92 4.52 ;
      RECT 84.71 4.915 86.885 5.08 ;
      RECT 86.74 3.795 86.885 5.08 ;
      RECT 83.63 4.71 83.91 5.08 ;
      RECT 83.63 4.825 84.85 4.965 ;
      RECT 86.46 3.795 86.885 3.935 ;
      RECT 86.46 3.615 86.72 3.935 ;
      RECT 79.8 5.195 83.46 5.335 ;
      RECT 83.32 4.38 83.46 5.335 ;
      RECT 79.8 4.265 79.94 5.335 ;
      RECT 86.34 4.455 86.6 4.775 ;
      RECT 83.32 4.38 85.85 4.52 ;
      RECT 85.57 4.15 85.85 4.52 ;
      RECT 79.8 4.265 80.25 4.52 ;
      RECT 79.97 4.15 80.25 4.52 ;
      RECT 86.34 4.265 86.54 4.775 ;
      RECT 85.57 4.265 86.54 4.405 ;
      RECT 86.14 3.055 86.28 4.405 ;
      RECT 86.08 3.055 86.34 3.375 ;
      RECT 77.4 8.94 77.75 9.29 ;
      RECT 85.955 8.895 86.305 9.245 ;
      RECT 77.4 8.97 86.305 9.17 ;
      RECT 79.98 3.615 80.24 3.935 ;
      RECT 79.98 3.705 81.02 3.845 ;
      RECT 80.88 2.915 81.02 3.845 ;
      RECT 83.64 3.055 83.9 3.375 ;
      RECT 80.88 2.915 83.84 3.055 ;
      RECT 83.02 3.895 83.28 4.215 ;
      RECT 83.02 3.895 83.34 4.125 ;
      RECT 83.13 3.59 83.41 3.96 ;
      RECT 82.72 4.455 83.04 4.775 ;
      RECT 82.72 3.335 82.86 4.775 ;
      RECT 82.66 3.335 82.92 3.655 ;
      RECT 80.22 4.735 80.48 5.055 ;
      RECT 80.22 4.825 81.9 4.965 ;
      RECT 81.76 4.545 81.9 4.965 ;
      RECT 81.76 4.545 82.2 4.775 ;
      RECT 81.94 4.455 82.2 4.775 ;
      RECT 81.26 3.615 81.66 4.125 ;
      RECT 81.45 3.59 81.73 3.96 ;
      RECT 81.2 3.615 81.73 3.935 ;
      RECT 74.265 8.505 74.585 8.83 ;
      RECT 74.295 7.98 74.465 8.83 ;
      RECT 74.295 7.98 74.47 8.33 ;
      RECT 74.295 7.98 75.27 8.155 ;
      RECT 75.095 3.26 75.27 8.155 ;
      RECT 75.04 3.26 75.39 3.61 ;
      RECT 75.065 8.94 75.39 9.265 ;
      RECT 73.95 9.03 75.39 9.2 ;
      RECT 73.95 3.69 74.11 9.2 ;
      RECT 74.265 3.66 74.585 3.98 ;
      RECT 73.95 3.69 74.585 3.86 ;
      RECT 62.685 4.15 62.965 4.52 ;
      RECT 62.74 2.585 62.91 4.52 ;
      RECT 72.735 2.585 72.905 3.11 ;
      RECT 72.645 2.755 72.985 3.105 ;
      RECT 62.74 2.585 72.905 2.755 ;
      RECT 69.365 3.59 69.645 3.96 ;
      RECT 68.295 3.615 68.555 3.935 ;
      RECT 70.845 3.425 71.125 3.795 ;
      RECT 71.455 3.335 71.715 3.655 ;
      RECT 68.355 2.775 68.495 3.935 ;
      RECT 69.435 2.775 69.575 3.96 ;
      RECT 70.555 3.425 71.715 3.565 ;
      RECT 70.555 2.775 70.695 3.565 ;
      RECT 68.355 2.775 70.695 2.915 ;
      RECT 71.325 4.15 71.605 4.52 ;
      RECT 71.335 3.895 71.595 4.52 ;
      RECT 68.385 4.915 70.56 5.08 ;
      RECT 70.415 3.795 70.56 5.08 ;
      RECT 67.305 4.71 67.585 5.08 ;
      RECT 67.305 4.825 68.525 4.965 ;
      RECT 70.135 3.795 70.56 3.935 ;
      RECT 70.135 3.615 70.395 3.935 ;
      RECT 63.475 5.195 67.135 5.335 ;
      RECT 66.995 4.38 67.135 5.335 ;
      RECT 63.475 4.265 63.615 5.335 ;
      RECT 70.015 4.455 70.275 4.775 ;
      RECT 66.995 4.38 69.525 4.52 ;
      RECT 69.245 4.15 69.525 4.52 ;
      RECT 63.475 4.265 63.925 4.52 ;
      RECT 63.645 4.15 63.925 4.52 ;
      RECT 70.015 4.265 70.215 4.775 ;
      RECT 69.245 4.265 70.215 4.405 ;
      RECT 69.815 3.055 69.955 4.405 ;
      RECT 69.755 3.055 70.015 3.375 ;
      RECT 61.075 8.94 61.425 9.29 ;
      RECT 69.625 8.895 69.975 9.245 ;
      RECT 61.075 8.97 69.975 9.17 ;
      RECT 63.655 3.615 63.915 3.935 ;
      RECT 63.655 3.705 64.695 3.845 ;
      RECT 64.555 2.915 64.695 3.845 ;
      RECT 67.315 3.055 67.575 3.375 ;
      RECT 64.555 2.915 67.515 3.055 ;
      RECT 66.695 3.895 66.955 4.215 ;
      RECT 66.695 3.895 67.015 4.125 ;
      RECT 66.805 3.59 67.085 3.96 ;
      RECT 66.395 4.455 66.715 4.775 ;
      RECT 66.395 3.335 66.535 4.775 ;
      RECT 66.335 3.335 66.595 3.655 ;
      RECT 63.895 4.735 64.155 5.055 ;
      RECT 63.895 4.825 65.575 4.965 ;
      RECT 65.435 4.545 65.575 4.965 ;
      RECT 65.435 4.545 65.875 4.775 ;
      RECT 65.615 4.455 65.875 4.775 ;
      RECT 64.935 3.615 65.335 4.125 ;
      RECT 65.125 3.59 65.405 3.96 ;
      RECT 64.875 3.615 65.405 3.935 ;
      RECT 57.94 8.505 58.26 8.83 ;
      RECT 57.97 7.98 58.14 8.83 ;
      RECT 57.97 7.98 58.145 8.33 ;
      RECT 57.97 7.98 58.945 8.155 ;
      RECT 58.77 3.26 58.945 8.155 ;
      RECT 58.715 3.26 59.065 3.61 ;
      RECT 58.74 8.94 59.065 9.265 ;
      RECT 57.625 9.03 59.065 9.2 ;
      RECT 57.625 3.69 57.785 9.2 ;
      RECT 57.94 3.66 58.26 3.98 ;
      RECT 57.625 3.69 58.26 3.86 ;
      RECT 46.36 4.15 46.64 4.52 ;
      RECT 46.415 2.585 46.585 4.52 ;
      RECT 56.41 2.585 56.58 3.11 ;
      RECT 56.32 2.755 56.66 3.105 ;
      RECT 46.415 2.585 56.58 2.755 ;
      RECT 53.04 3.59 53.32 3.96 ;
      RECT 51.97 3.615 52.23 3.935 ;
      RECT 54.52 3.425 54.8 3.795 ;
      RECT 55.13 3.335 55.39 3.655 ;
      RECT 52.03 2.775 52.17 3.935 ;
      RECT 53.11 2.775 53.25 3.96 ;
      RECT 54.23 3.425 55.39 3.565 ;
      RECT 54.23 2.775 54.37 3.565 ;
      RECT 52.03 2.775 54.37 2.915 ;
      RECT 55 4.15 55.28 4.52 ;
      RECT 55.01 3.895 55.27 4.52 ;
      RECT 52.06 4.915 54.235 5.08 ;
      RECT 54.09 3.795 54.235 5.08 ;
      RECT 50.98 4.71 51.26 5.08 ;
      RECT 50.98 4.825 52.2 4.965 ;
      RECT 53.81 3.795 54.235 3.935 ;
      RECT 53.81 3.615 54.07 3.935 ;
      RECT 47.15 5.195 50.81 5.335 ;
      RECT 50.67 4.38 50.81 5.335 ;
      RECT 47.15 4.265 47.29 5.335 ;
      RECT 53.69 4.455 53.95 4.775 ;
      RECT 50.67 4.38 53.2 4.52 ;
      RECT 52.92 4.15 53.2 4.52 ;
      RECT 47.15 4.265 47.6 4.52 ;
      RECT 47.32 4.15 47.6 4.52 ;
      RECT 53.69 4.265 53.89 4.775 ;
      RECT 52.92 4.265 53.89 4.405 ;
      RECT 53.49 3.055 53.63 4.405 ;
      RECT 53.43 3.055 53.69 3.375 ;
      RECT 44.795 8.945 45.145 9.295 ;
      RECT 53.3 8.9 53.65 9.25 ;
      RECT 44.795 8.975 53.65 9.175 ;
      RECT 47.33 3.615 47.59 3.935 ;
      RECT 47.33 3.705 48.37 3.845 ;
      RECT 48.23 2.915 48.37 3.845 ;
      RECT 50.99 3.055 51.25 3.375 ;
      RECT 48.23 2.915 51.19 3.055 ;
      RECT 50.37 3.895 50.63 4.215 ;
      RECT 50.37 3.895 50.69 4.125 ;
      RECT 50.48 3.59 50.76 3.96 ;
      RECT 50.07 4.455 50.39 4.775 ;
      RECT 50.07 3.335 50.21 4.775 ;
      RECT 50.01 3.335 50.27 3.655 ;
      RECT 47.57 4.735 47.83 5.055 ;
      RECT 47.57 4.825 49.25 4.965 ;
      RECT 49.11 4.545 49.25 4.965 ;
      RECT 49.11 4.545 49.55 4.775 ;
      RECT 49.29 4.455 49.55 4.775 ;
      RECT 48.61 3.615 49.01 4.125 ;
      RECT 48.8 3.59 49.08 3.96 ;
      RECT 48.55 3.615 49.08 3.935 ;
      RECT 41.615 8.505 41.935 8.83 ;
      RECT 41.645 7.98 41.815 8.83 ;
      RECT 41.645 7.98 41.82 8.33 ;
      RECT 41.645 7.98 42.62 8.155 ;
      RECT 42.445 3.26 42.62 8.155 ;
      RECT 42.39 3.26 42.74 3.61 ;
      RECT 42.415 8.94 42.74 9.265 ;
      RECT 41.3 9.03 42.74 9.2 ;
      RECT 41.3 3.69 41.46 9.2 ;
      RECT 41.615 3.66 41.935 3.98 ;
      RECT 41.3 3.69 41.935 3.86 ;
      RECT 30.035 4.15 30.315 4.52 ;
      RECT 30.09 2.585 30.26 4.52 ;
      RECT 40.085 2.585 40.255 3.11 ;
      RECT 39.995 2.755 40.335 3.105 ;
      RECT 30.09 2.585 40.255 2.755 ;
      RECT 36.715 3.59 36.995 3.96 ;
      RECT 35.645 3.615 35.905 3.935 ;
      RECT 38.195 3.425 38.475 3.795 ;
      RECT 38.805 3.335 39.065 3.655 ;
      RECT 35.705 2.775 35.845 3.935 ;
      RECT 36.785 2.775 36.925 3.96 ;
      RECT 37.905 3.425 39.065 3.565 ;
      RECT 37.905 2.775 38.045 3.565 ;
      RECT 35.705 2.775 38.045 2.915 ;
      RECT 38.675 4.15 38.955 4.52 ;
      RECT 38.685 3.895 38.945 4.52 ;
      RECT 35.735 4.915 37.91 5.08 ;
      RECT 37.765 3.795 37.91 5.08 ;
      RECT 34.655 4.71 34.935 5.08 ;
      RECT 34.655 4.825 35.875 4.965 ;
      RECT 37.485 3.795 37.91 3.935 ;
      RECT 37.485 3.615 37.745 3.935 ;
      RECT 30.825 5.195 34.485 5.335 ;
      RECT 34.345 4.38 34.485 5.335 ;
      RECT 30.825 4.265 30.965 5.335 ;
      RECT 37.365 4.455 37.625 4.775 ;
      RECT 34.345 4.38 36.875 4.52 ;
      RECT 36.595 4.15 36.875 4.52 ;
      RECT 30.825 4.265 31.275 4.52 ;
      RECT 30.995 4.15 31.275 4.52 ;
      RECT 37.365 4.265 37.565 4.775 ;
      RECT 36.595 4.265 37.565 4.405 ;
      RECT 37.165 3.055 37.305 4.405 ;
      RECT 37.105 3.055 37.365 3.375 ;
      RECT 28.47 8.94 28.82 9.29 ;
      RECT 36.975 8.895 37.325 9.245 ;
      RECT 28.47 8.97 37.325 9.17 ;
      RECT 31.005 3.615 31.265 3.935 ;
      RECT 31.005 3.705 32.045 3.845 ;
      RECT 31.905 2.915 32.045 3.845 ;
      RECT 34.665 3.055 34.925 3.375 ;
      RECT 31.905 2.915 34.865 3.055 ;
      RECT 34.045 3.895 34.305 4.215 ;
      RECT 34.045 3.895 34.365 4.125 ;
      RECT 34.155 3.59 34.435 3.96 ;
      RECT 33.745 4.455 34.065 4.775 ;
      RECT 33.745 3.335 33.885 4.775 ;
      RECT 33.685 3.335 33.945 3.655 ;
      RECT 31.245 4.735 31.505 5.055 ;
      RECT 31.245 4.825 32.925 4.965 ;
      RECT 32.785 4.545 32.925 4.965 ;
      RECT 32.785 4.545 33.225 4.775 ;
      RECT 32.965 4.455 33.225 4.775 ;
      RECT 32.285 3.615 32.685 4.125 ;
      RECT 32.475 3.59 32.755 3.96 ;
      RECT 32.225 3.615 32.755 3.935 ;
      RECT 25.29 8.505 25.61 8.83 ;
      RECT 25.32 7.98 25.49 8.83 ;
      RECT 25.32 7.98 25.495 8.33 ;
      RECT 25.32 7.98 26.295 8.155 ;
      RECT 26.12 3.26 26.295 8.155 ;
      RECT 26.065 3.26 26.415 3.61 ;
      RECT 26.09 8.94 26.415 9.265 ;
      RECT 24.975 9.03 26.415 9.2 ;
      RECT 24.975 3.69 25.135 9.2 ;
      RECT 25.29 3.66 25.61 3.98 ;
      RECT 24.975 3.69 25.61 3.86 ;
      RECT 13.71 4.15 13.99 4.52 ;
      RECT 13.765 2.585 13.935 4.52 ;
      RECT 23.76 2.585 23.93 3.11 ;
      RECT 23.67 2.755 24.01 3.105 ;
      RECT 13.765 2.585 23.93 2.755 ;
      RECT 20.39 3.59 20.67 3.96 ;
      RECT 19.32 3.615 19.58 3.935 ;
      RECT 21.87 3.425 22.15 3.795 ;
      RECT 22.48 3.335 22.74 3.655 ;
      RECT 19.38 2.775 19.52 3.935 ;
      RECT 20.46 2.775 20.6 3.96 ;
      RECT 21.58 3.425 22.74 3.565 ;
      RECT 21.58 2.775 21.72 3.565 ;
      RECT 19.38 2.775 21.72 2.915 ;
      RECT 22.35 4.15 22.63 4.52 ;
      RECT 22.36 3.895 22.62 4.52 ;
      RECT 11.44 9.28 11.73 9.63 ;
      RECT 11.44 9.335 12.78 9.505 ;
      RECT 12.61 8.97 12.78 9.505 ;
      RECT 21.485 8.89 21.835 9.24 ;
      RECT 12.61 8.97 21.835 9.14 ;
      RECT 19.41 4.915 21.585 5.08 ;
      RECT 21.44 3.795 21.585 5.08 ;
      RECT 18.33 4.71 18.61 5.08 ;
      RECT 18.33 4.825 19.55 4.965 ;
      RECT 21.16 3.795 21.585 3.935 ;
      RECT 21.16 3.615 21.42 3.935 ;
      RECT 14.5 5.195 18.16 5.335 ;
      RECT 18.02 4.38 18.16 5.335 ;
      RECT 14.5 4.265 14.64 5.335 ;
      RECT 21.04 4.455 21.3 4.775 ;
      RECT 18.02 4.38 20.55 4.52 ;
      RECT 20.27 4.15 20.55 4.52 ;
      RECT 14.5 4.265 14.95 4.52 ;
      RECT 14.67 4.15 14.95 4.52 ;
      RECT 21.04 4.265 21.24 4.775 ;
      RECT 20.27 4.265 21.24 4.405 ;
      RECT 20.84 3.055 20.98 4.405 ;
      RECT 20.78 3.055 21.04 3.375 ;
      RECT 14.68 3.615 14.94 3.935 ;
      RECT 14.68 3.705 15.72 3.845 ;
      RECT 15.58 2.915 15.72 3.845 ;
      RECT 18.34 3.055 18.6 3.375 ;
      RECT 15.58 2.915 18.54 3.055 ;
      RECT 17.72 3.895 17.98 4.215 ;
      RECT 17.72 3.895 18.04 4.125 ;
      RECT 17.83 3.59 18.11 3.96 ;
      RECT 17.42 4.455 17.74 4.775 ;
      RECT 17.42 3.335 17.56 4.775 ;
      RECT 17.36 3.335 17.62 3.655 ;
      RECT 14.92 4.735 15.18 5.055 ;
      RECT 14.92 4.825 16.6 4.965 ;
      RECT 16.46 4.545 16.6 4.965 ;
      RECT 16.46 4.545 16.9 4.775 ;
      RECT 16.64 4.455 16.9 4.775 ;
      RECT 15.96 3.615 16.36 4.125 ;
      RECT 16.15 3.59 16.43 3.96 ;
      RECT 15.9 3.615 16.43 3.935 ;
      RECT 10.095 10.785 10.475 11.165 ;
      RECT 10.135 0 10.275 11.165 ;
      RECT 10.09 0 10.47 0.38 ;
      RECT 85.3 9.34 85.67 9.71 ;
      RECT 84.01 3.59 84.29 3.96 ;
      RECT 82.17 3.59 82.45 3.96 ;
      RECT 80.45 3.03 80.73 3.4 ;
      RECT 68.975 9.34 69.345 9.71 ;
      RECT 67.685 3.59 67.965 3.96 ;
      RECT 65.845 3.59 66.125 3.96 ;
      RECT 64.125 3.03 64.405 3.4 ;
      RECT 52.65 9.34 53.02 9.71 ;
      RECT 51.36 3.59 51.64 3.96 ;
      RECT 49.52 3.59 49.8 3.96 ;
      RECT 47.8 3.03 48.08 3.4 ;
      RECT 36.325 9.34 36.695 9.71 ;
      RECT 35.035 3.59 35.315 3.96 ;
      RECT 33.195 3.59 33.475 3.96 ;
      RECT 31.475 3.03 31.755 3.4 ;
      RECT 20 9.34 20.37 9.71 ;
      RECT 18.71 3.59 18.99 3.96 ;
      RECT 16.87 3.59 17.15 3.96 ;
      RECT 15.15 3.03 15.43 3.4 ;
    LAYER via1 ;
      RECT 93.85 9.66 94 9.81 ;
      RECT 91.48 9.025 91.63 9.175 ;
      RECT 91.465 3.36 91.615 3.51 ;
      RECT 90.675 3.745 90.825 3.895 ;
      RECT 90.675 8.61 90.825 8.76 ;
      RECT 89.07 2.855 89.22 3.005 ;
      RECT 87.835 3.42 87.985 3.57 ;
      RECT 87.715 3.98 87.865 4.13 ;
      RECT 86.515 3.7 86.665 3.85 ;
      RECT 86.395 4.54 86.545 4.69 ;
      RECT 86.135 3.14 86.285 3.29 ;
      RECT 86.055 8.995 86.205 9.145 ;
      RECT 85.41 9.45 85.56 9.6 ;
      RECT 84.675 3.7 84.825 3.85 ;
      RECT 84.075 3.7 84.225 3.85 ;
      RECT 83.695 3.14 83.845 3.29 ;
      RECT 83.075 3.98 83.225 4.13 ;
      RECT 82.835 4.54 82.985 4.69 ;
      RECT 82.715 3.42 82.865 3.57 ;
      RECT 82.235 3.7 82.385 3.85 ;
      RECT 81.995 4.54 82.145 4.69 ;
      RECT 81.255 3.7 81.405 3.85 ;
      RECT 80.515 3.14 80.665 3.29 ;
      RECT 80.275 4.82 80.425 4.97 ;
      RECT 80.035 3.7 80.185 3.85 ;
      RECT 80.035 4.26 80.185 4.41 ;
      RECT 79.075 4.26 79.225 4.41 ;
      RECT 77.5 9.04 77.65 9.19 ;
      RECT 75.155 9.025 75.305 9.175 ;
      RECT 75.14 3.36 75.29 3.51 ;
      RECT 74.35 3.745 74.5 3.895 ;
      RECT 74.35 8.61 74.5 8.76 ;
      RECT 72.745 2.855 72.895 3.005 ;
      RECT 71.51 3.42 71.66 3.57 ;
      RECT 71.39 3.98 71.54 4.13 ;
      RECT 70.19 3.7 70.34 3.85 ;
      RECT 70.07 4.54 70.22 4.69 ;
      RECT 69.81 3.14 69.96 3.29 ;
      RECT 69.725 8.995 69.875 9.145 ;
      RECT 69.085 9.45 69.235 9.6 ;
      RECT 68.35 3.7 68.5 3.85 ;
      RECT 67.75 3.7 67.9 3.85 ;
      RECT 67.37 3.14 67.52 3.29 ;
      RECT 66.75 3.98 66.9 4.13 ;
      RECT 66.51 4.54 66.66 4.69 ;
      RECT 66.39 3.42 66.54 3.57 ;
      RECT 65.91 3.7 66.06 3.85 ;
      RECT 65.67 4.54 65.82 4.69 ;
      RECT 64.93 3.7 65.08 3.85 ;
      RECT 64.19 3.14 64.34 3.29 ;
      RECT 63.95 4.82 64.1 4.97 ;
      RECT 63.71 3.7 63.86 3.85 ;
      RECT 63.71 4.26 63.86 4.41 ;
      RECT 62.75 4.26 62.9 4.41 ;
      RECT 61.175 9.04 61.325 9.19 ;
      RECT 58.83 9.025 58.98 9.175 ;
      RECT 58.815 3.36 58.965 3.51 ;
      RECT 58.025 3.745 58.175 3.895 ;
      RECT 58.025 8.61 58.175 8.76 ;
      RECT 56.42 2.855 56.57 3.005 ;
      RECT 55.185 3.42 55.335 3.57 ;
      RECT 55.065 3.98 55.215 4.13 ;
      RECT 53.865 3.7 54.015 3.85 ;
      RECT 53.745 4.54 53.895 4.69 ;
      RECT 53.485 3.14 53.635 3.29 ;
      RECT 53.4 9 53.55 9.15 ;
      RECT 52.76 9.45 52.91 9.6 ;
      RECT 52.025 3.7 52.175 3.85 ;
      RECT 51.425 3.7 51.575 3.85 ;
      RECT 51.045 3.14 51.195 3.29 ;
      RECT 50.425 3.98 50.575 4.13 ;
      RECT 50.185 4.54 50.335 4.69 ;
      RECT 50.065 3.42 50.215 3.57 ;
      RECT 49.585 3.7 49.735 3.85 ;
      RECT 49.345 4.54 49.495 4.69 ;
      RECT 48.605 3.7 48.755 3.85 ;
      RECT 47.865 3.14 48.015 3.29 ;
      RECT 47.625 4.82 47.775 4.97 ;
      RECT 47.385 3.7 47.535 3.85 ;
      RECT 47.385 4.26 47.535 4.41 ;
      RECT 46.425 4.26 46.575 4.41 ;
      RECT 44.895 9.045 45.045 9.195 ;
      RECT 42.505 9.025 42.655 9.175 ;
      RECT 42.49 3.36 42.64 3.51 ;
      RECT 41.7 3.745 41.85 3.895 ;
      RECT 41.7 8.61 41.85 8.76 ;
      RECT 40.095 2.855 40.245 3.005 ;
      RECT 38.86 3.42 39.01 3.57 ;
      RECT 38.74 3.98 38.89 4.13 ;
      RECT 37.54 3.7 37.69 3.85 ;
      RECT 37.42 4.54 37.57 4.69 ;
      RECT 37.16 3.14 37.31 3.29 ;
      RECT 37.075 8.995 37.225 9.145 ;
      RECT 36.435 9.45 36.585 9.6 ;
      RECT 35.7 3.7 35.85 3.85 ;
      RECT 35.1 3.7 35.25 3.85 ;
      RECT 34.72 3.14 34.87 3.29 ;
      RECT 34.1 3.98 34.25 4.13 ;
      RECT 33.86 4.54 34.01 4.69 ;
      RECT 33.74 3.42 33.89 3.57 ;
      RECT 33.26 3.7 33.41 3.85 ;
      RECT 33.02 4.54 33.17 4.69 ;
      RECT 32.28 3.7 32.43 3.85 ;
      RECT 31.54 3.14 31.69 3.29 ;
      RECT 31.3 4.82 31.45 4.97 ;
      RECT 31.06 3.7 31.21 3.85 ;
      RECT 31.06 4.26 31.21 4.41 ;
      RECT 30.1 4.26 30.25 4.41 ;
      RECT 28.57 9.04 28.72 9.19 ;
      RECT 26.18 9.025 26.33 9.175 ;
      RECT 26.165 3.36 26.315 3.51 ;
      RECT 25.375 3.745 25.525 3.895 ;
      RECT 25.375 8.61 25.525 8.76 ;
      RECT 23.77 2.855 23.92 3.005 ;
      RECT 22.535 3.42 22.685 3.57 ;
      RECT 22.415 3.98 22.565 4.13 ;
      RECT 21.585 8.99 21.735 9.14 ;
      RECT 21.215 3.7 21.365 3.85 ;
      RECT 21.095 4.54 21.245 4.69 ;
      RECT 20.835 3.14 20.985 3.29 ;
      RECT 20.11 9.45 20.26 9.6 ;
      RECT 19.375 3.7 19.525 3.85 ;
      RECT 18.775 3.7 18.925 3.85 ;
      RECT 18.395 3.14 18.545 3.29 ;
      RECT 17.775 3.98 17.925 4.13 ;
      RECT 17.535 4.54 17.685 4.69 ;
      RECT 17.415 3.42 17.565 3.57 ;
      RECT 16.935 3.7 17.085 3.85 ;
      RECT 16.695 4.54 16.845 4.69 ;
      RECT 15.955 3.7 16.105 3.85 ;
      RECT 15.215 3.14 15.365 3.29 ;
      RECT 14.975 4.82 15.125 4.97 ;
      RECT 14.735 3.7 14.885 3.85 ;
      RECT 14.735 4.26 14.885 4.41 ;
      RECT 13.775 4.26 13.925 4.41 ;
      RECT 11.51 9.38 11.66 9.53 ;
      RECT 11.135 8.64 11.285 8.79 ;
      RECT 10.21 10.9 10.36 11.05 ;
      RECT 10.205 0.115 10.355 0.265 ;
    LAYER met1 ;
      RECT 9.9 10.86 94.325 12.46 ;
      RECT 84.57 8.6 84.745 12.46 ;
      RECT 68.245 8.6 68.42 12.46 ;
      RECT 51.92 8.6 52.095 12.46 ;
      RECT 35.595 8.6 35.77 12.46 ;
      RECT 19.27 8.6 19.445 12.46 ;
      RECT 9.905 10.85 10.71 12.46 ;
      RECT 10.11 10.83 10.46 12.46 ;
      RECT 84.945 8.57 85.235 8.8 ;
      RECT 68.62 8.57 68.91 8.8 ;
      RECT 52.295 8.57 52.585 8.8 ;
      RECT 35.97 8.57 36.26 8.8 ;
      RECT 19.645 8.57 19.935 8.8 ;
      RECT 84.57 8.6 85.235 8.77 ;
      RECT 68.245 8.6 68.91 8.77 ;
      RECT 51.92 8.6 52.585 8.77 ;
      RECT 35.595 8.6 36.26 8.77 ;
      RECT 19.27 8.6 19.935 8.77 ;
      RECT 87.585 4.305 87.905 4.35 ;
      RECT 87.665 3.925 87.905 4.35 ;
      RECT 71.26 4.305 71.58 4.35 ;
      RECT 71.34 3.925 71.58 4.35 ;
      RECT 54.935 4.305 55.255 4.35 ;
      RECT 55.015 3.925 55.255 4.35 ;
      RECT 38.61 4.305 38.93 4.35 ;
      RECT 38.69 3.925 38.93 4.35 ;
      RECT 22.285 4.305 22.605 4.35 ;
      RECT 22.365 3.925 22.605 4.35 ;
      RECT 86.14 4.125 87.905 4.265 ;
      RECT 69.815 4.125 71.58 4.265 ;
      RECT 53.49 4.125 55.255 4.265 ;
      RECT 37.165 4.125 38.93 4.265 ;
      RECT 20.84 4.125 22.605 4.265 ;
      RECT 88.365 0 88.55 4.24 ;
      RECT 72.04 0 72.225 4.24 ;
      RECT 55.715 0 55.9 4.24 ;
      RECT 39.39 0 39.575 4.24 ;
      RECT 23.065 0 23.25 4.24 ;
      RECT 85.805 3.985 86.28 4.17 ;
      RECT 69.48 3.985 69.955 4.17 ;
      RECT 53.155 3.985 53.63 4.17 ;
      RECT 36.83 3.985 37.305 4.17 ;
      RECT 20.505 3.985 20.98 4.17 ;
      RECT 87.6 4.055 88.55 4.24 ;
      RECT 71.275 4.055 72.225 4.24 ;
      RECT 54.95 4.055 55.9 4.24 ;
      RECT 38.625 4.055 39.575 4.24 ;
      RECT 22.3 4.055 23.25 4.24 ;
      RECT 87.6 3.985 88.055 4.24 ;
      RECT 87.63 3.94 88.055 4.24 ;
      RECT 71.275 3.985 71.73 4.24 ;
      RECT 71.305 3.94 71.73 4.24 ;
      RECT 54.95 3.985 55.405 4.24 ;
      RECT 54.98 3.94 55.405 4.24 ;
      RECT 38.625 3.985 39.08 4.24 ;
      RECT 38.655 3.94 39.08 4.24 ;
      RECT 22.3 3.985 22.755 4.24 ;
      RECT 22.33 3.94 22.755 4.24 ;
      RECT 85.805 3.94 86.095 4.17 ;
      RECT 69.48 3.94 69.77 4.17 ;
      RECT 53.155 3.94 53.445 4.17 ;
      RECT 36.83 3.94 37.12 4.17 ;
      RECT 20.505 3.94 20.795 4.17 ;
      RECT 87.63 3.925 87.95 4.24 ;
      RECT 71.305 3.925 71.625 4.24 ;
      RECT 54.98 3.925 55.3 4.24 ;
      RECT 38.655 3.925 38.975 4.24 ;
      RECT 22.33 3.925 22.65 4.24 ;
      RECT 78.735 0 88.55 2.935 ;
      RECT 62.41 0 72.225 2.935 ;
      RECT 46.085 0 55.9 2.935 ;
      RECT 29.76 0 39.575 2.935 ;
      RECT 13.435 0 23.25 2.935 ;
      RECT 9.9 0 94.32 1.6 ;
      RECT 93.715 10.055 94.005 10.285 ;
      RECT 93.775 8.575 93.945 10.285 ;
      RECT 93.75 9.56 94.1 9.91 ;
      RECT 93.715 8.575 94.005 8.805 ;
      RECT 93.31 3.69 93.415 4.26 ;
      RECT 93.31 4.025 93.635 4.255 ;
      RECT 93.31 4.055 93.805 4.225 ;
      RECT 93.31 3.69 93.5 4.255 ;
      RECT 92.725 3.655 93.015 3.885 ;
      RECT 92.725 3.69 93.5 3.86 ;
      RECT 92.785 2.175 92.955 3.885 ;
      RECT 92.725 2.175 93.015 2.405 ;
      RECT 92.725 10.055 93.015 10.285 ;
      RECT 92.785 8.575 92.955 10.285 ;
      RECT 92.725 8.575 93.015 8.805 ;
      RECT 92.725 8.61 93.58 8.77 ;
      RECT 93.41 8.205 93.58 8.77 ;
      RECT 92.725 8.605 93.12 8.77 ;
      RECT 93.345 8.205 93.635 8.435 ;
      RECT 93.345 8.235 93.805 8.405 ;
      RECT 92.355 4.025 92.645 4.255 ;
      RECT 92.355 4.055 92.815 4.225 ;
      RECT 92.42 2.95 92.585 4.255 ;
      RECT 90.935 2.92 91.225 3.15 ;
      RECT 90.935 2.95 92.585 3.12 ;
      RECT 90.995 2.18 91.165 3.15 ;
      RECT 90.935 2.18 91.225 2.41 ;
      RECT 90.935 10.05 91.225 10.28 ;
      RECT 90.995 9.31 91.165 10.28 ;
      RECT 90.995 9.405 92.585 9.575 ;
      RECT 92.415 8.205 92.585 9.575 ;
      RECT 90.935 9.31 91.225 9.54 ;
      RECT 92.355 8.205 92.645 8.435 ;
      RECT 92.355 8.235 92.815 8.405 ;
      RECT 91.365 3.26 91.715 3.61 ;
      RECT 89.06 3.32 91.715 3.49 ;
      RECT 89.06 2.755 89.23 3.49 ;
      RECT 88.97 2.755 89.31 3.105 ;
      RECT 91.39 8.94 91.715 9.265 ;
      RECT 85.955 8.895 86.305 9.245 ;
      RECT 91.365 8.94 91.715 9.17 ;
      RECT 85.75 8.94 86.305 9.17 ;
      RECT 85.58 8.97 91.715 9.14 ;
      RECT 90.59 3.66 90.91 3.98 ;
      RECT 90.56 3.66 90.91 3.89 ;
      RECT 90.39 3.69 90.91 3.86 ;
      RECT 90.59 8.54 90.91 8.83 ;
      RECT 90.56 8.57 90.91 8.8 ;
      RECT 90.39 8.6 90.91 8.77 ;
      RECT 87.045 3.66 87.335 3.89 ;
      RECT 87.045 3.66 87.5 3.845 ;
      RECT 87.36 3.565 87.98 3.705 ;
      RECT 87.75 3.365 88.07 3.625 ;
      RECT 86.43 3.645 86.75 3.905 ;
      RECT 86.43 3.645 86.895 3.89 ;
      RECT 86.755 3.265 86.895 3.89 ;
      RECT 86.755 3.265 87.02 3.405 ;
      RECT 87.285 3.1 87.575 3.33 ;
      RECT 86.88 3.145 87.575 3.285 ;
      RECT 86.325 4.485 86.615 5.01 ;
      RECT 86.31 4.485 86.63 4.745 ;
      RECT 86.05 3.085 86.37 3.345 ;
      RECT 86.05 3.1 86.615 3.33 ;
      RECT 85.325 4.78 85.615 5.01 ;
      RECT 85.52 3.425 85.66 4.965 ;
      RECT 85.565 3.38 85.855 3.61 ;
      RECT 85.16 3.425 85.855 3.565 ;
      RECT 85.16 3.265 85.3 3.565 ;
      RECT 83.7 3.265 85.3 3.405 ;
      RECT 83.61 3.085 83.93 3.345 ;
      RECT 83.61 3.1 84.175 3.345 ;
      RECT 85.32 10.05 85.61 10.28 ;
      RECT 85.38 9.31 85.55 10.28 ;
      RECT 85.3 9.36 85.67 9.71 ;
      RECT 85.3 9.34 85.61 9.71 ;
      RECT 85.32 9.31 85.61 9.71 ;
      RECT 82.72 4.125 85.3 4.265 ;
      RECT 85.085 3.94 85.375 4.17 ;
      RECT 82.645 3.94 83.31 4.17 ;
      RECT 82.99 3.925 83.31 4.265 ;
      RECT 83.99 3.645 84.31 3.905 ;
      RECT 83.99 3.66 84.415 3.89 ;
      RECT 82.63 3.365 82.95 3.625 ;
      RECT 83.125 3.38 83.415 3.61 ;
      RECT 82.63 3.425 83.415 3.565 ;
      RECT 82.75 4.485 83.07 4.745 ;
      RECT 81.91 4.485 82.23 4.745 ;
      RECT 82.75 4.5 83.175 4.73 ;
      RECT 81.91 4.545 83.175 4.685 ;
      RECT 81.445 4.22 81.735 4.45 ;
      RECT 81.52 3.145 81.66 4.45 ;
      RECT 81.17 3.645 81.66 3.905 ;
      RECT 80.925 3.66 81.66 3.89 ;
      RECT 81.925 3.1 82.215 3.33 ;
      RECT 81.52 3.145 82.215 3.285 ;
      RECT 80.685 4.5 80.975 4.73 ;
      RECT 80.685 4.5 81.14 4.685 ;
      RECT 81 4.125 81.14 4.685 ;
      RECT 80.64 4.125 81.14 4.265 ;
      RECT 80.64 3.145 80.78 4.265 ;
      RECT 80.43 3.085 80.75 3.345 ;
      RECT 80.19 4.765 80.51 5.025 ;
      RECT 79.485 4.78 79.775 5.01 ;
      RECT 79.485 4.825 80.51 4.965 ;
      RECT 79.56 4.775 79.82 4.965 ;
      RECT 79.95 3.645 80.27 3.905 ;
      RECT 79.95 3.66 80.495 3.89 ;
      RECT 79.95 4.205 80.27 4.465 ;
      RECT 79.95 4.22 80.495 4.45 ;
      RECT 78.99 4.205 79.31 4.465 ;
      RECT 79.08 3.145 79.22 4.465 ;
      RECT 79.485 3.1 79.775 3.33 ;
      RECT 79.08 3.145 79.775 3.285 ;
      RECT 77.39 10.055 77.68 10.285 ;
      RECT 77.45 8.575 77.62 10.285 ;
      RECT 77.4 8.94 77.75 9.29 ;
      RECT 77.39 8.575 77.68 8.805 ;
      RECT 76.985 3.69 77.09 4.26 ;
      RECT 76.985 4.025 77.31 4.255 ;
      RECT 76.985 4.055 77.48 4.225 ;
      RECT 76.985 3.69 77.175 4.255 ;
      RECT 76.4 3.655 76.69 3.885 ;
      RECT 76.4 3.69 77.175 3.86 ;
      RECT 76.46 2.175 76.63 3.885 ;
      RECT 76.4 2.175 76.69 2.405 ;
      RECT 76.4 10.055 76.69 10.285 ;
      RECT 76.46 8.575 76.63 10.285 ;
      RECT 76.4 8.575 76.69 8.805 ;
      RECT 76.4 8.61 77.255 8.77 ;
      RECT 77.085 8.205 77.255 8.77 ;
      RECT 76.4 8.605 76.795 8.77 ;
      RECT 77.02 8.205 77.31 8.435 ;
      RECT 77.02 8.235 77.48 8.405 ;
      RECT 76.03 4.025 76.32 4.255 ;
      RECT 76.03 4.055 76.49 4.225 ;
      RECT 76.095 2.95 76.26 4.255 ;
      RECT 74.61 2.92 74.9 3.15 ;
      RECT 74.61 2.95 76.26 3.12 ;
      RECT 74.67 2.18 74.84 3.15 ;
      RECT 74.61 2.18 74.9 2.41 ;
      RECT 74.61 10.05 74.9 10.28 ;
      RECT 74.67 9.31 74.84 10.28 ;
      RECT 74.67 9.405 76.26 9.575 ;
      RECT 76.09 8.205 76.26 9.575 ;
      RECT 74.61 9.31 74.9 9.54 ;
      RECT 76.03 8.205 76.32 8.435 ;
      RECT 76.03 8.235 76.49 8.405 ;
      RECT 75.04 3.26 75.39 3.61 ;
      RECT 72.735 3.32 75.39 3.49 ;
      RECT 72.735 2.755 72.905 3.49 ;
      RECT 72.645 2.755 72.985 3.105 ;
      RECT 75.065 8.94 75.39 9.265 ;
      RECT 69.625 8.895 69.975 9.245 ;
      RECT 75.04 8.94 75.39 9.17 ;
      RECT 69.425 8.94 69.975 9.17 ;
      RECT 69.255 8.97 75.39 9.14 ;
      RECT 74.265 3.66 74.585 3.98 ;
      RECT 74.235 3.66 74.585 3.89 ;
      RECT 74.065 3.69 74.585 3.86 ;
      RECT 74.265 8.54 74.585 8.83 ;
      RECT 74.235 8.57 74.585 8.8 ;
      RECT 74.065 8.6 74.585 8.77 ;
      RECT 70.72 3.66 71.01 3.89 ;
      RECT 70.72 3.66 71.175 3.845 ;
      RECT 71.035 3.565 71.655 3.705 ;
      RECT 71.425 3.365 71.745 3.625 ;
      RECT 70.105 3.645 70.425 3.905 ;
      RECT 70.105 3.645 70.57 3.89 ;
      RECT 70.43 3.265 70.57 3.89 ;
      RECT 70.43 3.265 70.695 3.405 ;
      RECT 70.96 3.1 71.25 3.33 ;
      RECT 70.555 3.145 71.25 3.285 ;
      RECT 70 4.485 70.29 5.01 ;
      RECT 69.985 4.485 70.305 4.745 ;
      RECT 69.725 3.085 70.045 3.345 ;
      RECT 69.725 3.1 70.29 3.33 ;
      RECT 69 4.78 69.29 5.01 ;
      RECT 69.195 3.425 69.335 4.965 ;
      RECT 69.24 3.38 69.53 3.61 ;
      RECT 68.835 3.425 69.53 3.565 ;
      RECT 68.835 3.265 68.975 3.565 ;
      RECT 67.375 3.265 68.975 3.405 ;
      RECT 67.285 3.085 67.605 3.345 ;
      RECT 67.285 3.1 67.85 3.345 ;
      RECT 68.995 10.05 69.285 10.28 ;
      RECT 69.055 9.31 69.225 10.28 ;
      RECT 68.975 9.36 69.345 9.71 ;
      RECT 68.975 9.34 69.285 9.71 ;
      RECT 68.995 9.31 69.285 9.71 ;
      RECT 66.395 4.125 68.975 4.265 ;
      RECT 68.76 3.94 69.05 4.17 ;
      RECT 66.32 3.94 66.985 4.17 ;
      RECT 66.665 3.925 66.985 4.265 ;
      RECT 67.665 3.645 67.985 3.905 ;
      RECT 67.665 3.66 68.09 3.89 ;
      RECT 66.305 3.365 66.625 3.625 ;
      RECT 66.8 3.38 67.09 3.61 ;
      RECT 66.305 3.425 67.09 3.565 ;
      RECT 66.425 4.485 66.745 4.745 ;
      RECT 65.585 4.485 65.905 4.745 ;
      RECT 66.425 4.5 66.85 4.73 ;
      RECT 65.585 4.545 66.85 4.685 ;
      RECT 65.12 4.22 65.41 4.45 ;
      RECT 65.195 3.145 65.335 4.45 ;
      RECT 64.845 3.645 65.335 3.905 ;
      RECT 64.6 3.66 65.335 3.89 ;
      RECT 65.6 3.1 65.89 3.33 ;
      RECT 65.195 3.145 65.89 3.285 ;
      RECT 64.36 4.5 64.65 4.73 ;
      RECT 64.36 4.5 64.815 4.685 ;
      RECT 64.675 4.125 64.815 4.685 ;
      RECT 64.315 4.125 64.815 4.265 ;
      RECT 64.315 3.145 64.455 4.265 ;
      RECT 64.105 3.085 64.425 3.345 ;
      RECT 63.865 4.765 64.185 5.025 ;
      RECT 63.16 4.78 63.45 5.01 ;
      RECT 63.16 4.825 64.185 4.965 ;
      RECT 63.235 4.775 63.495 4.965 ;
      RECT 63.625 3.645 63.945 3.905 ;
      RECT 63.625 3.66 64.17 3.89 ;
      RECT 63.625 4.205 63.945 4.465 ;
      RECT 63.625 4.22 64.17 4.45 ;
      RECT 62.665 4.205 62.985 4.465 ;
      RECT 62.755 3.145 62.895 4.465 ;
      RECT 63.16 3.1 63.45 3.33 ;
      RECT 62.755 3.145 63.45 3.285 ;
      RECT 61.065 10.055 61.355 10.285 ;
      RECT 61.125 8.575 61.295 10.285 ;
      RECT 61.075 8.94 61.425 9.29 ;
      RECT 61.065 8.575 61.355 8.805 ;
      RECT 60.66 3.69 60.765 4.26 ;
      RECT 60.66 4.025 60.985 4.255 ;
      RECT 60.66 4.055 61.155 4.225 ;
      RECT 60.66 3.69 60.85 4.255 ;
      RECT 60.075 3.655 60.365 3.885 ;
      RECT 60.075 3.69 60.85 3.86 ;
      RECT 60.135 2.175 60.305 3.885 ;
      RECT 60.075 2.175 60.365 2.405 ;
      RECT 60.075 10.055 60.365 10.285 ;
      RECT 60.135 8.575 60.305 10.285 ;
      RECT 60.075 8.575 60.365 8.805 ;
      RECT 60.075 8.61 60.93 8.77 ;
      RECT 60.76 8.205 60.93 8.77 ;
      RECT 60.075 8.605 60.47 8.77 ;
      RECT 60.695 8.205 60.985 8.435 ;
      RECT 60.695 8.235 61.155 8.405 ;
      RECT 59.705 4.025 59.995 4.255 ;
      RECT 59.705 4.055 60.165 4.225 ;
      RECT 59.77 2.95 59.935 4.255 ;
      RECT 58.285 2.92 58.575 3.15 ;
      RECT 58.285 2.95 59.935 3.12 ;
      RECT 58.345 2.18 58.515 3.15 ;
      RECT 58.285 2.18 58.575 2.41 ;
      RECT 58.285 10.05 58.575 10.28 ;
      RECT 58.345 9.31 58.515 10.28 ;
      RECT 58.345 9.405 59.935 9.575 ;
      RECT 59.765 8.205 59.935 9.575 ;
      RECT 58.285 9.31 58.575 9.54 ;
      RECT 59.705 8.205 59.995 8.435 ;
      RECT 59.705 8.235 60.165 8.405 ;
      RECT 58.715 3.26 59.065 3.61 ;
      RECT 56.41 3.32 59.065 3.49 ;
      RECT 56.41 2.755 56.58 3.49 ;
      RECT 56.32 2.755 56.66 3.105 ;
      RECT 58.74 8.94 59.065 9.265 ;
      RECT 53.3 8.9 53.65 9.25 ;
      RECT 58.715 8.94 59.065 9.17 ;
      RECT 53.1 8.94 53.65 9.17 ;
      RECT 52.93 8.97 59.065 9.14 ;
      RECT 57.94 3.66 58.26 3.98 ;
      RECT 57.91 3.66 58.26 3.89 ;
      RECT 57.74 3.69 58.26 3.86 ;
      RECT 57.94 8.54 58.26 8.83 ;
      RECT 57.91 8.57 58.26 8.8 ;
      RECT 57.74 8.6 58.26 8.77 ;
      RECT 54.395 3.66 54.685 3.89 ;
      RECT 54.395 3.66 54.85 3.845 ;
      RECT 54.71 3.565 55.33 3.705 ;
      RECT 55.1 3.365 55.42 3.625 ;
      RECT 53.78 3.645 54.1 3.905 ;
      RECT 53.78 3.645 54.245 3.89 ;
      RECT 54.105 3.265 54.245 3.89 ;
      RECT 54.105 3.265 54.37 3.405 ;
      RECT 54.635 3.1 54.925 3.33 ;
      RECT 54.23 3.145 54.925 3.285 ;
      RECT 53.675 4.485 53.965 5.01 ;
      RECT 53.66 4.485 53.98 4.745 ;
      RECT 53.4 3.085 53.72 3.345 ;
      RECT 53.4 3.1 53.965 3.33 ;
      RECT 52.675 4.78 52.965 5.01 ;
      RECT 52.87 3.425 53.01 4.965 ;
      RECT 52.915 3.38 53.205 3.61 ;
      RECT 52.51 3.425 53.205 3.565 ;
      RECT 52.51 3.265 52.65 3.565 ;
      RECT 51.05 3.265 52.65 3.405 ;
      RECT 50.96 3.085 51.28 3.345 ;
      RECT 50.96 3.1 51.525 3.345 ;
      RECT 52.67 10.05 52.96 10.28 ;
      RECT 52.73 9.31 52.9 10.28 ;
      RECT 52.65 9.36 53.02 9.71 ;
      RECT 52.65 9.34 52.96 9.71 ;
      RECT 52.67 9.31 52.96 9.71 ;
      RECT 50.07 4.125 52.65 4.265 ;
      RECT 52.435 3.94 52.725 4.17 ;
      RECT 49.995 3.94 50.66 4.17 ;
      RECT 50.34 3.925 50.66 4.265 ;
      RECT 51.34 3.645 51.66 3.905 ;
      RECT 51.34 3.66 51.765 3.89 ;
      RECT 49.98 3.365 50.3 3.625 ;
      RECT 50.475 3.38 50.765 3.61 ;
      RECT 49.98 3.425 50.765 3.565 ;
      RECT 50.1 4.485 50.42 4.745 ;
      RECT 49.26 4.485 49.58 4.745 ;
      RECT 50.1 4.5 50.525 4.73 ;
      RECT 49.26 4.545 50.525 4.685 ;
      RECT 48.795 4.22 49.085 4.45 ;
      RECT 48.87 3.145 49.01 4.45 ;
      RECT 48.52 3.645 49.01 3.905 ;
      RECT 48.275 3.66 49.01 3.89 ;
      RECT 49.275 3.1 49.565 3.33 ;
      RECT 48.87 3.145 49.565 3.285 ;
      RECT 48.035 4.5 48.325 4.73 ;
      RECT 48.035 4.5 48.49 4.685 ;
      RECT 48.35 4.125 48.49 4.685 ;
      RECT 47.99 4.125 48.49 4.265 ;
      RECT 47.99 3.145 48.13 4.265 ;
      RECT 47.78 3.085 48.1 3.345 ;
      RECT 47.54 4.765 47.86 5.025 ;
      RECT 46.835 4.78 47.125 5.01 ;
      RECT 46.835 4.825 47.86 4.965 ;
      RECT 46.91 4.775 47.17 4.965 ;
      RECT 47.3 3.645 47.62 3.905 ;
      RECT 47.3 3.66 47.845 3.89 ;
      RECT 47.3 4.205 47.62 4.465 ;
      RECT 47.3 4.22 47.845 4.45 ;
      RECT 46.34 4.205 46.66 4.465 ;
      RECT 46.43 3.145 46.57 4.465 ;
      RECT 46.835 3.1 47.125 3.33 ;
      RECT 46.43 3.145 47.125 3.285 ;
      RECT 44.74 10.055 45.03 10.285 ;
      RECT 44.8 8.575 44.97 10.285 ;
      RECT 44.79 8.945 45.145 9.3 ;
      RECT 44.74 8.575 45.03 8.805 ;
      RECT 44.335 3.69 44.44 4.26 ;
      RECT 44.335 4.025 44.66 4.255 ;
      RECT 44.335 4.055 44.83 4.225 ;
      RECT 44.335 3.69 44.525 4.255 ;
      RECT 43.75 3.655 44.04 3.885 ;
      RECT 43.75 3.69 44.525 3.86 ;
      RECT 43.81 2.175 43.98 3.885 ;
      RECT 43.75 2.175 44.04 2.405 ;
      RECT 43.75 10.055 44.04 10.285 ;
      RECT 43.81 8.575 43.98 10.285 ;
      RECT 43.75 8.575 44.04 8.805 ;
      RECT 43.75 8.61 44.605 8.77 ;
      RECT 44.435 8.205 44.605 8.77 ;
      RECT 43.75 8.605 44.145 8.77 ;
      RECT 44.37 8.205 44.66 8.435 ;
      RECT 44.37 8.235 44.83 8.405 ;
      RECT 43.38 4.025 43.67 4.255 ;
      RECT 43.38 4.055 43.84 4.225 ;
      RECT 43.445 2.95 43.61 4.255 ;
      RECT 41.96 2.92 42.25 3.15 ;
      RECT 41.96 2.95 43.61 3.12 ;
      RECT 42.02 2.18 42.19 3.15 ;
      RECT 41.96 2.18 42.25 2.41 ;
      RECT 41.96 10.05 42.25 10.28 ;
      RECT 42.02 9.31 42.19 10.28 ;
      RECT 42.02 9.405 43.61 9.575 ;
      RECT 43.44 8.205 43.61 9.575 ;
      RECT 41.96 9.31 42.25 9.54 ;
      RECT 43.38 8.205 43.67 8.435 ;
      RECT 43.38 8.235 43.84 8.405 ;
      RECT 42.39 3.26 42.74 3.61 ;
      RECT 40.085 3.32 42.74 3.49 ;
      RECT 40.085 2.755 40.255 3.49 ;
      RECT 39.995 2.755 40.335 3.105 ;
      RECT 42.415 8.94 42.74 9.265 ;
      RECT 36.975 8.895 37.325 9.245 ;
      RECT 42.39 8.94 42.74 9.17 ;
      RECT 36.775 8.94 37.325 9.17 ;
      RECT 36.605 8.97 42.74 9.14 ;
      RECT 41.615 3.66 41.935 3.98 ;
      RECT 41.585 3.66 41.935 3.89 ;
      RECT 41.415 3.69 41.935 3.86 ;
      RECT 41.615 8.54 41.935 8.83 ;
      RECT 41.585 8.57 41.935 8.8 ;
      RECT 41.415 8.6 41.935 8.77 ;
      RECT 38.07 3.66 38.36 3.89 ;
      RECT 38.07 3.66 38.525 3.845 ;
      RECT 38.385 3.565 39.005 3.705 ;
      RECT 38.775 3.365 39.095 3.625 ;
      RECT 37.455 3.645 37.775 3.905 ;
      RECT 37.455 3.645 37.92 3.89 ;
      RECT 37.78 3.265 37.92 3.89 ;
      RECT 37.78 3.265 38.045 3.405 ;
      RECT 38.31 3.1 38.6 3.33 ;
      RECT 37.905 3.145 38.6 3.285 ;
      RECT 37.35 4.485 37.64 5.01 ;
      RECT 37.335 4.485 37.655 4.745 ;
      RECT 37.075 3.085 37.395 3.345 ;
      RECT 37.075 3.1 37.64 3.33 ;
      RECT 36.35 4.78 36.64 5.01 ;
      RECT 36.545 3.425 36.685 4.965 ;
      RECT 36.59 3.38 36.88 3.61 ;
      RECT 36.185 3.425 36.88 3.565 ;
      RECT 36.185 3.265 36.325 3.565 ;
      RECT 34.725 3.265 36.325 3.405 ;
      RECT 34.635 3.085 34.955 3.345 ;
      RECT 34.635 3.1 35.2 3.345 ;
      RECT 36.345 10.05 36.635 10.28 ;
      RECT 36.405 9.31 36.575 10.28 ;
      RECT 36.325 9.36 36.695 9.71 ;
      RECT 36.325 9.34 36.635 9.71 ;
      RECT 36.345 9.31 36.635 9.71 ;
      RECT 33.745 4.125 36.325 4.265 ;
      RECT 36.11 3.94 36.4 4.17 ;
      RECT 33.67 3.94 34.335 4.17 ;
      RECT 34.015 3.925 34.335 4.265 ;
      RECT 35.015 3.645 35.335 3.905 ;
      RECT 35.015 3.66 35.44 3.89 ;
      RECT 33.655 3.365 33.975 3.625 ;
      RECT 34.15 3.38 34.44 3.61 ;
      RECT 33.655 3.425 34.44 3.565 ;
      RECT 33.775 4.485 34.095 4.745 ;
      RECT 32.935 4.485 33.255 4.745 ;
      RECT 33.775 4.5 34.2 4.73 ;
      RECT 32.935 4.545 34.2 4.685 ;
      RECT 32.47 4.22 32.76 4.45 ;
      RECT 32.545 3.145 32.685 4.45 ;
      RECT 32.195 3.645 32.685 3.905 ;
      RECT 31.95 3.66 32.685 3.89 ;
      RECT 32.95 3.1 33.24 3.33 ;
      RECT 32.545 3.145 33.24 3.285 ;
      RECT 31.71 4.5 32 4.73 ;
      RECT 31.71 4.5 32.165 4.685 ;
      RECT 32.025 4.125 32.165 4.685 ;
      RECT 31.665 4.125 32.165 4.265 ;
      RECT 31.665 3.145 31.805 4.265 ;
      RECT 31.455 3.085 31.775 3.345 ;
      RECT 31.215 4.765 31.535 5.025 ;
      RECT 30.51 4.78 30.8 5.01 ;
      RECT 30.51 4.825 31.535 4.965 ;
      RECT 30.585 4.775 30.845 4.965 ;
      RECT 30.975 3.645 31.295 3.905 ;
      RECT 30.975 3.66 31.52 3.89 ;
      RECT 30.975 4.205 31.295 4.465 ;
      RECT 30.975 4.22 31.52 4.45 ;
      RECT 30.015 4.205 30.335 4.465 ;
      RECT 30.105 3.145 30.245 4.465 ;
      RECT 30.51 3.1 30.8 3.33 ;
      RECT 30.105 3.145 30.8 3.285 ;
      RECT 28.415 10.055 28.705 10.285 ;
      RECT 28.475 8.575 28.645 10.285 ;
      RECT 28.47 8.94 28.82 9.29 ;
      RECT 28.415 8.575 28.705 8.805 ;
      RECT 28.01 3.69 28.115 4.26 ;
      RECT 28.01 4.025 28.335 4.255 ;
      RECT 28.01 4.055 28.505 4.225 ;
      RECT 28.01 3.69 28.2 4.255 ;
      RECT 27.425 3.655 27.715 3.885 ;
      RECT 27.425 3.69 28.2 3.86 ;
      RECT 27.485 2.175 27.655 3.885 ;
      RECT 27.425 2.175 27.715 2.405 ;
      RECT 27.425 10.055 27.715 10.285 ;
      RECT 27.485 8.575 27.655 10.285 ;
      RECT 27.425 8.575 27.715 8.805 ;
      RECT 27.425 8.61 28.28 8.77 ;
      RECT 28.11 8.205 28.28 8.77 ;
      RECT 27.425 8.605 27.82 8.77 ;
      RECT 28.045 8.205 28.335 8.435 ;
      RECT 28.045 8.235 28.505 8.405 ;
      RECT 27.055 4.025 27.345 4.255 ;
      RECT 27.055 4.055 27.515 4.225 ;
      RECT 27.12 2.95 27.285 4.255 ;
      RECT 25.635 2.92 25.925 3.15 ;
      RECT 25.635 2.95 27.285 3.12 ;
      RECT 25.695 2.18 25.865 3.15 ;
      RECT 25.635 2.18 25.925 2.41 ;
      RECT 25.635 10.05 25.925 10.28 ;
      RECT 25.695 9.31 25.865 10.28 ;
      RECT 25.695 9.405 27.285 9.575 ;
      RECT 27.115 8.205 27.285 9.575 ;
      RECT 25.635 9.31 25.925 9.54 ;
      RECT 27.055 8.205 27.345 8.435 ;
      RECT 27.055 8.235 27.515 8.405 ;
      RECT 26.065 3.26 26.415 3.61 ;
      RECT 23.76 3.32 26.415 3.49 ;
      RECT 23.76 2.755 23.93 3.49 ;
      RECT 23.67 2.755 24.01 3.105 ;
      RECT 26.09 8.94 26.415 9.265 ;
      RECT 21.485 8.89 21.835 9.24 ;
      RECT 26.065 8.94 26.415 9.17 ;
      RECT 20.45 8.94 20.74 9.17 ;
      RECT 20.28 8.97 26.415 9.14 ;
      RECT 25.29 3.66 25.61 3.98 ;
      RECT 25.26 3.66 25.61 3.89 ;
      RECT 25.09 3.69 25.61 3.86 ;
      RECT 25.29 8.54 25.61 8.83 ;
      RECT 25.26 8.57 25.61 8.8 ;
      RECT 25.09 8.6 25.61 8.77 ;
      RECT 21.745 3.66 22.035 3.89 ;
      RECT 21.745 3.66 22.2 3.845 ;
      RECT 22.06 3.565 22.68 3.705 ;
      RECT 22.45 3.365 22.77 3.625 ;
      RECT 21.13 3.645 21.45 3.905 ;
      RECT 21.13 3.645 21.595 3.89 ;
      RECT 21.455 3.265 21.595 3.89 ;
      RECT 21.455 3.265 21.72 3.405 ;
      RECT 21.985 3.1 22.275 3.33 ;
      RECT 21.58 3.145 22.275 3.285 ;
      RECT 21.025 4.485 21.315 5.01 ;
      RECT 21.01 4.485 21.33 4.745 ;
      RECT 20.75 3.085 21.07 3.345 ;
      RECT 20.75 3.1 21.315 3.33 ;
      RECT 20.025 4.78 20.315 5.01 ;
      RECT 20.22 3.425 20.36 4.965 ;
      RECT 20.265 3.38 20.555 3.61 ;
      RECT 19.86 3.425 20.555 3.565 ;
      RECT 19.86 3.265 20 3.565 ;
      RECT 18.4 3.265 20 3.405 ;
      RECT 18.31 3.085 18.63 3.345 ;
      RECT 18.31 3.1 18.875 3.345 ;
      RECT 20.02 10.05 20.31 10.28 ;
      RECT 20.08 9.31 20.25 10.28 ;
      RECT 20 9.36 20.37 9.71 ;
      RECT 20 9.34 20.31 9.71 ;
      RECT 20.02 9.31 20.31 9.71 ;
      RECT 17.42 4.125 20 4.265 ;
      RECT 19.785 3.94 20.075 4.17 ;
      RECT 17.345 3.94 18.01 4.17 ;
      RECT 17.69 3.925 18.01 4.265 ;
      RECT 18.69 3.645 19.01 3.905 ;
      RECT 18.69 3.66 19.115 3.89 ;
      RECT 17.33 3.365 17.65 3.625 ;
      RECT 17.825 3.38 18.115 3.61 ;
      RECT 17.33 3.425 18.115 3.565 ;
      RECT 17.45 4.485 17.77 4.745 ;
      RECT 16.61 4.485 16.93 4.745 ;
      RECT 17.45 4.5 17.875 4.73 ;
      RECT 16.61 4.545 17.875 4.685 ;
      RECT 16.145 4.22 16.435 4.45 ;
      RECT 16.22 3.145 16.36 4.45 ;
      RECT 15.87 3.645 16.36 3.905 ;
      RECT 15.625 3.66 16.36 3.89 ;
      RECT 16.625 3.1 16.915 3.33 ;
      RECT 16.22 3.145 16.915 3.285 ;
      RECT 15.385 4.5 15.675 4.73 ;
      RECT 15.385 4.5 15.84 4.685 ;
      RECT 15.7 4.125 15.84 4.685 ;
      RECT 15.34 4.125 15.84 4.265 ;
      RECT 15.34 3.145 15.48 4.265 ;
      RECT 15.13 3.085 15.45 3.345 ;
      RECT 14.89 4.765 15.21 5.025 ;
      RECT 14.185 4.78 14.475 5.01 ;
      RECT 14.185 4.825 15.21 4.965 ;
      RECT 14.26 4.775 14.52 4.965 ;
      RECT 14.65 3.645 14.97 3.905 ;
      RECT 14.65 3.66 15.195 3.89 ;
      RECT 14.65 4.205 14.97 4.465 ;
      RECT 14.65 4.22 15.195 4.45 ;
      RECT 13.69 4.205 14.01 4.465 ;
      RECT 13.78 3.145 13.92 4.465 ;
      RECT 14.185 3.1 14.475 3.33 ;
      RECT 13.78 3.145 14.475 3.285 ;
      RECT 11.44 10.05 11.73 10.28 ;
      RECT 11.5 9.31 11.67 10.28 ;
      RECT 11.41 9.31 11.76 9.6 ;
      RECT 11.035 8.57 11.385 8.86 ;
      RECT 10.895 8.6 11.385 8.77 ;
      RECT 84.59 3.645 84.91 3.905 ;
      RECT 82.15 3.645 82.47 3.905 ;
      RECT 68.265 3.645 68.585 3.905 ;
      RECT 65.825 3.645 66.145 3.905 ;
      RECT 51.94 3.645 52.26 3.905 ;
      RECT 49.5 3.645 49.82 3.905 ;
      RECT 35.615 3.645 35.935 3.905 ;
      RECT 33.175 3.645 33.495 3.905 ;
      RECT 19.29 3.645 19.61 3.905 ;
      RECT 16.85 3.645 17.17 3.905 ;
    LAYER mcon ;
      RECT 93.775 8.605 93.945 8.775 ;
      RECT 93.78 8.6 93.95 8.77 ;
      RECT 77.45 8.605 77.62 8.775 ;
      RECT 77.455 8.6 77.625 8.77 ;
      RECT 61.125 8.605 61.295 8.775 ;
      RECT 61.13 8.6 61.3 8.77 ;
      RECT 44.8 8.605 44.97 8.775 ;
      RECT 44.805 8.6 44.975 8.77 ;
      RECT 28.475 8.605 28.645 8.775 ;
      RECT 28.48 8.6 28.65 8.77 ;
      RECT 93.775 10.085 93.945 10.255 ;
      RECT 93.425 1.395 93.595 1.565 ;
      RECT 93.425 10.895 93.595 11.065 ;
      RECT 93.405 4.055 93.575 4.225 ;
      RECT 93.405 8.235 93.575 8.405 ;
      RECT 92.785 2.205 92.955 2.375 ;
      RECT 92.785 3.685 92.955 3.855 ;
      RECT 92.785 8.605 92.955 8.775 ;
      RECT 92.785 10.085 92.955 10.255 ;
      RECT 92.435 1.395 92.605 1.565 ;
      RECT 92.435 10.895 92.605 11.065 ;
      RECT 92.415 4.055 92.585 4.225 ;
      RECT 92.415 8.235 92.585 8.405 ;
      RECT 91.735 1.4 91.905 1.57 ;
      RECT 91.735 10.89 91.905 11.06 ;
      RECT 91.425 3.32 91.595 3.49 ;
      RECT 91.425 8.97 91.595 9.14 ;
      RECT 91.055 1.4 91.225 1.57 ;
      RECT 91.055 10.89 91.225 11.06 ;
      RECT 90.995 2.21 91.165 2.38 ;
      RECT 90.995 2.95 91.165 3.12 ;
      RECT 90.995 9.34 91.165 9.51 ;
      RECT 90.995 10.08 91.165 10.25 ;
      RECT 90.62 3.69 90.79 3.86 ;
      RECT 90.62 8.6 90.79 8.77 ;
      RECT 90.375 1.4 90.545 1.57 ;
      RECT 90.375 10.89 90.545 11.06 ;
      RECT 89.695 1.4 89.865 1.57 ;
      RECT 89.695 10.89 89.865 11.06 ;
      RECT 88.08 2.61 88.25 2.78 ;
      RECT 87.825 3.97 87.995 4.14 ;
      RECT 87.62 2.61 87.79 2.78 ;
      RECT 87.345 3.13 87.515 3.3 ;
      RECT 87.16 2.61 87.33 2.78 ;
      RECT 87.105 3.69 87.275 3.86 ;
      RECT 86.7 2.61 86.87 2.78 ;
      RECT 86.625 3.69 86.795 3.86 ;
      RECT 86.385 3.13 86.555 3.3 ;
      RECT 86.385 4.81 86.555 4.98 ;
      RECT 86.24 2.61 86.41 2.78 ;
      RECT 86.12 10.89 86.29 11.06 ;
      RECT 85.865 3.97 86.035 4.14 ;
      RECT 85.81 8.97 85.98 9.14 ;
      RECT 85.78 2.61 85.95 2.78 ;
      RECT 85.625 3.41 85.795 3.58 ;
      RECT 85.44 10.89 85.61 11.06 ;
      RECT 85.385 4.81 85.555 4.98 ;
      RECT 85.38 9.34 85.55 9.51 ;
      RECT 85.38 10.08 85.55 10.25 ;
      RECT 85.32 2.61 85.49 2.78 ;
      RECT 85.145 3.97 85.315 4.14 ;
      RECT 85.005 8.6 85.175 8.77 ;
      RECT 84.86 2.61 85.03 2.78 ;
      RECT 84.76 10.89 84.93 11.06 ;
      RECT 84.665 3.69 84.835 3.86 ;
      RECT 84.4 2.61 84.57 2.78 ;
      RECT 84.185 3.69 84.355 3.86 ;
      RECT 84.08 10.89 84.25 11.06 ;
      RECT 83.945 3.13 84.115 3.3 ;
      RECT 83.94 2.61 84.11 2.78 ;
      RECT 83.48 2.61 83.65 2.78 ;
      RECT 83.185 3.41 83.355 3.58 ;
      RECT 83.02 2.61 83.19 2.78 ;
      RECT 82.945 4.53 83.115 4.7 ;
      RECT 82.705 3.97 82.875 4.14 ;
      RECT 82.56 2.61 82.73 2.78 ;
      RECT 82.225 3.69 82.395 3.86 ;
      RECT 82.1 2.61 82.27 2.78 ;
      RECT 81.985 3.13 82.155 3.3 ;
      RECT 81.985 4.53 82.155 4.7 ;
      RECT 81.64 2.61 81.81 2.78 ;
      RECT 81.505 4.25 81.675 4.42 ;
      RECT 81.18 2.61 81.35 2.78 ;
      RECT 80.985 3.69 81.155 3.86 ;
      RECT 80.745 4.53 80.915 4.7 ;
      RECT 80.72 2.61 80.89 2.78 ;
      RECT 80.505 3.13 80.675 3.3 ;
      RECT 80.265 3.69 80.435 3.86 ;
      RECT 80.265 4.25 80.435 4.42 ;
      RECT 80.26 2.61 80.43 2.78 ;
      RECT 79.8 2.61 79.97 2.78 ;
      RECT 79.545 3.13 79.715 3.3 ;
      RECT 79.545 4.81 79.715 4.98 ;
      RECT 79.34 2.61 79.51 2.78 ;
      RECT 79.065 4.25 79.235 4.42 ;
      RECT 78.88 2.61 79.05 2.78 ;
      RECT 77.45 10.085 77.62 10.255 ;
      RECT 77.1 1.395 77.27 1.565 ;
      RECT 77.1 10.895 77.27 11.065 ;
      RECT 77.08 4.055 77.25 4.225 ;
      RECT 77.08 8.235 77.25 8.405 ;
      RECT 76.46 2.205 76.63 2.375 ;
      RECT 76.46 3.685 76.63 3.855 ;
      RECT 76.46 8.605 76.63 8.775 ;
      RECT 76.46 10.085 76.63 10.255 ;
      RECT 76.11 1.395 76.28 1.565 ;
      RECT 76.11 10.895 76.28 11.065 ;
      RECT 76.09 4.055 76.26 4.225 ;
      RECT 76.09 8.235 76.26 8.405 ;
      RECT 75.41 1.4 75.58 1.57 ;
      RECT 75.41 10.89 75.58 11.06 ;
      RECT 75.1 3.32 75.27 3.49 ;
      RECT 75.1 8.97 75.27 9.14 ;
      RECT 74.73 1.4 74.9 1.57 ;
      RECT 74.73 10.89 74.9 11.06 ;
      RECT 74.67 2.21 74.84 2.38 ;
      RECT 74.67 2.95 74.84 3.12 ;
      RECT 74.67 9.34 74.84 9.51 ;
      RECT 74.67 10.08 74.84 10.25 ;
      RECT 74.295 3.69 74.465 3.86 ;
      RECT 74.295 8.6 74.465 8.77 ;
      RECT 74.05 1.4 74.22 1.57 ;
      RECT 74.05 10.89 74.22 11.06 ;
      RECT 73.37 1.4 73.54 1.57 ;
      RECT 73.37 10.89 73.54 11.06 ;
      RECT 71.755 2.61 71.925 2.78 ;
      RECT 71.5 3.97 71.67 4.14 ;
      RECT 71.295 2.61 71.465 2.78 ;
      RECT 71.02 3.13 71.19 3.3 ;
      RECT 70.835 2.61 71.005 2.78 ;
      RECT 70.78 3.69 70.95 3.86 ;
      RECT 70.375 2.61 70.545 2.78 ;
      RECT 70.3 3.69 70.47 3.86 ;
      RECT 70.06 3.13 70.23 3.3 ;
      RECT 70.06 4.81 70.23 4.98 ;
      RECT 69.915 2.61 70.085 2.78 ;
      RECT 69.795 10.89 69.965 11.06 ;
      RECT 69.54 3.97 69.71 4.14 ;
      RECT 69.485 8.97 69.655 9.14 ;
      RECT 69.455 2.61 69.625 2.78 ;
      RECT 69.3 3.41 69.47 3.58 ;
      RECT 69.115 10.89 69.285 11.06 ;
      RECT 69.06 4.81 69.23 4.98 ;
      RECT 69.055 9.34 69.225 9.51 ;
      RECT 69.055 10.08 69.225 10.25 ;
      RECT 68.995 2.61 69.165 2.78 ;
      RECT 68.82 3.97 68.99 4.14 ;
      RECT 68.68 8.6 68.85 8.77 ;
      RECT 68.535 2.61 68.705 2.78 ;
      RECT 68.435 10.89 68.605 11.06 ;
      RECT 68.34 3.69 68.51 3.86 ;
      RECT 68.075 2.61 68.245 2.78 ;
      RECT 67.86 3.69 68.03 3.86 ;
      RECT 67.755 10.89 67.925 11.06 ;
      RECT 67.62 3.13 67.79 3.3 ;
      RECT 67.615 2.61 67.785 2.78 ;
      RECT 67.155 2.61 67.325 2.78 ;
      RECT 66.86 3.41 67.03 3.58 ;
      RECT 66.695 2.61 66.865 2.78 ;
      RECT 66.62 4.53 66.79 4.7 ;
      RECT 66.38 3.97 66.55 4.14 ;
      RECT 66.235 2.61 66.405 2.78 ;
      RECT 65.9 3.69 66.07 3.86 ;
      RECT 65.775 2.61 65.945 2.78 ;
      RECT 65.66 3.13 65.83 3.3 ;
      RECT 65.66 4.53 65.83 4.7 ;
      RECT 65.315 2.61 65.485 2.78 ;
      RECT 65.18 4.25 65.35 4.42 ;
      RECT 64.855 2.61 65.025 2.78 ;
      RECT 64.66 3.69 64.83 3.86 ;
      RECT 64.42 4.53 64.59 4.7 ;
      RECT 64.395 2.61 64.565 2.78 ;
      RECT 64.18 3.13 64.35 3.3 ;
      RECT 63.94 3.69 64.11 3.86 ;
      RECT 63.94 4.25 64.11 4.42 ;
      RECT 63.935 2.61 64.105 2.78 ;
      RECT 63.475 2.61 63.645 2.78 ;
      RECT 63.22 3.13 63.39 3.3 ;
      RECT 63.22 4.81 63.39 4.98 ;
      RECT 63.015 2.61 63.185 2.78 ;
      RECT 62.74 4.25 62.91 4.42 ;
      RECT 62.555 2.61 62.725 2.78 ;
      RECT 61.125 10.085 61.295 10.255 ;
      RECT 60.775 1.395 60.945 1.565 ;
      RECT 60.775 10.895 60.945 11.065 ;
      RECT 60.755 4.055 60.925 4.225 ;
      RECT 60.755 8.235 60.925 8.405 ;
      RECT 60.135 2.205 60.305 2.375 ;
      RECT 60.135 3.685 60.305 3.855 ;
      RECT 60.135 8.605 60.305 8.775 ;
      RECT 60.135 10.085 60.305 10.255 ;
      RECT 59.785 1.395 59.955 1.565 ;
      RECT 59.785 10.895 59.955 11.065 ;
      RECT 59.765 4.055 59.935 4.225 ;
      RECT 59.765 8.235 59.935 8.405 ;
      RECT 59.085 1.4 59.255 1.57 ;
      RECT 59.085 10.89 59.255 11.06 ;
      RECT 58.775 3.32 58.945 3.49 ;
      RECT 58.775 8.97 58.945 9.14 ;
      RECT 58.405 1.4 58.575 1.57 ;
      RECT 58.405 10.89 58.575 11.06 ;
      RECT 58.345 2.21 58.515 2.38 ;
      RECT 58.345 2.95 58.515 3.12 ;
      RECT 58.345 9.34 58.515 9.51 ;
      RECT 58.345 10.08 58.515 10.25 ;
      RECT 57.97 3.69 58.14 3.86 ;
      RECT 57.97 8.6 58.14 8.77 ;
      RECT 57.725 1.4 57.895 1.57 ;
      RECT 57.725 10.89 57.895 11.06 ;
      RECT 57.045 1.4 57.215 1.57 ;
      RECT 57.045 10.89 57.215 11.06 ;
      RECT 55.43 2.61 55.6 2.78 ;
      RECT 55.175 3.97 55.345 4.14 ;
      RECT 54.97 2.61 55.14 2.78 ;
      RECT 54.695 3.13 54.865 3.3 ;
      RECT 54.51 2.61 54.68 2.78 ;
      RECT 54.455 3.69 54.625 3.86 ;
      RECT 54.05 2.61 54.22 2.78 ;
      RECT 53.975 3.69 54.145 3.86 ;
      RECT 53.735 3.13 53.905 3.3 ;
      RECT 53.735 4.81 53.905 4.98 ;
      RECT 53.59 2.61 53.76 2.78 ;
      RECT 53.47 10.89 53.64 11.06 ;
      RECT 53.215 3.97 53.385 4.14 ;
      RECT 53.16 8.97 53.33 9.14 ;
      RECT 53.13 2.61 53.3 2.78 ;
      RECT 52.975 3.41 53.145 3.58 ;
      RECT 52.79 10.89 52.96 11.06 ;
      RECT 52.735 4.81 52.905 4.98 ;
      RECT 52.73 9.34 52.9 9.51 ;
      RECT 52.73 10.08 52.9 10.25 ;
      RECT 52.67 2.61 52.84 2.78 ;
      RECT 52.495 3.97 52.665 4.14 ;
      RECT 52.355 8.6 52.525 8.77 ;
      RECT 52.21 2.61 52.38 2.78 ;
      RECT 52.11 10.89 52.28 11.06 ;
      RECT 52.015 3.69 52.185 3.86 ;
      RECT 51.75 2.61 51.92 2.78 ;
      RECT 51.535 3.69 51.705 3.86 ;
      RECT 51.43 10.89 51.6 11.06 ;
      RECT 51.295 3.13 51.465 3.3 ;
      RECT 51.29 2.61 51.46 2.78 ;
      RECT 50.83 2.61 51 2.78 ;
      RECT 50.535 3.41 50.705 3.58 ;
      RECT 50.37 2.61 50.54 2.78 ;
      RECT 50.295 4.53 50.465 4.7 ;
      RECT 50.055 3.97 50.225 4.14 ;
      RECT 49.91 2.61 50.08 2.78 ;
      RECT 49.575 3.69 49.745 3.86 ;
      RECT 49.45 2.61 49.62 2.78 ;
      RECT 49.335 3.13 49.505 3.3 ;
      RECT 49.335 4.53 49.505 4.7 ;
      RECT 48.99 2.61 49.16 2.78 ;
      RECT 48.855 4.25 49.025 4.42 ;
      RECT 48.53 2.61 48.7 2.78 ;
      RECT 48.335 3.69 48.505 3.86 ;
      RECT 48.095 4.53 48.265 4.7 ;
      RECT 48.07 2.61 48.24 2.78 ;
      RECT 47.855 3.13 48.025 3.3 ;
      RECT 47.615 3.69 47.785 3.86 ;
      RECT 47.615 4.25 47.785 4.42 ;
      RECT 47.61 2.61 47.78 2.78 ;
      RECT 47.15 2.61 47.32 2.78 ;
      RECT 46.895 3.13 47.065 3.3 ;
      RECT 46.895 4.81 47.065 4.98 ;
      RECT 46.69 2.61 46.86 2.78 ;
      RECT 46.415 4.25 46.585 4.42 ;
      RECT 46.23 2.61 46.4 2.78 ;
      RECT 44.8 10.085 44.97 10.255 ;
      RECT 44.45 1.395 44.62 1.565 ;
      RECT 44.45 10.895 44.62 11.065 ;
      RECT 44.43 4.055 44.6 4.225 ;
      RECT 44.43 8.235 44.6 8.405 ;
      RECT 43.81 2.205 43.98 2.375 ;
      RECT 43.81 3.685 43.98 3.855 ;
      RECT 43.81 8.605 43.98 8.775 ;
      RECT 43.81 10.085 43.98 10.255 ;
      RECT 43.46 1.395 43.63 1.565 ;
      RECT 43.46 10.895 43.63 11.065 ;
      RECT 43.44 4.055 43.61 4.225 ;
      RECT 43.44 8.235 43.61 8.405 ;
      RECT 42.76 1.4 42.93 1.57 ;
      RECT 42.76 10.89 42.93 11.06 ;
      RECT 42.45 3.32 42.62 3.49 ;
      RECT 42.45 8.97 42.62 9.14 ;
      RECT 42.08 1.4 42.25 1.57 ;
      RECT 42.08 10.89 42.25 11.06 ;
      RECT 42.02 2.21 42.19 2.38 ;
      RECT 42.02 2.95 42.19 3.12 ;
      RECT 42.02 9.34 42.19 9.51 ;
      RECT 42.02 10.08 42.19 10.25 ;
      RECT 41.645 3.69 41.815 3.86 ;
      RECT 41.645 8.6 41.815 8.77 ;
      RECT 41.4 1.4 41.57 1.57 ;
      RECT 41.4 10.89 41.57 11.06 ;
      RECT 40.72 1.4 40.89 1.57 ;
      RECT 40.72 10.89 40.89 11.06 ;
      RECT 39.105 2.61 39.275 2.78 ;
      RECT 38.85 3.97 39.02 4.14 ;
      RECT 38.645 2.61 38.815 2.78 ;
      RECT 38.37 3.13 38.54 3.3 ;
      RECT 38.185 2.61 38.355 2.78 ;
      RECT 38.13 3.69 38.3 3.86 ;
      RECT 37.725 2.61 37.895 2.78 ;
      RECT 37.65 3.69 37.82 3.86 ;
      RECT 37.41 3.13 37.58 3.3 ;
      RECT 37.41 4.81 37.58 4.98 ;
      RECT 37.265 2.61 37.435 2.78 ;
      RECT 37.145 10.89 37.315 11.06 ;
      RECT 36.89 3.97 37.06 4.14 ;
      RECT 36.835 8.97 37.005 9.14 ;
      RECT 36.805 2.61 36.975 2.78 ;
      RECT 36.65 3.41 36.82 3.58 ;
      RECT 36.465 10.89 36.635 11.06 ;
      RECT 36.41 4.81 36.58 4.98 ;
      RECT 36.405 9.34 36.575 9.51 ;
      RECT 36.405 10.08 36.575 10.25 ;
      RECT 36.345 2.61 36.515 2.78 ;
      RECT 36.17 3.97 36.34 4.14 ;
      RECT 36.03 8.6 36.2 8.77 ;
      RECT 35.885 2.61 36.055 2.78 ;
      RECT 35.785 10.89 35.955 11.06 ;
      RECT 35.69 3.69 35.86 3.86 ;
      RECT 35.425 2.61 35.595 2.78 ;
      RECT 35.21 3.69 35.38 3.86 ;
      RECT 35.105 10.89 35.275 11.06 ;
      RECT 34.97 3.13 35.14 3.3 ;
      RECT 34.965 2.61 35.135 2.78 ;
      RECT 34.505 2.61 34.675 2.78 ;
      RECT 34.21 3.41 34.38 3.58 ;
      RECT 34.045 2.61 34.215 2.78 ;
      RECT 33.97 4.53 34.14 4.7 ;
      RECT 33.73 3.97 33.9 4.14 ;
      RECT 33.585 2.61 33.755 2.78 ;
      RECT 33.25 3.69 33.42 3.86 ;
      RECT 33.125 2.61 33.295 2.78 ;
      RECT 33.01 3.13 33.18 3.3 ;
      RECT 33.01 4.53 33.18 4.7 ;
      RECT 32.665 2.61 32.835 2.78 ;
      RECT 32.53 4.25 32.7 4.42 ;
      RECT 32.205 2.61 32.375 2.78 ;
      RECT 32.01 3.69 32.18 3.86 ;
      RECT 31.77 4.53 31.94 4.7 ;
      RECT 31.745 2.61 31.915 2.78 ;
      RECT 31.53 3.13 31.7 3.3 ;
      RECT 31.29 3.69 31.46 3.86 ;
      RECT 31.29 4.25 31.46 4.42 ;
      RECT 31.285 2.61 31.455 2.78 ;
      RECT 30.825 2.61 30.995 2.78 ;
      RECT 30.57 3.13 30.74 3.3 ;
      RECT 30.57 4.81 30.74 4.98 ;
      RECT 30.365 2.61 30.535 2.78 ;
      RECT 30.09 4.25 30.26 4.42 ;
      RECT 29.905 2.61 30.075 2.78 ;
      RECT 28.475 10.085 28.645 10.255 ;
      RECT 28.125 1.395 28.295 1.565 ;
      RECT 28.125 10.895 28.295 11.065 ;
      RECT 28.105 4.055 28.275 4.225 ;
      RECT 28.105 8.235 28.275 8.405 ;
      RECT 27.485 2.205 27.655 2.375 ;
      RECT 27.485 3.685 27.655 3.855 ;
      RECT 27.485 8.605 27.655 8.775 ;
      RECT 27.485 10.085 27.655 10.255 ;
      RECT 27.135 1.395 27.305 1.565 ;
      RECT 27.135 10.895 27.305 11.065 ;
      RECT 27.115 4.055 27.285 4.225 ;
      RECT 27.115 8.235 27.285 8.405 ;
      RECT 26.435 1.4 26.605 1.57 ;
      RECT 26.435 10.89 26.605 11.06 ;
      RECT 26.125 3.32 26.295 3.49 ;
      RECT 26.125 8.97 26.295 9.14 ;
      RECT 25.755 1.4 25.925 1.57 ;
      RECT 25.755 10.89 25.925 11.06 ;
      RECT 25.695 2.21 25.865 2.38 ;
      RECT 25.695 2.95 25.865 3.12 ;
      RECT 25.695 9.34 25.865 9.51 ;
      RECT 25.695 10.08 25.865 10.25 ;
      RECT 25.32 3.69 25.49 3.86 ;
      RECT 25.32 8.6 25.49 8.77 ;
      RECT 25.075 1.4 25.245 1.57 ;
      RECT 25.075 10.89 25.245 11.06 ;
      RECT 24.395 1.4 24.565 1.57 ;
      RECT 24.395 10.89 24.565 11.06 ;
      RECT 22.78 2.61 22.95 2.78 ;
      RECT 22.525 3.97 22.695 4.14 ;
      RECT 22.32 2.61 22.49 2.78 ;
      RECT 22.045 3.13 22.215 3.3 ;
      RECT 21.86 2.61 22.03 2.78 ;
      RECT 21.805 3.69 21.975 3.86 ;
      RECT 21.4 2.61 21.57 2.78 ;
      RECT 21.325 3.69 21.495 3.86 ;
      RECT 21.085 3.13 21.255 3.3 ;
      RECT 21.085 4.81 21.255 4.98 ;
      RECT 20.94 2.61 21.11 2.78 ;
      RECT 20.82 10.89 20.99 11.06 ;
      RECT 20.565 3.97 20.735 4.14 ;
      RECT 20.51 8.97 20.68 9.14 ;
      RECT 20.48 2.61 20.65 2.78 ;
      RECT 20.325 3.41 20.495 3.58 ;
      RECT 20.14 10.89 20.31 11.06 ;
      RECT 20.085 4.81 20.255 4.98 ;
      RECT 20.08 9.34 20.25 9.51 ;
      RECT 20.08 10.08 20.25 10.25 ;
      RECT 20.02 2.61 20.19 2.78 ;
      RECT 19.845 3.97 20.015 4.14 ;
      RECT 19.705 8.6 19.875 8.77 ;
      RECT 19.56 2.61 19.73 2.78 ;
      RECT 19.46 10.89 19.63 11.06 ;
      RECT 19.365 3.69 19.535 3.86 ;
      RECT 19.1 2.61 19.27 2.78 ;
      RECT 18.885 3.69 19.055 3.86 ;
      RECT 18.78 10.89 18.95 11.06 ;
      RECT 18.645 3.13 18.815 3.3 ;
      RECT 18.64 2.61 18.81 2.78 ;
      RECT 18.18 2.61 18.35 2.78 ;
      RECT 17.885 3.41 18.055 3.58 ;
      RECT 17.72 2.61 17.89 2.78 ;
      RECT 17.645 4.53 17.815 4.7 ;
      RECT 17.405 3.97 17.575 4.14 ;
      RECT 17.26 2.61 17.43 2.78 ;
      RECT 16.925 3.69 17.095 3.86 ;
      RECT 16.8 2.61 16.97 2.78 ;
      RECT 16.685 3.13 16.855 3.3 ;
      RECT 16.685 4.53 16.855 4.7 ;
      RECT 16.34 2.61 16.51 2.78 ;
      RECT 16.205 4.25 16.375 4.42 ;
      RECT 15.88 2.61 16.05 2.78 ;
      RECT 15.685 3.69 15.855 3.86 ;
      RECT 15.445 4.53 15.615 4.7 ;
      RECT 15.42 2.61 15.59 2.78 ;
      RECT 15.205 3.13 15.375 3.3 ;
      RECT 14.965 3.69 15.135 3.86 ;
      RECT 14.965 4.25 15.135 4.42 ;
      RECT 14.96 2.61 15.13 2.78 ;
      RECT 14.5 2.61 14.67 2.78 ;
      RECT 14.245 3.13 14.415 3.3 ;
      RECT 14.245 4.81 14.415 4.98 ;
      RECT 14.04 2.61 14.21 2.78 ;
      RECT 13.765 4.25 13.935 4.42 ;
      RECT 13.58 2.61 13.75 2.78 ;
      RECT 12.24 10.89 12.41 11.06 ;
      RECT 11.56 10.89 11.73 11.06 ;
      RECT 11.5 9.34 11.67 9.51 ;
      RECT 11.5 10.08 11.67 10.25 ;
      RECT 11.125 8.6 11.295 8.77 ;
      RECT 10.88 10.89 11.05 11.06 ;
      RECT 10.2 10.89 10.37 11.06 ;
    LAYER li1 ;
      RECT 9.9 10.86 94.325 12.46 ;
      RECT 93.345 10.235 93.515 12.46 ;
      RECT 92.355 10.235 92.525 12.46 ;
      RECT 89.615 10.23 89.785 12.46 ;
      RECT 84 10.23 84.17 12.46 ;
      RECT 77.02 10.235 77.19 12.46 ;
      RECT 76.03 10.235 76.2 12.46 ;
      RECT 73.29 10.23 73.46 12.46 ;
      RECT 67.675 10.23 67.845 12.46 ;
      RECT 60.695 10.235 60.865 12.46 ;
      RECT 59.705 10.235 59.875 12.46 ;
      RECT 56.965 10.23 57.135 12.46 ;
      RECT 51.35 10.23 51.52 12.46 ;
      RECT 44.37 10.235 44.54 12.46 ;
      RECT 43.38 10.235 43.55 12.46 ;
      RECT 40.64 10.23 40.81 12.46 ;
      RECT 35.025 10.23 35.195 12.46 ;
      RECT 28.045 10.235 28.215 12.46 ;
      RECT 27.055 10.235 27.225 12.46 ;
      RECT 24.315 10.23 24.485 12.46 ;
      RECT 18.7 10.23 18.87 12.46 ;
      RECT 9.905 10.85 10.71 12.46 ;
      RECT 10.12 10.83 10.37 12.46 ;
      RECT 10.12 10.23 10.29 12.46 ;
      RECT 86.865 0 87.035 3.28 ;
      RECT 84.905 0 85.075 3.28 ;
      RECT 82.465 0 82.635 3.28 ;
      RECT 81.505 0 81.675 3.28 ;
      RECT 80.985 0 81.155 3.28 ;
      RECT 80.025 0 80.195 3.28 ;
      RECT 79.065 0 79.235 3.28 ;
      RECT 70.54 0 70.71 3.28 ;
      RECT 68.58 0 68.75 3.28 ;
      RECT 66.14 0 66.31 3.28 ;
      RECT 65.18 0 65.35 3.28 ;
      RECT 64.66 0 64.83 3.28 ;
      RECT 63.7 0 63.87 3.28 ;
      RECT 62.74 0 62.91 3.28 ;
      RECT 54.215 0 54.385 3.28 ;
      RECT 52.255 0 52.425 3.28 ;
      RECT 49.815 0 49.985 3.28 ;
      RECT 48.855 0 49.025 3.28 ;
      RECT 48.335 0 48.505 3.28 ;
      RECT 47.375 0 47.545 3.28 ;
      RECT 46.415 0 46.585 3.28 ;
      RECT 37.89 0 38.06 3.28 ;
      RECT 35.93 0 36.1 3.28 ;
      RECT 33.49 0 33.66 3.28 ;
      RECT 32.53 0 32.7 3.28 ;
      RECT 32.01 0 32.18 3.28 ;
      RECT 31.05 0 31.22 3.28 ;
      RECT 30.09 0 30.26 3.28 ;
      RECT 21.565 0 21.735 3.28 ;
      RECT 19.605 0 19.775 3.28 ;
      RECT 17.165 0 17.335 3.28 ;
      RECT 16.205 0 16.375 3.28 ;
      RECT 15.685 0 15.855 3.28 ;
      RECT 14.725 0 14.895 3.28 ;
      RECT 13.765 0 13.935 3.28 ;
      RECT 84.835 0 85.075 2.89 ;
      RECT 81.16 0 81.355 2.89 ;
      RECT 78.86 0 79.055 2.89 ;
      RECT 68.51 0 68.75 2.89 ;
      RECT 64.835 0 65.03 2.89 ;
      RECT 62.535 0 62.73 2.89 ;
      RECT 52.185 0 52.425 2.89 ;
      RECT 48.51 0 48.705 2.89 ;
      RECT 46.21 0 46.405 2.89 ;
      RECT 35.86 0 36.1 2.89 ;
      RECT 32.185 0 32.38 2.89 ;
      RECT 29.885 0 30.08 2.89 ;
      RECT 19.535 0 19.775 2.89 ;
      RECT 15.86 0 16.055 2.89 ;
      RECT 13.56 0 13.755 2.89 ;
      RECT 88.36 0 88.55 2.88 ;
      RECT 72.035 0 72.225 2.88 ;
      RECT 55.71 0 55.9 2.88 ;
      RECT 39.385 0 39.575 2.88 ;
      RECT 23.06 0 23.25 2.88 ;
      RECT 86.685 0 87.035 2.865 ;
      RECT 70.36 0 70.71 2.865 ;
      RECT 54.035 0 54.385 2.865 ;
      RECT 37.71 0 38.06 2.865 ;
      RECT 21.385 0 21.735 2.865 ;
      RECT 88.355 0 88.55 2.86 ;
      RECT 82.995 0 83.19 2.86 ;
      RECT 72.03 0 72.225 2.86 ;
      RECT 66.67 0 66.865 2.86 ;
      RECT 55.705 0 55.9 2.86 ;
      RECT 50.345 0 50.54 2.86 ;
      RECT 39.38 0 39.575 2.86 ;
      RECT 34.02 0 34.215 2.86 ;
      RECT 23.055 0 23.25 2.86 ;
      RECT 17.695 0 17.89 2.86 ;
      RECT 78.735 0 88.55 2.78 ;
      RECT 62.41 0 72.225 2.78 ;
      RECT 46.085 0 55.9 2.78 ;
      RECT 29.76 0 39.575 2.78 ;
      RECT 13.435 0 23.25 2.78 ;
      RECT 89.615 0 89.785 2.23 ;
      RECT 73.29 0 73.46 2.23 ;
      RECT 56.965 0 57.135 2.23 ;
      RECT 40.64 0 40.81 2.23 ;
      RECT 24.315 0 24.485 2.23 ;
      RECT 93.345 0 93.515 2.225 ;
      RECT 92.355 0 92.525 2.225 ;
      RECT 77.02 0 77.19 2.225 ;
      RECT 76.03 0 76.2 2.225 ;
      RECT 60.695 0 60.865 2.225 ;
      RECT 59.705 0 59.875 2.225 ;
      RECT 44.37 0 44.54 2.225 ;
      RECT 43.38 0 43.55 2.225 ;
      RECT 28.045 0 28.215 2.225 ;
      RECT 27.055 0 27.225 2.225 ;
      RECT 9.9 0 94.32 1.6 ;
      RECT 93.775 7.305 93.945 8.775 ;
      RECT 93.775 8.6 93.95 8.77 ;
      RECT 93.405 3.035 93.575 4.225 ;
      RECT 93.405 3.035 93.875 3.205 ;
      RECT 93.405 9.255 93.875 9.425 ;
      RECT 93.405 8.235 93.575 9.425 ;
      RECT 92.415 3.035 92.585 4.225 ;
      RECT 92.415 3.035 92.885 3.205 ;
      RECT 92.415 9.255 92.885 9.425 ;
      RECT 92.415 8.235 92.585 9.425 ;
      RECT 90.565 3.93 90.735 5.16 ;
      RECT 90.62 2.15 90.79 4.1 ;
      RECT 90.565 1.87 90.735 2.32 ;
      RECT 90.565 10.14 90.735 10.59 ;
      RECT 90.62 8.36 90.79 10.31 ;
      RECT 90.565 7.3 90.735 8.53 ;
      RECT 90.045 1.87 90.215 5.16 ;
      RECT 90.045 3.37 90.45 3.7 ;
      RECT 90.045 2.53 90.45 2.86 ;
      RECT 90.045 7.3 90.215 10.59 ;
      RECT 90.045 9.6 90.45 9.93 ;
      RECT 90.045 8.76 90.45 9.09 ;
      RECT 87.345 3.03 87.515 3.3 ;
      RECT 87.345 3.03 88.075 3.2 ;
      RECT 87.825 3.77 87.995 4.14 ;
      RECT 87.505 3.77 87.995 3.94 ;
      RECT 87.265 4.42 87.595 4.59 ;
      RECT 86.505 4.25 87.515 4.42 ;
      RECT 86.505 3.77 86.675 4.42 ;
      RECT 86.625 3.69 86.795 4.02 ;
      RECT 85.785 4.42 86.115 4.59 ;
      RECT 83.865 4.42 85.155 4.59 ;
      RECT 84.905 4.335 86.035 4.505 ;
      RECT 85.625 3.41 86.035 3.58 ;
      RECT 85.865 2.95 86.035 3.58 ;
      RECT 85.865 3.77 86.035 4.14 ;
      RECT 85.545 3.77 86.035 3.94 ;
      RECT 84.95 10.14 85.12 10.59 ;
      RECT 85.005 8.36 85.175 10.31 ;
      RECT 84.95 7.3 85.12 8.53 ;
      RECT 84.43 7.3 84.6 10.59 ;
      RECT 84.43 9.6 84.835 9.93 ;
      RECT 84.43 8.76 84.835 9.09 ;
      RECT 83.105 3.77 84.435 3.94 ;
      RECT 84.185 3.69 84.355 3.94 ;
      RECT 83.185 3.37 83.355 3.58 ;
      RECT 83.185 3.37 83.675 3.54 ;
      RECT 81.865 4.53 82.155 4.7 ;
      RECT 81.865 3.77 82.035 4.7 ;
      RECT 81.665 3.77 82.035 3.94 ;
      RECT 80.665 3.77 81.155 3.94 ;
      RECT 80.985 3.69 81.155 3.94 ;
      RECT 80.745 4.53 81.155 4.7 ;
      RECT 80.985 4.34 81.155 4.7 ;
      RECT 79.785 4.25 80.435 4.42 ;
      RECT 79.785 3.69 79.955 4.42 ;
      RECT 79.425 4.81 79.715 4.98 ;
      RECT 79.425 3.77 79.595 4.98 ;
      RECT 79.225 3.77 79.595 3.94 ;
      RECT 77.45 7.305 77.62 8.775 ;
      RECT 77.45 8.6 77.625 8.77 ;
      RECT 77.08 3.035 77.25 4.225 ;
      RECT 77.08 3.035 77.55 3.205 ;
      RECT 77.08 9.255 77.55 9.425 ;
      RECT 77.08 8.235 77.25 9.425 ;
      RECT 76.09 3.035 76.26 4.225 ;
      RECT 76.09 3.035 76.56 3.205 ;
      RECT 76.09 9.255 76.56 9.425 ;
      RECT 76.09 8.235 76.26 9.425 ;
      RECT 74.24 3.93 74.41 5.16 ;
      RECT 74.295 2.15 74.465 4.1 ;
      RECT 74.24 1.87 74.41 2.32 ;
      RECT 74.24 10.14 74.41 10.59 ;
      RECT 74.295 8.36 74.465 10.31 ;
      RECT 74.24 7.3 74.41 8.53 ;
      RECT 73.72 1.87 73.89 5.16 ;
      RECT 73.72 3.37 74.125 3.7 ;
      RECT 73.72 2.53 74.125 2.86 ;
      RECT 73.72 7.3 73.89 10.59 ;
      RECT 73.72 9.6 74.125 9.93 ;
      RECT 73.72 8.76 74.125 9.09 ;
      RECT 71.02 3.03 71.19 3.3 ;
      RECT 71.02 3.03 71.75 3.2 ;
      RECT 71.5 3.77 71.67 4.14 ;
      RECT 71.18 3.77 71.67 3.94 ;
      RECT 70.94 4.42 71.27 4.59 ;
      RECT 70.18 4.25 71.19 4.42 ;
      RECT 70.18 3.77 70.35 4.42 ;
      RECT 70.3 3.69 70.47 4.02 ;
      RECT 69.46 4.42 69.79 4.59 ;
      RECT 67.54 4.42 68.83 4.59 ;
      RECT 68.58 4.335 69.71 4.505 ;
      RECT 69.3 3.41 69.71 3.58 ;
      RECT 69.54 2.95 69.71 3.58 ;
      RECT 69.54 3.77 69.71 4.14 ;
      RECT 69.22 3.77 69.71 3.94 ;
      RECT 68.625 10.14 68.795 10.59 ;
      RECT 68.68 8.36 68.85 10.31 ;
      RECT 68.625 7.3 68.795 8.53 ;
      RECT 68.105 7.3 68.275 10.59 ;
      RECT 68.105 9.6 68.51 9.93 ;
      RECT 68.105 8.76 68.51 9.09 ;
      RECT 66.78 3.77 68.11 3.94 ;
      RECT 67.86 3.69 68.03 3.94 ;
      RECT 66.86 3.37 67.03 3.58 ;
      RECT 66.86 3.37 67.35 3.54 ;
      RECT 65.54 4.53 65.83 4.7 ;
      RECT 65.54 3.77 65.71 4.7 ;
      RECT 65.34 3.77 65.71 3.94 ;
      RECT 64.34 3.77 64.83 3.94 ;
      RECT 64.66 3.69 64.83 3.94 ;
      RECT 64.42 4.53 64.83 4.7 ;
      RECT 64.66 4.34 64.83 4.7 ;
      RECT 63.46 4.25 64.11 4.42 ;
      RECT 63.46 3.69 63.63 4.42 ;
      RECT 63.1 4.81 63.39 4.98 ;
      RECT 63.1 3.77 63.27 4.98 ;
      RECT 62.9 3.77 63.27 3.94 ;
      RECT 61.125 7.305 61.295 8.775 ;
      RECT 61.125 8.6 61.3 8.77 ;
      RECT 60.755 3.035 60.925 4.225 ;
      RECT 60.755 3.035 61.225 3.205 ;
      RECT 60.755 9.255 61.225 9.425 ;
      RECT 60.755 8.235 60.925 9.425 ;
      RECT 59.765 3.035 59.935 4.225 ;
      RECT 59.765 3.035 60.235 3.205 ;
      RECT 59.765 9.255 60.235 9.425 ;
      RECT 59.765 8.235 59.935 9.425 ;
      RECT 57.915 3.93 58.085 5.16 ;
      RECT 57.97 2.15 58.14 4.1 ;
      RECT 57.915 1.87 58.085 2.32 ;
      RECT 57.915 10.14 58.085 10.59 ;
      RECT 57.97 8.36 58.14 10.31 ;
      RECT 57.915 7.3 58.085 8.53 ;
      RECT 57.395 1.87 57.565 5.16 ;
      RECT 57.395 3.37 57.8 3.7 ;
      RECT 57.395 2.53 57.8 2.86 ;
      RECT 57.395 7.3 57.565 10.59 ;
      RECT 57.395 9.6 57.8 9.93 ;
      RECT 57.395 8.76 57.8 9.09 ;
      RECT 54.695 3.03 54.865 3.3 ;
      RECT 54.695 3.03 55.425 3.2 ;
      RECT 55.175 3.77 55.345 4.14 ;
      RECT 54.855 3.77 55.345 3.94 ;
      RECT 54.615 4.42 54.945 4.59 ;
      RECT 53.855 4.25 54.865 4.42 ;
      RECT 53.855 3.77 54.025 4.42 ;
      RECT 53.975 3.69 54.145 4.02 ;
      RECT 53.135 4.42 53.465 4.59 ;
      RECT 51.215 4.42 52.505 4.59 ;
      RECT 52.255 4.335 53.385 4.505 ;
      RECT 52.975 3.41 53.385 3.58 ;
      RECT 53.215 2.95 53.385 3.58 ;
      RECT 53.215 3.77 53.385 4.14 ;
      RECT 52.895 3.77 53.385 3.94 ;
      RECT 52.3 10.14 52.47 10.59 ;
      RECT 52.355 8.36 52.525 10.31 ;
      RECT 52.3 7.3 52.47 8.53 ;
      RECT 51.78 7.3 51.95 10.59 ;
      RECT 51.78 9.6 52.185 9.93 ;
      RECT 51.78 8.76 52.185 9.09 ;
      RECT 50.455 3.77 51.785 3.94 ;
      RECT 51.535 3.69 51.705 3.94 ;
      RECT 50.535 3.37 50.705 3.58 ;
      RECT 50.535 3.37 51.025 3.54 ;
      RECT 49.215 4.53 49.505 4.7 ;
      RECT 49.215 3.77 49.385 4.7 ;
      RECT 49.015 3.77 49.385 3.94 ;
      RECT 48.015 3.77 48.505 3.94 ;
      RECT 48.335 3.69 48.505 3.94 ;
      RECT 48.095 4.53 48.505 4.7 ;
      RECT 48.335 4.34 48.505 4.7 ;
      RECT 47.135 4.25 47.785 4.42 ;
      RECT 47.135 3.69 47.305 4.42 ;
      RECT 46.775 4.81 47.065 4.98 ;
      RECT 46.775 3.77 46.945 4.98 ;
      RECT 46.575 3.77 46.945 3.94 ;
      RECT 44.8 7.305 44.97 8.775 ;
      RECT 44.8 8.6 44.975 8.77 ;
      RECT 44.43 3.035 44.6 4.225 ;
      RECT 44.43 3.035 44.9 3.205 ;
      RECT 44.43 9.255 44.9 9.425 ;
      RECT 44.43 8.235 44.6 9.425 ;
      RECT 43.44 3.035 43.61 4.225 ;
      RECT 43.44 3.035 43.91 3.205 ;
      RECT 43.44 9.255 43.91 9.425 ;
      RECT 43.44 8.235 43.61 9.425 ;
      RECT 41.59 3.93 41.76 5.16 ;
      RECT 41.645 2.15 41.815 4.1 ;
      RECT 41.59 1.87 41.76 2.32 ;
      RECT 41.59 10.14 41.76 10.59 ;
      RECT 41.645 8.36 41.815 10.31 ;
      RECT 41.59 7.3 41.76 8.53 ;
      RECT 41.07 1.87 41.24 5.16 ;
      RECT 41.07 3.37 41.475 3.7 ;
      RECT 41.07 2.53 41.475 2.86 ;
      RECT 41.07 7.3 41.24 10.59 ;
      RECT 41.07 9.6 41.475 9.93 ;
      RECT 41.07 8.76 41.475 9.09 ;
      RECT 38.37 3.03 38.54 3.3 ;
      RECT 38.37 3.03 39.1 3.2 ;
      RECT 38.85 3.77 39.02 4.14 ;
      RECT 38.53 3.77 39.02 3.94 ;
      RECT 38.29 4.42 38.62 4.59 ;
      RECT 37.53 4.25 38.54 4.42 ;
      RECT 37.53 3.77 37.7 4.42 ;
      RECT 37.65 3.69 37.82 4.02 ;
      RECT 36.81 4.42 37.14 4.59 ;
      RECT 34.89 4.42 36.18 4.59 ;
      RECT 35.93 4.335 37.06 4.505 ;
      RECT 36.65 3.41 37.06 3.58 ;
      RECT 36.89 2.95 37.06 3.58 ;
      RECT 36.89 3.77 37.06 4.14 ;
      RECT 36.57 3.77 37.06 3.94 ;
      RECT 35.975 10.14 36.145 10.59 ;
      RECT 36.03 8.36 36.2 10.31 ;
      RECT 35.975 7.3 36.145 8.53 ;
      RECT 35.455 7.3 35.625 10.59 ;
      RECT 35.455 9.6 35.86 9.93 ;
      RECT 35.455 8.76 35.86 9.09 ;
      RECT 34.13 3.77 35.46 3.94 ;
      RECT 35.21 3.69 35.38 3.94 ;
      RECT 34.21 3.37 34.38 3.58 ;
      RECT 34.21 3.37 34.7 3.54 ;
      RECT 32.89 4.53 33.18 4.7 ;
      RECT 32.89 3.77 33.06 4.7 ;
      RECT 32.69 3.77 33.06 3.94 ;
      RECT 31.69 3.77 32.18 3.94 ;
      RECT 32.01 3.69 32.18 3.94 ;
      RECT 31.77 4.53 32.18 4.7 ;
      RECT 32.01 4.34 32.18 4.7 ;
      RECT 30.81 4.25 31.46 4.42 ;
      RECT 30.81 3.69 30.98 4.42 ;
      RECT 30.45 4.81 30.74 4.98 ;
      RECT 30.45 3.77 30.62 4.98 ;
      RECT 30.25 3.77 30.62 3.94 ;
      RECT 28.475 7.305 28.645 8.775 ;
      RECT 28.475 8.6 28.65 8.77 ;
      RECT 28.105 3.035 28.275 4.225 ;
      RECT 28.105 3.035 28.575 3.205 ;
      RECT 28.105 9.255 28.575 9.425 ;
      RECT 28.105 8.235 28.275 9.425 ;
      RECT 27.115 3.035 27.285 4.225 ;
      RECT 27.115 3.035 27.585 3.205 ;
      RECT 27.115 9.255 27.585 9.425 ;
      RECT 27.115 8.235 27.285 9.425 ;
      RECT 25.265 3.93 25.435 5.16 ;
      RECT 25.32 2.15 25.49 4.1 ;
      RECT 25.265 1.87 25.435 2.32 ;
      RECT 25.265 10.14 25.435 10.59 ;
      RECT 25.32 8.36 25.49 10.31 ;
      RECT 25.265 7.3 25.435 8.53 ;
      RECT 24.745 1.87 24.915 5.16 ;
      RECT 24.745 3.37 25.15 3.7 ;
      RECT 24.745 2.53 25.15 2.86 ;
      RECT 24.745 7.3 24.915 10.59 ;
      RECT 24.745 9.6 25.15 9.93 ;
      RECT 24.745 8.76 25.15 9.09 ;
      RECT 22.045 3.03 22.215 3.3 ;
      RECT 22.045 3.03 22.775 3.2 ;
      RECT 22.525 3.77 22.695 4.14 ;
      RECT 22.205 3.77 22.695 3.94 ;
      RECT 21.965 4.42 22.295 4.59 ;
      RECT 21.205 4.25 22.215 4.42 ;
      RECT 21.205 3.77 21.375 4.42 ;
      RECT 21.325 3.69 21.495 4.02 ;
      RECT 20.485 4.42 20.815 4.59 ;
      RECT 18.565 4.42 19.855 4.59 ;
      RECT 19.605 4.335 20.735 4.505 ;
      RECT 20.325 3.41 20.735 3.58 ;
      RECT 20.565 2.95 20.735 3.58 ;
      RECT 20.565 3.77 20.735 4.14 ;
      RECT 20.245 3.77 20.735 3.94 ;
      RECT 19.65 10.14 19.82 10.59 ;
      RECT 19.705 8.36 19.875 10.31 ;
      RECT 19.65 7.3 19.82 8.53 ;
      RECT 19.13 7.3 19.3 10.59 ;
      RECT 19.13 9.6 19.535 9.93 ;
      RECT 19.13 8.76 19.535 9.09 ;
      RECT 17.805 3.77 19.135 3.94 ;
      RECT 18.885 3.69 19.055 3.94 ;
      RECT 17.885 3.37 18.055 3.58 ;
      RECT 17.885 3.37 18.375 3.54 ;
      RECT 16.565 4.53 16.855 4.7 ;
      RECT 16.565 3.77 16.735 4.7 ;
      RECT 16.365 3.77 16.735 3.94 ;
      RECT 15.365 3.77 15.855 3.94 ;
      RECT 15.685 3.69 15.855 3.94 ;
      RECT 15.445 4.53 15.855 4.7 ;
      RECT 15.685 4.34 15.855 4.7 ;
      RECT 14.485 4.25 15.135 4.42 ;
      RECT 14.485 3.69 14.655 4.42 ;
      RECT 14.125 4.81 14.415 4.98 ;
      RECT 14.125 3.77 14.295 4.98 ;
      RECT 13.925 3.77 14.295 3.94 ;
      RECT 11.07 10.14 11.24 10.59 ;
      RECT 11.125 8.36 11.295 10.31 ;
      RECT 11.07 7.3 11.24 8.53 ;
      RECT 10.55 7.3 10.72 10.59 ;
      RECT 10.55 9.6 10.955 9.93 ;
      RECT 10.55 8.76 10.955 9.09 ;
      RECT 93.775 10.085 93.945 10.595 ;
      RECT 92.785 1.865 92.955 2.375 ;
      RECT 92.785 3.685 92.955 5.155 ;
      RECT 92.785 7.305 92.955 8.775 ;
      RECT 92.785 10.085 92.955 10.595 ;
      RECT 91.425 1.87 91.595 5.16 ;
      RECT 91.425 7.3 91.595 10.59 ;
      RECT 90.995 1.87 91.165 2.38 ;
      RECT 90.995 2.95 91.165 5.16 ;
      RECT 90.995 7.3 91.165 9.51 ;
      RECT 90.995 10.08 91.165 10.59 ;
      RECT 87.105 3.69 87.275 4.02 ;
      RECT 86.385 2.95 86.555 3.3 ;
      RECT 86.385 4.68 86.555 5.01 ;
      RECT 85.81 7.3 85.98 10.59 ;
      RECT 85.385 4.68 85.555 5.01 ;
      RECT 85.38 7.3 85.55 9.51 ;
      RECT 85.38 10.08 85.55 10.59 ;
      RECT 85.145 3.69 85.315 4.14 ;
      RECT 84.665 3.69 84.835 4.02 ;
      RECT 83.945 2.95 84.115 3.3 ;
      RECT 83.285 2.86 83.48 2.89 ;
      RECT 82.945 4.34 83.115 4.7 ;
      RECT 82.705 3.69 82.875 4.14 ;
      RECT 82.225 3.69 82.395 4.02 ;
      RECT 81.985 2.95 82.155 3.3 ;
      RECT 81.505 4.25 81.675 4.67 ;
      RECT 80.505 2.95 80.675 3.3 ;
      RECT 80.265 3.69 80.435 4.02 ;
      RECT 79.545 2.95 79.715 3.3 ;
      RECT 79.065 4.25 79.235 4.67 ;
      RECT 77.45 10.085 77.62 10.595 ;
      RECT 76.46 1.865 76.63 2.375 ;
      RECT 76.46 3.685 76.63 5.155 ;
      RECT 76.46 7.305 76.63 8.775 ;
      RECT 76.46 10.085 76.63 10.595 ;
      RECT 75.1 1.87 75.27 5.16 ;
      RECT 75.1 7.3 75.27 10.59 ;
      RECT 74.67 1.87 74.84 2.38 ;
      RECT 74.67 2.95 74.84 5.16 ;
      RECT 74.67 7.3 74.84 9.51 ;
      RECT 74.67 10.08 74.84 10.59 ;
      RECT 70.78 3.69 70.95 4.02 ;
      RECT 70.06 2.95 70.23 3.3 ;
      RECT 70.06 4.68 70.23 5.01 ;
      RECT 69.485 7.3 69.655 10.59 ;
      RECT 69.06 4.68 69.23 5.01 ;
      RECT 69.055 7.3 69.225 9.51 ;
      RECT 69.055 10.08 69.225 10.59 ;
      RECT 68.82 3.69 68.99 4.14 ;
      RECT 68.34 3.69 68.51 4.02 ;
      RECT 67.62 2.95 67.79 3.3 ;
      RECT 66.96 2.86 67.155 2.89 ;
      RECT 66.62 4.34 66.79 4.7 ;
      RECT 66.38 3.69 66.55 4.14 ;
      RECT 65.9 3.69 66.07 4.02 ;
      RECT 65.66 2.95 65.83 3.3 ;
      RECT 65.18 4.25 65.35 4.67 ;
      RECT 64.18 2.95 64.35 3.3 ;
      RECT 63.94 3.69 64.11 4.02 ;
      RECT 63.22 2.95 63.39 3.3 ;
      RECT 62.74 4.25 62.91 4.67 ;
      RECT 61.125 10.085 61.295 10.595 ;
      RECT 60.135 1.865 60.305 2.375 ;
      RECT 60.135 3.685 60.305 5.155 ;
      RECT 60.135 7.305 60.305 8.775 ;
      RECT 60.135 10.085 60.305 10.595 ;
      RECT 58.775 1.87 58.945 5.16 ;
      RECT 58.775 7.3 58.945 10.59 ;
      RECT 58.345 1.87 58.515 2.38 ;
      RECT 58.345 2.95 58.515 5.16 ;
      RECT 58.345 7.3 58.515 9.51 ;
      RECT 58.345 10.08 58.515 10.59 ;
      RECT 54.455 3.69 54.625 4.02 ;
      RECT 53.735 2.95 53.905 3.3 ;
      RECT 53.735 4.68 53.905 5.01 ;
      RECT 53.16 7.3 53.33 10.59 ;
      RECT 52.735 4.68 52.905 5.01 ;
      RECT 52.73 7.3 52.9 9.51 ;
      RECT 52.73 10.08 52.9 10.59 ;
      RECT 52.495 3.69 52.665 4.14 ;
      RECT 52.015 3.69 52.185 4.02 ;
      RECT 51.295 2.95 51.465 3.3 ;
      RECT 50.635 2.86 50.83 2.89 ;
      RECT 50.295 4.34 50.465 4.7 ;
      RECT 50.055 3.69 50.225 4.14 ;
      RECT 49.575 3.69 49.745 4.02 ;
      RECT 49.335 2.95 49.505 3.3 ;
      RECT 48.855 4.25 49.025 4.67 ;
      RECT 47.855 2.95 48.025 3.3 ;
      RECT 47.615 3.69 47.785 4.02 ;
      RECT 46.895 2.95 47.065 3.3 ;
      RECT 46.415 4.25 46.585 4.67 ;
      RECT 44.8 10.085 44.97 10.595 ;
      RECT 43.81 1.865 43.98 2.375 ;
      RECT 43.81 3.685 43.98 5.155 ;
      RECT 43.81 7.305 43.98 8.775 ;
      RECT 43.81 10.085 43.98 10.595 ;
      RECT 42.45 1.87 42.62 5.16 ;
      RECT 42.45 7.3 42.62 10.59 ;
      RECT 42.02 1.87 42.19 2.38 ;
      RECT 42.02 2.95 42.19 5.16 ;
      RECT 42.02 7.3 42.19 9.51 ;
      RECT 42.02 10.08 42.19 10.59 ;
      RECT 38.13 3.69 38.3 4.02 ;
      RECT 37.41 2.95 37.58 3.3 ;
      RECT 37.41 4.68 37.58 5.01 ;
      RECT 36.835 7.3 37.005 10.59 ;
      RECT 36.41 4.68 36.58 5.01 ;
      RECT 36.405 7.3 36.575 9.51 ;
      RECT 36.405 10.08 36.575 10.59 ;
      RECT 36.17 3.69 36.34 4.14 ;
      RECT 35.69 3.69 35.86 4.02 ;
      RECT 34.97 2.95 35.14 3.3 ;
      RECT 34.31 2.86 34.505 2.89 ;
      RECT 33.97 4.34 34.14 4.7 ;
      RECT 33.73 3.69 33.9 4.14 ;
      RECT 33.25 3.69 33.42 4.02 ;
      RECT 33.01 2.95 33.18 3.3 ;
      RECT 32.53 4.25 32.7 4.67 ;
      RECT 31.53 2.95 31.7 3.3 ;
      RECT 31.29 3.69 31.46 4.02 ;
      RECT 30.57 2.95 30.74 3.3 ;
      RECT 30.09 4.25 30.26 4.67 ;
      RECT 28.475 10.085 28.645 10.595 ;
      RECT 27.485 1.865 27.655 2.375 ;
      RECT 27.485 3.685 27.655 5.155 ;
      RECT 27.485 7.305 27.655 8.775 ;
      RECT 27.485 10.085 27.655 10.595 ;
      RECT 26.125 1.87 26.295 5.16 ;
      RECT 26.125 7.3 26.295 10.59 ;
      RECT 25.695 1.87 25.865 2.38 ;
      RECT 25.695 2.95 25.865 5.16 ;
      RECT 25.695 7.3 25.865 9.51 ;
      RECT 25.695 10.08 25.865 10.59 ;
      RECT 21.805 3.69 21.975 4.02 ;
      RECT 21.085 2.95 21.255 3.3 ;
      RECT 21.085 4.68 21.255 5.01 ;
      RECT 20.51 7.3 20.68 10.59 ;
      RECT 20.085 4.68 20.255 5.01 ;
      RECT 20.08 7.3 20.25 9.51 ;
      RECT 20.08 10.08 20.25 10.59 ;
      RECT 19.845 3.69 20.015 4.14 ;
      RECT 19.365 3.69 19.535 4.02 ;
      RECT 18.645 2.95 18.815 3.3 ;
      RECT 17.985 2.86 18.18 2.89 ;
      RECT 17.645 4.34 17.815 4.7 ;
      RECT 17.405 3.69 17.575 4.14 ;
      RECT 16.925 3.69 17.095 4.02 ;
      RECT 16.685 2.95 16.855 3.3 ;
      RECT 16.205 4.25 16.375 4.67 ;
      RECT 15.205 2.95 15.375 3.3 ;
      RECT 14.965 3.69 15.135 4.02 ;
      RECT 14.245 2.95 14.415 3.3 ;
      RECT 13.765 4.25 13.935 4.67 ;
      RECT 11.5 7.3 11.67 9.51 ;
      RECT 11.5 10.08 11.67 10.59 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  ORIGIN -12.125 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r1 ;
  SIZE 95.615 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 32.94 1.87 33.11 2.38 ;
        RECT 32.94 3.69 33.11 5.16 ;
      LAYER met1 ;
        RECT 32.88 3.66 33.17 3.89 ;
        RECT 32.88 2.18 33.17 2.41 ;
        RECT 32.94 2.18 33.11 3.89 ;
      LAYER mcon ;
        RECT 32.94 3.69 33.11 3.86 ;
        RECT 32.94 2.21 33.11 2.38 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 51.5 1.87 51.67 2.38 ;
        RECT 51.5 3.69 51.67 5.16 ;
      LAYER met1 ;
        RECT 51.44 3.66 51.73 3.89 ;
        RECT 51.44 2.18 51.73 2.41 ;
        RECT 51.5 2.18 51.67 3.89 ;
      LAYER mcon ;
        RECT 51.5 3.69 51.67 3.86 ;
        RECT 51.5 2.21 51.67 2.38 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 70.06 1.87 70.23 2.38 ;
        RECT 70.06 3.69 70.23 5.16 ;
      LAYER met1 ;
        RECT 70 3.66 70.29 3.89 ;
        RECT 70 2.18 70.29 2.41 ;
        RECT 70.06 2.18 70.23 3.89 ;
      LAYER mcon ;
        RECT 70.06 3.69 70.23 3.86 ;
        RECT 70.06 2.21 70.23 2.38 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 88.62 1.87 88.79 2.38 ;
        RECT 88.62 3.69 88.79 5.16 ;
      LAYER met1 ;
        RECT 88.56 3.66 88.85 3.89 ;
        RECT 88.56 2.18 88.85 2.41 ;
        RECT 88.62 2.18 88.79 3.89 ;
      LAYER mcon ;
        RECT 88.62 3.69 88.79 3.86 ;
        RECT 88.62 2.21 88.79 2.38 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 107.18 1.87 107.35 2.38 ;
        RECT 107.18 3.69 107.35 5.16 ;
      LAYER met1 ;
        RECT 107.12 3.66 107.41 3.89 ;
        RECT 107.12 2.18 107.41 2.41 ;
        RECT 107.18 2.18 107.35 3.89 ;
      LAYER mcon ;
        RECT 107.18 3.69 107.35 3.86 ;
        RECT 107.18 2.21 107.35 2.38 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 28.79 2.955 28.96 4.23 ;
        RECT 28.79 8.235 28.96 9.51 ;
        RECT 23.175 8.235 23.345 9.51 ;
      LAYER met2 ;
        RECT 28.715 4 29.055 4.35 ;
        RECT 28.705 8.135 29.045 8.485 ;
        RECT 28.79 4 28.96 8.485 ;
      LAYER met1 ;
        RECT 28.715 4.06 29.19 4.23 ;
        RECT 28.715 4 29.055 4.35 ;
        RECT 23.115 8.235 29.19 8.405 ;
        RECT 28.705 8.135 29.045 8.485 ;
        RECT 23.115 8.205 23.405 8.435 ;
      LAYER via1 ;
        RECT 28.805 8.235 28.955 8.385 ;
        RECT 28.815 4.1 28.965 4.25 ;
      LAYER mcon ;
        RECT 23.175 8.235 23.345 8.405 ;
        RECT 28.79 8.235 28.96 8.405 ;
        RECT 28.79 4.06 28.96 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 47.35 2.955 47.52 4.23 ;
        RECT 47.35 8.235 47.52 9.51 ;
        RECT 41.735 8.235 41.905 9.51 ;
      LAYER met2 ;
        RECT 47.275 4 47.615 4.35 ;
        RECT 47.265 8.135 47.605 8.485 ;
        RECT 47.35 4 47.52 8.485 ;
      LAYER met1 ;
        RECT 47.275 4.06 47.75 4.23 ;
        RECT 47.275 4 47.615 4.35 ;
        RECT 41.675 8.235 47.75 8.405 ;
        RECT 47.265 8.135 47.605 8.485 ;
        RECT 41.675 8.205 41.965 8.435 ;
      LAYER via1 ;
        RECT 47.365 8.235 47.515 8.385 ;
        RECT 47.375 4.1 47.525 4.25 ;
      LAYER mcon ;
        RECT 41.735 8.235 41.905 8.405 ;
        RECT 47.35 8.235 47.52 8.405 ;
        RECT 47.35 4.06 47.52 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 65.91 2.955 66.08 4.23 ;
        RECT 65.91 8.235 66.08 9.51 ;
        RECT 60.295 8.235 60.465 9.51 ;
      LAYER met2 ;
        RECT 65.835 4 66.175 4.35 ;
        RECT 65.825 8.135 66.165 8.485 ;
        RECT 65.91 4 66.08 8.485 ;
      LAYER met1 ;
        RECT 65.835 4.06 66.31 4.23 ;
        RECT 65.835 4 66.175 4.35 ;
        RECT 60.235 8.235 66.31 8.405 ;
        RECT 65.825 8.135 66.165 8.485 ;
        RECT 60.235 8.205 60.525 8.435 ;
      LAYER via1 ;
        RECT 65.925 8.235 66.075 8.385 ;
        RECT 65.935 4.1 66.085 4.25 ;
      LAYER mcon ;
        RECT 60.295 8.235 60.465 8.405 ;
        RECT 65.91 8.235 66.08 8.405 ;
        RECT 65.91 4.06 66.08 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 84.47 2.955 84.64 4.23 ;
        RECT 84.47 8.235 84.64 9.51 ;
        RECT 78.855 8.235 79.025 9.51 ;
      LAYER met2 ;
        RECT 84.395 4 84.735 4.35 ;
        RECT 84.385 8.135 84.725 8.485 ;
        RECT 84.47 4 84.64 8.485 ;
      LAYER met1 ;
        RECT 84.395 4.06 84.87 4.23 ;
        RECT 84.395 4 84.735 4.35 ;
        RECT 78.795 8.235 84.87 8.405 ;
        RECT 84.385 8.135 84.725 8.485 ;
        RECT 78.795 8.205 79.085 8.435 ;
      LAYER via1 ;
        RECT 84.485 8.235 84.635 8.385 ;
        RECT 84.495 4.1 84.645 4.25 ;
      LAYER mcon ;
        RECT 78.855 8.235 79.025 8.405 ;
        RECT 84.47 8.235 84.64 8.405 ;
        RECT 84.47 4.06 84.64 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 103.03 2.955 103.2 4.23 ;
        RECT 103.03 8.235 103.2 9.51 ;
        RECT 97.415 8.235 97.585 9.51 ;
      LAYER met2 ;
        RECT 102.955 4 103.295 4.35 ;
        RECT 102.945 8.135 103.285 8.485 ;
        RECT 103.03 4 103.2 8.485 ;
      LAYER met1 ;
        RECT 102.955 4.06 103.43 4.23 ;
        RECT 102.955 4 103.295 4.35 ;
        RECT 97.355 8.235 103.43 8.405 ;
        RECT 102.945 8.135 103.285 8.485 ;
        RECT 97.355 8.205 97.645 8.435 ;
      LAYER via1 ;
        RECT 103.045 8.235 103.195 8.385 ;
        RECT 103.055 4.1 103.205 4.25 ;
      LAYER mcon ;
        RECT 97.415 8.235 97.585 8.405 ;
        RECT 103.03 8.235 103.2 8.405 ;
        RECT 103.03 4.06 103.2 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 12.36 8.235 12.53 9.51 ;
      LAYER met1 ;
        RECT 12.3 8.235 12.76 8.405 ;
        RECT 12.3 8.205 12.59 8.435 ;
      LAYER mcon ;
        RECT 12.36 8.235 12.53 8.405 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 91.525 3.71 92.255 4.04 ;
        RECT 72.965 3.71 73.695 4.04 ;
        RECT 54.405 3.71 55.135 4.04 ;
        RECT 35.845 3.71 36.575 4.04 ;
        RECT 17.285 3.71 18.015 4.04 ;
        RECT 12.135 10.79 12.94 11.17 ;
        RECT 12.13 0 12.935 0.38 ;
      LAYER li1 ;
        RECT 12.13 10.865 107.73 12.465 ;
        RECT 106.75 10.235 106.92 12.465 ;
        RECT 105.76 10.235 105.93 12.465 ;
        RECT 103.02 10.235 103.19 12.465 ;
        RECT 97.405 10.235 97.575 12.465 ;
        RECT 88.19 10.235 88.36 12.465 ;
        RECT 87.2 10.235 87.37 12.465 ;
        RECT 84.46 10.235 84.63 12.465 ;
        RECT 78.845 10.235 79.015 12.465 ;
        RECT 69.63 10.235 69.8 12.465 ;
        RECT 68.64 10.235 68.81 12.465 ;
        RECT 65.9 10.235 66.07 12.465 ;
        RECT 60.285 10.235 60.455 12.465 ;
        RECT 51.07 10.235 51.24 12.465 ;
        RECT 50.08 10.235 50.25 12.465 ;
        RECT 47.34 10.235 47.51 12.465 ;
        RECT 41.725 10.235 41.895 12.465 ;
        RECT 32.51 10.235 32.68 12.465 ;
        RECT 31.52 10.235 31.69 12.465 ;
        RECT 28.78 10.235 28.95 12.465 ;
        RECT 23.165 10.235 23.335 12.465 ;
        RECT 12.135 10.855 12.94 12.465 ;
        RECT 12.35 10.835 12.6 12.465 ;
        RECT 12.35 10.235 12.52 12.465 ;
        RECT 12.13 0 107.725 1.6 ;
        RECT 106.75 0 106.92 2.23 ;
        RECT 105.76 0 105.93 2.23 ;
        RECT 103.02 0 103.19 2.23 ;
        RECT 89.91 0 101.955 2.88 ;
        RECT 100.96 0 101.13 3.38 ;
        RECT 100 0 100.17 3.38 ;
        RECT 99.04 0 99.21 3.38 ;
        RECT 98.52 0 98.69 3.38 ;
        RECT 98.24 0 98.435 2.89 ;
        RECT 97.56 0 97.73 3.38 ;
        RECT 96.56 0 96.73 3.38 ;
        RECT 95.6 0 95.77 3.38 ;
        RECT 94.565 0 94.76 2.89 ;
        RECT 94.12 0 94.29 3.38 ;
        RECT 92.2 0 92.46 2.89 ;
        RECT 92.2 0 92.37 3.38 ;
        RECT 90.72 0 90.89 3.38 ;
        RECT 88.19 0 88.36 2.23 ;
        RECT 87.2 0 87.37 2.23 ;
        RECT 84.46 0 84.63 2.23 ;
        RECT 71.35 0 83.395 2.88 ;
        RECT 82.4 0 82.57 3.38 ;
        RECT 81.44 0 81.61 3.38 ;
        RECT 80.48 0 80.65 3.38 ;
        RECT 79.96 0 80.13 3.38 ;
        RECT 79.68 0 79.875 2.89 ;
        RECT 79 0 79.17 3.38 ;
        RECT 78 0 78.17 3.38 ;
        RECT 77.04 0 77.21 3.38 ;
        RECT 76.005 0 76.2 2.89 ;
        RECT 75.56 0 75.73 3.38 ;
        RECT 73.64 0 73.9 2.89 ;
        RECT 73.64 0 73.81 3.38 ;
        RECT 72.16 0 72.33 3.38 ;
        RECT 69.63 0 69.8 2.23 ;
        RECT 68.64 0 68.81 2.23 ;
        RECT 65.9 0 66.07 2.23 ;
        RECT 52.79 0 64.835 2.88 ;
        RECT 63.84 0 64.01 3.38 ;
        RECT 62.88 0 63.05 3.38 ;
        RECT 61.92 0 62.09 3.38 ;
        RECT 61.4 0 61.57 3.38 ;
        RECT 61.12 0 61.315 2.89 ;
        RECT 60.44 0 60.61 3.38 ;
        RECT 59.44 0 59.61 3.38 ;
        RECT 58.48 0 58.65 3.38 ;
        RECT 57.445 0 57.64 2.89 ;
        RECT 57 0 57.17 3.38 ;
        RECT 55.08 0 55.34 2.89 ;
        RECT 55.08 0 55.25 3.38 ;
        RECT 53.6 0 53.77 3.38 ;
        RECT 51.07 0 51.24 2.23 ;
        RECT 50.08 0 50.25 2.23 ;
        RECT 47.34 0 47.51 2.23 ;
        RECT 34.23 0 46.275 2.88 ;
        RECT 45.28 0 45.45 3.38 ;
        RECT 44.32 0 44.49 3.38 ;
        RECT 43.36 0 43.53 3.38 ;
        RECT 42.84 0 43.01 3.38 ;
        RECT 42.56 0 42.755 2.89 ;
        RECT 41.88 0 42.05 3.38 ;
        RECT 40.88 0 41.05 3.38 ;
        RECT 39.92 0 40.09 3.38 ;
        RECT 38.885 0 39.08 2.89 ;
        RECT 38.44 0 38.61 3.38 ;
        RECT 36.52 0 36.78 2.89 ;
        RECT 36.52 0 36.69 3.38 ;
        RECT 35.04 0 35.21 3.38 ;
        RECT 32.51 0 32.68 2.23 ;
        RECT 31.52 0 31.69 2.23 ;
        RECT 28.78 0 28.95 2.23 ;
        RECT 15.67 0 27.715 2.88 ;
        RECT 26.72 0 26.89 3.38 ;
        RECT 25.76 0 25.93 3.38 ;
        RECT 24.8 0 24.97 3.38 ;
        RECT 24.28 0 24.45 3.38 ;
        RECT 24 0 24.195 2.89 ;
        RECT 23.32 0 23.49 3.38 ;
        RECT 22.32 0 22.49 3.38 ;
        RECT 21.36 0 21.53 3.38 ;
        RECT 20.325 0 20.52 2.89 ;
        RECT 19.88 0 20.05 3.38 ;
        RECT 17.96 0 18.22 2.89 ;
        RECT 17.96 0 18.13 3.38 ;
        RECT 16.48 0 16.65 3.38 ;
        RECT 98.41 8.365 98.58 10.315 ;
        RECT 98.355 10.145 98.525 10.595 ;
        RECT 98.355 7.305 98.525 8.535 ;
        RECT 93.4 3.79 93.57 4.12 ;
        RECT 91.56 4.35 91.85 4.52 ;
        RECT 91.56 3.87 91.73 4.52 ;
        RECT 91.36 3.87 91.73 4.04 ;
        RECT 79.85 8.365 80.02 10.315 ;
        RECT 79.795 10.145 79.965 10.595 ;
        RECT 79.795 7.305 79.965 8.535 ;
        RECT 74.84 3.79 75.01 4.12 ;
        RECT 73 4.35 73.29 4.52 ;
        RECT 73 3.87 73.17 4.52 ;
        RECT 72.8 3.87 73.17 4.04 ;
        RECT 61.29 8.365 61.46 10.315 ;
        RECT 61.235 10.145 61.405 10.595 ;
        RECT 61.235 7.305 61.405 8.535 ;
        RECT 56.28 3.79 56.45 4.12 ;
        RECT 54.44 4.35 54.73 4.52 ;
        RECT 54.44 3.87 54.61 4.52 ;
        RECT 54.24 3.87 54.61 4.04 ;
        RECT 42.73 8.365 42.9 10.315 ;
        RECT 42.675 10.145 42.845 10.595 ;
        RECT 42.675 7.305 42.845 8.535 ;
        RECT 37.72 3.79 37.89 4.12 ;
        RECT 35.88 4.35 36.17 4.52 ;
        RECT 35.88 3.87 36.05 4.52 ;
        RECT 35.68 3.87 36.05 4.04 ;
        RECT 24.17 8.365 24.34 10.315 ;
        RECT 24.115 10.145 24.285 10.595 ;
        RECT 24.115 7.305 24.285 8.535 ;
        RECT 19.16 3.79 19.33 4.12 ;
        RECT 17.32 4.35 17.61 4.52 ;
        RECT 17.32 3.87 17.49 4.52 ;
        RECT 17.12 3.87 17.49 4.04 ;
      LAYER met2 ;
        RECT 93.355 3.715 93.615 4.035 ;
        RECT 91.575 3.805 93.615 3.945 ;
        RECT 91.955 2.295 92.295 2.635 ;
        RECT 91.885 3.69 92.165 4.06 ;
        RECT 91.98 2.295 92.15 4.06 ;
        RECT 91.635 4.275 91.895 4.595 ;
        RECT 91.575 3.805 91.715 4.505 ;
        RECT 74.795 3.715 75.055 4.035 ;
        RECT 73.015 3.805 75.055 3.945 ;
        RECT 73.395 2.295 73.735 2.635 ;
        RECT 73.325 3.69 73.605 4.06 ;
        RECT 73.42 2.295 73.59 4.06 ;
        RECT 73.075 4.275 73.335 4.595 ;
        RECT 73.015 3.805 73.155 4.505 ;
        RECT 56.235 3.715 56.495 4.035 ;
        RECT 54.455 3.805 56.495 3.945 ;
        RECT 54.835 2.295 55.175 2.635 ;
        RECT 54.765 3.69 55.045 4.06 ;
        RECT 54.86 2.295 55.03 4.06 ;
        RECT 54.515 4.275 54.775 4.595 ;
        RECT 54.455 3.805 54.595 4.505 ;
        RECT 37.675 3.715 37.935 4.035 ;
        RECT 35.895 3.805 37.935 3.945 ;
        RECT 36.275 2.295 36.615 2.635 ;
        RECT 36.205 3.69 36.485 4.06 ;
        RECT 36.3 2.295 36.47 4.06 ;
        RECT 35.955 4.275 36.215 4.595 ;
        RECT 35.895 3.805 36.035 4.505 ;
        RECT 19.115 3.715 19.375 4.035 ;
        RECT 17.335 3.805 19.375 3.945 ;
        RECT 17.715 2.295 18.055 2.635 ;
        RECT 17.645 3.69 17.925 4.06 ;
        RECT 17.74 2.295 17.91 4.06 ;
        RECT 17.395 4.275 17.655 4.595 ;
        RECT 17.335 3.805 17.475 4.505 ;
        RECT 12.325 10.79 12.705 11.17 ;
        RECT 12.32 0 12.7 0.38 ;
        RECT 12.365 0 12.535 11.17 ;
      LAYER met1 ;
        RECT 12.13 0 107.73 1.6 ;
        RECT 89.91 0 101.955 2.88 ;
        RECT 89.91 0 101.87 3.035 ;
        RECT 71.35 0 83.395 2.88 ;
        RECT 71.35 0 83.31 3.035 ;
        RECT 52.79 0 64.835 2.88 ;
        RECT 52.79 0 64.75 3.035 ;
        RECT 34.23 0 46.275 2.88 ;
        RECT 34.23 0 46.19 3.035 ;
        RECT 15.67 0 27.715 2.88 ;
        RECT 15.67 0 27.63 3.035 ;
        RECT 12.13 10.865 107.73 12.465 ;
        RECT 98.35 8.575 98.64 8.805 ;
        RECT 97.915 8.605 98.64 8.775 ;
        RECT 97.915 8.605 98.085 12.465 ;
        RECT 79.79 8.575 80.08 8.805 ;
        RECT 79.355 8.605 80.08 8.775 ;
        RECT 79.355 8.605 79.525 12.465 ;
        RECT 61.23 8.575 61.52 8.805 ;
        RECT 60.795 8.605 61.52 8.775 ;
        RECT 60.795 8.605 60.965 12.465 ;
        RECT 42.67 8.575 42.96 8.805 ;
        RECT 42.235 8.605 42.96 8.775 ;
        RECT 42.235 8.605 42.405 12.465 ;
        RECT 24.11 8.575 24.4 8.805 ;
        RECT 23.675 8.605 24.4 8.775 ;
        RECT 23.675 8.605 23.845 12.465 ;
        RECT 12.135 10.855 12.94 12.465 ;
        RECT 12.34 10.835 12.69 12.465 ;
        RECT 93.34 3.665 93.63 4.035 ;
        RECT 92.575 3.665 93.63 3.805 ;
        RECT 91.605 4.305 91.925 4.565 ;
        RECT 74.78 3.665 75.07 4.035 ;
        RECT 74.015 3.665 75.07 3.805 ;
        RECT 73.045 4.305 73.365 4.565 ;
        RECT 56.22 3.665 56.51 4.035 ;
        RECT 55.455 3.665 56.51 3.805 ;
        RECT 54.485 4.305 54.805 4.565 ;
        RECT 37.66 3.665 37.95 4.035 ;
        RECT 36.895 3.665 37.95 3.805 ;
        RECT 35.925 4.305 36.245 4.565 ;
        RECT 19.1 3.665 19.39 4.035 ;
        RECT 18.335 3.665 19.39 3.805 ;
        RECT 17.365 4.305 17.685 4.565 ;
      LAYER via2 ;
        RECT 12.41 0.09 12.61 0.29 ;
        RECT 12.415 10.88 12.615 11.08 ;
        RECT 17.685 3.775 17.885 3.975 ;
        RECT 36.245 3.775 36.445 3.975 ;
        RECT 54.805 3.775 55.005 3.975 ;
        RECT 73.365 3.775 73.565 3.975 ;
        RECT 91.925 3.775 92.125 3.975 ;
      LAYER via1 ;
        RECT 12.435 0.115 12.585 0.265 ;
        RECT 12.44 10.905 12.59 11.055 ;
        RECT 17.45 4.36 17.6 4.51 ;
        RECT 17.81 2.39 17.96 2.54 ;
        RECT 19.17 3.8 19.32 3.95 ;
        RECT 36.01 4.36 36.16 4.51 ;
        RECT 36.37 2.39 36.52 2.54 ;
        RECT 37.73 3.8 37.88 3.95 ;
        RECT 54.57 4.36 54.72 4.51 ;
        RECT 54.93 2.39 55.08 2.54 ;
        RECT 56.29 3.8 56.44 3.95 ;
        RECT 73.13 4.36 73.28 4.51 ;
        RECT 73.49 2.39 73.64 2.54 ;
        RECT 74.85 3.8 75 3.95 ;
        RECT 91.69 4.36 91.84 4.51 ;
        RECT 92.05 2.39 92.2 2.54 ;
        RECT 93.41 3.8 93.56 3.95 ;
      LAYER mcon ;
        RECT 12.43 10.895 12.6 11.065 ;
        RECT 13.11 10.895 13.28 11.065 ;
        RECT 13.79 10.895 13.96 11.065 ;
        RECT 14.47 10.895 14.64 11.065 ;
        RECT 15.815 2.71 15.985 2.88 ;
        RECT 16.275 2.71 16.445 2.88 ;
        RECT 16.735 2.71 16.905 2.88 ;
        RECT 17.195 2.71 17.365 2.88 ;
        RECT 17.44 4.35 17.61 4.52 ;
        RECT 17.655 2.71 17.825 2.88 ;
        RECT 18.115 2.71 18.285 2.88 ;
        RECT 18.575 2.71 18.745 2.88 ;
        RECT 19.035 2.71 19.205 2.88 ;
        RECT 19.16 3.79 19.33 3.96 ;
        RECT 19.495 2.71 19.665 2.88 ;
        RECT 19.955 2.71 20.125 2.88 ;
        RECT 20.415 2.71 20.585 2.88 ;
        RECT 20.875 2.71 21.045 2.88 ;
        RECT 21.335 2.71 21.505 2.88 ;
        RECT 21.795 2.71 21.965 2.88 ;
        RECT 22.255 2.71 22.425 2.88 ;
        RECT 22.715 2.71 22.885 2.88 ;
        RECT 23.175 2.71 23.345 2.88 ;
        RECT 23.245 10.895 23.415 11.065 ;
        RECT 23.635 2.71 23.805 2.88 ;
        RECT 23.925 10.895 24.095 11.065 ;
        RECT 24.095 2.71 24.265 2.88 ;
        RECT 24.17 8.605 24.34 8.775 ;
        RECT 24.555 2.71 24.725 2.88 ;
        RECT 24.605 10.895 24.775 11.065 ;
        RECT 25.015 2.71 25.185 2.88 ;
        RECT 25.285 10.895 25.455 11.065 ;
        RECT 25.475 2.71 25.645 2.88 ;
        RECT 25.935 2.71 26.105 2.88 ;
        RECT 26.395 2.71 26.565 2.88 ;
        RECT 26.855 2.71 27.025 2.88 ;
        RECT 27.315 2.71 27.485 2.88 ;
        RECT 28.86 10.895 29.03 11.065 ;
        RECT 28.86 1.4 29.03 1.57 ;
        RECT 29.54 10.895 29.71 11.065 ;
        RECT 29.54 1.4 29.71 1.57 ;
        RECT 30.22 10.895 30.39 11.065 ;
        RECT 30.22 1.4 30.39 1.57 ;
        RECT 30.9 10.895 31.07 11.065 ;
        RECT 30.9 1.4 31.07 1.57 ;
        RECT 31.6 10.895 31.77 11.065 ;
        RECT 31.6 1.4 31.77 1.57 ;
        RECT 32.59 10.895 32.76 11.065 ;
        RECT 32.59 1.4 32.76 1.57 ;
        RECT 34.375 2.71 34.545 2.88 ;
        RECT 34.835 2.71 35.005 2.88 ;
        RECT 35.295 2.71 35.465 2.88 ;
        RECT 35.755 2.71 35.925 2.88 ;
        RECT 36 4.35 36.17 4.52 ;
        RECT 36.215 2.71 36.385 2.88 ;
        RECT 36.675 2.71 36.845 2.88 ;
        RECT 37.135 2.71 37.305 2.88 ;
        RECT 37.595 2.71 37.765 2.88 ;
        RECT 37.72 3.79 37.89 3.96 ;
        RECT 38.055 2.71 38.225 2.88 ;
        RECT 38.515 2.71 38.685 2.88 ;
        RECT 38.975 2.71 39.145 2.88 ;
        RECT 39.435 2.71 39.605 2.88 ;
        RECT 39.895 2.71 40.065 2.88 ;
        RECT 40.355 2.71 40.525 2.88 ;
        RECT 40.815 2.71 40.985 2.88 ;
        RECT 41.275 2.71 41.445 2.88 ;
        RECT 41.735 2.71 41.905 2.88 ;
        RECT 41.805 10.895 41.975 11.065 ;
        RECT 42.195 2.71 42.365 2.88 ;
        RECT 42.485 10.895 42.655 11.065 ;
        RECT 42.655 2.71 42.825 2.88 ;
        RECT 42.73 8.605 42.9 8.775 ;
        RECT 43.115 2.71 43.285 2.88 ;
        RECT 43.165 10.895 43.335 11.065 ;
        RECT 43.575 2.71 43.745 2.88 ;
        RECT 43.845 10.895 44.015 11.065 ;
        RECT 44.035 2.71 44.205 2.88 ;
        RECT 44.495 2.71 44.665 2.88 ;
        RECT 44.955 2.71 45.125 2.88 ;
        RECT 45.415 2.71 45.585 2.88 ;
        RECT 45.875 2.71 46.045 2.88 ;
        RECT 47.42 10.895 47.59 11.065 ;
        RECT 47.42 1.4 47.59 1.57 ;
        RECT 48.1 10.895 48.27 11.065 ;
        RECT 48.1 1.4 48.27 1.57 ;
        RECT 48.78 10.895 48.95 11.065 ;
        RECT 48.78 1.4 48.95 1.57 ;
        RECT 49.46 10.895 49.63 11.065 ;
        RECT 49.46 1.4 49.63 1.57 ;
        RECT 50.16 10.895 50.33 11.065 ;
        RECT 50.16 1.4 50.33 1.57 ;
        RECT 51.15 10.895 51.32 11.065 ;
        RECT 51.15 1.4 51.32 1.57 ;
        RECT 52.935 2.71 53.105 2.88 ;
        RECT 53.395 2.71 53.565 2.88 ;
        RECT 53.855 2.71 54.025 2.88 ;
        RECT 54.315 2.71 54.485 2.88 ;
        RECT 54.56 4.35 54.73 4.52 ;
        RECT 54.775 2.71 54.945 2.88 ;
        RECT 55.235 2.71 55.405 2.88 ;
        RECT 55.695 2.71 55.865 2.88 ;
        RECT 56.155 2.71 56.325 2.88 ;
        RECT 56.28 3.79 56.45 3.96 ;
        RECT 56.615 2.71 56.785 2.88 ;
        RECT 57.075 2.71 57.245 2.88 ;
        RECT 57.535 2.71 57.705 2.88 ;
        RECT 57.995 2.71 58.165 2.88 ;
        RECT 58.455 2.71 58.625 2.88 ;
        RECT 58.915 2.71 59.085 2.88 ;
        RECT 59.375 2.71 59.545 2.88 ;
        RECT 59.835 2.71 60.005 2.88 ;
        RECT 60.295 2.71 60.465 2.88 ;
        RECT 60.365 10.895 60.535 11.065 ;
        RECT 60.755 2.71 60.925 2.88 ;
        RECT 61.045 10.895 61.215 11.065 ;
        RECT 61.215 2.71 61.385 2.88 ;
        RECT 61.29 8.605 61.46 8.775 ;
        RECT 61.675 2.71 61.845 2.88 ;
        RECT 61.725 10.895 61.895 11.065 ;
        RECT 62.135 2.71 62.305 2.88 ;
        RECT 62.405 10.895 62.575 11.065 ;
        RECT 62.595 2.71 62.765 2.88 ;
        RECT 63.055 2.71 63.225 2.88 ;
        RECT 63.515 2.71 63.685 2.88 ;
        RECT 63.975 2.71 64.145 2.88 ;
        RECT 64.435 2.71 64.605 2.88 ;
        RECT 65.98 10.895 66.15 11.065 ;
        RECT 65.98 1.4 66.15 1.57 ;
        RECT 66.66 10.895 66.83 11.065 ;
        RECT 66.66 1.4 66.83 1.57 ;
        RECT 67.34 10.895 67.51 11.065 ;
        RECT 67.34 1.4 67.51 1.57 ;
        RECT 68.02 10.895 68.19 11.065 ;
        RECT 68.02 1.4 68.19 1.57 ;
        RECT 68.72 10.895 68.89 11.065 ;
        RECT 68.72 1.4 68.89 1.57 ;
        RECT 69.71 10.895 69.88 11.065 ;
        RECT 69.71 1.4 69.88 1.57 ;
        RECT 71.495 2.71 71.665 2.88 ;
        RECT 71.955 2.71 72.125 2.88 ;
        RECT 72.415 2.71 72.585 2.88 ;
        RECT 72.875 2.71 73.045 2.88 ;
        RECT 73.12 4.35 73.29 4.52 ;
        RECT 73.335 2.71 73.505 2.88 ;
        RECT 73.795 2.71 73.965 2.88 ;
        RECT 74.255 2.71 74.425 2.88 ;
        RECT 74.715 2.71 74.885 2.88 ;
        RECT 74.84 3.79 75.01 3.96 ;
        RECT 75.175 2.71 75.345 2.88 ;
        RECT 75.635 2.71 75.805 2.88 ;
        RECT 76.095 2.71 76.265 2.88 ;
        RECT 76.555 2.71 76.725 2.88 ;
        RECT 77.015 2.71 77.185 2.88 ;
        RECT 77.475 2.71 77.645 2.88 ;
        RECT 77.935 2.71 78.105 2.88 ;
        RECT 78.395 2.71 78.565 2.88 ;
        RECT 78.855 2.71 79.025 2.88 ;
        RECT 78.925 10.895 79.095 11.065 ;
        RECT 79.315 2.71 79.485 2.88 ;
        RECT 79.605 10.895 79.775 11.065 ;
        RECT 79.775 2.71 79.945 2.88 ;
        RECT 79.85 8.605 80.02 8.775 ;
        RECT 80.235 2.71 80.405 2.88 ;
        RECT 80.285 10.895 80.455 11.065 ;
        RECT 80.695 2.71 80.865 2.88 ;
        RECT 80.965 10.895 81.135 11.065 ;
        RECT 81.155 2.71 81.325 2.88 ;
        RECT 81.615 2.71 81.785 2.88 ;
        RECT 82.075 2.71 82.245 2.88 ;
        RECT 82.535 2.71 82.705 2.88 ;
        RECT 82.995 2.71 83.165 2.88 ;
        RECT 84.54 10.895 84.71 11.065 ;
        RECT 84.54 1.4 84.71 1.57 ;
        RECT 85.22 10.895 85.39 11.065 ;
        RECT 85.22 1.4 85.39 1.57 ;
        RECT 85.9 10.895 86.07 11.065 ;
        RECT 85.9 1.4 86.07 1.57 ;
        RECT 86.58 10.895 86.75 11.065 ;
        RECT 86.58 1.4 86.75 1.57 ;
        RECT 87.28 10.895 87.45 11.065 ;
        RECT 87.28 1.4 87.45 1.57 ;
        RECT 88.27 10.895 88.44 11.065 ;
        RECT 88.27 1.4 88.44 1.57 ;
        RECT 90.055 2.71 90.225 2.88 ;
        RECT 90.515 2.71 90.685 2.88 ;
        RECT 90.975 2.71 91.145 2.88 ;
        RECT 91.435 2.71 91.605 2.88 ;
        RECT 91.68 4.35 91.85 4.52 ;
        RECT 91.895 2.71 92.065 2.88 ;
        RECT 92.355 2.71 92.525 2.88 ;
        RECT 92.815 2.71 92.985 2.88 ;
        RECT 93.275 2.71 93.445 2.88 ;
        RECT 93.4 3.79 93.57 3.96 ;
        RECT 93.735 2.71 93.905 2.88 ;
        RECT 94.195 2.71 94.365 2.88 ;
        RECT 94.655 2.71 94.825 2.88 ;
        RECT 95.115 2.71 95.285 2.88 ;
        RECT 95.575 2.71 95.745 2.88 ;
        RECT 96.035 2.71 96.205 2.88 ;
        RECT 96.495 2.71 96.665 2.88 ;
        RECT 96.955 2.71 97.125 2.88 ;
        RECT 97.415 2.71 97.585 2.88 ;
        RECT 97.485 10.895 97.655 11.065 ;
        RECT 97.875 2.71 98.045 2.88 ;
        RECT 98.165 10.895 98.335 11.065 ;
        RECT 98.335 2.71 98.505 2.88 ;
        RECT 98.41 8.605 98.58 8.775 ;
        RECT 98.795 2.71 98.965 2.88 ;
        RECT 98.845 10.895 99.015 11.065 ;
        RECT 99.255 2.71 99.425 2.88 ;
        RECT 99.525 10.895 99.695 11.065 ;
        RECT 99.715 2.71 99.885 2.88 ;
        RECT 100.175 2.71 100.345 2.88 ;
        RECT 100.635 2.71 100.805 2.88 ;
        RECT 101.095 2.71 101.265 2.88 ;
        RECT 101.555 2.71 101.725 2.88 ;
        RECT 103.1 10.895 103.27 11.065 ;
        RECT 103.1 1.4 103.27 1.57 ;
        RECT 103.78 10.895 103.95 11.065 ;
        RECT 103.78 1.4 103.95 1.57 ;
        RECT 104.46 10.895 104.63 11.065 ;
        RECT 104.46 1.4 104.63 1.57 ;
        RECT 105.14 10.895 105.31 11.065 ;
        RECT 105.14 1.4 105.31 1.57 ;
        RECT 105.84 10.895 106.01 11.065 ;
        RECT 105.84 1.4 106.01 1.57 ;
        RECT 106.83 10.895 107 11.065 ;
        RECT 106.83 1.4 107 1.57 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 98.685 9.345 99.06 9.715 ;
      RECT 80.125 9.345 80.5 9.715 ;
      RECT 61.565 9.345 61.94 9.715 ;
      RECT 43.005 9.345 43.38 9.715 ;
      RECT 24.445 9.345 24.82 9.715 ;
      RECT 98.685 9.385 99.69 9.685 ;
      RECT 99.39 5.45 99.69 9.685 ;
      RECT 80.125 9.385 81.13 9.685 ;
      RECT 80.83 5.45 81.13 9.685 ;
      RECT 61.565 9.385 62.57 9.685 ;
      RECT 62.27 5.45 62.57 9.685 ;
      RECT 43.005 9.385 44.01 9.685 ;
      RECT 43.71 5.45 44.01 9.685 ;
      RECT 24.445 9.385 25.45 9.685 ;
      RECT 25.15 5.45 25.45 9.685 ;
      RECT 12.125 5.45 107.725 7.05 ;
      RECT 94.065 3.71 94.365 7.05 ;
      RECT 92.63 4.27 92.93 7.05 ;
      RECT 89.165 5.435 90.005 7.05 ;
      RECT 75.505 3.71 75.805 7.05 ;
      RECT 74.07 4.27 74.37 7.05 ;
      RECT 70.605 5.435 71.445 7.05 ;
      RECT 56.945 3.71 57.245 7.05 ;
      RECT 55.51 4.27 55.81 7.05 ;
      RECT 52.045 5.435 52.885 7.05 ;
      RECT 38.385 3.71 38.685 7.05 ;
      RECT 36.95 4.27 37.25 7.05 ;
      RECT 33.485 5.435 34.325 7.05 ;
      RECT 19.825 3.71 20.125 7.05 ;
      RECT 18.39 4.27 18.69 7.05 ;
      RECT 14.925 5.435 15.765 7.05 ;
      RECT 89.56 3.715 89.86 7.05 ;
      RECT 71 3.715 71.3 7.05 ;
      RECT 52.44 3.715 52.74 7.05 ;
      RECT 33.88 3.715 34.18 7.05 ;
      RECT 15.32 3.715 15.62 7.05 ;
      RECT 92.6 4.27 93.33 4.6 ;
      RECT 74.04 4.27 74.77 4.6 ;
      RECT 55.48 4.27 56.21 4.6 ;
      RECT 36.92 4.27 37.65 4.6 ;
      RECT 18.36 4.27 19.09 4.6 ;
      RECT 94.04 3.71 94.77 4.04 ;
      RECT 90.49 3.71 91.22 4.04 ;
      RECT 75.48 3.71 76.21 4.04 ;
      RECT 71.93 3.71 72.66 4.04 ;
      RECT 56.92 3.71 57.65 4.04 ;
      RECT 53.37 3.71 54.1 4.04 ;
      RECT 38.36 3.71 39.09 4.04 ;
      RECT 34.81 3.71 35.54 4.04 ;
      RECT 19.8 3.71 20.53 4.04 ;
      RECT 16.25 3.71 16.98 4.04 ;
      RECT 89.56 3.715 91.22 4.015 ;
      RECT 71 3.715 72.66 4.015 ;
      RECT 52.44 3.715 54.1 4.015 ;
      RECT 33.88 3.715 35.54 4.015 ;
      RECT 15.32 3.715 16.98 4.015 ;
      RECT 99.215 4.83 99.77 5.16 ;
      RECT 99.215 3.165 99.515 5.16 ;
      RECT 95.28 4.27 95.835 4.6 ;
      RECT 95.535 3.165 95.835 4.6 ;
      RECT 95.535 3.165 99.515 3.465 ;
      RECT 80.655 4.83 81.21 5.16 ;
      RECT 80.655 3.165 80.955 5.16 ;
      RECT 76.72 4.27 77.275 4.6 ;
      RECT 76.975 3.165 77.275 4.6 ;
      RECT 76.975 3.165 80.955 3.465 ;
      RECT 62.095 4.83 62.65 5.16 ;
      RECT 62.095 3.165 62.395 5.16 ;
      RECT 58.16 4.27 58.715 4.6 ;
      RECT 58.415 3.165 58.715 4.6 ;
      RECT 58.415 3.165 62.395 3.465 ;
      RECT 43.535 4.83 44.09 5.16 ;
      RECT 43.535 3.165 43.835 5.16 ;
      RECT 39.6 4.27 40.155 4.6 ;
      RECT 39.855 3.165 40.155 4.6 ;
      RECT 39.855 3.165 43.835 3.465 ;
      RECT 24.975 4.83 25.53 5.16 ;
      RECT 24.975 3.165 25.275 5.16 ;
      RECT 21.04 4.27 21.595 4.6 ;
      RECT 21.295 3.165 21.595 4.6 ;
      RECT 21.295 3.165 25.275 3.465 ;
      RECT 100.4 3.15 101.13 3.48 ;
      RECT 98.18 4.83 98.91 5.16 ;
      RECT 96.48 4.83 97.21 5.16 ;
      RECT 90.16 4.83 90.89 5.16 ;
      RECT 81.84 3.15 82.57 3.48 ;
      RECT 79.62 4.83 80.35 5.16 ;
      RECT 77.92 4.83 78.65 5.16 ;
      RECT 71.6 4.83 72.33 5.16 ;
      RECT 63.28 3.15 64.01 3.48 ;
      RECT 61.06 4.83 61.79 5.16 ;
      RECT 59.36 4.83 60.09 5.16 ;
      RECT 53.04 4.83 53.77 5.16 ;
      RECT 44.72 3.15 45.45 3.48 ;
      RECT 42.5 4.83 43.23 5.16 ;
      RECT 40.8 4.83 41.53 5.16 ;
      RECT 34.48 4.83 35.21 5.16 ;
      RECT 26.16 3.15 26.89 3.48 ;
      RECT 23.94 4.83 24.67 5.16 ;
      RECT 22.24 4.83 22.97 5.16 ;
      RECT 15.92 4.83 16.65 5.16 ;
    LAYER via2 ;
      RECT 100.465 3.215 100.665 3.415 ;
      RECT 99.505 4.895 99.705 5.095 ;
      RECT 98.77 9.43 98.97 9.63 ;
      RECT 98.505 4.895 98.705 5.095 ;
      RECT 96.545 4.895 96.745 5.095 ;
      RECT 95.345 4.335 95.545 4.535 ;
      RECT 94.105 3.775 94.305 3.975 ;
      RECT 92.665 4.335 92.865 4.535 ;
      RECT 90.705 3.775 90.905 3.975 ;
      RECT 90.225 4.895 90.425 5.095 ;
      RECT 81.905 3.215 82.105 3.415 ;
      RECT 80.945 4.895 81.145 5.095 ;
      RECT 80.21 9.43 80.41 9.63 ;
      RECT 79.945 4.895 80.145 5.095 ;
      RECT 77.985 4.895 78.185 5.095 ;
      RECT 76.785 4.335 76.985 4.535 ;
      RECT 75.545 3.775 75.745 3.975 ;
      RECT 74.105 4.335 74.305 4.535 ;
      RECT 72.145 3.775 72.345 3.975 ;
      RECT 71.665 4.895 71.865 5.095 ;
      RECT 63.345 3.215 63.545 3.415 ;
      RECT 62.385 4.895 62.585 5.095 ;
      RECT 61.65 9.43 61.85 9.63 ;
      RECT 61.385 4.895 61.585 5.095 ;
      RECT 59.425 4.895 59.625 5.095 ;
      RECT 58.225 4.335 58.425 4.535 ;
      RECT 56.985 3.775 57.185 3.975 ;
      RECT 55.545 4.335 55.745 4.535 ;
      RECT 53.585 3.775 53.785 3.975 ;
      RECT 53.105 4.895 53.305 5.095 ;
      RECT 44.785 3.215 44.985 3.415 ;
      RECT 43.825 4.895 44.025 5.095 ;
      RECT 43.09 9.43 43.29 9.63 ;
      RECT 42.825 4.895 43.025 5.095 ;
      RECT 40.865 4.895 41.065 5.095 ;
      RECT 39.665 4.335 39.865 4.535 ;
      RECT 38.425 3.775 38.625 3.975 ;
      RECT 36.985 4.335 37.185 4.535 ;
      RECT 35.025 3.775 35.225 3.975 ;
      RECT 34.545 4.895 34.745 5.095 ;
      RECT 26.225 3.215 26.425 3.415 ;
      RECT 25.265 4.895 25.465 5.095 ;
      RECT 24.53 9.43 24.73 9.63 ;
      RECT 24.265 4.895 24.465 5.095 ;
      RECT 22.305 4.895 22.505 5.095 ;
      RECT 21.105 4.335 21.305 4.535 ;
      RECT 19.865 3.775 20.065 3.975 ;
      RECT 18.425 4.335 18.625 4.535 ;
      RECT 16.465 3.775 16.665 3.975 ;
      RECT 15.985 4.895 16.185 5.095 ;
      RECT 13.9 6.645 14.1 6.845 ;
    LAYER met2 ;
      RECT 13.36 10.69 107.355 10.86 ;
      RECT 107.185 9.565 107.355 10.86 ;
      RECT 13.36 8.545 13.53 10.86 ;
      RECT 107.155 9.565 107.505 9.915 ;
      RECT 13.295 8.545 13.585 8.895 ;
      RECT 103.995 8.51 104.315 8.835 ;
      RECT 104.025 7.985 104.195 8.835 ;
      RECT 104.025 7.985 104.2 8.335 ;
      RECT 104.025 7.985 105 8.16 ;
      RECT 104.825 3.26 105 8.16 ;
      RECT 104.77 3.26 105.12 3.61 ;
      RECT 104.795 8.945 105.12 9.27 ;
      RECT 103.68 9.035 105.12 9.205 ;
      RECT 103.68 3.69 103.84 9.205 ;
      RECT 103.995 3.66 104.315 3.98 ;
      RECT 103.68 3.69 104.315 3.86 ;
      RECT 98.515 5.43 102.65 5.62 ;
      RECT 102.48 4.44 102.65 5.62 ;
      RECT 102.46 4.445 102.65 5.62 ;
      RECT 98.515 4.81 98.705 5.62 ;
      RECT 98.465 4.81 98.745 5.18 ;
      RECT 102.39 4.445 102.73 4.795 ;
      RECT 88.57 8.945 88.92 9.295 ;
      RECT 99.355 8.9 99.705 9.25 ;
      RECT 88.57 8.975 99.705 9.175 ;
      RECT 98.995 4.275 99.255 4.595 ;
      RECT 99.055 3.155 99.195 4.595 ;
      RECT 98.995 3.155 99.255 3.475 ;
      RECT 97.995 4.835 98.255 5.155 ;
      RECT 97.995 4.25 98.195 5.155 ;
      RECT 97.935 3.155 98.075 4.785 ;
      RECT 97.935 4.25 98.435 4.62 ;
      RECT 97.875 3.155 98.135 3.475 ;
      RECT 97.515 4.835 97.775 5.155 ;
      RECT 97.575 3.245 97.715 5.155 ;
      RECT 97.275 3.245 97.715 3.475 ;
      RECT 97.275 3.155 97.535 3.475 ;
      RECT 97.035 3.715 97.295 4.035 ;
      RECT 96.455 3.805 97.295 3.945 ;
      RECT 96.455 2.865 96.595 3.945 ;
      RECT 93.115 3.155 93.375 3.475 ;
      RECT 93.115 3.245 94.155 3.385 ;
      RECT 94.015 2.865 94.155 3.385 ;
      RECT 94.015 2.865 96.595 3.005 ;
      RECT 96.505 4.81 96.785 5.18 ;
      RECT 96.575 4.365 96.715 5.18 ;
      RECT 96.385 4.25 96.665 4.62 ;
      RECT 96.095 4.365 96.715 4.505 ;
      RECT 96.095 3.155 96.235 4.505 ;
      RECT 96.035 3.155 96.295 3.475 ;
      RECT 95.305 4.25 95.585 4.62 ;
      RECT 95.375 3.155 95.515 4.62 ;
      RECT 95.315 3.155 95.575 3.475 ;
      RECT 94.955 4.835 95.215 5.155 ;
      RECT 95.015 3.245 95.155 5.155 ;
      RECT 94.595 3.155 94.855 3.475 ;
      RECT 94.595 3.245 95.155 3.385 ;
      RECT 92.625 4.25 92.905 4.62 ;
      RECT 94.595 4.275 94.855 4.595 ;
      RECT 92.275 4.275 92.905 4.595 ;
      RECT 92.275 4.365 94.855 4.505 ;
      RECT 94.065 3.69 94.345 4.06 ;
      RECT 94.065 3.715 94.595 4.035 ;
      RECT 91.155 4.275 91.415 4.595 ;
      RECT 91.215 3.155 91.355 4.595 ;
      RECT 91.155 3.155 91.415 3.475 ;
      RECT 90.185 4.81 90.465 5.18 ;
      RECT 90.195 4.555 90.455 5.18 ;
      RECT 85.435 8.51 85.755 8.835 ;
      RECT 85.465 7.985 85.635 8.835 ;
      RECT 85.465 7.985 85.64 8.335 ;
      RECT 85.465 7.985 86.44 8.16 ;
      RECT 86.265 3.26 86.44 8.16 ;
      RECT 86.21 3.26 86.56 3.61 ;
      RECT 86.235 8.945 86.56 9.27 ;
      RECT 85.12 9.035 86.56 9.205 ;
      RECT 85.12 3.69 85.28 9.205 ;
      RECT 85.435 3.66 85.755 3.98 ;
      RECT 85.12 3.69 85.755 3.86 ;
      RECT 79.955 5.43 84.09 5.62 ;
      RECT 83.92 4.44 84.09 5.62 ;
      RECT 83.9 4.445 84.09 5.62 ;
      RECT 79.955 4.81 80.145 5.62 ;
      RECT 79.905 4.81 80.185 5.18 ;
      RECT 83.83 4.445 84.17 4.795 ;
      RECT 70.01 8.945 70.36 9.295 ;
      RECT 80.795 8.9 81.145 9.25 ;
      RECT 70.01 8.975 81.145 9.175 ;
      RECT 80.435 4.275 80.695 4.595 ;
      RECT 80.495 3.155 80.635 4.595 ;
      RECT 80.435 3.155 80.695 3.475 ;
      RECT 79.435 4.835 79.695 5.155 ;
      RECT 79.435 4.25 79.635 5.155 ;
      RECT 79.375 3.155 79.515 4.785 ;
      RECT 79.375 4.25 79.875 4.62 ;
      RECT 79.315 3.155 79.575 3.475 ;
      RECT 78.955 4.835 79.215 5.155 ;
      RECT 79.015 3.245 79.155 5.155 ;
      RECT 78.715 3.245 79.155 3.475 ;
      RECT 78.715 3.155 78.975 3.475 ;
      RECT 78.475 3.715 78.735 4.035 ;
      RECT 77.895 3.805 78.735 3.945 ;
      RECT 77.895 2.865 78.035 3.945 ;
      RECT 74.555 3.155 74.815 3.475 ;
      RECT 74.555 3.245 75.595 3.385 ;
      RECT 75.455 2.865 75.595 3.385 ;
      RECT 75.455 2.865 78.035 3.005 ;
      RECT 77.945 4.81 78.225 5.18 ;
      RECT 78.015 4.365 78.155 5.18 ;
      RECT 77.825 4.25 78.105 4.62 ;
      RECT 77.535 4.365 78.155 4.505 ;
      RECT 77.535 3.155 77.675 4.505 ;
      RECT 77.475 3.155 77.735 3.475 ;
      RECT 76.745 4.25 77.025 4.62 ;
      RECT 76.815 3.155 76.955 4.62 ;
      RECT 76.755 3.155 77.015 3.475 ;
      RECT 76.395 4.835 76.655 5.155 ;
      RECT 76.455 3.245 76.595 5.155 ;
      RECT 76.035 3.155 76.295 3.475 ;
      RECT 76.035 3.245 76.595 3.385 ;
      RECT 74.065 4.25 74.345 4.62 ;
      RECT 76.035 4.275 76.295 4.595 ;
      RECT 73.715 4.275 74.345 4.595 ;
      RECT 73.715 4.365 76.295 4.505 ;
      RECT 75.505 3.69 75.785 4.06 ;
      RECT 75.505 3.715 76.035 4.035 ;
      RECT 72.595 4.275 72.855 4.595 ;
      RECT 72.655 3.155 72.795 4.595 ;
      RECT 72.595 3.155 72.855 3.475 ;
      RECT 71.625 4.81 71.905 5.18 ;
      RECT 71.635 4.555 71.895 5.18 ;
      RECT 66.875 8.51 67.195 8.835 ;
      RECT 66.905 7.985 67.075 8.835 ;
      RECT 66.905 7.985 67.08 8.335 ;
      RECT 66.905 7.985 67.88 8.16 ;
      RECT 67.705 3.26 67.88 8.16 ;
      RECT 67.65 3.26 68 3.61 ;
      RECT 67.675 8.945 68 9.27 ;
      RECT 66.56 9.035 68 9.205 ;
      RECT 66.56 3.69 66.72 9.205 ;
      RECT 66.875 3.66 67.195 3.98 ;
      RECT 66.56 3.69 67.195 3.86 ;
      RECT 61.395 5.43 65.53 5.62 ;
      RECT 65.36 4.44 65.53 5.62 ;
      RECT 65.34 4.445 65.53 5.62 ;
      RECT 61.395 4.81 61.585 5.62 ;
      RECT 61.345 4.81 61.625 5.18 ;
      RECT 65.27 4.445 65.61 4.795 ;
      RECT 51.495 8.95 51.845 9.3 ;
      RECT 62.235 8.905 62.585 9.255 ;
      RECT 51.495 8.98 62.585 9.18 ;
      RECT 61.875 4.275 62.135 4.595 ;
      RECT 61.935 3.155 62.075 4.595 ;
      RECT 61.875 3.155 62.135 3.475 ;
      RECT 60.875 4.835 61.135 5.155 ;
      RECT 60.875 4.25 61.075 5.155 ;
      RECT 60.815 3.155 60.955 4.785 ;
      RECT 60.815 4.25 61.315 4.62 ;
      RECT 60.755 3.155 61.015 3.475 ;
      RECT 60.395 4.835 60.655 5.155 ;
      RECT 60.455 3.245 60.595 5.155 ;
      RECT 60.155 3.245 60.595 3.475 ;
      RECT 60.155 3.155 60.415 3.475 ;
      RECT 59.915 3.715 60.175 4.035 ;
      RECT 59.335 3.805 60.175 3.945 ;
      RECT 59.335 2.865 59.475 3.945 ;
      RECT 55.995 3.155 56.255 3.475 ;
      RECT 55.995 3.245 57.035 3.385 ;
      RECT 56.895 2.865 57.035 3.385 ;
      RECT 56.895 2.865 59.475 3.005 ;
      RECT 59.385 4.81 59.665 5.18 ;
      RECT 59.455 4.365 59.595 5.18 ;
      RECT 59.265 4.25 59.545 4.62 ;
      RECT 58.975 4.365 59.595 4.505 ;
      RECT 58.975 3.155 59.115 4.505 ;
      RECT 58.915 3.155 59.175 3.475 ;
      RECT 58.185 4.25 58.465 4.62 ;
      RECT 58.255 3.155 58.395 4.62 ;
      RECT 58.195 3.155 58.455 3.475 ;
      RECT 57.835 4.835 58.095 5.155 ;
      RECT 57.895 3.245 58.035 5.155 ;
      RECT 57.475 3.155 57.735 3.475 ;
      RECT 57.475 3.245 58.035 3.385 ;
      RECT 55.505 4.25 55.785 4.62 ;
      RECT 57.475 4.275 57.735 4.595 ;
      RECT 55.155 4.275 55.785 4.595 ;
      RECT 55.155 4.365 57.735 4.505 ;
      RECT 56.945 3.69 57.225 4.06 ;
      RECT 56.945 3.715 57.475 4.035 ;
      RECT 54.035 4.275 54.295 4.595 ;
      RECT 54.095 3.155 54.235 4.595 ;
      RECT 54.035 3.155 54.295 3.475 ;
      RECT 53.065 4.81 53.345 5.18 ;
      RECT 53.075 4.555 53.335 5.18 ;
      RECT 48.315 8.51 48.635 8.835 ;
      RECT 48.345 7.985 48.515 8.835 ;
      RECT 48.345 7.985 48.52 8.335 ;
      RECT 48.345 7.985 49.32 8.16 ;
      RECT 49.145 3.26 49.32 8.16 ;
      RECT 49.09 3.26 49.44 3.61 ;
      RECT 49.115 8.945 49.44 9.27 ;
      RECT 48 9.035 49.44 9.205 ;
      RECT 48 3.69 48.16 9.205 ;
      RECT 48.315 3.66 48.635 3.98 ;
      RECT 48 3.69 48.635 3.86 ;
      RECT 42.835 5.43 46.97 5.62 ;
      RECT 46.8 4.44 46.97 5.62 ;
      RECT 46.78 4.445 46.97 5.62 ;
      RECT 42.835 4.81 43.025 5.62 ;
      RECT 42.785 4.81 43.065 5.18 ;
      RECT 46.71 4.445 47.05 4.795 ;
      RECT 32.935 8.945 33.285 9.295 ;
      RECT 43.68 8.9 44.03 9.25 ;
      RECT 32.935 8.975 44.03 9.175 ;
      RECT 43.315 4.275 43.575 4.595 ;
      RECT 43.375 3.155 43.515 4.595 ;
      RECT 43.315 3.155 43.575 3.475 ;
      RECT 42.315 4.835 42.575 5.155 ;
      RECT 42.315 4.25 42.515 5.155 ;
      RECT 42.255 3.155 42.395 4.785 ;
      RECT 42.255 4.25 42.755 4.62 ;
      RECT 42.195 3.155 42.455 3.475 ;
      RECT 41.835 4.835 42.095 5.155 ;
      RECT 41.895 3.245 42.035 5.155 ;
      RECT 41.595 3.245 42.035 3.475 ;
      RECT 41.595 3.155 41.855 3.475 ;
      RECT 41.355 3.715 41.615 4.035 ;
      RECT 40.775 3.805 41.615 3.945 ;
      RECT 40.775 2.865 40.915 3.945 ;
      RECT 37.435 3.155 37.695 3.475 ;
      RECT 37.435 3.245 38.475 3.385 ;
      RECT 38.335 2.865 38.475 3.385 ;
      RECT 38.335 2.865 40.915 3.005 ;
      RECT 40.825 4.81 41.105 5.18 ;
      RECT 40.895 4.365 41.035 5.18 ;
      RECT 40.705 4.25 40.985 4.62 ;
      RECT 40.415 4.365 41.035 4.505 ;
      RECT 40.415 3.155 40.555 4.505 ;
      RECT 40.355 3.155 40.615 3.475 ;
      RECT 39.625 4.25 39.905 4.62 ;
      RECT 39.695 3.155 39.835 4.62 ;
      RECT 39.635 3.155 39.895 3.475 ;
      RECT 39.275 4.835 39.535 5.155 ;
      RECT 39.335 3.245 39.475 5.155 ;
      RECT 38.915 3.155 39.175 3.475 ;
      RECT 38.915 3.245 39.475 3.385 ;
      RECT 36.945 4.25 37.225 4.62 ;
      RECT 38.915 4.275 39.175 4.595 ;
      RECT 36.595 4.275 37.225 4.595 ;
      RECT 36.595 4.365 39.175 4.505 ;
      RECT 38.385 3.69 38.665 4.06 ;
      RECT 38.385 3.715 38.915 4.035 ;
      RECT 35.475 4.275 35.735 4.595 ;
      RECT 35.535 3.155 35.675 4.595 ;
      RECT 35.475 3.155 35.735 3.475 ;
      RECT 34.505 4.81 34.785 5.18 ;
      RECT 34.515 4.555 34.775 5.18 ;
      RECT 29.755 8.51 30.075 8.835 ;
      RECT 29.785 7.985 29.955 8.835 ;
      RECT 29.785 7.985 29.96 8.335 ;
      RECT 29.785 7.985 30.76 8.16 ;
      RECT 30.585 3.26 30.76 8.16 ;
      RECT 30.53 3.26 30.88 3.61 ;
      RECT 30.555 8.945 30.88 9.27 ;
      RECT 29.44 9.035 30.88 9.205 ;
      RECT 29.44 3.69 29.6 9.205 ;
      RECT 29.755 3.66 30.075 3.98 ;
      RECT 29.44 3.69 30.075 3.86 ;
      RECT 24.275 5.43 28.41 5.62 ;
      RECT 28.24 4.44 28.41 5.62 ;
      RECT 28.22 4.445 28.41 5.62 ;
      RECT 24.275 4.81 24.465 5.62 ;
      RECT 24.225 4.81 24.505 5.18 ;
      RECT 28.15 4.445 28.49 4.795 ;
      RECT 13.67 9.285 13.96 9.635 ;
      RECT 13.67 9.34 14.985 9.51 ;
      RECT 14.815 8.975 14.985 9.51 ;
      RECT 25.12 8.895 25.47 9.245 ;
      RECT 14.815 8.975 25.47 9.145 ;
      RECT 24.755 4.275 25.015 4.595 ;
      RECT 24.815 3.155 24.955 4.595 ;
      RECT 24.755 3.155 25.015 3.475 ;
      RECT 23.755 4.835 24.015 5.155 ;
      RECT 23.755 4.25 23.955 5.155 ;
      RECT 23.695 3.155 23.835 4.785 ;
      RECT 23.695 4.25 24.195 4.62 ;
      RECT 23.635 3.155 23.895 3.475 ;
      RECT 23.275 4.835 23.535 5.155 ;
      RECT 23.335 3.245 23.475 5.155 ;
      RECT 23.035 3.245 23.475 3.475 ;
      RECT 23.035 3.155 23.295 3.475 ;
      RECT 22.795 3.715 23.055 4.035 ;
      RECT 22.215 3.805 23.055 3.945 ;
      RECT 22.215 2.865 22.355 3.945 ;
      RECT 18.875 3.155 19.135 3.475 ;
      RECT 18.875 3.245 19.915 3.385 ;
      RECT 19.775 2.865 19.915 3.385 ;
      RECT 19.775 2.865 22.355 3.005 ;
      RECT 22.265 4.81 22.545 5.18 ;
      RECT 22.335 4.365 22.475 5.18 ;
      RECT 22.145 4.25 22.425 4.62 ;
      RECT 21.855 4.365 22.475 4.505 ;
      RECT 21.855 3.155 21.995 4.505 ;
      RECT 21.795 3.155 22.055 3.475 ;
      RECT 21.065 4.25 21.345 4.62 ;
      RECT 21.135 3.155 21.275 4.62 ;
      RECT 21.075 3.155 21.335 3.475 ;
      RECT 20.715 4.835 20.975 5.155 ;
      RECT 20.775 3.245 20.915 5.155 ;
      RECT 20.355 3.155 20.615 3.475 ;
      RECT 20.355 3.245 20.915 3.385 ;
      RECT 18.385 4.25 18.665 4.62 ;
      RECT 20.355 4.275 20.615 4.595 ;
      RECT 18.035 4.275 18.665 4.595 ;
      RECT 18.035 4.365 20.615 4.505 ;
      RECT 19.825 3.69 20.105 4.06 ;
      RECT 19.825 3.715 20.355 4.035 ;
      RECT 16.915 4.275 17.175 4.595 ;
      RECT 16.975 3.155 17.115 4.595 ;
      RECT 16.915 3.155 17.175 3.475 ;
      RECT 15.945 4.81 16.225 5.18 ;
      RECT 15.955 4.555 16.215 5.18 ;
      RECT 100.425 3.13 100.705 3.5 ;
      RECT 99.465 4.81 99.745 5.18 ;
      RECT 98.685 9.345 99.06 9.715 ;
      RECT 90.665 3.69 90.945 4.06 ;
      RECT 81.865 3.13 82.145 3.5 ;
      RECT 80.905 4.81 81.185 5.18 ;
      RECT 80.125 9.345 80.5 9.715 ;
      RECT 72.105 3.69 72.385 4.06 ;
      RECT 63.305 3.13 63.585 3.5 ;
      RECT 62.345 4.81 62.625 5.18 ;
      RECT 61.565 9.345 61.94 9.715 ;
      RECT 53.545 3.69 53.825 4.06 ;
      RECT 44.745 3.13 45.025 3.5 ;
      RECT 43.785 4.81 44.065 5.18 ;
      RECT 43.005 9.345 43.38 9.715 ;
      RECT 34.985 3.69 35.265 4.06 ;
      RECT 26.185 3.13 26.465 3.5 ;
      RECT 25.225 4.81 25.505 5.18 ;
      RECT 24.445 9.345 24.82 9.715 ;
      RECT 16.425 3.69 16.705 4.06 ;
      RECT 13.81 6.555 14.19 6.935 ;
    LAYER via1 ;
      RECT 107.255 9.665 107.405 9.815 ;
      RECT 104.885 9.03 105.035 9.18 ;
      RECT 104.87 3.36 105.02 3.51 ;
      RECT 104.08 3.745 104.23 3.895 ;
      RECT 104.08 8.615 104.23 8.765 ;
      RECT 102.49 4.545 102.64 4.695 ;
      RECT 100.49 3.24 100.64 3.39 ;
      RECT 99.53 4.92 99.68 5.07 ;
      RECT 99.455 9 99.605 9.15 ;
      RECT 99.05 3.24 99.2 3.39 ;
      RECT 99.05 4.36 99.2 4.51 ;
      RECT 98.795 9.455 98.945 9.605 ;
      RECT 98.53 4.92 98.68 5.07 ;
      RECT 98.05 4.92 98.2 5.07 ;
      RECT 97.93 3.24 98.08 3.39 ;
      RECT 97.57 4.92 97.72 5.07 ;
      RECT 97.33 3.24 97.48 3.39 ;
      RECT 97.09 3.8 97.24 3.95 ;
      RECT 96.57 4.92 96.72 5.07 ;
      RECT 96.09 3.24 96.24 3.39 ;
      RECT 95.37 3.24 95.52 3.39 ;
      RECT 95.37 4.36 95.52 4.51 ;
      RECT 95.01 4.92 95.16 5.07 ;
      RECT 94.65 3.24 94.8 3.39 ;
      RECT 94.65 4.36 94.8 4.51 ;
      RECT 94.39 3.8 94.54 3.95 ;
      RECT 93.17 3.24 93.32 3.39 ;
      RECT 92.33 4.36 92.48 4.51 ;
      RECT 91.21 3.24 91.36 3.39 ;
      RECT 91.21 4.36 91.36 4.51 ;
      RECT 90.73 3.8 90.88 3.95 ;
      RECT 90.25 4.64 90.4 4.79 ;
      RECT 88.67 9.045 88.82 9.195 ;
      RECT 86.325 9.03 86.475 9.18 ;
      RECT 86.31 3.36 86.46 3.51 ;
      RECT 85.52 3.745 85.67 3.895 ;
      RECT 85.52 8.615 85.67 8.765 ;
      RECT 83.93 4.545 84.08 4.695 ;
      RECT 81.93 3.24 82.08 3.39 ;
      RECT 80.97 4.92 81.12 5.07 ;
      RECT 80.895 9 81.045 9.15 ;
      RECT 80.49 3.24 80.64 3.39 ;
      RECT 80.49 4.36 80.64 4.51 ;
      RECT 80.235 9.455 80.385 9.605 ;
      RECT 79.97 4.92 80.12 5.07 ;
      RECT 79.49 4.92 79.64 5.07 ;
      RECT 79.37 3.24 79.52 3.39 ;
      RECT 79.01 4.92 79.16 5.07 ;
      RECT 78.77 3.24 78.92 3.39 ;
      RECT 78.53 3.8 78.68 3.95 ;
      RECT 78.01 4.92 78.16 5.07 ;
      RECT 77.53 3.24 77.68 3.39 ;
      RECT 76.81 3.24 76.96 3.39 ;
      RECT 76.81 4.36 76.96 4.51 ;
      RECT 76.45 4.92 76.6 5.07 ;
      RECT 76.09 3.24 76.24 3.39 ;
      RECT 76.09 4.36 76.24 4.51 ;
      RECT 75.83 3.8 75.98 3.95 ;
      RECT 74.61 3.24 74.76 3.39 ;
      RECT 73.77 4.36 73.92 4.51 ;
      RECT 72.65 3.24 72.8 3.39 ;
      RECT 72.65 4.36 72.8 4.51 ;
      RECT 72.17 3.8 72.32 3.95 ;
      RECT 71.69 4.64 71.84 4.79 ;
      RECT 70.11 9.045 70.26 9.195 ;
      RECT 67.765 9.03 67.915 9.18 ;
      RECT 67.75 3.36 67.9 3.51 ;
      RECT 66.96 3.745 67.11 3.895 ;
      RECT 66.96 8.615 67.11 8.765 ;
      RECT 65.37 4.545 65.52 4.695 ;
      RECT 63.37 3.24 63.52 3.39 ;
      RECT 62.41 4.92 62.56 5.07 ;
      RECT 62.335 9.005 62.485 9.155 ;
      RECT 61.93 3.24 62.08 3.39 ;
      RECT 61.93 4.36 62.08 4.51 ;
      RECT 61.675 9.455 61.825 9.605 ;
      RECT 61.41 4.92 61.56 5.07 ;
      RECT 60.93 4.92 61.08 5.07 ;
      RECT 60.81 3.24 60.96 3.39 ;
      RECT 60.45 4.92 60.6 5.07 ;
      RECT 60.21 3.24 60.36 3.39 ;
      RECT 59.97 3.8 60.12 3.95 ;
      RECT 59.45 4.92 59.6 5.07 ;
      RECT 58.97 3.24 59.12 3.39 ;
      RECT 58.25 3.24 58.4 3.39 ;
      RECT 58.25 4.36 58.4 4.51 ;
      RECT 57.89 4.92 58.04 5.07 ;
      RECT 57.53 3.24 57.68 3.39 ;
      RECT 57.53 4.36 57.68 4.51 ;
      RECT 57.27 3.8 57.42 3.95 ;
      RECT 56.05 3.24 56.2 3.39 ;
      RECT 55.21 4.36 55.36 4.51 ;
      RECT 54.09 3.24 54.24 3.39 ;
      RECT 54.09 4.36 54.24 4.51 ;
      RECT 53.61 3.8 53.76 3.95 ;
      RECT 53.13 4.64 53.28 4.79 ;
      RECT 51.595 9.05 51.745 9.2 ;
      RECT 49.205 9.03 49.355 9.18 ;
      RECT 49.19 3.36 49.34 3.51 ;
      RECT 48.4 3.745 48.55 3.895 ;
      RECT 48.4 8.615 48.55 8.765 ;
      RECT 46.81 4.545 46.96 4.695 ;
      RECT 44.81 3.24 44.96 3.39 ;
      RECT 43.85 4.92 44 5.07 ;
      RECT 43.78 9 43.93 9.15 ;
      RECT 43.37 3.24 43.52 3.39 ;
      RECT 43.37 4.36 43.52 4.51 ;
      RECT 43.115 9.455 43.265 9.605 ;
      RECT 42.85 4.92 43 5.07 ;
      RECT 42.37 4.92 42.52 5.07 ;
      RECT 42.25 3.24 42.4 3.39 ;
      RECT 41.89 4.92 42.04 5.07 ;
      RECT 41.65 3.24 41.8 3.39 ;
      RECT 41.41 3.8 41.56 3.95 ;
      RECT 40.89 4.92 41.04 5.07 ;
      RECT 40.41 3.24 40.56 3.39 ;
      RECT 39.69 3.24 39.84 3.39 ;
      RECT 39.69 4.36 39.84 4.51 ;
      RECT 39.33 4.92 39.48 5.07 ;
      RECT 38.97 3.24 39.12 3.39 ;
      RECT 38.97 4.36 39.12 4.51 ;
      RECT 38.71 3.8 38.86 3.95 ;
      RECT 37.49 3.24 37.64 3.39 ;
      RECT 36.65 4.36 36.8 4.51 ;
      RECT 35.53 3.24 35.68 3.39 ;
      RECT 35.53 4.36 35.68 4.51 ;
      RECT 35.05 3.8 35.2 3.95 ;
      RECT 34.57 4.64 34.72 4.79 ;
      RECT 33.035 9.045 33.185 9.195 ;
      RECT 30.645 9.03 30.795 9.18 ;
      RECT 30.63 3.36 30.78 3.51 ;
      RECT 29.84 3.745 29.99 3.895 ;
      RECT 29.84 8.615 29.99 8.765 ;
      RECT 28.25 4.545 28.4 4.695 ;
      RECT 26.25 3.24 26.4 3.39 ;
      RECT 25.29 4.92 25.44 5.07 ;
      RECT 25.22 8.995 25.37 9.145 ;
      RECT 24.81 3.24 24.96 3.39 ;
      RECT 24.81 4.36 24.96 4.51 ;
      RECT 24.555 9.455 24.705 9.605 ;
      RECT 24.29 4.92 24.44 5.07 ;
      RECT 23.81 4.92 23.96 5.07 ;
      RECT 23.69 3.24 23.84 3.39 ;
      RECT 23.33 4.92 23.48 5.07 ;
      RECT 23.09 3.24 23.24 3.39 ;
      RECT 22.85 3.8 23 3.95 ;
      RECT 22.33 4.92 22.48 5.07 ;
      RECT 21.85 3.24 22 3.39 ;
      RECT 21.13 3.24 21.28 3.39 ;
      RECT 21.13 4.36 21.28 4.51 ;
      RECT 20.77 4.92 20.92 5.07 ;
      RECT 20.41 3.24 20.56 3.39 ;
      RECT 20.41 4.36 20.56 4.51 ;
      RECT 20.15 3.8 20.3 3.95 ;
      RECT 18.93 3.24 19.08 3.39 ;
      RECT 18.09 4.36 18.24 4.51 ;
      RECT 16.97 3.24 17.12 3.39 ;
      RECT 16.97 4.36 17.12 4.51 ;
      RECT 16.49 3.8 16.64 3.95 ;
      RECT 16.01 4.64 16.16 4.79 ;
      RECT 13.925 6.67 14.075 6.82 ;
      RECT 13.74 9.385 13.89 9.535 ;
      RECT 13.365 8.645 13.515 8.795 ;
    LAYER met1 ;
      RECT 12.125 5.45 107.725 7.05 ;
      RECT 14.94 5.425 107.74 7.025 ;
      RECT 89.91 5.275 101.87 7.05 ;
      RECT 71.35 5.275 83.31 7.05 ;
      RECT 52.79 5.275 64.75 7.05 ;
      RECT 34.23 5.275 46.19 7.05 ;
      RECT 15.67 5.275 27.63 7.05 ;
      RECT 107.12 10.055 107.41 10.285 ;
      RECT 107.18 8.575 107.35 10.285 ;
      RECT 107.155 9.565 107.505 9.915 ;
      RECT 107.12 8.575 107.41 8.805 ;
      RECT 106.75 4.03 107.04 4.26 ;
      RECT 106.715 3.725 106.905 4.255 ;
      RECT 106.715 4.06 107.21 4.23 ;
      RECT 106.36 3.725 106.905 3.895 ;
      RECT 106.19 2.18 106.36 3.89 ;
      RECT 106.13 3.66 106.42 3.89 ;
      RECT 106.13 2.18 106.42 2.41 ;
      RECT 106.13 10.055 106.42 10.285 ;
      RECT 106.19 8.575 106.36 10.285 ;
      RECT 106.19 8.81 106.98 8.97 ;
      RECT 106.825 8.205 106.98 8.97 ;
      RECT 106.815 8.63 106.98 8.97 ;
      RECT 106.19 8.575 106.42 8.97 ;
      RECT 106.13 8.575 106.42 8.805 ;
      RECT 106.75 8.205 107.04 8.435 ;
      RECT 106.75 8.235 107.21 8.405 ;
      RECT 105.825 4.03 105.995 4.335 ;
      RECT 105.76 4.03 106.05 4.26 ;
      RECT 105.76 4.06 106.22 4.23 ;
      RECT 105.825 2.95 105.99 4.335 ;
      RECT 104.34 2.92 104.63 3.15 ;
      RECT 104.34 2.95 105.99 3.12 ;
      RECT 104.4 2.18 104.57 3.15 ;
      RECT 104.34 2.18 104.63 2.41 ;
      RECT 104.34 10.055 104.63 10.285 ;
      RECT 104.4 9.315 104.57 10.285 ;
      RECT 104.4 9.41 105.99 9.58 ;
      RECT 105.82 8.205 105.99 9.58 ;
      RECT 104.34 9.315 104.63 9.545 ;
      RECT 105.76 8.205 106.05 8.435 ;
      RECT 105.76 8.235 106.22 8.405 ;
      RECT 102.39 4.445 102.73 4.795 ;
      RECT 102.48 3.32 102.65 4.795 ;
      RECT 104.77 3.26 105.12 3.61 ;
      RECT 102.48 3.32 105.12 3.49 ;
      RECT 104.795 8.945 105.12 9.27 ;
      RECT 99.355 8.9 99.705 9.25 ;
      RECT 104.77 8.945 105.12 9.175 ;
      RECT 99.155 8.945 99.705 9.175 ;
      RECT 98.985 8.975 105.12 9.145 ;
      RECT 103.995 3.66 104.315 3.98 ;
      RECT 103.965 3.66 104.315 3.89 ;
      RECT 103.795 3.69 104.315 3.86 ;
      RECT 103.995 8.545 104.315 8.835 ;
      RECT 103.965 8.575 104.315 8.805 ;
      RECT 103.795 8.605 104.315 8.775 ;
      RECT 99.445 4.865 99.765 5.125 ;
      RECT 100.735 4.04 100.875 4.9 ;
      RECT 99.535 4.76 100.875 4.9 ;
      RECT 99.535 4.32 99.675 5.125 ;
      RECT 99.46 4.32 99.75 4.55 ;
      RECT 100.66 4.04 100.95 4.27 ;
      RECT 100.18 4.32 100.47 4.55 ;
      RECT 100.375 3.245 100.515 4.505 ;
      RECT 100.405 3.185 100.725 3.445 ;
      RECT 97.005 3.745 97.325 4.005 ;
      RECT 99.7 3.76 99.99 3.99 ;
      RECT 97.095 3.665 99.915 3.805 ;
      RECT 98.965 3.185 99.285 3.445 ;
      RECT 99.46 3.2 99.75 3.43 ;
      RECT 98.965 3.245 99.75 3.385 ;
      RECT 98.965 4.305 99.285 4.565 ;
      RECT 98.965 4.085 99.195 4.565 ;
      RECT 98.46 4.04 98.75 4.27 ;
      RECT 98.46 4.085 99.195 4.225 ;
      RECT 98.725 10.055 99.015 10.285 ;
      RECT 98.785 9.315 98.955 10.285 ;
      RECT 98.685 9.345 99.065 9.715 ;
      RECT 98.725 9.315 99.015 9.715 ;
      RECT 97.485 4.865 97.805 5.125 ;
      RECT 97.02 4.88 97.31 5.11 ;
      RECT 97.02 4.925 97.805 5.065 ;
      RECT 95.78 3.76 96.07 3.99 ;
      RECT 95.78 3.805 96.715 3.945 ;
      RECT 96.575 3.245 96.715 3.945 ;
      RECT 97.245 3.185 97.565 3.445 ;
      RECT 97.02 3.2 97.565 3.43 ;
      RECT 96.575 3.245 97.565 3.385 ;
      RECT 94.925 4.865 95.245 5.125 ;
      RECT 94.925 4.925 95.995 5.065 ;
      RECT 95.855 4.365 95.995 5.065 ;
      RECT 97.02 4.32 97.31 4.55 ;
      RECT 95.855 4.365 97.31 4.505 ;
      RECT 95.285 3.185 95.605 3.445 ;
      RECT 95.06 3.2 95.605 3.43 ;
      RECT 94.305 3.745 94.625 4.005 ;
      RECT 95.3 3.76 95.59 3.99 ;
      RECT 94.06 3.76 94.625 3.99 ;
      RECT 94.06 3.805 95.59 3.945 ;
      RECT 93.58 4.32 93.87 4.55 ;
      RECT 93.775 3.245 93.915 4.505 ;
      RECT 94.565 3.185 94.885 3.445 ;
      RECT 93.58 3.2 93.87 3.43 ;
      RECT 93.58 3.245 94.885 3.385 ;
      RECT 93.175 4.76 94.275 4.9 ;
      RECT 94.06 4.6 94.35 4.83 ;
      RECT 93.1 4.6 93.39 4.83 ;
      RECT 93.085 3.185 93.405 3.445 ;
      RECT 91.125 3.185 91.445 3.445 ;
      RECT 91.125 3.245 93.405 3.385 ;
      RECT 92.245 4.305 92.565 4.565 ;
      RECT 92.245 4.305 93.075 4.445 ;
      RECT 92.86 4.04 93.075 4.445 ;
      RECT 92.86 4.04 93.15 4.27 ;
      RECT 90.645 3.745 90.965 4.005 ;
      RECT 92.055 3.76 92.345 3.99 ;
      RECT 90.645 3.76 91.19 3.99 ;
      RECT 90.645 3.845 91.595 3.985 ;
      RECT 91.455 3.665 91.595 3.985 ;
      RECT 91.955 3.76 92.345 3.945 ;
      RECT 91.455 3.665 92.095 3.805 ;
      RECT 90.165 4.555 90.485 4.97 ;
      RECT 90.245 3.2 90.4 4.97 ;
      RECT 90.18 3.2 90.47 3.43 ;
      RECT 88.56 10.055 88.85 10.285 ;
      RECT 88.62 8.575 88.79 10.285 ;
      RECT 88.57 8.945 88.92 9.295 ;
      RECT 88.56 8.575 88.85 8.805 ;
      RECT 88.19 4.03 88.48 4.26 ;
      RECT 88.155 3.725 88.345 4.255 ;
      RECT 88.155 4.06 88.65 4.23 ;
      RECT 87.8 3.725 88.345 3.895 ;
      RECT 87.63 2.18 87.8 3.89 ;
      RECT 87.57 3.66 87.86 3.89 ;
      RECT 87.57 2.18 87.86 2.41 ;
      RECT 87.57 10.055 87.86 10.285 ;
      RECT 87.63 8.575 87.8 10.285 ;
      RECT 87.63 8.81 88.42 8.97 ;
      RECT 88.265 8.205 88.42 8.97 ;
      RECT 88.255 8.63 88.42 8.97 ;
      RECT 87.63 8.575 87.86 8.97 ;
      RECT 87.57 8.575 87.86 8.805 ;
      RECT 88.19 8.205 88.48 8.435 ;
      RECT 88.19 8.235 88.65 8.405 ;
      RECT 87.265 4.03 87.435 4.335 ;
      RECT 87.2 4.03 87.49 4.26 ;
      RECT 87.2 4.06 87.66 4.23 ;
      RECT 87.265 2.95 87.43 4.335 ;
      RECT 85.78 2.92 86.07 3.15 ;
      RECT 85.78 2.95 87.43 3.12 ;
      RECT 85.84 2.18 86.01 3.15 ;
      RECT 85.78 2.18 86.07 2.41 ;
      RECT 85.78 10.055 86.07 10.285 ;
      RECT 85.84 9.315 86.01 10.285 ;
      RECT 85.84 9.41 87.43 9.58 ;
      RECT 87.26 8.205 87.43 9.58 ;
      RECT 85.78 9.315 86.07 9.545 ;
      RECT 87.2 8.205 87.49 8.435 ;
      RECT 87.2 8.235 87.66 8.405 ;
      RECT 83.83 4.445 84.17 4.795 ;
      RECT 83.92 3.32 84.09 4.795 ;
      RECT 86.21 3.26 86.56 3.61 ;
      RECT 83.92 3.32 86.56 3.49 ;
      RECT 86.235 8.945 86.56 9.27 ;
      RECT 80.795 8.9 81.145 9.25 ;
      RECT 86.21 8.945 86.56 9.175 ;
      RECT 80.595 8.945 81.145 9.175 ;
      RECT 80.425 8.975 86.56 9.145 ;
      RECT 85.435 3.66 85.755 3.98 ;
      RECT 85.405 3.66 85.755 3.89 ;
      RECT 85.235 3.69 85.755 3.86 ;
      RECT 85.435 8.545 85.755 8.835 ;
      RECT 85.405 8.575 85.755 8.805 ;
      RECT 85.235 8.605 85.755 8.775 ;
      RECT 80.885 4.865 81.205 5.125 ;
      RECT 82.175 4.04 82.315 4.9 ;
      RECT 80.975 4.76 82.315 4.9 ;
      RECT 80.975 4.32 81.115 5.125 ;
      RECT 80.9 4.32 81.19 4.55 ;
      RECT 82.1 4.04 82.39 4.27 ;
      RECT 81.62 4.32 81.91 4.55 ;
      RECT 81.815 3.245 81.955 4.505 ;
      RECT 81.845 3.185 82.165 3.445 ;
      RECT 78.445 3.745 78.765 4.005 ;
      RECT 81.14 3.76 81.43 3.99 ;
      RECT 78.535 3.665 81.355 3.805 ;
      RECT 80.405 3.185 80.725 3.445 ;
      RECT 80.9 3.2 81.19 3.43 ;
      RECT 80.405 3.245 81.19 3.385 ;
      RECT 80.405 4.305 80.725 4.565 ;
      RECT 80.405 4.085 80.635 4.565 ;
      RECT 79.9 4.04 80.19 4.27 ;
      RECT 79.9 4.085 80.635 4.225 ;
      RECT 80.165 10.055 80.455 10.285 ;
      RECT 80.225 9.315 80.395 10.285 ;
      RECT 80.125 9.345 80.505 9.715 ;
      RECT 80.165 9.315 80.455 9.715 ;
      RECT 78.925 4.865 79.245 5.125 ;
      RECT 78.46 4.88 78.75 5.11 ;
      RECT 78.46 4.925 79.245 5.065 ;
      RECT 77.22 3.76 77.51 3.99 ;
      RECT 77.22 3.805 78.155 3.945 ;
      RECT 78.015 3.245 78.155 3.945 ;
      RECT 78.685 3.185 79.005 3.445 ;
      RECT 78.46 3.2 79.005 3.43 ;
      RECT 78.015 3.245 79.005 3.385 ;
      RECT 76.365 4.865 76.685 5.125 ;
      RECT 76.365 4.925 77.435 5.065 ;
      RECT 77.295 4.365 77.435 5.065 ;
      RECT 78.46 4.32 78.75 4.55 ;
      RECT 77.295 4.365 78.75 4.505 ;
      RECT 76.725 3.185 77.045 3.445 ;
      RECT 76.5 3.2 77.045 3.43 ;
      RECT 75.745 3.745 76.065 4.005 ;
      RECT 76.74 3.76 77.03 3.99 ;
      RECT 75.5 3.76 76.065 3.99 ;
      RECT 75.5 3.805 77.03 3.945 ;
      RECT 75.02 4.32 75.31 4.55 ;
      RECT 75.215 3.245 75.355 4.505 ;
      RECT 76.005 3.185 76.325 3.445 ;
      RECT 75.02 3.2 75.31 3.43 ;
      RECT 75.02 3.245 76.325 3.385 ;
      RECT 74.615 4.76 75.715 4.9 ;
      RECT 75.5 4.6 75.79 4.83 ;
      RECT 74.54 4.6 74.83 4.83 ;
      RECT 74.525 3.185 74.845 3.445 ;
      RECT 72.565 3.185 72.885 3.445 ;
      RECT 72.565 3.245 74.845 3.385 ;
      RECT 73.685 4.305 74.005 4.565 ;
      RECT 73.685 4.305 74.515 4.445 ;
      RECT 74.3 4.04 74.515 4.445 ;
      RECT 74.3 4.04 74.59 4.27 ;
      RECT 72.085 3.745 72.405 4.005 ;
      RECT 73.495 3.76 73.785 3.99 ;
      RECT 72.085 3.76 72.63 3.99 ;
      RECT 72.085 3.845 73.035 3.985 ;
      RECT 72.895 3.665 73.035 3.985 ;
      RECT 73.395 3.76 73.785 3.945 ;
      RECT 72.895 3.665 73.535 3.805 ;
      RECT 71.605 4.555 71.925 4.97 ;
      RECT 71.685 3.2 71.84 4.97 ;
      RECT 71.62 3.2 71.91 3.43 ;
      RECT 70 10.055 70.29 10.285 ;
      RECT 70.06 8.575 70.23 10.285 ;
      RECT 70.01 8.945 70.36 9.295 ;
      RECT 70 8.575 70.29 8.805 ;
      RECT 69.63 4.03 69.92 4.26 ;
      RECT 69.595 3.725 69.785 4.255 ;
      RECT 69.595 4.06 70.09 4.23 ;
      RECT 69.24 3.725 69.785 3.895 ;
      RECT 69.07 2.18 69.24 3.89 ;
      RECT 69.01 3.66 69.3 3.89 ;
      RECT 69.01 2.18 69.3 2.41 ;
      RECT 69.01 10.055 69.3 10.285 ;
      RECT 69.07 8.575 69.24 10.285 ;
      RECT 69.07 8.81 69.86 8.97 ;
      RECT 69.705 8.205 69.86 8.97 ;
      RECT 69.695 8.63 69.86 8.97 ;
      RECT 69.07 8.575 69.3 8.97 ;
      RECT 69.01 8.575 69.3 8.805 ;
      RECT 69.63 8.205 69.92 8.435 ;
      RECT 69.63 8.235 70.09 8.405 ;
      RECT 68.705 4.03 68.875 4.335 ;
      RECT 68.64 4.03 68.93 4.26 ;
      RECT 68.64 4.06 69.1 4.23 ;
      RECT 68.705 2.95 68.87 4.335 ;
      RECT 67.22 2.92 67.51 3.15 ;
      RECT 67.22 2.95 68.87 3.12 ;
      RECT 67.28 2.18 67.45 3.15 ;
      RECT 67.22 2.18 67.51 2.41 ;
      RECT 67.22 10.055 67.51 10.285 ;
      RECT 67.28 9.315 67.45 10.285 ;
      RECT 67.28 9.41 68.87 9.58 ;
      RECT 68.7 8.205 68.87 9.58 ;
      RECT 67.22 9.315 67.51 9.545 ;
      RECT 68.64 8.205 68.93 8.435 ;
      RECT 68.64 8.235 69.1 8.405 ;
      RECT 65.27 4.445 65.61 4.795 ;
      RECT 65.36 3.32 65.53 4.795 ;
      RECT 67.65 3.26 68 3.61 ;
      RECT 65.36 3.32 68 3.49 ;
      RECT 67.675 8.945 68 9.27 ;
      RECT 62.235 8.905 62.585 9.255 ;
      RECT 67.65 8.945 68 9.175 ;
      RECT 62.035 8.945 62.585 9.175 ;
      RECT 61.865 8.975 68 9.145 ;
      RECT 66.875 3.66 67.195 3.98 ;
      RECT 66.845 3.66 67.195 3.89 ;
      RECT 66.675 3.69 67.195 3.86 ;
      RECT 66.875 8.545 67.195 8.835 ;
      RECT 66.845 8.575 67.195 8.805 ;
      RECT 66.675 8.605 67.195 8.775 ;
      RECT 62.325 4.865 62.645 5.125 ;
      RECT 63.615 4.04 63.755 4.9 ;
      RECT 62.415 4.76 63.755 4.9 ;
      RECT 62.415 4.32 62.555 5.125 ;
      RECT 62.34 4.32 62.63 4.55 ;
      RECT 63.54 4.04 63.83 4.27 ;
      RECT 63.06 4.32 63.35 4.55 ;
      RECT 63.255 3.245 63.395 4.505 ;
      RECT 63.285 3.185 63.605 3.445 ;
      RECT 59.885 3.745 60.205 4.005 ;
      RECT 62.58 3.76 62.87 3.99 ;
      RECT 59.975 3.665 62.795 3.805 ;
      RECT 61.845 3.185 62.165 3.445 ;
      RECT 62.34 3.2 62.63 3.43 ;
      RECT 61.845 3.245 62.63 3.385 ;
      RECT 61.845 4.305 62.165 4.565 ;
      RECT 61.845 4.085 62.075 4.565 ;
      RECT 61.34 4.04 61.63 4.27 ;
      RECT 61.34 4.085 62.075 4.225 ;
      RECT 61.605 10.055 61.895 10.285 ;
      RECT 61.665 9.315 61.835 10.285 ;
      RECT 61.565 9.345 61.945 9.715 ;
      RECT 61.605 9.315 61.895 9.715 ;
      RECT 60.365 4.865 60.685 5.125 ;
      RECT 59.9 4.88 60.19 5.11 ;
      RECT 59.9 4.925 60.685 5.065 ;
      RECT 58.66 3.76 58.95 3.99 ;
      RECT 58.66 3.805 59.595 3.945 ;
      RECT 59.455 3.245 59.595 3.945 ;
      RECT 60.125 3.185 60.445 3.445 ;
      RECT 59.9 3.2 60.445 3.43 ;
      RECT 59.455 3.245 60.445 3.385 ;
      RECT 57.805 4.865 58.125 5.125 ;
      RECT 57.805 4.925 58.875 5.065 ;
      RECT 58.735 4.365 58.875 5.065 ;
      RECT 59.9 4.32 60.19 4.55 ;
      RECT 58.735 4.365 60.19 4.505 ;
      RECT 58.165 3.185 58.485 3.445 ;
      RECT 57.94 3.2 58.485 3.43 ;
      RECT 57.185 3.745 57.505 4.005 ;
      RECT 58.18 3.76 58.47 3.99 ;
      RECT 56.94 3.76 57.505 3.99 ;
      RECT 56.94 3.805 58.47 3.945 ;
      RECT 56.46 4.32 56.75 4.55 ;
      RECT 56.655 3.245 56.795 4.505 ;
      RECT 57.445 3.185 57.765 3.445 ;
      RECT 56.46 3.2 56.75 3.43 ;
      RECT 56.46 3.245 57.765 3.385 ;
      RECT 56.055 4.76 57.155 4.9 ;
      RECT 56.94 4.6 57.23 4.83 ;
      RECT 55.98 4.6 56.27 4.83 ;
      RECT 55.965 3.185 56.285 3.445 ;
      RECT 54.005 3.185 54.325 3.445 ;
      RECT 54.005 3.245 56.285 3.385 ;
      RECT 55.125 4.305 55.445 4.565 ;
      RECT 55.125 4.305 55.955 4.445 ;
      RECT 55.74 4.04 55.955 4.445 ;
      RECT 55.74 4.04 56.03 4.27 ;
      RECT 53.525 3.745 53.845 4.005 ;
      RECT 54.935 3.76 55.225 3.99 ;
      RECT 53.525 3.76 54.07 3.99 ;
      RECT 53.525 3.845 54.475 3.985 ;
      RECT 54.335 3.665 54.475 3.985 ;
      RECT 54.835 3.76 55.225 3.945 ;
      RECT 54.335 3.665 54.975 3.805 ;
      RECT 53.045 4.555 53.365 4.97 ;
      RECT 53.125 3.2 53.28 4.97 ;
      RECT 53.06 3.2 53.35 3.43 ;
      RECT 51.44 10.055 51.73 10.285 ;
      RECT 51.5 8.575 51.67 10.285 ;
      RECT 51.49 8.95 51.845 9.305 ;
      RECT 51.44 8.575 51.73 8.805 ;
      RECT 51.07 4.03 51.36 4.26 ;
      RECT 51.035 3.725 51.225 4.255 ;
      RECT 51.035 4.06 51.53 4.23 ;
      RECT 50.68 3.725 51.225 3.895 ;
      RECT 50.51 2.18 50.68 3.89 ;
      RECT 50.45 3.66 50.74 3.89 ;
      RECT 50.45 2.18 50.74 2.41 ;
      RECT 50.45 10.055 50.74 10.285 ;
      RECT 50.51 8.575 50.68 10.285 ;
      RECT 50.51 8.81 51.3 8.97 ;
      RECT 51.145 8.205 51.3 8.97 ;
      RECT 51.135 8.63 51.3 8.97 ;
      RECT 50.51 8.575 50.74 8.97 ;
      RECT 50.45 8.575 50.74 8.805 ;
      RECT 51.07 8.205 51.36 8.435 ;
      RECT 51.07 8.235 51.53 8.405 ;
      RECT 50.145 4.03 50.315 4.335 ;
      RECT 50.08 4.03 50.37 4.26 ;
      RECT 50.08 4.06 50.54 4.23 ;
      RECT 50.145 2.95 50.31 4.335 ;
      RECT 48.66 2.92 48.95 3.15 ;
      RECT 48.66 2.95 50.31 3.12 ;
      RECT 48.72 2.18 48.89 3.15 ;
      RECT 48.66 2.18 48.95 2.41 ;
      RECT 48.66 10.055 48.95 10.285 ;
      RECT 48.72 9.315 48.89 10.285 ;
      RECT 48.72 9.41 50.31 9.58 ;
      RECT 50.14 8.205 50.31 9.58 ;
      RECT 48.66 9.315 48.95 9.545 ;
      RECT 50.08 8.205 50.37 8.435 ;
      RECT 50.08 8.235 50.54 8.405 ;
      RECT 46.71 4.445 47.05 4.795 ;
      RECT 46.8 3.32 46.97 4.795 ;
      RECT 49.09 3.26 49.44 3.61 ;
      RECT 46.8 3.32 49.44 3.49 ;
      RECT 49.115 8.945 49.44 9.27 ;
      RECT 43.68 8.9 44.03 9.25 ;
      RECT 49.09 8.945 49.44 9.175 ;
      RECT 43.475 8.945 44.03 9.175 ;
      RECT 43.305 8.975 49.44 9.145 ;
      RECT 48.315 3.66 48.635 3.98 ;
      RECT 48.285 3.66 48.635 3.89 ;
      RECT 48.115 3.69 48.635 3.86 ;
      RECT 48.315 8.545 48.635 8.835 ;
      RECT 48.285 8.575 48.635 8.805 ;
      RECT 48.115 8.605 48.635 8.775 ;
      RECT 43.765 4.865 44.085 5.125 ;
      RECT 45.055 4.04 45.195 4.9 ;
      RECT 43.855 4.76 45.195 4.9 ;
      RECT 43.855 4.32 43.995 5.125 ;
      RECT 43.78 4.32 44.07 4.55 ;
      RECT 44.98 4.04 45.27 4.27 ;
      RECT 44.5 4.32 44.79 4.55 ;
      RECT 44.695 3.245 44.835 4.505 ;
      RECT 44.725 3.185 45.045 3.445 ;
      RECT 41.325 3.745 41.645 4.005 ;
      RECT 44.02 3.76 44.31 3.99 ;
      RECT 41.415 3.665 44.235 3.805 ;
      RECT 43.285 3.185 43.605 3.445 ;
      RECT 43.78 3.2 44.07 3.43 ;
      RECT 43.285 3.245 44.07 3.385 ;
      RECT 43.285 4.305 43.605 4.565 ;
      RECT 43.285 4.085 43.515 4.565 ;
      RECT 42.78 4.04 43.07 4.27 ;
      RECT 42.78 4.085 43.515 4.225 ;
      RECT 43.045 10.055 43.335 10.285 ;
      RECT 43.105 9.315 43.275 10.285 ;
      RECT 43.005 9.345 43.385 9.715 ;
      RECT 43.045 9.315 43.335 9.715 ;
      RECT 41.805 4.865 42.125 5.125 ;
      RECT 41.34 4.88 41.63 5.11 ;
      RECT 41.34 4.925 42.125 5.065 ;
      RECT 40.1 3.76 40.39 3.99 ;
      RECT 40.1 3.805 41.035 3.945 ;
      RECT 40.895 3.245 41.035 3.945 ;
      RECT 41.565 3.185 41.885 3.445 ;
      RECT 41.34 3.2 41.885 3.43 ;
      RECT 40.895 3.245 41.885 3.385 ;
      RECT 39.245 4.865 39.565 5.125 ;
      RECT 39.245 4.925 40.315 5.065 ;
      RECT 40.175 4.365 40.315 5.065 ;
      RECT 41.34 4.32 41.63 4.55 ;
      RECT 40.175 4.365 41.63 4.505 ;
      RECT 39.605 3.185 39.925 3.445 ;
      RECT 39.38 3.2 39.925 3.43 ;
      RECT 38.625 3.745 38.945 4.005 ;
      RECT 39.62 3.76 39.91 3.99 ;
      RECT 38.38 3.76 38.945 3.99 ;
      RECT 38.38 3.805 39.91 3.945 ;
      RECT 37.9 4.32 38.19 4.55 ;
      RECT 38.095 3.245 38.235 4.505 ;
      RECT 38.885 3.185 39.205 3.445 ;
      RECT 37.9 3.2 38.19 3.43 ;
      RECT 37.9 3.245 39.205 3.385 ;
      RECT 37.495 4.76 38.595 4.9 ;
      RECT 38.38 4.6 38.67 4.83 ;
      RECT 37.42 4.6 37.71 4.83 ;
      RECT 37.405 3.185 37.725 3.445 ;
      RECT 35.445 3.185 35.765 3.445 ;
      RECT 35.445 3.245 37.725 3.385 ;
      RECT 36.565 4.305 36.885 4.565 ;
      RECT 36.565 4.305 37.395 4.445 ;
      RECT 37.18 4.04 37.395 4.445 ;
      RECT 37.18 4.04 37.47 4.27 ;
      RECT 34.965 3.745 35.285 4.005 ;
      RECT 36.375 3.76 36.665 3.99 ;
      RECT 34.965 3.76 35.51 3.99 ;
      RECT 34.965 3.845 35.915 3.985 ;
      RECT 35.775 3.665 35.915 3.985 ;
      RECT 36.275 3.76 36.665 3.945 ;
      RECT 35.775 3.665 36.415 3.805 ;
      RECT 34.485 4.555 34.805 4.97 ;
      RECT 34.565 3.2 34.72 4.97 ;
      RECT 34.5 3.2 34.79 3.43 ;
      RECT 32.88 10.055 33.17 10.285 ;
      RECT 32.94 8.575 33.11 10.285 ;
      RECT 32.935 8.945 33.285 9.295 ;
      RECT 32.88 8.575 33.17 8.805 ;
      RECT 32.51 4.03 32.8 4.26 ;
      RECT 32.475 3.725 32.665 4.255 ;
      RECT 32.475 4.06 32.97 4.23 ;
      RECT 32.12 3.725 32.665 3.895 ;
      RECT 31.95 2.18 32.12 3.89 ;
      RECT 31.89 3.66 32.18 3.89 ;
      RECT 31.89 2.18 32.18 2.41 ;
      RECT 31.89 10.055 32.18 10.285 ;
      RECT 31.95 8.575 32.12 10.285 ;
      RECT 31.95 8.81 32.74 8.97 ;
      RECT 32.585 8.205 32.74 8.97 ;
      RECT 32.575 8.63 32.74 8.97 ;
      RECT 31.95 8.575 32.18 8.97 ;
      RECT 31.89 8.575 32.18 8.805 ;
      RECT 32.51 8.205 32.8 8.435 ;
      RECT 32.51 8.235 32.97 8.405 ;
      RECT 31.585 4.03 31.755 4.335 ;
      RECT 31.52 4.03 31.81 4.26 ;
      RECT 31.52 4.06 31.98 4.23 ;
      RECT 31.585 2.95 31.75 4.335 ;
      RECT 30.1 2.92 30.39 3.15 ;
      RECT 30.1 2.95 31.75 3.12 ;
      RECT 30.16 2.18 30.33 3.15 ;
      RECT 30.1 2.18 30.39 2.41 ;
      RECT 30.1 10.055 30.39 10.285 ;
      RECT 30.16 9.315 30.33 10.285 ;
      RECT 30.16 9.41 31.75 9.58 ;
      RECT 31.58 8.205 31.75 9.58 ;
      RECT 30.1 9.315 30.39 9.545 ;
      RECT 31.52 8.205 31.81 8.435 ;
      RECT 31.52 8.235 31.98 8.405 ;
      RECT 28.15 4.445 28.49 4.795 ;
      RECT 28.24 3.32 28.41 4.795 ;
      RECT 30.53 3.26 30.88 3.61 ;
      RECT 28.24 3.32 30.88 3.49 ;
      RECT 30.555 8.945 30.88 9.27 ;
      RECT 25.12 8.895 25.47 9.245 ;
      RECT 30.53 8.945 30.88 9.175 ;
      RECT 24.915 8.945 25.47 9.175 ;
      RECT 24.745 8.975 30.88 9.145 ;
      RECT 29.755 3.66 30.075 3.98 ;
      RECT 29.725 3.66 30.075 3.89 ;
      RECT 29.555 3.69 30.075 3.86 ;
      RECT 29.755 8.545 30.075 8.835 ;
      RECT 29.725 8.575 30.075 8.805 ;
      RECT 29.555 8.605 30.075 8.775 ;
      RECT 25.205 4.865 25.525 5.125 ;
      RECT 26.495 4.04 26.635 4.9 ;
      RECT 25.295 4.76 26.635 4.9 ;
      RECT 25.295 4.32 25.435 5.125 ;
      RECT 25.22 4.32 25.51 4.55 ;
      RECT 26.42 4.04 26.71 4.27 ;
      RECT 25.94 4.32 26.23 4.55 ;
      RECT 26.135 3.245 26.275 4.505 ;
      RECT 26.165 3.185 26.485 3.445 ;
      RECT 22.765 3.745 23.085 4.005 ;
      RECT 25.46 3.76 25.75 3.99 ;
      RECT 22.855 3.665 25.675 3.805 ;
      RECT 24.725 3.185 25.045 3.445 ;
      RECT 25.22 3.2 25.51 3.43 ;
      RECT 24.725 3.245 25.51 3.385 ;
      RECT 24.725 4.305 25.045 4.565 ;
      RECT 24.725 4.085 24.955 4.565 ;
      RECT 24.22 4.04 24.51 4.27 ;
      RECT 24.22 4.085 24.955 4.225 ;
      RECT 24.485 10.055 24.775 10.285 ;
      RECT 24.545 9.315 24.715 10.285 ;
      RECT 24.445 9.345 24.825 9.715 ;
      RECT 24.485 9.315 24.775 9.715 ;
      RECT 23.245 4.865 23.565 5.125 ;
      RECT 22.78 4.88 23.07 5.11 ;
      RECT 22.78 4.925 23.565 5.065 ;
      RECT 21.54 3.76 21.83 3.99 ;
      RECT 21.54 3.805 22.475 3.945 ;
      RECT 22.335 3.245 22.475 3.945 ;
      RECT 23.005 3.185 23.325 3.445 ;
      RECT 22.78 3.2 23.325 3.43 ;
      RECT 22.335 3.245 23.325 3.385 ;
      RECT 20.685 4.865 21.005 5.125 ;
      RECT 20.685 4.925 21.755 5.065 ;
      RECT 21.615 4.365 21.755 5.065 ;
      RECT 22.78 4.32 23.07 4.55 ;
      RECT 21.615 4.365 23.07 4.505 ;
      RECT 21.045 3.185 21.365 3.445 ;
      RECT 20.82 3.2 21.365 3.43 ;
      RECT 20.065 3.745 20.385 4.005 ;
      RECT 21.06 3.76 21.35 3.99 ;
      RECT 19.82 3.76 20.385 3.99 ;
      RECT 19.82 3.805 21.35 3.945 ;
      RECT 19.34 4.32 19.63 4.55 ;
      RECT 19.535 3.245 19.675 4.505 ;
      RECT 20.325 3.185 20.645 3.445 ;
      RECT 19.34 3.2 19.63 3.43 ;
      RECT 19.34 3.245 20.645 3.385 ;
      RECT 18.935 4.76 20.035 4.9 ;
      RECT 19.82 4.6 20.11 4.83 ;
      RECT 18.86 4.6 19.15 4.83 ;
      RECT 18.845 3.185 19.165 3.445 ;
      RECT 16.885 3.185 17.205 3.445 ;
      RECT 16.885 3.245 19.165 3.385 ;
      RECT 18.005 4.305 18.325 4.565 ;
      RECT 18.005 4.305 18.835 4.445 ;
      RECT 18.62 4.04 18.835 4.445 ;
      RECT 18.62 4.04 18.91 4.27 ;
      RECT 16.405 3.745 16.725 4.005 ;
      RECT 17.815 3.76 18.105 3.99 ;
      RECT 16.405 3.76 16.95 3.99 ;
      RECT 16.405 3.845 17.355 3.985 ;
      RECT 17.215 3.665 17.355 3.985 ;
      RECT 17.715 3.76 18.105 3.945 ;
      RECT 17.215 3.665 17.855 3.805 ;
      RECT 15.925 4.555 16.245 4.97 ;
      RECT 16.005 3.2 16.16 4.97 ;
      RECT 15.94 3.2 16.23 3.43 ;
      RECT 14.1 8.945 14.39 9.175 ;
      RECT 13.93 8.975 14.39 9.145 ;
      RECT 13.67 10.055 13.96 10.285 ;
      RECT 13.73 9.315 13.9 10.285 ;
      RECT 13.64 9.315 13.99 9.605 ;
      RECT 13.265 8.575 13.615 8.865 ;
      RECT 13.125 8.605 13.615 8.775 ;
      RECT 98.445 4.865 98.765 5.125 ;
      RECT 97.845 3.185 98.525 3.445 ;
      RECT 97.965 4.865 98.285 5.125 ;
      RECT 96.485 4.865 96.805 5.125 ;
      RECT 96.005 3.185 96.325 3.445 ;
      RECT 95.285 4.305 95.605 4.565 ;
      RECT 94.565 4.305 94.885 4.565 ;
      RECT 91.125 4.305 91.445 4.565 ;
      RECT 79.885 4.865 80.205 5.125 ;
      RECT 79.285 3.185 79.965 3.445 ;
      RECT 79.405 4.865 79.725 5.125 ;
      RECT 77.925 4.865 78.245 5.125 ;
      RECT 77.445 3.185 77.765 3.445 ;
      RECT 76.725 4.305 77.045 4.565 ;
      RECT 76.005 4.305 76.325 4.565 ;
      RECT 72.565 4.305 72.885 4.565 ;
      RECT 61.325 4.865 61.645 5.125 ;
      RECT 60.725 3.185 61.405 3.445 ;
      RECT 60.845 4.865 61.165 5.125 ;
      RECT 59.365 4.865 59.685 5.125 ;
      RECT 58.885 3.185 59.205 3.445 ;
      RECT 58.165 4.305 58.485 4.565 ;
      RECT 57.445 4.305 57.765 4.565 ;
      RECT 54.005 4.305 54.325 4.565 ;
      RECT 42.765 4.865 43.085 5.125 ;
      RECT 42.165 3.185 42.845 3.445 ;
      RECT 42.285 4.865 42.605 5.125 ;
      RECT 40.805 4.865 41.125 5.125 ;
      RECT 40.325 3.185 40.645 3.445 ;
      RECT 39.605 4.305 39.925 4.565 ;
      RECT 38.885 4.305 39.205 4.565 ;
      RECT 35.445 4.305 35.765 4.565 ;
      RECT 24.205 4.865 24.525 5.125 ;
      RECT 23.605 3.185 24.285 3.445 ;
      RECT 23.725 4.865 24.045 5.125 ;
      RECT 22.245 4.865 22.565 5.125 ;
      RECT 21.765 3.185 22.085 3.445 ;
      RECT 21.045 4.305 21.365 4.565 ;
      RECT 20.325 4.305 20.645 4.565 ;
      RECT 16.885 4.305 17.205 4.565 ;
    LAYER mcon ;
      RECT 107.18 8.605 107.35 8.775 ;
      RECT 107.18 10.085 107.35 10.255 ;
      RECT 106.83 5.46 107 5.63 ;
      RECT 106.83 6.835 107 7.005 ;
      RECT 106.81 4.06 106.98 4.23 ;
      RECT 106.81 8.235 106.98 8.405 ;
      RECT 106.19 2.21 106.36 2.38 ;
      RECT 106.19 3.69 106.36 3.86 ;
      RECT 106.19 8.605 106.36 8.775 ;
      RECT 106.19 10.085 106.36 10.255 ;
      RECT 105.84 5.46 106.01 5.63 ;
      RECT 105.84 6.835 106.01 7.005 ;
      RECT 105.82 4.06 105.99 4.23 ;
      RECT 105.82 8.235 105.99 8.405 ;
      RECT 105.14 5.46 105.31 5.63 ;
      RECT 105.14 6.835 105.31 7.005 ;
      RECT 104.83 3.32 105 3.49 ;
      RECT 104.83 8.975 105 9.145 ;
      RECT 104.4 2.21 104.57 2.38 ;
      RECT 104.4 2.95 104.57 3.12 ;
      RECT 104.4 9.345 104.57 9.515 ;
      RECT 104.4 10.085 104.57 10.255 ;
      RECT 104.025 3.69 104.195 3.86 ;
      RECT 104.025 8.605 104.195 8.775 ;
      RECT 101.555 5.43 101.725 5.6 ;
      RECT 101.095 5.43 101.265 5.6 ;
      RECT 100.72 4.07 100.89 4.24 ;
      RECT 100.635 5.43 100.805 5.6 ;
      RECT 100.48 3.23 100.65 3.4 ;
      RECT 100.24 4.35 100.41 4.52 ;
      RECT 100.175 5.43 100.345 5.6 ;
      RECT 99.76 3.79 99.93 3.96 ;
      RECT 99.715 5.43 99.885 5.6 ;
      RECT 99.525 6.835 99.695 7.005 ;
      RECT 99.52 3.23 99.69 3.4 ;
      RECT 99.52 4.35 99.69 4.52 ;
      RECT 99.52 4.91 99.69 5.08 ;
      RECT 99.255 5.43 99.425 5.6 ;
      RECT 99.215 8.975 99.385 9.145 ;
      RECT 99.04 4.35 99.21 4.52 ;
      RECT 98.795 5.43 98.965 5.6 ;
      RECT 98.785 9.345 98.955 9.515 ;
      RECT 98.785 10.085 98.955 10.255 ;
      RECT 98.52 4.07 98.69 4.24 ;
      RECT 98.52 4.91 98.69 5.08 ;
      RECT 98.335 5.43 98.505 5.6 ;
      RECT 98.04 3.23 98.21 3.4 ;
      RECT 98.04 4.91 98.21 5.08 ;
      RECT 97.875 5.43 98.045 5.6 ;
      RECT 97.415 5.43 97.585 5.6 ;
      RECT 97.08 3.23 97.25 3.4 ;
      RECT 97.08 3.79 97.25 3.96 ;
      RECT 97.08 4.35 97.25 4.52 ;
      RECT 97.08 4.91 97.25 5.08 ;
      RECT 96.955 5.43 97.125 5.6 ;
      RECT 96.56 4.91 96.73 5.08 ;
      RECT 96.495 5.43 96.665 5.6 ;
      RECT 96.08 3.23 96.25 3.4 ;
      RECT 96.035 5.43 96.205 5.6 ;
      RECT 95.84 3.79 96.01 3.96 ;
      RECT 95.575 5.43 95.745 5.6 ;
      RECT 95.36 3.79 95.53 3.96 ;
      RECT 95.36 4.35 95.53 4.52 ;
      RECT 95.12 3.23 95.29 3.4 ;
      RECT 95.115 5.43 95.285 5.6 ;
      RECT 94.655 5.43 94.825 5.6 ;
      RECT 94.64 4.35 94.81 4.52 ;
      RECT 94.195 5.43 94.365 5.6 ;
      RECT 94.12 3.79 94.29 3.96 ;
      RECT 94.12 4.63 94.29 4.8 ;
      RECT 93.735 5.43 93.905 5.6 ;
      RECT 93.64 3.23 93.81 3.4 ;
      RECT 93.64 4.35 93.81 4.52 ;
      RECT 93.275 5.43 93.445 5.6 ;
      RECT 93.16 4.63 93.33 4.8 ;
      RECT 92.92 4.07 93.09 4.24 ;
      RECT 92.815 5.43 92.985 5.6 ;
      RECT 92.355 5.43 92.525 5.6 ;
      RECT 92.115 3.79 92.285 3.96 ;
      RECT 91.895 5.43 92.065 5.6 ;
      RECT 91.435 5.43 91.605 5.6 ;
      RECT 91.2 3.23 91.37 3.4 ;
      RECT 91.2 4.35 91.37 4.52 ;
      RECT 90.975 5.43 91.145 5.6 ;
      RECT 90.96 3.79 91.13 3.96 ;
      RECT 90.515 5.43 90.685 5.6 ;
      RECT 90.24 3.23 90.41 3.4 ;
      RECT 90.24 4.77 90.41 4.94 ;
      RECT 90.055 5.43 90.225 5.6 ;
      RECT 88.62 8.605 88.79 8.775 ;
      RECT 88.62 10.085 88.79 10.255 ;
      RECT 88.27 5.46 88.44 5.63 ;
      RECT 88.27 6.835 88.44 7.005 ;
      RECT 88.25 4.06 88.42 4.23 ;
      RECT 88.25 8.235 88.42 8.405 ;
      RECT 87.63 2.21 87.8 2.38 ;
      RECT 87.63 3.69 87.8 3.86 ;
      RECT 87.63 8.605 87.8 8.775 ;
      RECT 87.63 10.085 87.8 10.255 ;
      RECT 87.28 5.46 87.45 5.63 ;
      RECT 87.28 6.835 87.45 7.005 ;
      RECT 87.26 4.06 87.43 4.23 ;
      RECT 87.26 8.235 87.43 8.405 ;
      RECT 86.58 5.46 86.75 5.63 ;
      RECT 86.58 6.835 86.75 7.005 ;
      RECT 86.27 3.32 86.44 3.49 ;
      RECT 86.27 8.975 86.44 9.145 ;
      RECT 85.84 2.21 86.01 2.38 ;
      RECT 85.84 2.95 86.01 3.12 ;
      RECT 85.84 9.345 86.01 9.515 ;
      RECT 85.84 10.085 86.01 10.255 ;
      RECT 85.465 3.69 85.635 3.86 ;
      RECT 85.465 8.605 85.635 8.775 ;
      RECT 82.995 5.43 83.165 5.6 ;
      RECT 82.535 5.43 82.705 5.6 ;
      RECT 82.16 4.07 82.33 4.24 ;
      RECT 82.075 5.43 82.245 5.6 ;
      RECT 81.92 3.23 82.09 3.4 ;
      RECT 81.68 4.35 81.85 4.52 ;
      RECT 81.615 5.43 81.785 5.6 ;
      RECT 81.2 3.79 81.37 3.96 ;
      RECT 81.155 5.43 81.325 5.6 ;
      RECT 80.965 6.835 81.135 7.005 ;
      RECT 80.96 3.23 81.13 3.4 ;
      RECT 80.96 4.35 81.13 4.52 ;
      RECT 80.96 4.91 81.13 5.08 ;
      RECT 80.695 5.43 80.865 5.6 ;
      RECT 80.655 8.975 80.825 9.145 ;
      RECT 80.48 4.35 80.65 4.52 ;
      RECT 80.235 5.43 80.405 5.6 ;
      RECT 80.225 9.345 80.395 9.515 ;
      RECT 80.225 10.085 80.395 10.255 ;
      RECT 79.96 4.07 80.13 4.24 ;
      RECT 79.96 4.91 80.13 5.08 ;
      RECT 79.775 5.43 79.945 5.6 ;
      RECT 79.48 3.23 79.65 3.4 ;
      RECT 79.48 4.91 79.65 5.08 ;
      RECT 79.315 5.43 79.485 5.6 ;
      RECT 78.855 5.43 79.025 5.6 ;
      RECT 78.52 3.23 78.69 3.4 ;
      RECT 78.52 3.79 78.69 3.96 ;
      RECT 78.52 4.35 78.69 4.52 ;
      RECT 78.52 4.91 78.69 5.08 ;
      RECT 78.395 5.43 78.565 5.6 ;
      RECT 78 4.91 78.17 5.08 ;
      RECT 77.935 5.43 78.105 5.6 ;
      RECT 77.52 3.23 77.69 3.4 ;
      RECT 77.475 5.43 77.645 5.6 ;
      RECT 77.28 3.79 77.45 3.96 ;
      RECT 77.015 5.43 77.185 5.6 ;
      RECT 76.8 3.79 76.97 3.96 ;
      RECT 76.8 4.35 76.97 4.52 ;
      RECT 76.56 3.23 76.73 3.4 ;
      RECT 76.555 5.43 76.725 5.6 ;
      RECT 76.095 5.43 76.265 5.6 ;
      RECT 76.08 4.35 76.25 4.52 ;
      RECT 75.635 5.43 75.805 5.6 ;
      RECT 75.56 3.79 75.73 3.96 ;
      RECT 75.56 4.63 75.73 4.8 ;
      RECT 75.175 5.43 75.345 5.6 ;
      RECT 75.08 3.23 75.25 3.4 ;
      RECT 75.08 4.35 75.25 4.52 ;
      RECT 74.715 5.43 74.885 5.6 ;
      RECT 74.6 4.63 74.77 4.8 ;
      RECT 74.36 4.07 74.53 4.24 ;
      RECT 74.255 5.43 74.425 5.6 ;
      RECT 73.795 5.43 73.965 5.6 ;
      RECT 73.555 3.79 73.725 3.96 ;
      RECT 73.335 5.43 73.505 5.6 ;
      RECT 72.875 5.43 73.045 5.6 ;
      RECT 72.64 3.23 72.81 3.4 ;
      RECT 72.64 4.35 72.81 4.52 ;
      RECT 72.415 5.43 72.585 5.6 ;
      RECT 72.4 3.79 72.57 3.96 ;
      RECT 71.955 5.43 72.125 5.6 ;
      RECT 71.68 3.23 71.85 3.4 ;
      RECT 71.68 4.77 71.85 4.94 ;
      RECT 71.495 5.43 71.665 5.6 ;
      RECT 70.06 8.605 70.23 8.775 ;
      RECT 70.06 10.085 70.23 10.255 ;
      RECT 69.71 5.46 69.88 5.63 ;
      RECT 69.71 6.835 69.88 7.005 ;
      RECT 69.69 4.06 69.86 4.23 ;
      RECT 69.69 8.235 69.86 8.405 ;
      RECT 69.07 2.21 69.24 2.38 ;
      RECT 69.07 3.69 69.24 3.86 ;
      RECT 69.07 8.605 69.24 8.775 ;
      RECT 69.07 10.085 69.24 10.255 ;
      RECT 68.72 5.46 68.89 5.63 ;
      RECT 68.72 6.835 68.89 7.005 ;
      RECT 68.7 4.06 68.87 4.23 ;
      RECT 68.7 8.235 68.87 8.405 ;
      RECT 68.02 5.46 68.19 5.63 ;
      RECT 68.02 6.835 68.19 7.005 ;
      RECT 67.71 3.32 67.88 3.49 ;
      RECT 67.71 8.975 67.88 9.145 ;
      RECT 67.28 2.21 67.45 2.38 ;
      RECT 67.28 2.95 67.45 3.12 ;
      RECT 67.28 9.345 67.45 9.515 ;
      RECT 67.28 10.085 67.45 10.255 ;
      RECT 66.905 3.69 67.075 3.86 ;
      RECT 66.905 8.605 67.075 8.775 ;
      RECT 64.435 5.43 64.605 5.6 ;
      RECT 63.975 5.43 64.145 5.6 ;
      RECT 63.6 4.07 63.77 4.24 ;
      RECT 63.515 5.43 63.685 5.6 ;
      RECT 63.36 3.23 63.53 3.4 ;
      RECT 63.12 4.35 63.29 4.52 ;
      RECT 63.055 5.43 63.225 5.6 ;
      RECT 62.64 3.79 62.81 3.96 ;
      RECT 62.595 5.43 62.765 5.6 ;
      RECT 62.405 6.835 62.575 7.005 ;
      RECT 62.4 3.23 62.57 3.4 ;
      RECT 62.4 4.35 62.57 4.52 ;
      RECT 62.4 4.91 62.57 5.08 ;
      RECT 62.135 5.43 62.305 5.6 ;
      RECT 62.095 8.975 62.265 9.145 ;
      RECT 61.92 4.35 62.09 4.52 ;
      RECT 61.675 5.43 61.845 5.6 ;
      RECT 61.665 9.345 61.835 9.515 ;
      RECT 61.665 10.085 61.835 10.255 ;
      RECT 61.4 4.07 61.57 4.24 ;
      RECT 61.4 4.91 61.57 5.08 ;
      RECT 61.215 5.43 61.385 5.6 ;
      RECT 60.92 3.23 61.09 3.4 ;
      RECT 60.92 4.91 61.09 5.08 ;
      RECT 60.755 5.43 60.925 5.6 ;
      RECT 60.295 5.43 60.465 5.6 ;
      RECT 59.96 3.23 60.13 3.4 ;
      RECT 59.96 3.79 60.13 3.96 ;
      RECT 59.96 4.35 60.13 4.52 ;
      RECT 59.96 4.91 60.13 5.08 ;
      RECT 59.835 5.43 60.005 5.6 ;
      RECT 59.44 4.91 59.61 5.08 ;
      RECT 59.375 5.43 59.545 5.6 ;
      RECT 58.96 3.23 59.13 3.4 ;
      RECT 58.915 5.43 59.085 5.6 ;
      RECT 58.72 3.79 58.89 3.96 ;
      RECT 58.455 5.43 58.625 5.6 ;
      RECT 58.24 3.79 58.41 3.96 ;
      RECT 58.24 4.35 58.41 4.52 ;
      RECT 58 3.23 58.17 3.4 ;
      RECT 57.995 5.43 58.165 5.6 ;
      RECT 57.535 5.43 57.705 5.6 ;
      RECT 57.52 4.35 57.69 4.52 ;
      RECT 57.075 5.43 57.245 5.6 ;
      RECT 57 3.79 57.17 3.96 ;
      RECT 57 4.63 57.17 4.8 ;
      RECT 56.615 5.43 56.785 5.6 ;
      RECT 56.52 3.23 56.69 3.4 ;
      RECT 56.52 4.35 56.69 4.52 ;
      RECT 56.155 5.43 56.325 5.6 ;
      RECT 56.04 4.63 56.21 4.8 ;
      RECT 55.8 4.07 55.97 4.24 ;
      RECT 55.695 5.43 55.865 5.6 ;
      RECT 55.235 5.43 55.405 5.6 ;
      RECT 54.995 3.79 55.165 3.96 ;
      RECT 54.775 5.43 54.945 5.6 ;
      RECT 54.315 5.43 54.485 5.6 ;
      RECT 54.08 3.23 54.25 3.4 ;
      RECT 54.08 4.35 54.25 4.52 ;
      RECT 53.855 5.43 54.025 5.6 ;
      RECT 53.84 3.79 54.01 3.96 ;
      RECT 53.395 5.43 53.565 5.6 ;
      RECT 53.12 3.23 53.29 3.4 ;
      RECT 53.12 4.77 53.29 4.94 ;
      RECT 52.935 5.43 53.105 5.6 ;
      RECT 51.5 8.605 51.67 8.775 ;
      RECT 51.5 10.085 51.67 10.255 ;
      RECT 51.15 5.46 51.32 5.63 ;
      RECT 51.15 6.835 51.32 7.005 ;
      RECT 51.13 4.06 51.3 4.23 ;
      RECT 51.13 8.235 51.3 8.405 ;
      RECT 50.51 2.21 50.68 2.38 ;
      RECT 50.51 3.69 50.68 3.86 ;
      RECT 50.51 8.605 50.68 8.775 ;
      RECT 50.51 10.085 50.68 10.255 ;
      RECT 50.16 5.46 50.33 5.63 ;
      RECT 50.16 6.835 50.33 7.005 ;
      RECT 50.14 4.06 50.31 4.23 ;
      RECT 50.14 8.235 50.31 8.405 ;
      RECT 49.46 5.46 49.63 5.63 ;
      RECT 49.46 6.835 49.63 7.005 ;
      RECT 49.15 3.32 49.32 3.49 ;
      RECT 49.15 8.975 49.32 9.145 ;
      RECT 48.72 2.21 48.89 2.38 ;
      RECT 48.72 2.95 48.89 3.12 ;
      RECT 48.72 9.345 48.89 9.515 ;
      RECT 48.72 10.085 48.89 10.255 ;
      RECT 48.345 3.69 48.515 3.86 ;
      RECT 48.345 8.605 48.515 8.775 ;
      RECT 45.875 5.43 46.045 5.6 ;
      RECT 45.415 5.43 45.585 5.6 ;
      RECT 45.04 4.07 45.21 4.24 ;
      RECT 44.955 5.43 45.125 5.6 ;
      RECT 44.8 3.23 44.97 3.4 ;
      RECT 44.56 4.35 44.73 4.52 ;
      RECT 44.495 5.43 44.665 5.6 ;
      RECT 44.08 3.79 44.25 3.96 ;
      RECT 44.035 5.43 44.205 5.6 ;
      RECT 43.845 6.835 44.015 7.005 ;
      RECT 43.84 3.23 44.01 3.4 ;
      RECT 43.84 4.35 44.01 4.52 ;
      RECT 43.84 4.91 44.01 5.08 ;
      RECT 43.575 5.43 43.745 5.6 ;
      RECT 43.535 8.975 43.705 9.145 ;
      RECT 43.36 4.35 43.53 4.52 ;
      RECT 43.115 5.43 43.285 5.6 ;
      RECT 43.105 9.345 43.275 9.515 ;
      RECT 43.105 10.085 43.275 10.255 ;
      RECT 42.84 4.07 43.01 4.24 ;
      RECT 42.84 4.91 43.01 5.08 ;
      RECT 42.655 5.43 42.825 5.6 ;
      RECT 42.36 3.23 42.53 3.4 ;
      RECT 42.36 4.91 42.53 5.08 ;
      RECT 42.195 5.43 42.365 5.6 ;
      RECT 41.735 5.43 41.905 5.6 ;
      RECT 41.4 3.23 41.57 3.4 ;
      RECT 41.4 3.79 41.57 3.96 ;
      RECT 41.4 4.35 41.57 4.52 ;
      RECT 41.4 4.91 41.57 5.08 ;
      RECT 41.275 5.43 41.445 5.6 ;
      RECT 40.88 4.91 41.05 5.08 ;
      RECT 40.815 5.43 40.985 5.6 ;
      RECT 40.4 3.23 40.57 3.4 ;
      RECT 40.355 5.43 40.525 5.6 ;
      RECT 40.16 3.79 40.33 3.96 ;
      RECT 39.895 5.43 40.065 5.6 ;
      RECT 39.68 3.79 39.85 3.96 ;
      RECT 39.68 4.35 39.85 4.52 ;
      RECT 39.44 3.23 39.61 3.4 ;
      RECT 39.435 5.43 39.605 5.6 ;
      RECT 38.975 5.43 39.145 5.6 ;
      RECT 38.96 4.35 39.13 4.52 ;
      RECT 38.515 5.43 38.685 5.6 ;
      RECT 38.44 3.79 38.61 3.96 ;
      RECT 38.44 4.63 38.61 4.8 ;
      RECT 38.055 5.43 38.225 5.6 ;
      RECT 37.96 3.23 38.13 3.4 ;
      RECT 37.96 4.35 38.13 4.52 ;
      RECT 37.595 5.43 37.765 5.6 ;
      RECT 37.48 4.63 37.65 4.8 ;
      RECT 37.24 4.07 37.41 4.24 ;
      RECT 37.135 5.43 37.305 5.6 ;
      RECT 36.675 5.43 36.845 5.6 ;
      RECT 36.435 3.79 36.605 3.96 ;
      RECT 36.215 5.43 36.385 5.6 ;
      RECT 35.755 5.43 35.925 5.6 ;
      RECT 35.52 3.23 35.69 3.4 ;
      RECT 35.52 4.35 35.69 4.52 ;
      RECT 35.295 5.43 35.465 5.6 ;
      RECT 35.28 3.79 35.45 3.96 ;
      RECT 34.835 5.43 35.005 5.6 ;
      RECT 34.56 3.23 34.73 3.4 ;
      RECT 34.56 4.77 34.73 4.94 ;
      RECT 34.375 5.43 34.545 5.6 ;
      RECT 32.94 8.605 33.11 8.775 ;
      RECT 32.94 10.085 33.11 10.255 ;
      RECT 32.59 5.46 32.76 5.63 ;
      RECT 32.59 6.835 32.76 7.005 ;
      RECT 32.57 4.06 32.74 4.23 ;
      RECT 32.57 8.235 32.74 8.405 ;
      RECT 31.95 2.21 32.12 2.38 ;
      RECT 31.95 3.69 32.12 3.86 ;
      RECT 31.95 8.605 32.12 8.775 ;
      RECT 31.95 10.085 32.12 10.255 ;
      RECT 31.6 5.46 31.77 5.63 ;
      RECT 31.6 6.835 31.77 7.005 ;
      RECT 31.58 4.06 31.75 4.23 ;
      RECT 31.58 8.235 31.75 8.405 ;
      RECT 30.9 5.46 31.07 5.63 ;
      RECT 30.9 6.835 31.07 7.005 ;
      RECT 30.59 3.32 30.76 3.49 ;
      RECT 30.59 8.975 30.76 9.145 ;
      RECT 30.16 2.21 30.33 2.38 ;
      RECT 30.16 2.95 30.33 3.12 ;
      RECT 30.16 9.345 30.33 9.515 ;
      RECT 30.16 10.085 30.33 10.255 ;
      RECT 29.785 3.69 29.955 3.86 ;
      RECT 29.785 8.605 29.955 8.775 ;
      RECT 27.315 5.43 27.485 5.6 ;
      RECT 26.855 5.43 27.025 5.6 ;
      RECT 26.48 4.07 26.65 4.24 ;
      RECT 26.395 5.43 26.565 5.6 ;
      RECT 26.24 3.23 26.41 3.4 ;
      RECT 26 4.35 26.17 4.52 ;
      RECT 25.935 5.43 26.105 5.6 ;
      RECT 25.52 3.79 25.69 3.96 ;
      RECT 25.475 5.43 25.645 5.6 ;
      RECT 25.285 6.835 25.455 7.005 ;
      RECT 25.28 3.23 25.45 3.4 ;
      RECT 25.28 4.35 25.45 4.52 ;
      RECT 25.28 4.91 25.45 5.08 ;
      RECT 25.015 5.43 25.185 5.6 ;
      RECT 24.975 8.975 25.145 9.145 ;
      RECT 24.8 4.35 24.97 4.52 ;
      RECT 24.555 5.43 24.725 5.6 ;
      RECT 24.545 9.345 24.715 9.515 ;
      RECT 24.545 10.085 24.715 10.255 ;
      RECT 24.28 4.07 24.45 4.24 ;
      RECT 24.28 4.91 24.45 5.08 ;
      RECT 24.095 5.43 24.265 5.6 ;
      RECT 23.8 3.23 23.97 3.4 ;
      RECT 23.8 4.91 23.97 5.08 ;
      RECT 23.635 5.43 23.805 5.6 ;
      RECT 23.175 5.43 23.345 5.6 ;
      RECT 22.84 3.23 23.01 3.4 ;
      RECT 22.84 3.79 23.01 3.96 ;
      RECT 22.84 4.35 23.01 4.52 ;
      RECT 22.84 4.91 23.01 5.08 ;
      RECT 22.715 5.43 22.885 5.6 ;
      RECT 22.32 4.91 22.49 5.08 ;
      RECT 22.255 5.43 22.425 5.6 ;
      RECT 21.84 3.23 22.01 3.4 ;
      RECT 21.795 5.43 21.965 5.6 ;
      RECT 21.6 3.79 21.77 3.96 ;
      RECT 21.335 5.43 21.505 5.6 ;
      RECT 21.12 3.79 21.29 3.96 ;
      RECT 21.12 4.35 21.29 4.52 ;
      RECT 20.88 3.23 21.05 3.4 ;
      RECT 20.875 5.43 21.045 5.6 ;
      RECT 20.415 5.43 20.585 5.6 ;
      RECT 20.4 4.35 20.57 4.52 ;
      RECT 19.955 5.43 20.125 5.6 ;
      RECT 19.88 3.79 20.05 3.96 ;
      RECT 19.88 4.63 20.05 4.8 ;
      RECT 19.495 5.43 19.665 5.6 ;
      RECT 19.4 3.23 19.57 3.4 ;
      RECT 19.4 4.35 19.57 4.52 ;
      RECT 19.035 5.43 19.205 5.6 ;
      RECT 18.92 4.63 19.09 4.8 ;
      RECT 18.68 4.07 18.85 4.24 ;
      RECT 18.575 5.43 18.745 5.6 ;
      RECT 18.115 5.43 18.285 5.6 ;
      RECT 17.875 3.79 18.045 3.96 ;
      RECT 17.655 5.43 17.825 5.6 ;
      RECT 17.195 5.43 17.365 5.6 ;
      RECT 16.96 3.23 17.13 3.4 ;
      RECT 16.96 4.35 17.13 4.52 ;
      RECT 16.735 5.43 16.905 5.6 ;
      RECT 16.72 3.79 16.89 3.96 ;
      RECT 16.275 5.43 16.445 5.6 ;
      RECT 16 3.23 16.17 3.4 ;
      RECT 16 4.77 16.17 4.94 ;
      RECT 15.815 5.43 15.985 5.6 ;
      RECT 14.47 6.835 14.64 7.005 ;
      RECT 14.16 8.975 14.33 9.145 ;
      RECT 13.73 9.345 13.9 9.515 ;
      RECT 13.73 10.085 13.9 10.255 ;
      RECT 13.355 8.605 13.525 8.775 ;
    LAYER li1 ;
      RECT 14.16 5.45 14.33 10.595 ;
      RECT 106.75 4.7 106.92 7.765 ;
      RECT 105.76 4.7 105.93 7.765 ;
      RECT 103.02 4.7 103.19 7.765 ;
      RECT 97.405 5.43 97.575 7.765 ;
      RECT 88.19 4.7 88.36 7.765 ;
      RECT 87.2 4.7 87.37 7.765 ;
      RECT 84.46 4.7 84.63 7.765 ;
      RECT 78.845 5.43 79.015 7.765 ;
      RECT 69.63 4.7 69.8 7.765 ;
      RECT 68.64 4.7 68.81 7.765 ;
      RECT 65.9 4.7 66.07 7.765 ;
      RECT 60.285 5.43 60.455 7.765 ;
      RECT 51.07 4.7 51.24 7.765 ;
      RECT 50.08 4.7 50.25 7.765 ;
      RECT 47.34 4.7 47.51 7.765 ;
      RECT 41.725 5.43 41.895 7.765 ;
      RECT 32.51 4.7 32.68 7.765 ;
      RECT 31.52 4.7 31.69 7.765 ;
      RECT 28.78 4.7 28.95 7.765 ;
      RECT 23.165 5.43 23.335 7.765 ;
      RECT 12.35 5.45 12.52 7.765 ;
      RECT 12.125 5.45 107.725 7.05 ;
      RECT 89.91 5.43 107.725 7.05 ;
      RECT 14.925 5.435 107.725 7.05 ;
      RECT 71.35 5.43 89.165 7.05 ;
      RECT 52.79 5.43 70.605 7.05 ;
      RECT 34.23 5.43 52.045 7.05 ;
      RECT 15.67 5.43 33.485 7.05 ;
      RECT 100 4.93 100.17 7.05 ;
      RECT 97.56 4.93 97.73 7.05 ;
      RECT 95.6 4.93 95.77 7.05 ;
      RECT 94.64 4.93 94.81 7.05 ;
      RECT 92.68 4.93 92.85 7.05 ;
      RECT 91.68 4.93 91.85 7.05 ;
      RECT 90.72 4.93 90.89 7.05 ;
      RECT 81.44 4.93 81.61 7.05 ;
      RECT 79 4.93 79.17 7.05 ;
      RECT 77.04 4.93 77.21 7.05 ;
      RECT 76.08 4.93 76.25 7.05 ;
      RECT 74.12 4.93 74.29 7.05 ;
      RECT 73.12 4.93 73.29 7.05 ;
      RECT 72.16 4.93 72.33 7.05 ;
      RECT 62.88 4.93 63.05 7.05 ;
      RECT 60.44 4.93 60.61 7.05 ;
      RECT 58.48 4.93 58.65 7.05 ;
      RECT 57.52 4.93 57.69 7.05 ;
      RECT 55.56 4.93 55.73 7.05 ;
      RECT 54.56 4.93 54.73 7.05 ;
      RECT 53.6 4.93 53.77 7.05 ;
      RECT 44.32 4.93 44.49 7.05 ;
      RECT 41.88 4.93 42.05 7.05 ;
      RECT 39.92 4.93 40.09 7.05 ;
      RECT 38.96 4.93 39.13 7.05 ;
      RECT 37 4.93 37.17 7.05 ;
      RECT 36 4.93 36.17 7.05 ;
      RECT 35.04 4.93 35.21 7.05 ;
      RECT 25.76 4.93 25.93 7.05 ;
      RECT 23.32 4.93 23.49 7.05 ;
      RECT 21.36 4.93 21.53 7.05 ;
      RECT 20.4 4.93 20.57 7.05 ;
      RECT 18.44 4.93 18.61 7.05 ;
      RECT 17.44 4.93 17.61 7.05 ;
      RECT 16.48 4.93 16.65 7.05 ;
      RECT 106.81 3.04 106.98 4.23 ;
      RECT 106.81 3.04 107.28 3.21 ;
      RECT 106.81 9.255 107.28 9.425 ;
      RECT 106.81 8.235 106.98 9.425 ;
      RECT 105.82 3.04 105.99 4.23 ;
      RECT 105.82 3.04 106.29 3.21 ;
      RECT 105.82 9.255 106.29 9.425 ;
      RECT 105.82 8.235 105.99 9.425 ;
      RECT 103.97 3.93 104.14 5.16 ;
      RECT 104.025 2.15 104.195 4.1 ;
      RECT 103.97 1.87 104.14 2.32 ;
      RECT 103.97 10.145 104.14 10.595 ;
      RECT 104.025 8.365 104.195 10.315 ;
      RECT 103.97 7.305 104.14 8.535 ;
      RECT 103.45 1.87 103.62 5.16 ;
      RECT 103.45 3.37 103.855 3.7 ;
      RECT 103.45 2.53 103.855 2.86 ;
      RECT 103.45 7.305 103.62 10.595 ;
      RECT 103.45 9.605 103.855 9.935 ;
      RECT 103.45 8.765 103.855 9.095 ;
      RECT 100.24 4.52 101.21 4.69 ;
      RECT 100.24 4.35 100.41 4.69 ;
      RECT 99.76 3.79 99.93 4.12 ;
      RECT 99.76 3.87 100.49 4.04 ;
      RECT 99.4 4.91 99.69 5.08 ;
      RECT 99.4 3.87 99.57 5.08 ;
      RECT 99.4 4.35 99.69 4.52 ;
      RECT 99.2 3.87 99.57 4.04 ;
      RECT 98.52 3.97 98.69 4.24 ;
      RECT 98.28 3.97 98.69 4.14 ;
      RECT 98.2 3.87 98.53 4.04 ;
      RECT 98.04 4.91 98.69 5.08 ;
      RECT 98.52 4.44 98.69 5.08 ;
      RECT 98.4 4.52 98.69 5.08 ;
      RECT 97.835 7.305 98.005 10.595 ;
      RECT 97.835 9.605 98.24 9.935 ;
      RECT 97.835 8.765 98.24 9.095 ;
      RECT 97.08 4.21 97.25 4.52 ;
      RECT 97.08 4.21 97.97 4.38 ;
      RECT 97.8 3.79 97.97 4.38 ;
      RECT 97.08 3.87 97.57 4.04 ;
      RECT 97.08 3.79 97.25 4.04 ;
      RECT 95.04 4.52 95.53 4.69 ;
      RECT 96.2 3.87 96.37 4.52 ;
      RECT 95.36 4.35 96.37 4.52 ;
      RECT 96.32 3.79 96.49 4.12 ;
      RECT 95.12 3.13 95.29 3.4 ;
      RECT 94.56 3.13 95.29 3.3 ;
      RECT 94.64 3.87 94.81 4.52 ;
      RECT 94.64 3.87 95.13 4.04 ;
      RECT 93.8 3.87 94.29 4.04 ;
      RECT 94.12 3.79 94.29 4.04 ;
      RECT 93.64 3.13 93.81 3.4 ;
      RECT 93.08 3.13 93.81 3.3 ;
      RECT 93.16 4.52 93.33 4.8 ;
      RECT 92.12 4.52 93.41 4.69 ;
      RECT 92.115 3.87 92.69 4.04 ;
      RECT 92.115 3.79 92.285 4.04 ;
      RECT 91.2 3.13 91.37 3.4 ;
      RECT 91.2 3.13 91.93 3.3 ;
      RECT 91.2 4.35 91.37 4.77 ;
      RECT 90.58 4.435 91.37 4.605 ;
      RECT 90.58 4.21 90.75 4.605 ;
      RECT 90.48 3.79 90.65 4.38 ;
      RECT 90.24 3.87 90.65 4.14 ;
      RECT 88.25 3.04 88.42 4.23 ;
      RECT 88.25 3.04 88.72 3.21 ;
      RECT 88.25 9.255 88.72 9.425 ;
      RECT 88.25 8.235 88.42 9.425 ;
      RECT 87.26 3.04 87.43 4.23 ;
      RECT 87.26 3.04 87.73 3.21 ;
      RECT 87.26 9.255 87.73 9.425 ;
      RECT 87.26 8.235 87.43 9.425 ;
      RECT 85.41 3.93 85.58 5.16 ;
      RECT 85.465 2.15 85.635 4.1 ;
      RECT 85.41 1.87 85.58 2.32 ;
      RECT 85.41 10.145 85.58 10.595 ;
      RECT 85.465 8.365 85.635 10.315 ;
      RECT 85.41 7.305 85.58 8.535 ;
      RECT 84.89 1.87 85.06 5.16 ;
      RECT 84.89 3.37 85.295 3.7 ;
      RECT 84.89 2.53 85.295 2.86 ;
      RECT 84.89 7.305 85.06 10.595 ;
      RECT 84.89 9.605 85.295 9.935 ;
      RECT 84.89 8.765 85.295 9.095 ;
      RECT 81.68 4.52 82.65 4.69 ;
      RECT 81.68 4.35 81.85 4.69 ;
      RECT 81.2 3.79 81.37 4.12 ;
      RECT 81.2 3.87 81.93 4.04 ;
      RECT 80.84 4.91 81.13 5.08 ;
      RECT 80.84 3.87 81.01 5.08 ;
      RECT 80.84 4.35 81.13 4.52 ;
      RECT 80.64 3.87 81.01 4.04 ;
      RECT 79.96 3.97 80.13 4.24 ;
      RECT 79.72 3.97 80.13 4.14 ;
      RECT 79.64 3.87 79.97 4.04 ;
      RECT 79.48 4.91 80.13 5.08 ;
      RECT 79.96 4.44 80.13 5.08 ;
      RECT 79.84 4.52 80.13 5.08 ;
      RECT 79.275 7.305 79.445 10.595 ;
      RECT 79.275 9.605 79.68 9.935 ;
      RECT 79.275 8.765 79.68 9.095 ;
      RECT 78.52 4.21 78.69 4.52 ;
      RECT 78.52 4.21 79.41 4.38 ;
      RECT 79.24 3.79 79.41 4.38 ;
      RECT 78.52 3.87 79.01 4.04 ;
      RECT 78.52 3.79 78.69 4.04 ;
      RECT 76.48 4.52 76.97 4.69 ;
      RECT 77.64 3.87 77.81 4.52 ;
      RECT 76.8 4.35 77.81 4.52 ;
      RECT 77.76 3.79 77.93 4.12 ;
      RECT 76.56 3.13 76.73 3.4 ;
      RECT 76 3.13 76.73 3.3 ;
      RECT 76.08 3.87 76.25 4.52 ;
      RECT 76.08 3.87 76.57 4.04 ;
      RECT 75.24 3.87 75.73 4.04 ;
      RECT 75.56 3.79 75.73 4.04 ;
      RECT 75.08 3.13 75.25 3.4 ;
      RECT 74.52 3.13 75.25 3.3 ;
      RECT 74.6 4.52 74.77 4.8 ;
      RECT 73.56 4.52 74.85 4.69 ;
      RECT 73.555 3.87 74.13 4.04 ;
      RECT 73.555 3.79 73.725 4.04 ;
      RECT 72.64 3.13 72.81 3.4 ;
      RECT 72.64 3.13 73.37 3.3 ;
      RECT 72.64 4.35 72.81 4.77 ;
      RECT 72.02 4.435 72.81 4.605 ;
      RECT 72.02 4.21 72.19 4.605 ;
      RECT 71.92 3.79 72.09 4.38 ;
      RECT 71.68 3.87 72.09 4.14 ;
      RECT 69.69 3.04 69.86 4.23 ;
      RECT 69.69 3.04 70.16 3.21 ;
      RECT 69.69 9.255 70.16 9.425 ;
      RECT 69.69 8.235 69.86 9.425 ;
      RECT 68.7 3.04 68.87 4.23 ;
      RECT 68.7 3.04 69.17 3.21 ;
      RECT 68.7 9.255 69.17 9.425 ;
      RECT 68.7 8.235 68.87 9.425 ;
      RECT 66.85 3.93 67.02 5.16 ;
      RECT 66.905 2.15 67.075 4.1 ;
      RECT 66.85 1.87 67.02 2.32 ;
      RECT 66.85 10.145 67.02 10.595 ;
      RECT 66.905 8.365 67.075 10.315 ;
      RECT 66.85 7.305 67.02 8.535 ;
      RECT 66.33 1.87 66.5 5.16 ;
      RECT 66.33 3.37 66.735 3.7 ;
      RECT 66.33 2.53 66.735 2.86 ;
      RECT 66.33 7.305 66.5 10.595 ;
      RECT 66.33 9.605 66.735 9.935 ;
      RECT 66.33 8.765 66.735 9.095 ;
      RECT 63.12 4.52 64.09 4.69 ;
      RECT 63.12 4.35 63.29 4.69 ;
      RECT 62.64 3.79 62.81 4.12 ;
      RECT 62.64 3.87 63.37 4.04 ;
      RECT 62.28 4.91 62.57 5.08 ;
      RECT 62.28 3.87 62.45 5.08 ;
      RECT 62.28 4.35 62.57 4.52 ;
      RECT 62.08 3.87 62.45 4.04 ;
      RECT 61.4 3.97 61.57 4.24 ;
      RECT 61.16 3.97 61.57 4.14 ;
      RECT 61.08 3.87 61.41 4.04 ;
      RECT 60.92 4.91 61.57 5.08 ;
      RECT 61.4 4.44 61.57 5.08 ;
      RECT 61.28 4.52 61.57 5.08 ;
      RECT 60.715 7.305 60.885 10.595 ;
      RECT 60.715 9.605 61.12 9.935 ;
      RECT 60.715 8.765 61.12 9.095 ;
      RECT 59.96 4.21 60.13 4.52 ;
      RECT 59.96 4.21 60.85 4.38 ;
      RECT 60.68 3.79 60.85 4.38 ;
      RECT 59.96 3.87 60.45 4.04 ;
      RECT 59.96 3.79 60.13 4.04 ;
      RECT 57.92 4.52 58.41 4.69 ;
      RECT 59.08 3.87 59.25 4.52 ;
      RECT 58.24 4.35 59.25 4.52 ;
      RECT 59.2 3.79 59.37 4.12 ;
      RECT 58 3.13 58.17 3.4 ;
      RECT 57.44 3.13 58.17 3.3 ;
      RECT 57.52 3.87 57.69 4.52 ;
      RECT 57.52 3.87 58.01 4.04 ;
      RECT 56.68 3.87 57.17 4.04 ;
      RECT 57 3.79 57.17 4.04 ;
      RECT 56.52 3.13 56.69 3.4 ;
      RECT 55.96 3.13 56.69 3.3 ;
      RECT 56.04 4.52 56.21 4.8 ;
      RECT 55 4.52 56.29 4.69 ;
      RECT 54.995 3.87 55.57 4.04 ;
      RECT 54.995 3.79 55.165 4.04 ;
      RECT 54.08 3.13 54.25 3.4 ;
      RECT 54.08 3.13 54.81 3.3 ;
      RECT 54.08 4.35 54.25 4.77 ;
      RECT 53.46 4.435 54.25 4.605 ;
      RECT 53.46 4.21 53.63 4.605 ;
      RECT 53.36 3.79 53.53 4.38 ;
      RECT 53.12 3.87 53.53 4.14 ;
      RECT 51.13 3.04 51.3 4.23 ;
      RECT 51.13 3.04 51.6 3.21 ;
      RECT 51.13 9.255 51.6 9.425 ;
      RECT 51.13 8.235 51.3 9.425 ;
      RECT 50.14 3.04 50.31 4.23 ;
      RECT 50.14 3.04 50.61 3.21 ;
      RECT 50.14 9.255 50.61 9.425 ;
      RECT 50.14 8.235 50.31 9.425 ;
      RECT 48.29 3.93 48.46 5.16 ;
      RECT 48.345 2.15 48.515 4.1 ;
      RECT 48.29 1.87 48.46 2.32 ;
      RECT 48.29 10.145 48.46 10.595 ;
      RECT 48.345 8.365 48.515 10.315 ;
      RECT 48.29 7.305 48.46 8.535 ;
      RECT 47.77 1.87 47.94 5.16 ;
      RECT 47.77 3.37 48.175 3.7 ;
      RECT 47.77 2.53 48.175 2.86 ;
      RECT 47.77 7.305 47.94 10.595 ;
      RECT 47.77 9.605 48.175 9.935 ;
      RECT 47.77 8.765 48.175 9.095 ;
      RECT 44.56 4.52 45.53 4.69 ;
      RECT 44.56 4.35 44.73 4.69 ;
      RECT 44.08 3.79 44.25 4.12 ;
      RECT 44.08 3.87 44.81 4.04 ;
      RECT 43.72 4.91 44.01 5.08 ;
      RECT 43.72 3.87 43.89 5.08 ;
      RECT 43.72 4.35 44.01 4.52 ;
      RECT 43.52 3.87 43.89 4.04 ;
      RECT 42.84 3.97 43.01 4.24 ;
      RECT 42.6 3.97 43.01 4.14 ;
      RECT 42.52 3.87 42.85 4.04 ;
      RECT 42.36 4.91 43.01 5.08 ;
      RECT 42.84 4.44 43.01 5.08 ;
      RECT 42.72 4.52 43.01 5.08 ;
      RECT 42.155 7.305 42.325 10.595 ;
      RECT 42.155 9.605 42.56 9.935 ;
      RECT 42.155 8.765 42.56 9.095 ;
      RECT 41.4 4.21 41.57 4.52 ;
      RECT 41.4 4.21 42.29 4.38 ;
      RECT 42.12 3.79 42.29 4.38 ;
      RECT 41.4 3.87 41.89 4.04 ;
      RECT 41.4 3.79 41.57 4.04 ;
      RECT 39.36 4.52 39.85 4.69 ;
      RECT 40.52 3.87 40.69 4.52 ;
      RECT 39.68 4.35 40.69 4.52 ;
      RECT 40.64 3.79 40.81 4.12 ;
      RECT 39.44 3.13 39.61 3.4 ;
      RECT 38.88 3.13 39.61 3.3 ;
      RECT 38.96 3.87 39.13 4.52 ;
      RECT 38.96 3.87 39.45 4.04 ;
      RECT 38.12 3.87 38.61 4.04 ;
      RECT 38.44 3.79 38.61 4.04 ;
      RECT 37.96 3.13 38.13 3.4 ;
      RECT 37.4 3.13 38.13 3.3 ;
      RECT 37.48 4.52 37.65 4.8 ;
      RECT 36.44 4.52 37.73 4.69 ;
      RECT 36.435 3.87 37.01 4.04 ;
      RECT 36.435 3.79 36.605 4.04 ;
      RECT 35.52 3.13 35.69 3.4 ;
      RECT 35.52 3.13 36.25 3.3 ;
      RECT 35.52 4.35 35.69 4.77 ;
      RECT 34.9 4.435 35.69 4.605 ;
      RECT 34.9 4.21 35.07 4.605 ;
      RECT 34.8 3.79 34.97 4.38 ;
      RECT 34.56 3.87 34.97 4.14 ;
      RECT 32.57 3.04 32.74 4.23 ;
      RECT 32.57 3.04 33.04 3.21 ;
      RECT 32.57 9.255 33.04 9.425 ;
      RECT 32.57 8.235 32.74 9.425 ;
      RECT 31.58 3.04 31.75 4.23 ;
      RECT 31.58 3.04 32.05 3.21 ;
      RECT 31.58 9.255 32.05 9.425 ;
      RECT 31.58 8.235 31.75 9.425 ;
      RECT 29.73 3.93 29.9 5.16 ;
      RECT 29.785 2.15 29.955 4.1 ;
      RECT 29.73 1.87 29.9 2.32 ;
      RECT 29.73 10.145 29.9 10.595 ;
      RECT 29.785 8.365 29.955 10.315 ;
      RECT 29.73 7.305 29.9 8.535 ;
      RECT 29.21 1.87 29.38 5.16 ;
      RECT 29.21 3.37 29.615 3.7 ;
      RECT 29.21 2.53 29.615 2.86 ;
      RECT 29.21 7.305 29.38 10.595 ;
      RECT 29.21 9.605 29.615 9.935 ;
      RECT 29.21 8.765 29.615 9.095 ;
      RECT 26 4.52 26.97 4.69 ;
      RECT 26 4.35 26.17 4.69 ;
      RECT 25.52 3.79 25.69 4.12 ;
      RECT 25.52 3.87 26.25 4.04 ;
      RECT 25.16 4.91 25.45 5.08 ;
      RECT 25.16 3.87 25.33 5.08 ;
      RECT 25.16 4.35 25.45 4.52 ;
      RECT 24.96 3.87 25.33 4.04 ;
      RECT 24.28 3.97 24.45 4.24 ;
      RECT 24.04 3.97 24.45 4.14 ;
      RECT 23.96 3.87 24.29 4.04 ;
      RECT 23.8 4.91 24.45 5.08 ;
      RECT 24.28 4.44 24.45 5.08 ;
      RECT 24.16 4.52 24.45 5.08 ;
      RECT 23.595 7.305 23.765 10.595 ;
      RECT 23.595 9.605 24 9.935 ;
      RECT 23.595 8.765 24 9.095 ;
      RECT 22.84 4.21 23.01 4.52 ;
      RECT 22.84 4.21 23.73 4.38 ;
      RECT 23.56 3.79 23.73 4.38 ;
      RECT 22.84 3.87 23.33 4.04 ;
      RECT 22.84 3.79 23.01 4.04 ;
      RECT 20.8 4.52 21.29 4.69 ;
      RECT 21.96 3.87 22.13 4.52 ;
      RECT 21.12 4.35 22.13 4.52 ;
      RECT 22.08 3.79 22.25 4.12 ;
      RECT 20.88 3.13 21.05 3.4 ;
      RECT 20.32 3.13 21.05 3.3 ;
      RECT 20.4 3.87 20.57 4.52 ;
      RECT 20.4 3.87 20.89 4.04 ;
      RECT 19.56 3.87 20.05 4.04 ;
      RECT 19.88 3.79 20.05 4.04 ;
      RECT 19.4 3.13 19.57 3.4 ;
      RECT 18.84 3.13 19.57 3.3 ;
      RECT 18.92 4.52 19.09 4.8 ;
      RECT 17.88 4.52 19.17 4.69 ;
      RECT 17.875 3.87 18.45 4.04 ;
      RECT 17.875 3.79 18.045 4.04 ;
      RECT 16.96 3.13 17.13 3.4 ;
      RECT 16.96 3.13 17.69 3.3 ;
      RECT 16.96 4.35 17.13 4.77 ;
      RECT 16.34 4.435 17.13 4.605 ;
      RECT 16.34 4.21 16.51 4.605 ;
      RECT 16.24 3.79 16.41 4.38 ;
      RECT 16 3.87 16.41 4.14 ;
      RECT 13.3 10.145 13.47 10.595 ;
      RECT 13.355 8.365 13.525 10.315 ;
      RECT 13.3 7.305 13.47 8.535 ;
      RECT 12.78 7.305 12.95 10.595 ;
      RECT 12.78 9.605 13.185 9.935 ;
      RECT 12.78 8.765 13.185 9.095 ;
      RECT 107.18 7.305 107.35 8.775 ;
      RECT 107.18 10.085 107.35 10.595 ;
      RECT 106.19 1.87 106.36 2.38 ;
      RECT 106.19 3.69 106.36 5.16 ;
      RECT 106.19 7.305 106.36 8.775 ;
      RECT 106.19 10.085 106.36 10.595 ;
      RECT 104.83 1.87 105 5.16 ;
      RECT 104.83 7.305 105 10.595 ;
      RECT 104.4 1.87 104.57 2.38 ;
      RECT 104.4 2.95 104.57 5.16 ;
      RECT 104.4 7.305 104.57 9.515 ;
      RECT 104.4 10.085 104.57 10.595 ;
      RECT 100.72 3.79 100.89 4.24 ;
      RECT 100.48 3.05 100.65 3.4 ;
      RECT 99.52 3.05 99.69 3.4 ;
      RECT 99.215 7.305 99.385 10.595 ;
      RECT 99.04 4.35 99.21 4.77 ;
      RECT 98.785 7.305 98.955 9.515 ;
      RECT 98.785 10.085 98.955 10.595 ;
      RECT 98.04 3.05 98.21 3.4 ;
      RECT 97.08 3.05 97.25 3.4 ;
      RECT 97.08 4.78 97.25 5.11 ;
      RECT 96.56 4.44 96.73 5.08 ;
      RECT 96.08 3.05 96.25 3.4 ;
      RECT 95.84 3.79 96.01 4.12 ;
      RECT 95.36 3.79 95.53 4.12 ;
      RECT 94.12 4.44 94.29 4.8 ;
      RECT 93.64 4.35 93.81 4.77 ;
      RECT 92.92 3.79 93.09 4.24 ;
      RECT 90.96 3.79 91.13 4.12 ;
      RECT 90.24 3.05 90.41 3.4 ;
      RECT 90.24 4.58 90.41 4.94 ;
      RECT 88.62 7.305 88.79 8.775 ;
      RECT 88.62 10.085 88.79 10.595 ;
      RECT 87.63 1.87 87.8 2.38 ;
      RECT 87.63 3.69 87.8 5.16 ;
      RECT 87.63 7.305 87.8 8.775 ;
      RECT 87.63 10.085 87.8 10.595 ;
      RECT 86.27 1.87 86.44 5.16 ;
      RECT 86.27 7.305 86.44 10.595 ;
      RECT 85.84 1.87 86.01 2.38 ;
      RECT 85.84 2.95 86.01 5.16 ;
      RECT 85.84 7.305 86.01 9.515 ;
      RECT 85.84 10.085 86.01 10.595 ;
      RECT 82.16 3.79 82.33 4.24 ;
      RECT 81.92 3.05 82.09 3.4 ;
      RECT 80.96 3.05 81.13 3.4 ;
      RECT 80.655 7.305 80.825 10.595 ;
      RECT 80.48 4.35 80.65 4.77 ;
      RECT 80.225 7.305 80.395 9.515 ;
      RECT 80.225 10.085 80.395 10.595 ;
      RECT 79.48 3.05 79.65 3.4 ;
      RECT 78.52 3.05 78.69 3.4 ;
      RECT 78.52 4.78 78.69 5.11 ;
      RECT 78 4.44 78.17 5.08 ;
      RECT 77.52 3.05 77.69 3.4 ;
      RECT 77.28 3.79 77.45 4.12 ;
      RECT 76.8 3.79 76.97 4.12 ;
      RECT 75.56 4.44 75.73 4.8 ;
      RECT 75.08 4.35 75.25 4.77 ;
      RECT 74.36 3.79 74.53 4.24 ;
      RECT 72.4 3.79 72.57 4.12 ;
      RECT 71.68 3.05 71.85 3.4 ;
      RECT 71.68 4.58 71.85 4.94 ;
      RECT 70.06 7.305 70.23 8.775 ;
      RECT 70.06 10.085 70.23 10.595 ;
      RECT 69.07 1.87 69.24 2.38 ;
      RECT 69.07 3.69 69.24 5.16 ;
      RECT 69.07 7.305 69.24 8.775 ;
      RECT 69.07 10.085 69.24 10.595 ;
      RECT 67.71 1.87 67.88 5.16 ;
      RECT 67.71 7.305 67.88 10.595 ;
      RECT 67.28 1.87 67.45 2.38 ;
      RECT 67.28 2.95 67.45 5.16 ;
      RECT 67.28 7.305 67.45 9.515 ;
      RECT 67.28 10.085 67.45 10.595 ;
      RECT 63.6 3.79 63.77 4.24 ;
      RECT 63.36 3.05 63.53 3.4 ;
      RECT 62.4 3.05 62.57 3.4 ;
      RECT 62.095 7.305 62.265 10.595 ;
      RECT 61.92 4.35 62.09 4.77 ;
      RECT 61.665 7.305 61.835 9.515 ;
      RECT 61.665 10.085 61.835 10.595 ;
      RECT 60.92 3.05 61.09 3.4 ;
      RECT 59.96 3.05 60.13 3.4 ;
      RECT 59.96 4.78 60.13 5.11 ;
      RECT 59.44 4.44 59.61 5.08 ;
      RECT 58.96 3.05 59.13 3.4 ;
      RECT 58.72 3.79 58.89 4.12 ;
      RECT 58.24 3.79 58.41 4.12 ;
      RECT 57 4.44 57.17 4.8 ;
      RECT 56.52 4.35 56.69 4.77 ;
      RECT 55.8 3.79 55.97 4.24 ;
      RECT 53.84 3.79 54.01 4.12 ;
      RECT 53.12 3.05 53.29 3.4 ;
      RECT 53.12 4.58 53.29 4.94 ;
      RECT 51.5 7.305 51.67 8.775 ;
      RECT 51.5 10.085 51.67 10.595 ;
      RECT 50.51 1.87 50.68 2.38 ;
      RECT 50.51 3.69 50.68 5.16 ;
      RECT 50.51 7.305 50.68 8.775 ;
      RECT 50.51 10.085 50.68 10.595 ;
      RECT 49.15 1.87 49.32 5.16 ;
      RECT 49.15 7.305 49.32 10.595 ;
      RECT 48.72 1.87 48.89 2.38 ;
      RECT 48.72 2.95 48.89 5.16 ;
      RECT 48.72 7.305 48.89 9.515 ;
      RECT 48.72 10.085 48.89 10.595 ;
      RECT 45.04 3.79 45.21 4.24 ;
      RECT 44.8 3.05 44.97 3.4 ;
      RECT 43.84 3.05 44.01 3.4 ;
      RECT 43.535 7.305 43.705 10.595 ;
      RECT 43.36 4.35 43.53 4.77 ;
      RECT 43.105 7.305 43.275 9.515 ;
      RECT 43.105 10.085 43.275 10.595 ;
      RECT 42.36 3.05 42.53 3.4 ;
      RECT 41.4 3.05 41.57 3.4 ;
      RECT 41.4 4.78 41.57 5.11 ;
      RECT 40.88 4.44 41.05 5.08 ;
      RECT 40.4 3.05 40.57 3.4 ;
      RECT 40.16 3.79 40.33 4.12 ;
      RECT 39.68 3.79 39.85 4.12 ;
      RECT 38.44 4.44 38.61 4.8 ;
      RECT 37.96 4.35 38.13 4.77 ;
      RECT 37.24 3.79 37.41 4.24 ;
      RECT 35.28 3.79 35.45 4.12 ;
      RECT 34.56 3.05 34.73 3.4 ;
      RECT 34.56 4.58 34.73 4.94 ;
      RECT 32.94 7.305 33.11 8.775 ;
      RECT 32.94 10.085 33.11 10.595 ;
      RECT 31.95 1.87 32.12 2.38 ;
      RECT 31.95 3.69 32.12 5.16 ;
      RECT 31.95 7.305 32.12 8.775 ;
      RECT 31.95 10.085 32.12 10.595 ;
      RECT 30.59 1.87 30.76 5.16 ;
      RECT 30.59 7.305 30.76 10.595 ;
      RECT 30.16 1.87 30.33 2.38 ;
      RECT 30.16 2.95 30.33 5.16 ;
      RECT 30.16 7.305 30.33 9.515 ;
      RECT 30.16 10.085 30.33 10.595 ;
      RECT 26.48 3.79 26.65 4.24 ;
      RECT 26.24 3.05 26.41 3.4 ;
      RECT 25.28 3.05 25.45 3.4 ;
      RECT 24.975 7.305 25.145 10.595 ;
      RECT 24.8 4.35 24.97 4.77 ;
      RECT 24.545 7.305 24.715 9.515 ;
      RECT 24.545 10.085 24.715 10.595 ;
      RECT 23.8 3.05 23.97 3.4 ;
      RECT 22.84 3.05 23.01 3.4 ;
      RECT 22.84 4.78 23.01 5.11 ;
      RECT 22.32 4.44 22.49 5.08 ;
      RECT 21.84 3.05 22.01 3.4 ;
      RECT 21.6 3.79 21.77 4.12 ;
      RECT 21.12 3.79 21.29 4.12 ;
      RECT 19.88 4.44 20.05 4.8 ;
      RECT 19.4 4.35 19.57 4.77 ;
      RECT 18.68 3.79 18.85 4.24 ;
      RECT 16.72 3.79 16.89 4.12 ;
      RECT 16 3.05 16.17 3.4 ;
      RECT 16 4.58 16.17 4.94 ;
      RECT 13.73 7.305 13.9 9.515 ;
      RECT 13.73 10.085 13.9 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  ORIGIN -12.13 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r2 ;
  SIZE 95.6 BY 12.475 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 32.945 2.21 33.115 2.38 ;
        RECT 32.94 2.205 33.11 2.375 ;
        RECT 32.94 3.685 33.11 3.855 ;
      LAYER li1 ;
        RECT 32.945 2.21 33.115 2.38 ;
        RECT 32.94 1.865 33.11 2.375 ;
        RECT 32.94 3.685 33.11 5.155 ;
      LAYER met1 ;
        RECT 32.88 3.655 33.17 3.885 ;
        RECT 32.88 2.175 33.17 2.405 ;
        RECT 32.94 2.175 33.11 3.885 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 51.505 2.21 51.675 2.38 ;
        RECT 51.5 2.205 51.67 2.375 ;
        RECT 51.5 3.685 51.67 3.855 ;
      LAYER li1 ;
        RECT 51.505 2.21 51.675 2.38 ;
        RECT 51.5 1.865 51.67 2.375 ;
        RECT 51.5 3.685 51.67 5.155 ;
      LAYER met1 ;
        RECT 51.44 3.655 51.73 3.885 ;
        RECT 51.44 2.175 51.73 2.405 ;
        RECT 51.5 2.175 51.67 3.885 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 70.065 2.21 70.235 2.38 ;
        RECT 70.06 2.205 70.23 2.375 ;
        RECT 70.06 3.685 70.23 3.855 ;
      LAYER li1 ;
        RECT 70.065 2.21 70.235 2.38 ;
        RECT 70.06 1.865 70.23 2.375 ;
        RECT 70.06 3.685 70.23 5.155 ;
      LAYER met1 ;
        RECT 70 3.655 70.29 3.885 ;
        RECT 70 2.175 70.29 2.405 ;
        RECT 70.06 2.175 70.23 3.885 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 88.625 2.21 88.795 2.38 ;
        RECT 88.62 2.205 88.79 2.375 ;
        RECT 88.62 3.685 88.79 3.855 ;
      LAYER li1 ;
        RECT 88.625 2.21 88.795 2.38 ;
        RECT 88.62 1.865 88.79 2.375 ;
        RECT 88.62 3.685 88.79 5.155 ;
      LAYER met1 ;
        RECT 88.56 3.655 88.85 3.885 ;
        RECT 88.56 2.175 88.85 2.405 ;
        RECT 88.62 2.175 88.79 3.885 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER mcon ;
        RECT 107.185 2.21 107.355 2.38 ;
        RECT 107.18 2.205 107.35 2.375 ;
        RECT 107.18 3.685 107.35 3.855 ;
      LAYER li1 ;
        RECT 107.185 2.21 107.355 2.38 ;
        RECT 107.18 1.865 107.35 2.375 ;
        RECT 107.18 3.685 107.35 5.155 ;
      LAYER met1 ;
        RECT 107.12 3.655 107.41 3.885 ;
        RECT 107.12 2.175 107.41 2.405 ;
        RECT 107.18 2.175 107.35 3.885 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 28.79 2.955 28.96 4.23 ;
        RECT 28.79 8.235 28.96 9.51 ;
        RECT 23.175 8.235 23.345 9.51 ;
      LAYER met2 ;
        RECT 28.715 4 29.055 4.35 ;
        RECT 28.705 8.135 29.045 8.485 ;
        RECT 28.79 4 28.96 8.485 ;
      LAYER met1 ;
        RECT 28.715 4.06 29.19 4.23 ;
        RECT 28.715 4 29.055 4.35 ;
        RECT 23.115 8.235 29.19 8.405 ;
        RECT 28.705 8.135 29.045 8.485 ;
        RECT 23.115 8.205 23.405 8.435 ;
      LAYER via1 ;
        RECT 28.805 8.235 28.955 8.385 ;
        RECT 28.815 4.1 28.965 4.25 ;
      LAYER mcon ;
        RECT 23.175 8.235 23.345 8.405 ;
        RECT 28.79 8.235 28.96 8.405 ;
        RECT 28.79 4.06 28.96 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 47.35 2.955 47.52 4.23 ;
        RECT 47.35 8.235 47.52 9.51 ;
        RECT 41.735 8.235 41.905 9.51 ;
      LAYER met2 ;
        RECT 47.275 4 47.615 4.35 ;
        RECT 47.265 8.135 47.605 8.485 ;
        RECT 47.35 4 47.52 8.485 ;
      LAYER met1 ;
        RECT 47.275 4.06 47.75 4.23 ;
        RECT 47.275 4 47.615 4.35 ;
        RECT 41.675 8.235 47.75 8.405 ;
        RECT 47.265 8.135 47.605 8.485 ;
        RECT 41.675 8.205 41.965 8.435 ;
      LAYER via1 ;
        RECT 47.365 8.235 47.515 8.385 ;
        RECT 47.375 4.1 47.525 4.25 ;
      LAYER mcon ;
        RECT 41.735 8.235 41.905 8.405 ;
        RECT 47.35 8.235 47.52 8.405 ;
        RECT 47.35 4.06 47.52 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 65.91 2.955 66.08 4.23 ;
        RECT 65.91 8.235 66.08 9.51 ;
        RECT 60.295 8.235 60.465 9.51 ;
      LAYER met2 ;
        RECT 65.835 4 66.175 4.35 ;
        RECT 65.825 8.135 66.165 8.485 ;
        RECT 65.91 4 66.08 8.485 ;
      LAYER met1 ;
        RECT 65.835 4.06 66.31 4.23 ;
        RECT 65.835 4 66.175 4.35 ;
        RECT 60.235 8.235 66.31 8.405 ;
        RECT 65.825 8.135 66.165 8.485 ;
        RECT 60.235 8.205 60.525 8.435 ;
      LAYER via1 ;
        RECT 65.925 8.235 66.075 8.385 ;
        RECT 65.935 4.1 66.085 4.25 ;
      LAYER mcon ;
        RECT 60.295 8.235 60.465 8.405 ;
        RECT 65.91 8.235 66.08 8.405 ;
        RECT 65.91 4.06 66.08 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 84.47 2.955 84.64 4.23 ;
        RECT 84.47 8.235 84.64 9.51 ;
        RECT 78.855 8.235 79.025 9.51 ;
      LAYER met2 ;
        RECT 84.395 4 84.735 4.35 ;
        RECT 84.385 8.135 84.725 8.485 ;
        RECT 84.47 4 84.64 8.485 ;
      LAYER met1 ;
        RECT 84.395 4.06 84.87 4.23 ;
        RECT 84.395 4 84.735 4.35 ;
        RECT 78.795 8.235 84.87 8.405 ;
        RECT 84.385 8.135 84.725 8.485 ;
        RECT 78.795 8.205 79.085 8.435 ;
      LAYER via1 ;
        RECT 84.485 8.235 84.635 8.385 ;
        RECT 84.495 4.1 84.645 4.25 ;
      LAYER mcon ;
        RECT 78.855 8.235 79.025 8.405 ;
        RECT 84.47 8.235 84.64 8.405 ;
        RECT 84.47 4.06 84.64 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 103.03 2.955 103.2 4.23 ;
        RECT 103.03 8.235 103.2 9.51 ;
        RECT 97.415 8.235 97.585 9.51 ;
      LAYER met2 ;
        RECT 102.955 4 103.295 4.35 ;
        RECT 102.945 8.135 103.285 8.485 ;
        RECT 103.03 4 103.2 8.485 ;
      LAYER met1 ;
        RECT 102.955 4.06 103.43 4.23 ;
        RECT 102.955 4 103.295 4.35 ;
        RECT 97.355 8.235 103.43 8.405 ;
        RECT 102.945 8.135 103.285 8.485 ;
        RECT 97.355 8.205 97.645 8.435 ;
      LAYER via1 ;
        RECT 103.045 8.235 103.195 8.385 ;
        RECT 103.055 4.1 103.205 4.25 ;
      LAYER mcon ;
        RECT 97.415 8.235 97.585 8.405 ;
        RECT 103.03 8.235 103.2 8.405 ;
        RECT 103.03 4.06 103.2 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 12.36 8.235 12.53 9.51 ;
      LAYER met1 ;
        RECT 12.27 8.235 12.76 8.405 ;
        RECT 12.27 8.195 12.61 8.455 ;
      LAYER mcon ;
        RECT 12.36 8.235 12.53 8.405 ;
    END
  END start
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 91.525 3.71 92.255 4.04 ;
        RECT 72.965 3.71 73.695 4.04 ;
        RECT 54.405 3.71 55.135 4.04 ;
        RECT 35.845 3.71 36.575 4.04 ;
        RECT 17.285 3.71 18.015 4.04 ;
        RECT 12.135 10.79 12.94 11.17 ;
        RECT 12.13 0 12.935 0.38 ;
      LAYER li1 ;
        RECT 12.13 10.865 107.73 12.465 ;
        RECT 106.75 10.24 106.92 12.465 ;
        RECT 105.76 10.24 105.93 12.465 ;
        RECT 103.02 10.235 103.19 12.465 ;
        RECT 97.405 10.235 97.575 12.465 ;
        RECT 88.19 10.24 88.36 12.465 ;
        RECT 87.2 10.24 87.37 12.465 ;
        RECT 84.46 10.235 84.63 12.465 ;
        RECT 78.845 10.235 79.015 12.465 ;
        RECT 69.63 10.24 69.8 12.465 ;
        RECT 68.64 10.24 68.81 12.465 ;
        RECT 65.9 10.235 66.07 12.465 ;
        RECT 60.285 10.235 60.455 12.465 ;
        RECT 51.07 10.24 51.24 12.465 ;
        RECT 50.08 10.24 50.25 12.465 ;
        RECT 47.34 10.235 47.51 12.465 ;
        RECT 41.725 10.235 41.895 12.465 ;
        RECT 32.51 10.24 32.68 12.465 ;
        RECT 31.52 10.24 31.69 12.465 ;
        RECT 28.78 10.235 28.95 12.465 ;
        RECT 23.165 10.235 23.335 12.465 ;
        RECT 12.13 10.865 15.53 12.475 ;
        RECT 12.135 10.855 12.94 12.475 ;
        RECT 12.35 10.835 12.6 12.475 ;
        RECT 12.35 10.235 12.52 12.475 ;
        RECT 12.13 0 107.725 1.6 ;
        RECT 106.75 0 106.92 2.225 ;
        RECT 105.76 0 105.93 2.225 ;
        RECT 103.02 0 103.19 2.23 ;
        RECT 89.91 0 101.955 2.88 ;
        RECT 100.96 0 101.13 3.38 ;
        RECT 100 0 100.17 3.38 ;
        RECT 99.04 0 99.21 3.38 ;
        RECT 98.52 0 98.69 3.38 ;
        RECT 98.24 0 98.435 2.89 ;
        RECT 97.56 0 97.73 3.38 ;
        RECT 96.56 0 96.73 3.38 ;
        RECT 95.6 0 95.77 3.38 ;
        RECT 94.565 0 94.76 2.89 ;
        RECT 94.12 0 94.29 3.38 ;
        RECT 92.2 0 92.46 2.89 ;
        RECT 92.2 0 92.37 3.38 ;
        RECT 90.72 0 90.89 3.38 ;
        RECT 88.19 0 88.36 2.225 ;
        RECT 87.2 0 87.37 2.225 ;
        RECT 84.46 0 84.63 2.23 ;
        RECT 71.35 0 83.395 2.88 ;
        RECT 82.4 0 82.57 3.38 ;
        RECT 81.44 0 81.61 3.38 ;
        RECT 80.48 0 80.65 3.38 ;
        RECT 79.96 0 80.13 3.38 ;
        RECT 79.68 0 79.875 2.89 ;
        RECT 79 0 79.17 3.38 ;
        RECT 78 0 78.17 3.38 ;
        RECT 77.04 0 77.21 3.38 ;
        RECT 76.005 0 76.2 2.89 ;
        RECT 75.56 0 75.73 3.38 ;
        RECT 73.64 0 73.9 2.89 ;
        RECT 73.64 0 73.81 3.38 ;
        RECT 72.16 0 72.33 3.38 ;
        RECT 69.63 0 69.8 2.225 ;
        RECT 68.64 0 68.81 2.225 ;
        RECT 65.9 0 66.07 2.23 ;
        RECT 52.79 0 64.835 2.88 ;
        RECT 63.84 0 64.01 3.38 ;
        RECT 62.88 0 63.05 3.38 ;
        RECT 61.92 0 62.09 3.38 ;
        RECT 61.4 0 61.57 3.38 ;
        RECT 61.12 0 61.315 2.89 ;
        RECT 60.44 0 60.61 3.38 ;
        RECT 59.44 0 59.61 3.38 ;
        RECT 58.48 0 58.65 3.38 ;
        RECT 57.445 0 57.64 2.89 ;
        RECT 57 0 57.17 3.38 ;
        RECT 55.08 0 55.34 2.89 ;
        RECT 55.08 0 55.25 3.38 ;
        RECT 53.6 0 53.77 3.38 ;
        RECT 51.07 0 51.24 2.225 ;
        RECT 50.08 0 50.25 2.225 ;
        RECT 47.34 0 47.51 2.23 ;
        RECT 34.23 0 46.275 2.88 ;
        RECT 45.28 0 45.45 3.38 ;
        RECT 44.32 0 44.49 3.38 ;
        RECT 43.36 0 43.53 3.38 ;
        RECT 42.84 0 43.01 3.38 ;
        RECT 42.56 0 42.755 2.89 ;
        RECT 41.88 0 42.05 3.38 ;
        RECT 40.88 0 41.05 3.38 ;
        RECT 39.92 0 40.09 3.38 ;
        RECT 38.885 0 39.08 2.89 ;
        RECT 38.44 0 38.61 3.38 ;
        RECT 36.52 0 36.78 2.89 ;
        RECT 36.52 0 36.69 3.38 ;
        RECT 35.04 0 35.21 3.38 ;
        RECT 32.51 0 32.68 2.225 ;
        RECT 31.52 0 31.69 2.225 ;
        RECT 28.78 0 28.95 2.23 ;
        RECT 15.67 0 27.715 2.88 ;
        RECT 26.72 0 26.89 3.38 ;
        RECT 25.76 0 25.93 3.38 ;
        RECT 24.8 0 24.97 3.38 ;
        RECT 24.28 0 24.45 3.38 ;
        RECT 24 0 24.195 2.89 ;
        RECT 23.32 0 23.49 3.38 ;
        RECT 22.32 0 22.49 3.38 ;
        RECT 21.36 0 21.53 3.38 ;
        RECT 20.325 0 20.52 2.89 ;
        RECT 19.88 0 20.05 3.38 ;
        RECT 17.96 0 18.22 2.89 ;
        RECT 17.96 0 18.13 3.38 ;
        RECT 16.48 0 16.65 3.38 ;
        RECT 98.41 8.365 98.58 10.315 ;
        RECT 98.355 10.145 98.525 10.595 ;
        RECT 98.355 7.305 98.525 8.535 ;
        RECT 93.4 3.79 93.57 4.12 ;
        RECT 91.56 4.35 91.85 4.52 ;
        RECT 91.56 3.87 91.73 4.52 ;
        RECT 91.36 3.87 91.73 4.04 ;
        RECT 79.85 8.365 80.02 10.315 ;
        RECT 79.795 10.145 79.965 10.595 ;
        RECT 79.795 7.305 79.965 8.535 ;
        RECT 74.84 3.79 75.01 4.12 ;
        RECT 73 4.35 73.29 4.52 ;
        RECT 73 3.87 73.17 4.52 ;
        RECT 72.8 3.87 73.17 4.04 ;
        RECT 61.29 8.365 61.46 10.315 ;
        RECT 61.235 10.145 61.405 10.595 ;
        RECT 61.235 7.305 61.405 8.535 ;
        RECT 56.28 3.79 56.45 4.12 ;
        RECT 54.44 4.35 54.73 4.52 ;
        RECT 54.44 3.87 54.61 4.52 ;
        RECT 54.24 3.87 54.61 4.04 ;
        RECT 42.73 8.365 42.9 10.315 ;
        RECT 42.675 10.145 42.845 10.595 ;
        RECT 42.675 7.305 42.845 8.535 ;
        RECT 37.72 3.79 37.89 4.12 ;
        RECT 35.88 4.35 36.17 4.52 ;
        RECT 35.88 3.87 36.05 4.52 ;
        RECT 35.68 3.87 36.05 4.04 ;
        RECT 24.17 8.365 24.34 10.315 ;
        RECT 24.115 10.145 24.285 10.595 ;
        RECT 24.115 7.305 24.285 8.535 ;
        RECT 19.16 3.79 19.33 4.12 ;
        RECT 17.32 4.35 17.61 4.52 ;
        RECT 17.32 3.87 17.49 4.52 ;
        RECT 17.12 3.87 17.49 4.04 ;
      LAYER met2 ;
        RECT 93.355 3.715 93.615 4.035 ;
        RECT 91.575 3.805 93.615 3.945 ;
        RECT 91.955 2.295 92.295 2.635 ;
        RECT 91.885 3.69 92.165 4.06 ;
        RECT 91.98 2.295 92.15 4.06 ;
        RECT 91.635 4.275 91.895 4.595 ;
        RECT 91.575 3.805 91.715 4.505 ;
        RECT 74.795 3.715 75.055 4.035 ;
        RECT 73.015 3.805 75.055 3.945 ;
        RECT 73.395 2.295 73.735 2.635 ;
        RECT 73.325 3.69 73.605 4.06 ;
        RECT 73.42 2.295 73.59 4.06 ;
        RECT 73.075 4.275 73.335 4.595 ;
        RECT 73.015 3.805 73.155 4.505 ;
        RECT 56.235 3.715 56.495 4.035 ;
        RECT 54.455 3.805 56.495 3.945 ;
        RECT 54.835 2.295 55.175 2.635 ;
        RECT 54.765 3.69 55.045 4.06 ;
        RECT 54.86 2.295 55.03 4.06 ;
        RECT 54.515 4.275 54.775 4.595 ;
        RECT 54.455 3.805 54.595 4.505 ;
        RECT 37.675 3.715 37.935 4.035 ;
        RECT 35.895 3.805 37.935 3.945 ;
        RECT 36.275 2.295 36.615 2.635 ;
        RECT 36.205 3.69 36.485 4.06 ;
        RECT 36.3 2.295 36.47 4.06 ;
        RECT 35.955 4.275 36.215 4.595 ;
        RECT 35.895 3.805 36.035 4.505 ;
        RECT 19.115 3.715 19.375 4.035 ;
        RECT 17.335 3.805 19.375 3.945 ;
        RECT 17.715 2.295 18.055 2.635 ;
        RECT 17.645 3.69 17.925 4.06 ;
        RECT 17.74 2.295 17.91 4.06 ;
        RECT 17.395 4.275 17.655 4.595 ;
        RECT 17.335 3.805 17.475 4.505 ;
        RECT 12.325 10.79 12.705 11.17 ;
        RECT 12.32 0 12.7 0.38 ;
        RECT 12.365 0 12.525 11.17 ;
      LAYER met1 ;
        RECT 12.13 10.865 107.73 12.465 ;
        RECT 98.35 8.575 98.64 8.805 ;
        RECT 97.915 8.605 98.64 8.775 ;
        RECT 97.915 8.605 98.085 12.465 ;
        RECT 79.79 8.575 80.08 8.805 ;
        RECT 79.355 8.605 80.08 8.775 ;
        RECT 79.355 8.605 79.525 12.465 ;
        RECT 61.23 8.575 61.52 8.805 ;
        RECT 60.795 8.605 61.52 8.775 ;
        RECT 60.795 8.605 60.965 12.465 ;
        RECT 42.67 8.575 42.96 8.805 ;
        RECT 42.235 8.605 42.96 8.775 ;
        RECT 42.235 8.605 42.405 12.465 ;
        RECT 24.11 8.575 24.4 8.805 ;
        RECT 23.675 8.605 24.4 8.775 ;
        RECT 23.675 8.605 23.845 12.465 ;
        RECT 12.13 10.865 15.53 12.475 ;
        RECT 12.135 10.855 12.94 12.475 ;
        RECT 12.34 10.835 12.69 12.475 ;
        RECT 12.13 0 107.725 1.6 ;
        RECT 89.91 0 101.955 2.88 ;
        RECT 89.91 0 101.87 3.035 ;
        RECT 71.35 0 83.395 2.88 ;
        RECT 71.35 0 83.31 3.035 ;
        RECT 52.79 0 64.835 2.88 ;
        RECT 52.79 0 64.75 3.035 ;
        RECT 34.23 0 46.275 2.88 ;
        RECT 34.23 0 46.19 3.035 ;
        RECT 15.67 0 27.715 2.88 ;
        RECT 15.67 0 27.63 3.035 ;
        RECT 93.34 3.665 93.63 4.035 ;
        RECT 92.575 3.665 93.63 3.805 ;
        RECT 91.605 4.305 91.925 4.565 ;
        RECT 74.78 3.665 75.07 4.035 ;
        RECT 74.015 3.665 75.07 3.805 ;
        RECT 73.045 4.305 73.365 4.565 ;
        RECT 56.22 3.665 56.51 4.035 ;
        RECT 55.455 3.665 56.51 3.805 ;
        RECT 54.485 4.305 54.805 4.565 ;
        RECT 37.66 3.665 37.95 4.035 ;
        RECT 36.895 3.665 37.95 3.805 ;
        RECT 35.925 4.305 36.245 4.565 ;
        RECT 19.1 3.665 19.39 4.035 ;
        RECT 18.335 3.665 19.39 3.805 ;
        RECT 17.365 4.305 17.685 4.565 ;
      LAYER via2 ;
        RECT 12.41 0.09 12.61 0.29 ;
        RECT 12.415 10.88 12.615 11.08 ;
        RECT 17.685 3.775 17.885 3.975 ;
        RECT 36.245 3.775 36.445 3.975 ;
        RECT 54.805 3.775 55.005 3.975 ;
        RECT 73.365 3.775 73.565 3.975 ;
        RECT 91.925 3.775 92.125 3.975 ;
      LAYER via1 ;
        RECT 12.435 0.115 12.585 0.265 ;
        RECT 12.44 10.905 12.59 11.055 ;
        RECT 17.45 4.36 17.6 4.51 ;
        RECT 17.81 2.39 17.96 2.54 ;
        RECT 19.17 3.8 19.32 3.95 ;
        RECT 36.01 4.36 36.16 4.51 ;
        RECT 36.37 2.39 36.52 2.54 ;
        RECT 37.73 3.8 37.88 3.95 ;
        RECT 54.57 4.36 54.72 4.51 ;
        RECT 54.93 2.39 55.08 2.54 ;
        RECT 56.29 3.8 56.44 3.95 ;
        RECT 73.13 4.36 73.28 4.51 ;
        RECT 73.49 2.39 73.64 2.54 ;
        RECT 74.85 3.8 75 3.95 ;
        RECT 91.69 4.36 91.84 4.51 ;
        RECT 92.05 2.39 92.2 2.54 ;
        RECT 93.41 3.8 93.56 3.95 ;
      LAYER mcon ;
        RECT 12.43 10.895 12.6 11.065 ;
        RECT 13.11 10.895 13.28 11.065 ;
        RECT 13.79 10.895 13.96 11.065 ;
        RECT 14.47 10.895 14.64 11.065 ;
        RECT 15.815 2.71 15.985 2.88 ;
        RECT 16.275 2.71 16.445 2.88 ;
        RECT 16.735 2.71 16.905 2.88 ;
        RECT 17.195 2.71 17.365 2.88 ;
        RECT 17.44 4.35 17.61 4.52 ;
        RECT 17.655 2.71 17.825 2.88 ;
        RECT 18.115 2.71 18.285 2.88 ;
        RECT 18.575 2.71 18.745 2.88 ;
        RECT 19.035 2.71 19.205 2.88 ;
        RECT 19.16 3.79 19.33 3.96 ;
        RECT 19.495 2.71 19.665 2.88 ;
        RECT 19.955 2.71 20.125 2.88 ;
        RECT 20.415 2.71 20.585 2.88 ;
        RECT 20.875 2.71 21.045 2.88 ;
        RECT 21.335 2.71 21.505 2.88 ;
        RECT 21.795 2.71 21.965 2.88 ;
        RECT 22.255 2.71 22.425 2.88 ;
        RECT 22.715 2.71 22.885 2.88 ;
        RECT 23.175 2.71 23.345 2.88 ;
        RECT 23.245 10.895 23.415 11.065 ;
        RECT 23.635 2.71 23.805 2.88 ;
        RECT 23.925 10.895 24.095 11.065 ;
        RECT 24.095 2.71 24.265 2.88 ;
        RECT 24.17 8.605 24.34 8.775 ;
        RECT 24.555 2.71 24.725 2.88 ;
        RECT 24.605 10.895 24.775 11.065 ;
        RECT 25.015 2.71 25.185 2.88 ;
        RECT 25.285 10.895 25.455 11.065 ;
        RECT 25.475 2.71 25.645 2.88 ;
        RECT 25.935 2.71 26.105 2.88 ;
        RECT 26.395 2.71 26.565 2.88 ;
        RECT 26.855 2.71 27.025 2.88 ;
        RECT 27.315 2.71 27.485 2.88 ;
        RECT 28.86 10.895 29.03 11.065 ;
        RECT 28.86 1.4 29.03 1.57 ;
        RECT 29.54 10.895 29.71 11.065 ;
        RECT 29.54 1.4 29.71 1.57 ;
        RECT 30.22 10.895 30.39 11.065 ;
        RECT 30.22 1.4 30.39 1.57 ;
        RECT 30.9 10.895 31.07 11.065 ;
        RECT 30.9 1.4 31.07 1.57 ;
        RECT 31.6 10.9 31.77 11.07 ;
        RECT 31.6 1.395 31.77 1.565 ;
        RECT 32.59 10.9 32.76 11.07 ;
        RECT 32.59 1.395 32.76 1.565 ;
        RECT 34.375 2.71 34.545 2.88 ;
        RECT 34.835 2.71 35.005 2.88 ;
        RECT 35.295 2.71 35.465 2.88 ;
        RECT 35.755 2.71 35.925 2.88 ;
        RECT 36 4.35 36.17 4.52 ;
        RECT 36.215 2.71 36.385 2.88 ;
        RECT 36.675 2.71 36.845 2.88 ;
        RECT 37.135 2.71 37.305 2.88 ;
        RECT 37.595 2.71 37.765 2.88 ;
        RECT 37.72 3.79 37.89 3.96 ;
        RECT 38.055 2.71 38.225 2.88 ;
        RECT 38.515 2.71 38.685 2.88 ;
        RECT 38.975 2.71 39.145 2.88 ;
        RECT 39.435 2.71 39.605 2.88 ;
        RECT 39.895 2.71 40.065 2.88 ;
        RECT 40.355 2.71 40.525 2.88 ;
        RECT 40.815 2.71 40.985 2.88 ;
        RECT 41.275 2.71 41.445 2.88 ;
        RECT 41.735 2.71 41.905 2.88 ;
        RECT 41.805 10.895 41.975 11.065 ;
        RECT 42.195 2.71 42.365 2.88 ;
        RECT 42.485 10.895 42.655 11.065 ;
        RECT 42.655 2.71 42.825 2.88 ;
        RECT 42.73 8.605 42.9 8.775 ;
        RECT 43.115 2.71 43.285 2.88 ;
        RECT 43.165 10.895 43.335 11.065 ;
        RECT 43.575 2.71 43.745 2.88 ;
        RECT 43.845 10.895 44.015 11.065 ;
        RECT 44.035 2.71 44.205 2.88 ;
        RECT 44.495 2.71 44.665 2.88 ;
        RECT 44.955 2.71 45.125 2.88 ;
        RECT 45.415 2.71 45.585 2.88 ;
        RECT 45.875 2.71 46.045 2.88 ;
        RECT 47.42 10.895 47.59 11.065 ;
        RECT 47.42 1.4 47.59 1.57 ;
        RECT 48.1 10.895 48.27 11.065 ;
        RECT 48.1 1.4 48.27 1.57 ;
        RECT 48.78 10.895 48.95 11.065 ;
        RECT 48.78 1.4 48.95 1.57 ;
        RECT 49.46 10.895 49.63 11.065 ;
        RECT 49.46 1.4 49.63 1.57 ;
        RECT 50.16 10.9 50.33 11.07 ;
        RECT 50.16 1.395 50.33 1.565 ;
        RECT 51.15 10.9 51.32 11.07 ;
        RECT 51.15 1.395 51.32 1.565 ;
        RECT 52.935 2.71 53.105 2.88 ;
        RECT 53.395 2.71 53.565 2.88 ;
        RECT 53.855 2.71 54.025 2.88 ;
        RECT 54.315 2.71 54.485 2.88 ;
        RECT 54.56 4.35 54.73 4.52 ;
        RECT 54.775 2.71 54.945 2.88 ;
        RECT 55.235 2.71 55.405 2.88 ;
        RECT 55.695 2.71 55.865 2.88 ;
        RECT 56.155 2.71 56.325 2.88 ;
        RECT 56.28 3.79 56.45 3.96 ;
        RECT 56.615 2.71 56.785 2.88 ;
        RECT 57.075 2.71 57.245 2.88 ;
        RECT 57.535 2.71 57.705 2.88 ;
        RECT 57.995 2.71 58.165 2.88 ;
        RECT 58.455 2.71 58.625 2.88 ;
        RECT 58.915 2.71 59.085 2.88 ;
        RECT 59.375 2.71 59.545 2.88 ;
        RECT 59.835 2.71 60.005 2.88 ;
        RECT 60.295 2.71 60.465 2.88 ;
        RECT 60.365 10.895 60.535 11.065 ;
        RECT 60.755 2.71 60.925 2.88 ;
        RECT 61.045 10.895 61.215 11.065 ;
        RECT 61.215 2.71 61.385 2.88 ;
        RECT 61.29 8.605 61.46 8.775 ;
        RECT 61.675 2.71 61.845 2.88 ;
        RECT 61.725 10.895 61.895 11.065 ;
        RECT 62.135 2.71 62.305 2.88 ;
        RECT 62.405 10.895 62.575 11.065 ;
        RECT 62.595 2.71 62.765 2.88 ;
        RECT 63.055 2.71 63.225 2.88 ;
        RECT 63.515 2.71 63.685 2.88 ;
        RECT 63.975 2.71 64.145 2.88 ;
        RECT 64.435 2.71 64.605 2.88 ;
        RECT 65.98 10.895 66.15 11.065 ;
        RECT 65.98 1.4 66.15 1.57 ;
        RECT 66.66 10.895 66.83 11.065 ;
        RECT 66.66 1.4 66.83 1.57 ;
        RECT 67.34 10.895 67.51 11.065 ;
        RECT 67.34 1.4 67.51 1.57 ;
        RECT 68.02 10.895 68.19 11.065 ;
        RECT 68.02 1.4 68.19 1.57 ;
        RECT 68.72 10.9 68.89 11.07 ;
        RECT 68.72 1.395 68.89 1.565 ;
        RECT 69.71 10.9 69.88 11.07 ;
        RECT 69.71 1.395 69.88 1.565 ;
        RECT 71.495 2.71 71.665 2.88 ;
        RECT 71.955 2.71 72.125 2.88 ;
        RECT 72.415 2.71 72.585 2.88 ;
        RECT 72.875 2.71 73.045 2.88 ;
        RECT 73.12 4.35 73.29 4.52 ;
        RECT 73.335 2.71 73.505 2.88 ;
        RECT 73.795 2.71 73.965 2.88 ;
        RECT 74.255 2.71 74.425 2.88 ;
        RECT 74.715 2.71 74.885 2.88 ;
        RECT 74.84 3.79 75.01 3.96 ;
        RECT 75.175 2.71 75.345 2.88 ;
        RECT 75.635 2.71 75.805 2.88 ;
        RECT 76.095 2.71 76.265 2.88 ;
        RECT 76.555 2.71 76.725 2.88 ;
        RECT 77.015 2.71 77.185 2.88 ;
        RECT 77.475 2.71 77.645 2.88 ;
        RECT 77.935 2.71 78.105 2.88 ;
        RECT 78.395 2.71 78.565 2.88 ;
        RECT 78.855 2.71 79.025 2.88 ;
        RECT 78.925 10.895 79.095 11.065 ;
        RECT 79.315 2.71 79.485 2.88 ;
        RECT 79.605 10.895 79.775 11.065 ;
        RECT 79.775 2.71 79.945 2.88 ;
        RECT 79.85 8.605 80.02 8.775 ;
        RECT 80.235 2.71 80.405 2.88 ;
        RECT 80.285 10.895 80.455 11.065 ;
        RECT 80.695 2.71 80.865 2.88 ;
        RECT 80.965 10.895 81.135 11.065 ;
        RECT 81.155 2.71 81.325 2.88 ;
        RECT 81.615 2.71 81.785 2.88 ;
        RECT 82.075 2.71 82.245 2.88 ;
        RECT 82.535 2.71 82.705 2.88 ;
        RECT 82.995 2.71 83.165 2.88 ;
        RECT 84.54 10.895 84.71 11.065 ;
        RECT 84.54 1.4 84.71 1.57 ;
        RECT 85.22 10.895 85.39 11.065 ;
        RECT 85.22 1.4 85.39 1.57 ;
        RECT 85.9 10.895 86.07 11.065 ;
        RECT 85.9 1.4 86.07 1.57 ;
        RECT 86.58 10.895 86.75 11.065 ;
        RECT 86.58 1.4 86.75 1.57 ;
        RECT 87.28 10.9 87.45 11.07 ;
        RECT 87.28 1.395 87.45 1.565 ;
        RECT 88.27 10.9 88.44 11.07 ;
        RECT 88.27 1.395 88.44 1.565 ;
        RECT 90.055 2.71 90.225 2.88 ;
        RECT 90.515 2.71 90.685 2.88 ;
        RECT 90.975 2.71 91.145 2.88 ;
        RECT 91.435 2.71 91.605 2.88 ;
        RECT 91.68 4.35 91.85 4.52 ;
        RECT 91.895 2.71 92.065 2.88 ;
        RECT 92.355 2.71 92.525 2.88 ;
        RECT 92.815 2.71 92.985 2.88 ;
        RECT 93.275 2.71 93.445 2.88 ;
        RECT 93.4 3.79 93.57 3.96 ;
        RECT 93.735 2.71 93.905 2.88 ;
        RECT 94.195 2.71 94.365 2.88 ;
        RECT 94.655 2.71 94.825 2.88 ;
        RECT 95.115 2.71 95.285 2.88 ;
        RECT 95.575 2.71 95.745 2.88 ;
        RECT 96.035 2.71 96.205 2.88 ;
        RECT 96.495 2.71 96.665 2.88 ;
        RECT 96.955 2.71 97.125 2.88 ;
        RECT 97.415 2.71 97.585 2.88 ;
        RECT 97.485 10.895 97.655 11.065 ;
        RECT 97.875 2.71 98.045 2.88 ;
        RECT 98.165 10.895 98.335 11.065 ;
        RECT 98.335 2.71 98.505 2.88 ;
        RECT 98.41 8.605 98.58 8.775 ;
        RECT 98.795 2.71 98.965 2.88 ;
        RECT 98.845 10.895 99.015 11.065 ;
        RECT 99.255 2.71 99.425 2.88 ;
        RECT 99.525 10.895 99.695 11.065 ;
        RECT 99.715 2.71 99.885 2.88 ;
        RECT 100.175 2.71 100.345 2.88 ;
        RECT 100.635 2.71 100.805 2.88 ;
        RECT 101.095 2.71 101.265 2.88 ;
        RECT 101.555 2.71 101.725 2.88 ;
        RECT 103.1 10.895 103.27 11.065 ;
        RECT 103.1 1.4 103.27 1.57 ;
        RECT 103.78 10.895 103.95 11.065 ;
        RECT 103.78 1.4 103.95 1.57 ;
        RECT 104.46 10.895 104.63 11.065 ;
        RECT 104.46 1.4 104.63 1.57 ;
        RECT 105.14 10.895 105.31 11.065 ;
        RECT 105.14 1.4 105.31 1.57 ;
        RECT 105.84 10.9 106.01 11.07 ;
        RECT 105.84 1.395 106.01 1.565 ;
        RECT 106.83 10.9 107 11.07 ;
        RECT 106.83 1.395 107 1.565 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 99.215 4.83 99.77 5.16 ;
      RECT 99.215 3.165 99.515 5.16 ;
      RECT 95.28 4.27 95.835 4.6 ;
      RECT 95.535 3.165 95.835 4.6 ;
      RECT 95.535 3.165 99.515 3.465 ;
      RECT 98.685 9.345 99.06 9.715 ;
      RECT 98.685 9.385 99.69 9.685 ;
      RECT 99.39 6.695 99.69 9.685 ;
      RECT 89.56 6.695 99.69 6.995 ;
      RECT 94.065 3.71 94.365 6.995 ;
      RECT 92.63 4.27 92.93 6.995 ;
      RECT 89.56 3.715 89.86 6.995 ;
      RECT 92.6 4.27 93.33 4.6 ;
      RECT 94.04 3.71 94.77 4.04 ;
      RECT 90.49 3.71 91.22 4.04 ;
      RECT 89.56 3.715 91.22 4.015 ;
      RECT 80.655 4.83 81.21 5.16 ;
      RECT 80.655 3.165 80.955 5.16 ;
      RECT 76.72 4.27 77.275 4.6 ;
      RECT 76.975 3.165 77.275 4.6 ;
      RECT 76.975 3.165 80.955 3.465 ;
      RECT 80.125 9.345 80.5 9.715 ;
      RECT 80.125 9.385 81.13 9.685 ;
      RECT 80.83 6.695 81.13 9.685 ;
      RECT 71 6.695 81.13 6.995 ;
      RECT 75.505 3.71 75.805 6.995 ;
      RECT 74.07 4.27 74.37 6.995 ;
      RECT 71 3.715 71.3 6.995 ;
      RECT 74.04 4.27 74.77 4.6 ;
      RECT 75.48 3.71 76.21 4.04 ;
      RECT 71.93 3.71 72.66 4.04 ;
      RECT 71 3.715 72.66 4.015 ;
      RECT 62.095 4.83 62.65 5.16 ;
      RECT 62.095 3.165 62.395 5.16 ;
      RECT 58.16 4.27 58.715 4.6 ;
      RECT 58.415 3.165 58.715 4.6 ;
      RECT 58.415 3.165 62.395 3.465 ;
      RECT 61.565 9.345 61.94 9.715 ;
      RECT 61.565 9.385 62.57 9.685 ;
      RECT 62.27 6.695 62.57 9.685 ;
      RECT 52.44 6.695 62.57 6.995 ;
      RECT 56.945 3.71 57.245 6.995 ;
      RECT 55.51 4.27 55.81 6.995 ;
      RECT 52.44 3.715 52.74 6.995 ;
      RECT 55.48 4.27 56.21 4.6 ;
      RECT 56.92 3.71 57.65 4.04 ;
      RECT 53.37 3.71 54.1 4.04 ;
      RECT 52.44 3.715 54.1 4.015 ;
      RECT 43.535 4.83 44.09 5.16 ;
      RECT 43.535 3.165 43.835 5.16 ;
      RECT 39.6 4.27 40.155 4.6 ;
      RECT 39.855 3.165 40.155 4.6 ;
      RECT 39.855 3.165 43.835 3.465 ;
      RECT 43.005 9.345 43.38 9.715 ;
      RECT 43.005 9.385 44.01 9.685 ;
      RECT 43.71 6.695 44.01 9.685 ;
      RECT 33.88 6.695 44.01 6.995 ;
      RECT 38.385 3.71 38.685 6.995 ;
      RECT 36.95 4.27 37.25 6.995 ;
      RECT 33.88 3.715 34.18 6.995 ;
      RECT 36.92 4.27 37.65 4.6 ;
      RECT 38.36 3.71 39.09 4.04 ;
      RECT 34.81 3.71 35.54 4.04 ;
      RECT 33.88 3.715 35.54 4.015 ;
      RECT 24.975 4.83 25.53 5.16 ;
      RECT 24.975 3.165 25.275 5.16 ;
      RECT 21.04 4.27 21.595 4.6 ;
      RECT 21.295 3.165 21.595 4.6 ;
      RECT 21.295 3.165 25.275 3.465 ;
      RECT 24.445 9.345 24.82 9.715 ;
      RECT 24.445 9.385 25.45 9.685 ;
      RECT 25.15 6.695 25.45 9.685 ;
      RECT 15.32 6.695 25.45 6.995 ;
      RECT 19.825 3.71 20.125 6.995 ;
      RECT 18.39 4.27 18.69 6.995 ;
      RECT 15.32 3.715 15.62 6.995 ;
      RECT 18.36 4.27 19.09 4.6 ;
      RECT 19.8 3.71 20.53 4.04 ;
      RECT 16.25 3.71 16.98 4.04 ;
      RECT 15.32 3.715 16.98 4.015 ;
      RECT 100.4 3.15 101.13 3.48 ;
      RECT 98.18 4.83 98.91 5.16 ;
      RECT 96.48 4.83 97.21 5.16 ;
      RECT 90.16 4.83 90.89 5.16 ;
      RECT 81.84 3.15 82.57 3.48 ;
      RECT 79.62 4.83 80.35 5.16 ;
      RECT 77.92 4.83 78.65 5.16 ;
      RECT 71.6 4.83 72.33 5.16 ;
      RECT 63.28 3.15 64.01 3.48 ;
      RECT 61.06 4.83 61.79 5.16 ;
      RECT 59.36 4.83 60.09 5.16 ;
      RECT 53.04 4.83 53.77 5.16 ;
      RECT 44.72 3.15 45.45 3.48 ;
      RECT 42.5 4.83 43.23 5.16 ;
      RECT 40.8 4.83 41.53 5.16 ;
      RECT 34.48 4.83 35.21 5.16 ;
      RECT 26.16 3.15 26.89 3.48 ;
      RECT 23.94 4.83 24.67 5.16 ;
      RECT 22.24 4.83 22.97 5.16 ;
      RECT 15.92 4.83 16.65 5.16 ;
    LAYER via2 ;
      RECT 100.465 3.215 100.665 3.415 ;
      RECT 99.505 4.895 99.705 5.095 ;
      RECT 98.77 9.43 98.97 9.63 ;
      RECT 98.505 4.895 98.705 5.095 ;
      RECT 96.545 4.895 96.745 5.095 ;
      RECT 95.345 4.335 95.545 4.535 ;
      RECT 94.105 3.775 94.305 3.975 ;
      RECT 92.665 4.335 92.865 4.535 ;
      RECT 90.705 3.775 90.905 3.975 ;
      RECT 90.225 4.895 90.425 5.095 ;
      RECT 81.905 3.215 82.105 3.415 ;
      RECT 80.945 4.895 81.145 5.095 ;
      RECT 80.21 9.43 80.41 9.63 ;
      RECT 79.945 4.895 80.145 5.095 ;
      RECT 77.985 4.895 78.185 5.095 ;
      RECT 76.785 4.335 76.985 4.535 ;
      RECT 75.545 3.775 75.745 3.975 ;
      RECT 74.105 4.335 74.305 4.535 ;
      RECT 72.145 3.775 72.345 3.975 ;
      RECT 71.665 4.895 71.865 5.095 ;
      RECT 63.345 3.215 63.545 3.415 ;
      RECT 62.385 4.895 62.585 5.095 ;
      RECT 61.65 9.43 61.85 9.63 ;
      RECT 61.385 4.895 61.585 5.095 ;
      RECT 59.425 4.895 59.625 5.095 ;
      RECT 58.225 4.335 58.425 4.535 ;
      RECT 56.985 3.775 57.185 3.975 ;
      RECT 55.545 4.335 55.745 4.535 ;
      RECT 53.585 3.775 53.785 3.975 ;
      RECT 53.105 4.895 53.305 5.095 ;
      RECT 44.785 3.215 44.985 3.415 ;
      RECT 43.825 4.895 44.025 5.095 ;
      RECT 43.09 9.43 43.29 9.63 ;
      RECT 42.825 4.895 43.025 5.095 ;
      RECT 40.865 4.895 41.065 5.095 ;
      RECT 39.665 4.335 39.865 4.535 ;
      RECT 38.425 3.775 38.625 3.975 ;
      RECT 36.985 4.335 37.185 4.535 ;
      RECT 35.025 3.775 35.225 3.975 ;
      RECT 34.545 4.895 34.745 5.095 ;
      RECT 26.225 3.215 26.425 3.415 ;
      RECT 25.265 4.895 25.465 5.095 ;
      RECT 24.53 9.43 24.73 9.63 ;
      RECT 24.265 4.895 24.465 5.095 ;
      RECT 22.305 4.895 22.505 5.095 ;
      RECT 21.105 4.335 21.305 4.535 ;
      RECT 19.865 3.775 20.065 3.975 ;
      RECT 18.425 4.335 18.625 4.535 ;
      RECT 16.465 3.775 16.665 3.975 ;
      RECT 15.985 4.895 16.185 5.095 ;
    LAYER met2 ;
      RECT 13.355 10.69 107.355 10.86 ;
      RECT 107.185 9.565 107.355 10.86 ;
      RECT 13.355 8.545 13.525 10.86 ;
      RECT 107.155 9.565 107.505 9.915 ;
      RECT 13.295 8.545 13.585 8.895 ;
      RECT 103.995 8.51 104.315 8.835 ;
      RECT 104.025 7.985 104.195 8.835 ;
      RECT 104.025 7.985 104.2 8.335 ;
      RECT 104.025 7.985 105 8.16 ;
      RECT 104.825 3.26 105 8.16 ;
      RECT 104.77 3.26 105.12 3.61 ;
      RECT 104.795 8.945 105.12 9.27 ;
      RECT 103.68 9.035 105.12 9.205 ;
      RECT 103.68 3.69 103.84 9.205 ;
      RECT 103.995 3.66 104.315 3.98 ;
      RECT 103.68 3.69 104.315 3.86 ;
      RECT 96.56 5.43 102.65 5.62 ;
      RECT 102.48 4.44 102.65 5.62 ;
      RECT 102.46 4.445 102.65 5.62 ;
      RECT 96.56 4.81 96.73 5.62 ;
      RECT 96.505 4.81 96.785 5.18 ;
      RECT 96.575 4.365 96.715 5.62 ;
      RECT 102.39 4.445 102.73 4.795 ;
      RECT 96.385 4.25 96.665 4.62 ;
      RECT 96.095 4.365 96.715 4.505 ;
      RECT 96.095 3.155 96.235 4.505 ;
      RECT 96.035 3.155 96.295 3.475 ;
      RECT 88.57 8.945 88.92 9.295 ;
      RECT 99.355 8.9 99.705 9.25 ;
      RECT 88.57 8.975 99.705 9.175 ;
      RECT 98.995 4.275 99.255 4.595 ;
      RECT 99.055 3.155 99.195 4.595 ;
      RECT 98.995 3.155 99.255 3.475 ;
      RECT 97.995 4.835 98.255 5.155 ;
      RECT 97.995 4.25 98.195 5.155 ;
      RECT 97.935 3.155 98.075 4.785 ;
      RECT 97.935 4.25 98.435 4.62 ;
      RECT 97.875 3.155 98.135 3.475 ;
      RECT 97.515 4.835 97.775 5.155 ;
      RECT 97.575 3.245 97.715 5.155 ;
      RECT 97.275 3.245 97.715 3.475 ;
      RECT 97.275 3.155 97.535 3.475 ;
      RECT 97.035 3.715 97.295 4.035 ;
      RECT 96.455 3.805 97.295 3.945 ;
      RECT 96.455 2.865 96.595 3.945 ;
      RECT 93.115 3.155 93.375 3.475 ;
      RECT 93.115 3.245 94.155 3.385 ;
      RECT 94.015 2.865 94.155 3.385 ;
      RECT 94.015 2.865 96.595 3.005 ;
      RECT 95.305 4.25 95.585 4.62 ;
      RECT 95.375 3.155 95.515 4.62 ;
      RECT 95.315 3.155 95.575 3.475 ;
      RECT 94.955 4.835 95.215 5.155 ;
      RECT 95.015 3.245 95.155 5.155 ;
      RECT 94.595 3.155 94.855 3.475 ;
      RECT 94.595 3.245 95.155 3.385 ;
      RECT 92.625 4.25 92.905 4.62 ;
      RECT 94.595 4.275 94.855 4.595 ;
      RECT 92.275 4.275 92.905 4.595 ;
      RECT 92.275 4.365 94.855 4.505 ;
      RECT 94.065 3.69 94.345 4.06 ;
      RECT 94.065 3.715 94.595 4.035 ;
      RECT 91.155 4.275 91.415 4.595 ;
      RECT 91.215 3.155 91.355 4.595 ;
      RECT 91.155 3.155 91.415 3.475 ;
      RECT 90.185 4.81 90.465 5.18 ;
      RECT 90.195 4.555 90.455 5.18 ;
      RECT 85.435 8.51 85.755 8.835 ;
      RECT 85.465 7.985 85.635 8.835 ;
      RECT 85.465 7.985 85.64 8.335 ;
      RECT 85.465 7.985 86.44 8.16 ;
      RECT 86.265 3.26 86.44 8.16 ;
      RECT 86.21 3.26 86.56 3.61 ;
      RECT 86.235 8.945 86.56 9.27 ;
      RECT 85.12 9.035 86.56 9.205 ;
      RECT 85.12 3.69 85.28 9.205 ;
      RECT 85.435 3.66 85.755 3.98 ;
      RECT 85.12 3.69 85.755 3.86 ;
      RECT 78 5.43 84.09 5.62 ;
      RECT 83.92 4.44 84.09 5.62 ;
      RECT 83.9 4.445 84.09 5.62 ;
      RECT 78 4.81 78.17 5.62 ;
      RECT 77.945 4.81 78.225 5.18 ;
      RECT 78.015 4.365 78.155 5.62 ;
      RECT 83.83 4.445 84.17 4.795 ;
      RECT 77.825 4.25 78.105 4.62 ;
      RECT 77.535 4.365 78.155 4.505 ;
      RECT 77.535 3.155 77.675 4.505 ;
      RECT 77.475 3.155 77.735 3.475 ;
      RECT 70.01 8.945 70.36 9.295 ;
      RECT 80.795 8.9 81.145 9.25 ;
      RECT 70.01 8.975 81.145 9.175 ;
      RECT 80.435 4.275 80.695 4.595 ;
      RECT 80.495 3.155 80.635 4.595 ;
      RECT 80.435 3.155 80.695 3.475 ;
      RECT 79.435 4.835 79.695 5.155 ;
      RECT 79.435 4.25 79.635 5.155 ;
      RECT 79.375 3.155 79.515 4.785 ;
      RECT 79.375 4.25 79.875 4.62 ;
      RECT 79.315 3.155 79.575 3.475 ;
      RECT 78.955 4.835 79.215 5.155 ;
      RECT 79.015 3.245 79.155 5.155 ;
      RECT 78.715 3.245 79.155 3.475 ;
      RECT 78.715 3.155 78.975 3.475 ;
      RECT 78.475 3.715 78.735 4.035 ;
      RECT 77.895 3.805 78.735 3.945 ;
      RECT 77.895 2.865 78.035 3.945 ;
      RECT 74.555 3.155 74.815 3.475 ;
      RECT 74.555 3.245 75.595 3.385 ;
      RECT 75.455 2.865 75.595 3.385 ;
      RECT 75.455 2.865 78.035 3.005 ;
      RECT 76.745 4.25 77.025 4.62 ;
      RECT 76.815 3.155 76.955 4.62 ;
      RECT 76.755 3.155 77.015 3.475 ;
      RECT 76.395 4.835 76.655 5.155 ;
      RECT 76.455 3.245 76.595 5.155 ;
      RECT 76.035 3.155 76.295 3.475 ;
      RECT 76.035 3.245 76.595 3.385 ;
      RECT 74.065 4.25 74.345 4.62 ;
      RECT 76.035 4.275 76.295 4.595 ;
      RECT 73.715 4.275 74.345 4.595 ;
      RECT 73.715 4.365 76.295 4.505 ;
      RECT 75.505 3.69 75.785 4.06 ;
      RECT 75.505 3.715 76.035 4.035 ;
      RECT 72.595 4.275 72.855 4.595 ;
      RECT 72.655 3.155 72.795 4.595 ;
      RECT 72.595 3.155 72.855 3.475 ;
      RECT 71.625 4.81 71.905 5.18 ;
      RECT 71.635 4.555 71.895 5.18 ;
      RECT 66.875 8.51 67.195 8.835 ;
      RECT 66.905 7.985 67.075 8.835 ;
      RECT 66.905 7.985 67.08 8.335 ;
      RECT 66.905 7.985 67.88 8.16 ;
      RECT 67.705 3.26 67.88 8.16 ;
      RECT 67.65 3.26 68 3.61 ;
      RECT 67.675 8.945 68 9.27 ;
      RECT 66.56 9.035 68 9.205 ;
      RECT 66.56 3.69 66.72 9.205 ;
      RECT 66.875 3.66 67.195 3.98 ;
      RECT 66.56 3.69 67.195 3.86 ;
      RECT 59.44 5.43 65.53 5.62 ;
      RECT 65.36 4.44 65.53 5.62 ;
      RECT 65.34 4.445 65.53 5.62 ;
      RECT 59.44 4.81 59.61 5.62 ;
      RECT 59.385 4.81 59.665 5.18 ;
      RECT 59.455 4.365 59.595 5.62 ;
      RECT 65.27 4.445 65.61 4.795 ;
      RECT 59.265 4.25 59.545 4.62 ;
      RECT 58.975 4.365 59.595 4.505 ;
      RECT 58.975 3.155 59.115 4.505 ;
      RECT 58.915 3.155 59.175 3.475 ;
      RECT 51.495 8.95 51.845 9.3 ;
      RECT 62.235 8.905 62.585 9.255 ;
      RECT 51.495 8.98 62.585 9.18 ;
      RECT 61.875 4.275 62.135 4.595 ;
      RECT 61.935 3.155 62.075 4.595 ;
      RECT 61.875 3.155 62.135 3.475 ;
      RECT 60.875 4.835 61.135 5.155 ;
      RECT 60.875 4.25 61.075 5.155 ;
      RECT 60.815 3.155 60.955 4.785 ;
      RECT 60.815 4.25 61.315 4.62 ;
      RECT 60.755 3.155 61.015 3.475 ;
      RECT 60.395 4.835 60.655 5.155 ;
      RECT 60.455 3.245 60.595 5.155 ;
      RECT 60.155 3.245 60.595 3.475 ;
      RECT 60.155 3.155 60.415 3.475 ;
      RECT 59.915 3.715 60.175 4.035 ;
      RECT 59.335 3.805 60.175 3.945 ;
      RECT 59.335 2.865 59.475 3.945 ;
      RECT 55.995 3.155 56.255 3.475 ;
      RECT 55.995 3.245 57.035 3.385 ;
      RECT 56.895 2.865 57.035 3.385 ;
      RECT 56.895 2.865 59.475 3.005 ;
      RECT 58.185 4.25 58.465 4.62 ;
      RECT 58.255 3.155 58.395 4.62 ;
      RECT 58.195 3.155 58.455 3.475 ;
      RECT 57.835 4.835 58.095 5.155 ;
      RECT 57.895 3.245 58.035 5.155 ;
      RECT 57.475 3.155 57.735 3.475 ;
      RECT 57.475 3.245 58.035 3.385 ;
      RECT 55.505 4.25 55.785 4.62 ;
      RECT 57.475 4.275 57.735 4.595 ;
      RECT 55.155 4.275 55.785 4.595 ;
      RECT 55.155 4.365 57.735 4.505 ;
      RECT 56.945 3.69 57.225 4.06 ;
      RECT 56.945 3.715 57.475 4.035 ;
      RECT 54.035 4.275 54.295 4.595 ;
      RECT 54.095 3.155 54.235 4.595 ;
      RECT 54.035 3.155 54.295 3.475 ;
      RECT 53.065 4.81 53.345 5.18 ;
      RECT 53.075 4.555 53.335 5.18 ;
      RECT 48.315 8.51 48.635 8.835 ;
      RECT 48.345 7.985 48.515 8.835 ;
      RECT 48.345 7.985 48.52 8.335 ;
      RECT 48.345 7.985 49.32 8.16 ;
      RECT 49.145 3.26 49.32 8.16 ;
      RECT 49.09 3.26 49.44 3.61 ;
      RECT 49.115 8.945 49.44 9.27 ;
      RECT 48 9.035 49.44 9.205 ;
      RECT 48 3.69 48.16 9.205 ;
      RECT 48.315 3.66 48.635 3.98 ;
      RECT 48 3.69 48.635 3.86 ;
      RECT 40.88 5.43 46.97 5.62 ;
      RECT 46.8 4.44 46.97 5.62 ;
      RECT 46.78 4.445 46.97 5.62 ;
      RECT 40.88 4.81 41.05 5.62 ;
      RECT 40.825 4.81 41.105 5.18 ;
      RECT 40.895 4.365 41.035 5.62 ;
      RECT 46.71 4.445 47.05 4.795 ;
      RECT 40.705 4.25 40.985 4.62 ;
      RECT 40.415 4.365 41.035 4.505 ;
      RECT 40.415 3.155 40.555 4.505 ;
      RECT 40.355 3.155 40.615 3.475 ;
      RECT 32.935 8.945 33.285 9.295 ;
      RECT 43.68 8.9 44.03 9.25 ;
      RECT 32.935 8.975 44.03 9.175 ;
      RECT 43.315 4.275 43.575 4.595 ;
      RECT 43.375 3.155 43.515 4.595 ;
      RECT 43.315 3.155 43.575 3.475 ;
      RECT 42.315 4.835 42.575 5.155 ;
      RECT 42.315 4.25 42.515 5.155 ;
      RECT 42.255 3.155 42.395 4.785 ;
      RECT 42.255 4.25 42.755 4.62 ;
      RECT 42.195 3.155 42.455 3.475 ;
      RECT 41.835 4.835 42.095 5.155 ;
      RECT 41.895 3.245 42.035 5.155 ;
      RECT 41.595 3.245 42.035 3.475 ;
      RECT 41.595 3.155 41.855 3.475 ;
      RECT 41.355 3.715 41.615 4.035 ;
      RECT 40.775 3.805 41.615 3.945 ;
      RECT 40.775 2.865 40.915 3.945 ;
      RECT 37.435 3.155 37.695 3.475 ;
      RECT 37.435 3.245 38.475 3.385 ;
      RECT 38.335 2.865 38.475 3.385 ;
      RECT 38.335 2.865 40.915 3.005 ;
      RECT 39.625 4.25 39.905 4.62 ;
      RECT 39.695 3.155 39.835 4.62 ;
      RECT 39.635 3.155 39.895 3.475 ;
      RECT 39.275 4.835 39.535 5.155 ;
      RECT 39.335 3.245 39.475 5.155 ;
      RECT 38.915 3.155 39.175 3.475 ;
      RECT 38.915 3.245 39.475 3.385 ;
      RECT 36.945 4.25 37.225 4.62 ;
      RECT 38.915 4.275 39.175 4.595 ;
      RECT 36.595 4.275 37.225 4.595 ;
      RECT 36.595 4.365 39.175 4.505 ;
      RECT 38.385 3.69 38.665 4.06 ;
      RECT 38.385 3.715 38.915 4.035 ;
      RECT 35.475 4.275 35.735 4.595 ;
      RECT 35.535 3.155 35.675 4.595 ;
      RECT 35.475 3.155 35.735 3.475 ;
      RECT 34.505 4.81 34.785 5.18 ;
      RECT 34.515 4.555 34.775 5.18 ;
      RECT 29.755 8.51 30.075 8.835 ;
      RECT 29.785 7.985 29.955 8.835 ;
      RECT 29.785 7.985 29.96 8.335 ;
      RECT 29.785 7.985 30.76 8.16 ;
      RECT 30.585 3.26 30.76 8.16 ;
      RECT 30.53 3.26 30.88 3.61 ;
      RECT 30.555 8.945 30.88 9.27 ;
      RECT 29.44 9.035 30.88 9.205 ;
      RECT 29.44 3.69 29.6 9.205 ;
      RECT 29.755 3.66 30.075 3.98 ;
      RECT 29.44 3.69 30.075 3.86 ;
      RECT 22.32 5.43 28.41 5.62 ;
      RECT 28.24 4.44 28.41 5.62 ;
      RECT 28.22 4.445 28.41 5.62 ;
      RECT 22.32 4.81 22.49 5.62 ;
      RECT 22.265 4.81 22.545 5.18 ;
      RECT 22.335 4.365 22.475 5.62 ;
      RECT 28.15 4.445 28.49 4.795 ;
      RECT 22.145 4.25 22.425 4.62 ;
      RECT 21.855 4.365 22.475 4.505 ;
      RECT 21.855 3.155 21.995 4.505 ;
      RECT 21.795 3.155 22.055 3.475 ;
      RECT 13.67 9.285 13.96 9.635 ;
      RECT 13.67 9.345 14.86 9.515 ;
      RECT 14.69 8.975 14.86 9.515 ;
      RECT 25.12 8.895 25.47 9.245 ;
      RECT 14.69 8.975 25.47 9.145 ;
      RECT 24.755 4.275 25.015 4.595 ;
      RECT 24.815 3.155 24.955 4.595 ;
      RECT 24.755 3.155 25.015 3.475 ;
      RECT 23.755 4.835 24.015 5.155 ;
      RECT 23.755 4.25 23.955 5.155 ;
      RECT 23.695 3.155 23.835 4.785 ;
      RECT 23.695 4.25 24.195 4.62 ;
      RECT 23.635 3.155 23.895 3.475 ;
      RECT 23.275 4.835 23.535 5.155 ;
      RECT 23.335 3.245 23.475 5.155 ;
      RECT 23.035 3.245 23.475 3.475 ;
      RECT 23.035 3.155 23.295 3.475 ;
      RECT 22.795 3.715 23.055 4.035 ;
      RECT 22.215 3.805 23.055 3.945 ;
      RECT 22.215 2.865 22.355 3.945 ;
      RECT 18.875 3.155 19.135 3.475 ;
      RECT 18.875 3.245 19.915 3.385 ;
      RECT 19.775 2.865 19.915 3.385 ;
      RECT 19.775 2.865 22.355 3.005 ;
      RECT 21.065 4.25 21.345 4.62 ;
      RECT 21.135 3.155 21.275 4.62 ;
      RECT 21.075 3.155 21.335 3.475 ;
      RECT 20.715 4.835 20.975 5.155 ;
      RECT 20.775 3.245 20.915 5.155 ;
      RECT 20.355 3.155 20.615 3.475 ;
      RECT 20.355 3.245 20.915 3.385 ;
      RECT 18.385 4.25 18.665 4.62 ;
      RECT 20.355 4.275 20.615 4.595 ;
      RECT 18.035 4.275 18.665 4.595 ;
      RECT 18.035 4.365 20.615 4.505 ;
      RECT 19.825 3.69 20.105 4.06 ;
      RECT 19.825 3.715 20.355 4.035 ;
      RECT 16.915 4.275 17.175 4.595 ;
      RECT 16.975 3.155 17.115 4.595 ;
      RECT 16.915 3.155 17.175 3.475 ;
      RECT 15.945 4.81 16.225 5.18 ;
      RECT 15.955 4.555 16.215 5.18 ;
      RECT 100.425 3.13 100.705 3.5 ;
      RECT 99.465 4.81 99.745 5.18 ;
      RECT 98.685 9.345 99.06 9.715 ;
      RECT 98.465 4.81 98.745 5.18 ;
      RECT 90.665 3.69 90.945 4.06 ;
      RECT 81.865 3.13 82.145 3.5 ;
      RECT 80.905 4.81 81.185 5.18 ;
      RECT 80.125 9.345 80.5 9.715 ;
      RECT 79.905 4.81 80.185 5.18 ;
      RECT 72.105 3.69 72.385 4.06 ;
      RECT 63.305 3.13 63.585 3.5 ;
      RECT 62.345 4.81 62.625 5.18 ;
      RECT 61.565 9.345 61.94 9.715 ;
      RECT 61.345 4.81 61.625 5.18 ;
      RECT 53.545 3.69 53.825 4.06 ;
      RECT 44.745 3.13 45.025 3.5 ;
      RECT 43.785 4.81 44.065 5.18 ;
      RECT 43.005 9.345 43.38 9.715 ;
      RECT 42.785 4.81 43.065 5.18 ;
      RECT 34.985 3.69 35.265 4.06 ;
      RECT 26.185 3.13 26.465 3.5 ;
      RECT 25.225 4.81 25.505 5.18 ;
      RECT 24.445 9.345 24.82 9.715 ;
      RECT 24.225 4.81 24.505 5.18 ;
      RECT 16.425 3.69 16.705 4.06 ;
    LAYER via1 ;
      RECT 107.255 9.665 107.405 9.815 ;
      RECT 104.885 9.03 105.035 9.18 ;
      RECT 104.87 3.36 105.02 3.51 ;
      RECT 104.08 3.745 104.23 3.895 ;
      RECT 104.08 8.615 104.23 8.765 ;
      RECT 102.49 4.545 102.64 4.695 ;
      RECT 100.49 3.24 100.64 3.39 ;
      RECT 99.53 4.92 99.68 5.07 ;
      RECT 99.455 9 99.605 9.15 ;
      RECT 99.05 3.24 99.2 3.39 ;
      RECT 99.05 4.36 99.2 4.51 ;
      RECT 98.795 9.455 98.945 9.605 ;
      RECT 98.53 4.92 98.68 5.07 ;
      RECT 98.05 4.92 98.2 5.07 ;
      RECT 97.93 3.24 98.08 3.39 ;
      RECT 97.57 4.92 97.72 5.07 ;
      RECT 97.33 3.24 97.48 3.39 ;
      RECT 97.09 3.8 97.24 3.95 ;
      RECT 96.57 4.92 96.72 5.07 ;
      RECT 96.09 3.24 96.24 3.39 ;
      RECT 95.37 3.24 95.52 3.39 ;
      RECT 95.37 4.36 95.52 4.51 ;
      RECT 95.01 4.92 95.16 5.07 ;
      RECT 94.65 3.24 94.8 3.39 ;
      RECT 94.65 4.36 94.8 4.51 ;
      RECT 94.39 3.8 94.54 3.95 ;
      RECT 93.17 3.24 93.32 3.39 ;
      RECT 92.33 4.36 92.48 4.51 ;
      RECT 91.21 3.24 91.36 3.39 ;
      RECT 91.21 4.36 91.36 4.51 ;
      RECT 90.73 3.8 90.88 3.95 ;
      RECT 90.25 4.64 90.4 4.79 ;
      RECT 88.67 9.045 88.82 9.195 ;
      RECT 86.325 9.03 86.475 9.18 ;
      RECT 86.31 3.36 86.46 3.51 ;
      RECT 85.52 3.745 85.67 3.895 ;
      RECT 85.52 8.615 85.67 8.765 ;
      RECT 83.93 4.545 84.08 4.695 ;
      RECT 81.93 3.24 82.08 3.39 ;
      RECT 80.97 4.92 81.12 5.07 ;
      RECT 80.895 9 81.045 9.15 ;
      RECT 80.49 3.24 80.64 3.39 ;
      RECT 80.49 4.36 80.64 4.51 ;
      RECT 80.235 9.455 80.385 9.605 ;
      RECT 79.97 4.92 80.12 5.07 ;
      RECT 79.49 4.92 79.64 5.07 ;
      RECT 79.37 3.24 79.52 3.39 ;
      RECT 79.01 4.92 79.16 5.07 ;
      RECT 78.77 3.24 78.92 3.39 ;
      RECT 78.53 3.8 78.68 3.95 ;
      RECT 78.01 4.92 78.16 5.07 ;
      RECT 77.53 3.24 77.68 3.39 ;
      RECT 76.81 3.24 76.96 3.39 ;
      RECT 76.81 4.36 76.96 4.51 ;
      RECT 76.45 4.92 76.6 5.07 ;
      RECT 76.09 3.24 76.24 3.39 ;
      RECT 76.09 4.36 76.24 4.51 ;
      RECT 75.83 3.8 75.98 3.95 ;
      RECT 74.61 3.24 74.76 3.39 ;
      RECT 73.77 4.36 73.92 4.51 ;
      RECT 72.65 3.24 72.8 3.39 ;
      RECT 72.65 4.36 72.8 4.51 ;
      RECT 72.17 3.8 72.32 3.95 ;
      RECT 71.69 4.64 71.84 4.79 ;
      RECT 70.11 9.045 70.26 9.195 ;
      RECT 67.765 9.03 67.915 9.18 ;
      RECT 67.75 3.36 67.9 3.51 ;
      RECT 66.96 3.745 67.11 3.895 ;
      RECT 66.96 8.615 67.11 8.765 ;
      RECT 65.37 4.545 65.52 4.695 ;
      RECT 63.37 3.24 63.52 3.39 ;
      RECT 62.41 4.92 62.56 5.07 ;
      RECT 62.335 9.005 62.485 9.155 ;
      RECT 61.93 3.24 62.08 3.39 ;
      RECT 61.93 4.36 62.08 4.51 ;
      RECT 61.675 9.455 61.825 9.605 ;
      RECT 61.41 4.92 61.56 5.07 ;
      RECT 60.93 4.92 61.08 5.07 ;
      RECT 60.81 3.24 60.96 3.39 ;
      RECT 60.45 4.92 60.6 5.07 ;
      RECT 60.21 3.24 60.36 3.39 ;
      RECT 59.97 3.8 60.12 3.95 ;
      RECT 59.45 4.92 59.6 5.07 ;
      RECT 58.97 3.24 59.12 3.39 ;
      RECT 58.25 3.24 58.4 3.39 ;
      RECT 58.25 4.36 58.4 4.51 ;
      RECT 57.89 4.92 58.04 5.07 ;
      RECT 57.53 3.24 57.68 3.39 ;
      RECT 57.53 4.36 57.68 4.51 ;
      RECT 57.27 3.8 57.42 3.95 ;
      RECT 56.05 3.24 56.2 3.39 ;
      RECT 55.21 4.36 55.36 4.51 ;
      RECT 54.09 3.24 54.24 3.39 ;
      RECT 54.09 4.36 54.24 4.51 ;
      RECT 53.61 3.8 53.76 3.95 ;
      RECT 53.13 4.64 53.28 4.79 ;
      RECT 51.595 9.05 51.745 9.2 ;
      RECT 49.205 9.03 49.355 9.18 ;
      RECT 49.19 3.36 49.34 3.51 ;
      RECT 48.4 3.745 48.55 3.895 ;
      RECT 48.4 8.615 48.55 8.765 ;
      RECT 46.81 4.545 46.96 4.695 ;
      RECT 44.81 3.24 44.96 3.39 ;
      RECT 43.85 4.92 44 5.07 ;
      RECT 43.78 9 43.93 9.15 ;
      RECT 43.37 3.24 43.52 3.39 ;
      RECT 43.37 4.36 43.52 4.51 ;
      RECT 43.115 9.455 43.265 9.605 ;
      RECT 42.85 4.92 43 5.07 ;
      RECT 42.37 4.92 42.52 5.07 ;
      RECT 42.25 3.24 42.4 3.39 ;
      RECT 41.89 4.92 42.04 5.07 ;
      RECT 41.65 3.24 41.8 3.39 ;
      RECT 41.41 3.8 41.56 3.95 ;
      RECT 40.89 4.92 41.04 5.07 ;
      RECT 40.41 3.24 40.56 3.39 ;
      RECT 39.69 3.24 39.84 3.39 ;
      RECT 39.69 4.36 39.84 4.51 ;
      RECT 39.33 4.92 39.48 5.07 ;
      RECT 38.97 3.24 39.12 3.39 ;
      RECT 38.97 4.36 39.12 4.51 ;
      RECT 38.71 3.8 38.86 3.95 ;
      RECT 37.49 3.24 37.64 3.39 ;
      RECT 36.65 4.36 36.8 4.51 ;
      RECT 35.53 3.24 35.68 3.39 ;
      RECT 35.53 4.36 35.68 4.51 ;
      RECT 35.05 3.8 35.2 3.95 ;
      RECT 34.57 4.64 34.72 4.79 ;
      RECT 33.035 9.045 33.185 9.195 ;
      RECT 30.645 9.03 30.795 9.18 ;
      RECT 30.63 3.36 30.78 3.51 ;
      RECT 29.84 3.745 29.99 3.895 ;
      RECT 29.84 8.615 29.99 8.765 ;
      RECT 28.25 4.545 28.4 4.695 ;
      RECT 26.25 3.24 26.4 3.39 ;
      RECT 25.29 4.92 25.44 5.07 ;
      RECT 25.22 8.995 25.37 9.145 ;
      RECT 24.81 3.24 24.96 3.39 ;
      RECT 24.81 4.36 24.96 4.51 ;
      RECT 24.555 9.455 24.705 9.605 ;
      RECT 24.29 4.92 24.44 5.07 ;
      RECT 23.81 4.92 23.96 5.07 ;
      RECT 23.69 3.24 23.84 3.39 ;
      RECT 23.33 4.92 23.48 5.07 ;
      RECT 23.09 3.24 23.24 3.39 ;
      RECT 22.85 3.8 23 3.95 ;
      RECT 22.33 4.92 22.48 5.07 ;
      RECT 21.85 3.24 22 3.39 ;
      RECT 21.13 3.24 21.28 3.39 ;
      RECT 21.13 4.36 21.28 4.51 ;
      RECT 20.77 4.92 20.92 5.07 ;
      RECT 20.41 3.24 20.56 3.39 ;
      RECT 20.41 4.36 20.56 4.51 ;
      RECT 20.15 3.8 20.3 3.95 ;
      RECT 18.93 3.24 19.08 3.39 ;
      RECT 18.09 4.36 18.24 4.51 ;
      RECT 16.97 3.24 17.12 3.39 ;
      RECT 16.97 4.36 17.12 4.51 ;
      RECT 16.49 3.8 16.64 3.95 ;
      RECT 16.01 4.64 16.16 4.79 ;
      RECT 13.74 9.385 13.89 9.535 ;
      RECT 13.365 8.645 13.515 8.795 ;
    LAYER met1 ;
      RECT 12.13 5.44 107.625 7.04 ;
      RECT 89.91 5.43 107.725 7.035 ;
      RECT 71.35 5.43 89.165 7.04 ;
      RECT 52.79 5.43 70.605 7.04 ;
      RECT 34.23 5.43 52.045 7.04 ;
      RECT 15.67 5.43 33.485 7.04 ;
      RECT 105.59 5.425 107.57 7.04 ;
      RECT 89.91 5.275 101.87 7.04 ;
      RECT 87.03 5.425 89.01 7.04 ;
      RECT 71.35 5.275 83.31 7.04 ;
      RECT 68.47 5.425 70.45 7.04 ;
      RECT 52.79 5.275 64.75 7.04 ;
      RECT 49.91 5.425 51.89 7.04 ;
      RECT 34.23 5.275 46.19 7.04 ;
      RECT 31.35 5.425 33.33 7.04 ;
      RECT 15.67 5.275 27.63 7.04 ;
      RECT 107.12 10.06 107.41 10.29 ;
      RECT 107.18 8.58 107.35 10.29 ;
      RECT 107.155 9.565 107.505 9.915 ;
      RECT 107.12 8.58 107.41 8.81 ;
      RECT 106.715 3.69 106.82 4.26 ;
      RECT 106.715 4.025 107.04 4.255 ;
      RECT 106.715 4.055 107.21 4.225 ;
      RECT 106.715 3.69 106.905 4.255 ;
      RECT 106.13 3.655 106.42 3.885 ;
      RECT 106.13 3.69 106.905 3.86 ;
      RECT 106.19 2.175 106.36 3.885 ;
      RECT 106.13 2.175 106.42 2.405 ;
      RECT 106.13 10.06 106.42 10.29 ;
      RECT 106.19 8.58 106.36 10.29 ;
      RECT 106.13 8.58 106.42 8.81 ;
      RECT 106.13 8.615 106.985 8.775 ;
      RECT 106.815 8.21 106.985 8.775 ;
      RECT 106.13 8.61 106.525 8.775 ;
      RECT 106.75 8.21 107.04 8.44 ;
      RECT 106.75 8.24 107.21 8.41 ;
      RECT 105.76 4.025 106.05 4.255 ;
      RECT 105.76 4.055 106.22 4.225 ;
      RECT 105.825 2.95 105.99 4.255 ;
      RECT 104.34 2.92 104.63 3.15 ;
      RECT 104.34 2.95 105.99 3.12 ;
      RECT 104.4 2.18 104.57 3.15 ;
      RECT 104.34 2.18 104.63 2.41 ;
      RECT 104.34 10.055 104.63 10.285 ;
      RECT 104.4 9.315 104.57 10.285 ;
      RECT 104.4 9.41 105.99 9.58 ;
      RECT 105.82 8.21 105.99 9.58 ;
      RECT 104.34 9.315 104.63 9.545 ;
      RECT 105.76 8.21 106.05 8.44 ;
      RECT 105.76 8.24 106.22 8.41 ;
      RECT 102.39 4.445 102.73 4.795 ;
      RECT 102.48 3.32 102.65 4.795 ;
      RECT 104.77 3.26 105.12 3.61 ;
      RECT 102.48 3.32 105.12 3.49 ;
      RECT 104.795 8.945 105.12 9.27 ;
      RECT 99.355 8.9 99.705 9.25 ;
      RECT 104.77 8.945 105.12 9.175 ;
      RECT 99.155 8.945 99.705 9.175 ;
      RECT 98.985 8.975 105.12 9.145 ;
      RECT 103.995 3.66 104.315 3.98 ;
      RECT 103.965 3.66 104.315 3.89 ;
      RECT 103.795 3.69 104.315 3.86 ;
      RECT 103.995 8.545 104.315 8.835 ;
      RECT 103.965 8.575 104.315 8.805 ;
      RECT 103.795 8.605 104.315 8.775 ;
      RECT 99.445 4.865 99.765 5.125 ;
      RECT 100.735 4.04 100.875 4.9 ;
      RECT 99.535 4.76 100.875 4.9 ;
      RECT 99.535 4.32 99.675 5.125 ;
      RECT 99.46 4.32 99.75 4.55 ;
      RECT 100.66 4.04 100.95 4.27 ;
      RECT 100.18 4.32 100.47 4.55 ;
      RECT 100.375 3.245 100.515 4.505 ;
      RECT 100.405 3.185 100.725 3.445 ;
      RECT 97.005 3.745 97.325 4.005 ;
      RECT 99.7 3.76 99.99 3.99 ;
      RECT 97.095 3.665 99.915 3.805 ;
      RECT 98.965 3.185 99.285 3.445 ;
      RECT 99.46 3.2 99.75 3.43 ;
      RECT 98.965 3.245 99.75 3.385 ;
      RECT 98.965 4.305 99.285 4.565 ;
      RECT 98.965 4.085 99.195 4.565 ;
      RECT 98.46 4.04 98.75 4.27 ;
      RECT 98.46 4.085 99.195 4.225 ;
      RECT 98.725 10.055 99.015 10.285 ;
      RECT 98.785 9.315 98.955 10.285 ;
      RECT 98.685 9.345 99.065 9.715 ;
      RECT 98.725 9.315 99.015 9.715 ;
      RECT 97.485 4.865 97.805 5.125 ;
      RECT 97.02 4.88 97.31 5.11 ;
      RECT 97.02 4.925 97.805 5.065 ;
      RECT 95.78 3.76 96.07 3.99 ;
      RECT 95.78 3.805 96.715 3.945 ;
      RECT 96.575 3.245 96.715 3.945 ;
      RECT 97.245 3.185 97.565 3.445 ;
      RECT 97.02 3.2 97.565 3.43 ;
      RECT 96.575 3.245 97.565 3.385 ;
      RECT 94.925 4.865 95.245 5.125 ;
      RECT 94.925 4.925 95.995 5.065 ;
      RECT 95.855 4.365 95.995 5.065 ;
      RECT 97.02 4.32 97.31 4.55 ;
      RECT 95.855 4.365 97.31 4.505 ;
      RECT 95.285 3.185 95.605 3.445 ;
      RECT 95.06 3.2 95.605 3.43 ;
      RECT 94.305 3.745 94.625 4.005 ;
      RECT 95.3 3.76 95.59 3.99 ;
      RECT 94.06 3.76 94.625 3.99 ;
      RECT 94.06 3.805 95.59 3.945 ;
      RECT 93.58 4.32 93.87 4.55 ;
      RECT 93.775 3.245 93.915 4.505 ;
      RECT 94.565 3.185 94.885 3.445 ;
      RECT 93.58 3.2 93.87 3.43 ;
      RECT 93.58 3.245 94.885 3.385 ;
      RECT 93.175 4.76 94.275 4.9 ;
      RECT 94.06 4.6 94.35 4.83 ;
      RECT 93.1 4.6 93.39 4.83 ;
      RECT 93.085 3.185 93.405 3.445 ;
      RECT 91.125 3.185 91.445 3.445 ;
      RECT 91.125 3.245 93.405 3.385 ;
      RECT 92.245 4.305 92.565 4.565 ;
      RECT 92.245 4.305 93.075 4.445 ;
      RECT 92.86 4.04 93.075 4.445 ;
      RECT 92.86 4.04 93.15 4.27 ;
      RECT 90.645 3.745 90.965 4.005 ;
      RECT 92.055 3.76 92.345 3.99 ;
      RECT 90.645 3.76 91.19 3.99 ;
      RECT 90.645 3.845 91.595 3.985 ;
      RECT 91.455 3.665 91.595 3.985 ;
      RECT 91.955 3.76 92.345 3.945 ;
      RECT 91.455 3.665 92.095 3.805 ;
      RECT 90.165 4.555 90.485 4.97 ;
      RECT 90.245 3.2 90.4 4.97 ;
      RECT 90.18 3.2 90.47 3.43 ;
      RECT 88.56 10.06 88.85 10.29 ;
      RECT 88.62 8.58 88.79 10.29 ;
      RECT 88.57 8.945 88.92 9.295 ;
      RECT 88.56 8.58 88.85 8.81 ;
      RECT 88.155 3.69 88.26 4.26 ;
      RECT 88.155 4.025 88.48 4.255 ;
      RECT 88.155 4.055 88.65 4.225 ;
      RECT 88.155 3.69 88.345 4.255 ;
      RECT 87.57 3.655 87.86 3.885 ;
      RECT 87.57 3.69 88.345 3.86 ;
      RECT 87.63 2.175 87.8 3.885 ;
      RECT 87.57 2.175 87.86 2.405 ;
      RECT 87.57 10.06 87.86 10.29 ;
      RECT 87.63 8.58 87.8 10.29 ;
      RECT 87.57 8.58 87.86 8.81 ;
      RECT 87.57 8.615 88.425 8.775 ;
      RECT 88.255 8.21 88.425 8.775 ;
      RECT 87.57 8.61 87.965 8.775 ;
      RECT 88.19 8.21 88.48 8.44 ;
      RECT 88.19 8.24 88.65 8.41 ;
      RECT 87.2 4.025 87.49 4.255 ;
      RECT 87.2 4.055 87.66 4.225 ;
      RECT 87.265 2.95 87.43 4.255 ;
      RECT 85.78 2.92 86.07 3.15 ;
      RECT 85.78 2.95 87.43 3.12 ;
      RECT 85.84 2.18 86.01 3.15 ;
      RECT 85.78 2.18 86.07 2.41 ;
      RECT 85.78 10.055 86.07 10.285 ;
      RECT 85.84 9.315 86.01 10.285 ;
      RECT 85.84 9.41 87.43 9.58 ;
      RECT 87.26 8.21 87.43 9.58 ;
      RECT 85.78 9.315 86.07 9.545 ;
      RECT 87.2 8.21 87.49 8.44 ;
      RECT 87.2 8.24 87.66 8.41 ;
      RECT 83.83 4.445 84.17 4.795 ;
      RECT 83.92 3.32 84.09 4.795 ;
      RECT 86.21 3.26 86.56 3.61 ;
      RECT 83.92 3.32 86.56 3.49 ;
      RECT 86.235 8.945 86.56 9.27 ;
      RECT 80.795 8.9 81.145 9.25 ;
      RECT 86.21 8.945 86.56 9.175 ;
      RECT 80.595 8.945 81.145 9.175 ;
      RECT 80.425 8.975 86.56 9.145 ;
      RECT 85.435 3.66 85.755 3.98 ;
      RECT 85.405 3.66 85.755 3.89 ;
      RECT 85.235 3.69 85.755 3.86 ;
      RECT 85.435 8.545 85.755 8.835 ;
      RECT 85.405 8.575 85.755 8.805 ;
      RECT 85.235 8.605 85.755 8.775 ;
      RECT 80.885 4.865 81.205 5.125 ;
      RECT 82.175 4.04 82.315 4.9 ;
      RECT 80.975 4.76 82.315 4.9 ;
      RECT 80.975 4.32 81.115 5.125 ;
      RECT 80.9 4.32 81.19 4.55 ;
      RECT 82.1 4.04 82.39 4.27 ;
      RECT 81.62 4.32 81.91 4.55 ;
      RECT 81.815 3.245 81.955 4.505 ;
      RECT 81.845 3.185 82.165 3.445 ;
      RECT 78.445 3.745 78.765 4.005 ;
      RECT 81.14 3.76 81.43 3.99 ;
      RECT 78.535 3.665 81.355 3.805 ;
      RECT 80.405 3.185 80.725 3.445 ;
      RECT 80.9 3.2 81.19 3.43 ;
      RECT 80.405 3.245 81.19 3.385 ;
      RECT 80.405 4.305 80.725 4.565 ;
      RECT 80.405 4.085 80.635 4.565 ;
      RECT 79.9 4.04 80.19 4.27 ;
      RECT 79.9 4.085 80.635 4.225 ;
      RECT 80.165 10.055 80.455 10.285 ;
      RECT 80.225 9.315 80.395 10.285 ;
      RECT 80.125 9.345 80.505 9.715 ;
      RECT 80.165 9.315 80.455 9.715 ;
      RECT 78.925 4.865 79.245 5.125 ;
      RECT 78.46 4.88 78.75 5.11 ;
      RECT 78.46 4.925 79.245 5.065 ;
      RECT 77.22 3.76 77.51 3.99 ;
      RECT 77.22 3.805 78.155 3.945 ;
      RECT 78.015 3.245 78.155 3.945 ;
      RECT 78.685 3.185 79.005 3.445 ;
      RECT 78.46 3.2 79.005 3.43 ;
      RECT 78.015 3.245 79.005 3.385 ;
      RECT 76.365 4.865 76.685 5.125 ;
      RECT 76.365 4.925 77.435 5.065 ;
      RECT 77.295 4.365 77.435 5.065 ;
      RECT 78.46 4.32 78.75 4.55 ;
      RECT 77.295 4.365 78.75 4.505 ;
      RECT 76.725 3.185 77.045 3.445 ;
      RECT 76.5 3.2 77.045 3.43 ;
      RECT 75.745 3.745 76.065 4.005 ;
      RECT 76.74 3.76 77.03 3.99 ;
      RECT 75.5 3.76 76.065 3.99 ;
      RECT 75.5 3.805 77.03 3.945 ;
      RECT 75.02 4.32 75.31 4.55 ;
      RECT 75.215 3.245 75.355 4.505 ;
      RECT 76.005 3.185 76.325 3.445 ;
      RECT 75.02 3.2 75.31 3.43 ;
      RECT 75.02 3.245 76.325 3.385 ;
      RECT 74.615 4.76 75.715 4.9 ;
      RECT 75.5 4.6 75.79 4.83 ;
      RECT 74.54 4.6 74.83 4.83 ;
      RECT 74.525 3.185 74.845 3.445 ;
      RECT 72.565 3.185 72.885 3.445 ;
      RECT 72.565 3.245 74.845 3.385 ;
      RECT 73.685 4.305 74.005 4.565 ;
      RECT 73.685 4.305 74.515 4.445 ;
      RECT 74.3 4.04 74.515 4.445 ;
      RECT 74.3 4.04 74.59 4.27 ;
      RECT 72.085 3.745 72.405 4.005 ;
      RECT 73.495 3.76 73.785 3.99 ;
      RECT 72.085 3.76 72.63 3.99 ;
      RECT 72.085 3.845 73.035 3.985 ;
      RECT 72.895 3.665 73.035 3.985 ;
      RECT 73.395 3.76 73.785 3.945 ;
      RECT 72.895 3.665 73.535 3.805 ;
      RECT 71.605 4.555 71.925 4.97 ;
      RECT 71.685 3.2 71.84 4.97 ;
      RECT 71.62 3.2 71.91 3.43 ;
      RECT 70 10.06 70.29 10.29 ;
      RECT 70.06 8.58 70.23 10.29 ;
      RECT 70.01 8.945 70.36 9.295 ;
      RECT 70 8.58 70.29 8.81 ;
      RECT 69.595 3.69 69.7 4.26 ;
      RECT 69.595 4.025 69.92 4.255 ;
      RECT 69.595 4.055 70.09 4.225 ;
      RECT 69.595 3.69 69.785 4.255 ;
      RECT 69.01 3.655 69.3 3.885 ;
      RECT 69.01 3.69 69.785 3.86 ;
      RECT 69.07 2.175 69.24 3.885 ;
      RECT 69.01 2.175 69.3 2.405 ;
      RECT 69.01 10.06 69.3 10.29 ;
      RECT 69.07 8.58 69.24 10.29 ;
      RECT 69.01 8.58 69.3 8.81 ;
      RECT 69.01 8.615 69.865 8.775 ;
      RECT 69.695 8.21 69.865 8.775 ;
      RECT 69.01 8.61 69.405 8.775 ;
      RECT 69.63 8.21 69.92 8.44 ;
      RECT 69.63 8.24 70.09 8.41 ;
      RECT 68.64 4.025 68.93 4.255 ;
      RECT 68.64 4.055 69.1 4.225 ;
      RECT 68.705 2.95 68.87 4.255 ;
      RECT 67.22 2.92 67.51 3.15 ;
      RECT 67.22 2.95 68.87 3.12 ;
      RECT 67.28 2.18 67.45 3.15 ;
      RECT 67.22 2.18 67.51 2.41 ;
      RECT 67.22 10.055 67.51 10.285 ;
      RECT 67.28 9.315 67.45 10.285 ;
      RECT 67.28 9.41 68.87 9.58 ;
      RECT 68.7 8.21 68.87 9.58 ;
      RECT 67.22 9.315 67.51 9.545 ;
      RECT 68.64 8.21 68.93 8.44 ;
      RECT 68.64 8.24 69.1 8.41 ;
      RECT 65.27 4.445 65.61 4.795 ;
      RECT 65.36 3.32 65.53 4.795 ;
      RECT 67.65 3.26 68 3.61 ;
      RECT 65.36 3.32 68 3.49 ;
      RECT 67.675 8.945 68 9.27 ;
      RECT 62.235 8.905 62.585 9.255 ;
      RECT 67.65 8.945 68 9.175 ;
      RECT 62.035 8.945 62.585 9.175 ;
      RECT 61.865 8.975 68 9.145 ;
      RECT 66.875 3.66 67.195 3.98 ;
      RECT 66.845 3.66 67.195 3.89 ;
      RECT 66.675 3.69 67.195 3.86 ;
      RECT 66.875 8.545 67.195 8.835 ;
      RECT 66.845 8.575 67.195 8.805 ;
      RECT 66.675 8.605 67.195 8.775 ;
      RECT 62.325 4.865 62.645 5.125 ;
      RECT 63.615 4.04 63.755 4.9 ;
      RECT 62.415 4.76 63.755 4.9 ;
      RECT 62.415 4.32 62.555 5.125 ;
      RECT 62.34 4.32 62.63 4.55 ;
      RECT 63.54 4.04 63.83 4.27 ;
      RECT 63.06 4.32 63.35 4.55 ;
      RECT 63.255 3.245 63.395 4.505 ;
      RECT 63.285 3.185 63.605 3.445 ;
      RECT 59.885 3.745 60.205 4.005 ;
      RECT 62.58 3.76 62.87 3.99 ;
      RECT 59.975 3.665 62.795 3.805 ;
      RECT 61.845 3.185 62.165 3.445 ;
      RECT 62.34 3.2 62.63 3.43 ;
      RECT 61.845 3.245 62.63 3.385 ;
      RECT 61.845 4.305 62.165 4.565 ;
      RECT 61.845 4.085 62.075 4.565 ;
      RECT 61.34 4.04 61.63 4.27 ;
      RECT 61.34 4.085 62.075 4.225 ;
      RECT 61.605 10.055 61.895 10.285 ;
      RECT 61.665 9.315 61.835 10.285 ;
      RECT 61.565 9.345 61.945 9.715 ;
      RECT 61.605 9.315 61.895 9.715 ;
      RECT 60.365 4.865 60.685 5.125 ;
      RECT 59.9 4.88 60.19 5.11 ;
      RECT 59.9 4.925 60.685 5.065 ;
      RECT 58.66 3.76 58.95 3.99 ;
      RECT 58.66 3.805 59.595 3.945 ;
      RECT 59.455 3.245 59.595 3.945 ;
      RECT 60.125 3.185 60.445 3.445 ;
      RECT 59.9 3.2 60.445 3.43 ;
      RECT 59.455 3.245 60.445 3.385 ;
      RECT 57.805 4.865 58.125 5.125 ;
      RECT 57.805 4.925 58.875 5.065 ;
      RECT 58.735 4.365 58.875 5.065 ;
      RECT 59.9 4.32 60.19 4.55 ;
      RECT 58.735 4.365 60.19 4.505 ;
      RECT 58.165 3.185 58.485 3.445 ;
      RECT 57.94 3.2 58.485 3.43 ;
      RECT 57.185 3.745 57.505 4.005 ;
      RECT 58.18 3.76 58.47 3.99 ;
      RECT 56.94 3.76 57.505 3.99 ;
      RECT 56.94 3.805 58.47 3.945 ;
      RECT 56.46 4.32 56.75 4.55 ;
      RECT 56.655 3.245 56.795 4.505 ;
      RECT 57.445 3.185 57.765 3.445 ;
      RECT 56.46 3.2 56.75 3.43 ;
      RECT 56.46 3.245 57.765 3.385 ;
      RECT 56.055 4.76 57.155 4.9 ;
      RECT 56.94 4.6 57.23 4.83 ;
      RECT 55.98 4.6 56.27 4.83 ;
      RECT 55.965 3.185 56.285 3.445 ;
      RECT 54.005 3.185 54.325 3.445 ;
      RECT 54.005 3.245 56.285 3.385 ;
      RECT 55.125 4.305 55.445 4.565 ;
      RECT 55.125 4.305 55.955 4.445 ;
      RECT 55.74 4.04 55.955 4.445 ;
      RECT 55.74 4.04 56.03 4.27 ;
      RECT 53.525 3.745 53.845 4.005 ;
      RECT 54.935 3.76 55.225 3.99 ;
      RECT 53.525 3.76 54.07 3.99 ;
      RECT 53.525 3.845 54.475 3.985 ;
      RECT 54.335 3.665 54.475 3.985 ;
      RECT 54.835 3.76 55.225 3.945 ;
      RECT 54.335 3.665 54.975 3.805 ;
      RECT 53.045 4.555 53.365 4.97 ;
      RECT 53.125 3.2 53.28 4.97 ;
      RECT 53.06 3.2 53.35 3.43 ;
      RECT 51.44 10.06 51.73 10.29 ;
      RECT 51.5 8.58 51.67 10.29 ;
      RECT 51.49 8.95 51.845 9.305 ;
      RECT 51.44 8.58 51.73 8.81 ;
      RECT 51.035 3.69 51.14 4.26 ;
      RECT 51.035 4.025 51.36 4.255 ;
      RECT 51.035 4.055 51.53 4.225 ;
      RECT 51.035 3.69 51.225 4.255 ;
      RECT 50.45 3.655 50.74 3.885 ;
      RECT 50.45 3.69 51.225 3.86 ;
      RECT 50.51 2.175 50.68 3.885 ;
      RECT 50.45 2.175 50.74 2.405 ;
      RECT 50.45 10.06 50.74 10.29 ;
      RECT 50.51 8.58 50.68 10.29 ;
      RECT 50.45 8.58 50.74 8.81 ;
      RECT 50.45 8.615 51.305 8.775 ;
      RECT 51.135 8.21 51.305 8.775 ;
      RECT 50.45 8.61 50.845 8.775 ;
      RECT 51.07 8.21 51.36 8.44 ;
      RECT 51.07 8.24 51.53 8.41 ;
      RECT 50.08 4.025 50.37 4.255 ;
      RECT 50.08 4.055 50.54 4.225 ;
      RECT 50.145 2.95 50.31 4.255 ;
      RECT 48.66 2.92 48.95 3.15 ;
      RECT 48.66 2.95 50.31 3.12 ;
      RECT 48.72 2.18 48.89 3.15 ;
      RECT 48.66 2.18 48.95 2.41 ;
      RECT 48.66 10.055 48.95 10.285 ;
      RECT 48.72 9.315 48.89 10.285 ;
      RECT 48.72 9.41 50.31 9.58 ;
      RECT 50.14 8.21 50.31 9.58 ;
      RECT 48.66 9.315 48.95 9.545 ;
      RECT 50.08 8.21 50.37 8.44 ;
      RECT 50.08 8.24 50.54 8.41 ;
      RECT 46.71 4.445 47.05 4.795 ;
      RECT 46.8 3.32 46.97 4.795 ;
      RECT 49.09 3.26 49.44 3.61 ;
      RECT 46.8 3.32 49.44 3.49 ;
      RECT 49.115 8.945 49.44 9.27 ;
      RECT 43.68 8.9 44.03 9.25 ;
      RECT 49.09 8.945 49.44 9.175 ;
      RECT 43.475 8.945 44.03 9.175 ;
      RECT 43.305 8.975 49.44 9.145 ;
      RECT 48.315 3.66 48.635 3.98 ;
      RECT 48.285 3.66 48.635 3.89 ;
      RECT 48.115 3.69 48.635 3.86 ;
      RECT 48.315 8.545 48.635 8.835 ;
      RECT 48.285 8.575 48.635 8.805 ;
      RECT 48.115 8.605 48.635 8.775 ;
      RECT 43.765 4.865 44.085 5.125 ;
      RECT 45.055 4.04 45.195 4.9 ;
      RECT 43.855 4.76 45.195 4.9 ;
      RECT 43.855 4.32 43.995 5.125 ;
      RECT 43.78 4.32 44.07 4.55 ;
      RECT 44.98 4.04 45.27 4.27 ;
      RECT 44.5 4.32 44.79 4.55 ;
      RECT 44.695 3.245 44.835 4.505 ;
      RECT 44.725 3.185 45.045 3.445 ;
      RECT 41.325 3.745 41.645 4.005 ;
      RECT 44.02 3.76 44.31 3.99 ;
      RECT 41.415 3.665 44.235 3.805 ;
      RECT 43.285 3.185 43.605 3.445 ;
      RECT 43.78 3.2 44.07 3.43 ;
      RECT 43.285 3.245 44.07 3.385 ;
      RECT 43.285 4.305 43.605 4.565 ;
      RECT 43.285 4.085 43.515 4.565 ;
      RECT 42.78 4.04 43.07 4.27 ;
      RECT 42.78 4.085 43.515 4.225 ;
      RECT 43.045 10.055 43.335 10.285 ;
      RECT 43.105 9.315 43.275 10.285 ;
      RECT 43.005 9.345 43.385 9.715 ;
      RECT 43.045 9.315 43.335 9.715 ;
      RECT 41.805 4.865 42.125 5.125 ;
      RECT 41.34 4.88 41.63 5.11 ;
      RECT 41.34 4.925 42.125 5.065 ;
      RECT 40.1 3.76 40.39 3.99 ;
      RECT 40.1 3.805 41.035 3.945 ;
      RECT 40.895 3.245 41.035 3.945 ;
      RECT 41.565 3.185 41.885 3.445 ;
      RECT 41.34 3.2 41.885 3.43 ;
      RECT 40.895 3.245 41.885 3.385 ;
      RECT 39.245 4.865 39.565 5.125 ;
      RECT 39.245 4.925 40.315 5.065 ;
      RECT 40.175 4.365 40.315 5.065 ;
      RECT 41.34 4.32 41.63 4.55 ;
      RECT 40.175 4.365 41.63 4.505 ;
      RECT 39.605 3.185 39.925 3.445 ;
      RECT 39.38 3.2 39.925 3.43 ;
      RECT 38.625 3.745 38.945 4.005 ;
      RECT 39.62 3.76 39.91 3.99 ;
      RECT 38.38 3.76 38.945 3.99 ;
      RECT 38.38 3.805 39.91 3.945 ;
      RECT 37.9 4.32 38.19 4.55 ;
      RECT 38.095 3.245 38.235 4.505 ;
      RECT 38.885 3.185 39.205 3.445 ;
      RECT 37.9 3.2 38.19 3.43 ;
      RECT 37.9 3.245 39.205 3.385 ;
      RECT 37.495 4.76 38.595 4.9 ;
      RECT 38.38 4.6 38.67 4.83 ;
      RECT 37.42 4.6 37.71 4.83 ;
      RECT 37.405 3.185 37.725 3.445 ;
      RECT 35.445 3.185 35.765 3.445 ;
      RECT 35.445 3.245 37.725 3.385 ;
      RECT 36.565 4.305 36.885 4.565 ;
      RECT 36.565 4.305 37.395 4.445 ;
      RECT 37.18 4.04 37.395 4.445 ;
      RECT 37.18 4.04 37.47 4.27 ;
      RECT 34.965 3.745 35.285 4.005 ;
      RECT 36.375 3.76 36.665 3.99 ;
      RECT 34.965 3.76 35.51 3.99 ;
      RECT 34.965 3.845 35.915 3.985 ;
      RECT 35.775 3.665 35.915 3.985 ;
      RECT 36.275 3.76 36.665 3.945 ;
      RECT 35.775 3.665 36.415 3.805 ;
      RECT 34.485 4.555 34.805 4.97 ;
      RECT 34.565 3.2 34.72 4.97 ;
      RECT 34.5 3.2 34.79 3.43 ;
      RECT 32.88 10.06 33.17 10.29 ;
      RECT 32.94 8.58 33.11 10.29 ;
      RECT 32.935 8.945 33.285 9.295 ;
      RECT 32.88 8.58 33.17 8.81 ;
      RECT 32.475 3.69 32.58 4.26 ;
      RECT 32.475 4.025 32.8 4.255 ;
      RECT 32.475 4.055 32.97 4.225 ;
      RECT 32.475 3.69 32.665 4.255 ;
      RECT 31.89 3.655 32.18 3.885 ;
      RECT 31.89 3.69 32.665 3.86 ;
      RECT 31.95 2.175 32.12 3.885 ;
      RECT 31.89 2.175 32.18 2.405 ;
      RECT 31.89 10.06 32.18 10.29 ;
      RECT 31.95 8.58 32.12 10.29 ;
      RECT 31.89 8.58 32.18 8.81 ;
      RECT 31.89 8.615 32.745 8.775 ;
      RECT 32.575 8.21 32.745 8.775 ;
      RECT 31.89 8.61 32.285 8.775 ;
      RECT 32.51 8.21 32.8 8.44 ;
      RECT 32.51 8.24 32.97 8.41 ;
      RECT 31.52 4.025 31.81 4.255 ;
      RECT 31.52 4.055 31.98 4.225 ;
      RECT 31.585 2.95 31.75 4.255 ;
      RECT 30.1 2.92 30.39 3.15 ;
      RECT 30.1 2.95 31.75 3.12 ;
      RECT 30.16 2.18 30.33 3.15 ;
      RECT 30.1 2.18 30.39 2.41 ;
      RECT 30.1 10.055 30.39 10.285 ;
      RECT 30.16 9.315 30.33 10.285 ;
      RECT 30.16 9.41 31.75 9.58 ;
      RECT 31.58 8.21 31.75 9.58 ;
      RECT 30.1 9.315 30.39 9.545 ;
      RECT 31.52 8.21 31.81 8.44 ;
      RECT 31.52 8.24 31.98 8.41 ;
      RECT 28.15 4.445 28.49 4.795 ;
      RECT 28.24 3.32 28.41 4.795 ;
      RECT 30.53 3.26 30.88 3.61 ;
      RECT 28.24 3.32 30.88 3.49 ;
      RECT 30.555 8.945 30.88 9.27 ;
      RECT 25.12 8.895 25.47 9.245 ;
      RECT 30.53 8.945 30.88 9.175 ;
      RECT 24.915 8.945 25.47 9.175 ;
      RECT 24.745 8.975 30.88 9.145 ;
      RECT 29.755 3.66 30.075 3.98 ;
      RECT 29.725 3.66 30.075 3.89 ;
      RECT 29.555 3.69 30.075 3.86 ;
      RECT 29.755 8.545 30.075 8.835 ;
      RECT 29.725 8.575 30.075 8.805 ;
      RECT 29.555 8.605 30.075 8.775 ;
      RECT 25.205 4.865 25.525 5.125 ;
      RECT 26.495 4.04 26.635 4.9 ;
      RECT 25.295 4.76 26.635 4.9 ;
      RECT 25.295 4.32 25.435 5.125 ;
      RECT 25.22 4.32 25.51 4.55 ;
      RECT 26.42 4.04 26.71 4.27 ;
      RECT 25.94 4.32 26.23 4.55 ;
      RECT 26.135 3.245 26.275 4.505 ;
      RECT 26.165 3.185 26.485 3.445 ;
      RECT 22.765 3.745 23.085 4.005 ;
      RECT 25.46 3.76 25.75 3.99 ;
      RECT 22.855 3.665 25.675 3.805 ;
      RECT 24.725 3.185 25.045 3.445 ;
      RECT 25.22 3.2 25.51 3.43 ;
      RECT 24.725 3.245 25.51 3.385 ;
      RECT 24.725 4.305 25.045 4.565 ;
      RECT 24.725 4.085 24.955 4.565 ;
      RECT 24.22 4.04 24.51 4.27 ;
      RECT 24.22 4.085 24.955 4.225 ;
      RECT 24.485 10.055 24.775 10.285 ;
      RECT 24.545 9.315 24.715 10.285 ;
      RECT 24.445 9.345 24.825 9.715 ;
      RECT 24.485 9.315 24.775 9.715 ;
      RECT 23.245 4.865 23.565 5.125 ;
      RECT 22.78 4.88 23.07 5.11 ;
      RECT 22.78 4.925 23.565 5.065 ;
      RECT 21.54 3.76 21.83 3.99 ;
      RECT 21.54 3.805 22.475 3.945 ;
      RECT 22.335 3.245 22.475 3.945 ;
      RECT 23.005 3.185 23.325 3.445 ;
      RECT 22.78 3.2 23.325 3.43 ;
      RECT 22.335 3.245 23.325 3.385 ;
      RECT 20.685 4.865 21.005 5.125 ;
      RECT 20.685 4.925 21.755 5.065 ;
      RECT 21.615 4.365 21.755 5.065 ;
      RECT 22.78 4.32 23.07 4.55 ;
      RECT 21.615 4.365 23.07 4.505 ;
      RECT 21.045 3.185 21.365 3.445 ;
      RECT 20.82 3.2 21.365 3.43 ;
      RECT 20.065 3.745 20.385 4.005 ;
      RECT 21.06 3.76 21.35 3.99 ;
      RECT 19.82 3.76 20.385 3.99 ;
      RECT 19.82 3.805 21.35 3.945 ;
      RECT 19.34 4.32 19.63 4.55 ;
      RECT 19.535 3.245 19.675 4.505 ;
      RECT 20.325 3.185 20.645 3.445 ;
      RECT 19.34 3.2 19.63 3.43 ;
      RECT 19.34 3.245 20.645 3.385 ;
      RECT 18.935 4.76 20.035 4.9 ;
      RECT 19.82 4.6 20.11 4.83 ;
      RECT 18.86 4.6 19.15 4.83 ;
      RECT 18.845 3.185 19.165 3.445 ;
      RECT 16.885 3.185 17.205 3.445 ;
      RECT 16.885 3.245 19.165 3.385 ;
      RECT 18.005 4.305 18.325 4.565 ;
      RECT 18.005 4.305 18.835 4.445 ;
      RECT 18.62 4.04 18.835 4.445 ;
      RECT 18.62 4.04 18.91 4.27 ;
      RECT 16.405 3.745 16.725 4.005 ;
      RECT 17.815 3.76 18.105 3.99 ;
      RECT 16.405 3.76 16.95 3.99 ;
      RECT 16.405 3.845 17.355 3.985 ;
      RECT 17.215 3.665 17.355 3.985 ;
      RECT 17.715 3.76 18.105 3.945 ;
      RECT 17.215 3.665 17.855 3.805 ;
      RECT 15.925 4.555 16.245 4.97 ;
      RECT 16.005 3.2 16.16 4.97 ;
      RECT 15.94 3.2 16.23 3.43 ;
      RECT 14.1 8.945 14.39 9.175 ;
      RECT 13.93 8.975 14.39 9.145 ;
      RECT 13.67 10.055 13.96 10.285 ;
      RECT 13.73 9.315 13.9 10.285 ;
      RECT 13.64 9.315 13.99 9.605 ;
      RECT 13.265 8.575 13.615 8.865 ;
      RECT 13.125 8.605 13.615 8.775 ;
      RECT 98.445 4.865 98.765 5.125 ;
      RECT 97.845 3.185 98.525 3.445 ;
      RECT 97.965 4.865 98.285 5.125 ;
      RECT 96.485 4.865 96.805 5.125 ;
      RECT 96.005 3.185 96.325 3.445 ;
      RECT 95.285 4.305 95.605 4.565 ;
      RECT 94.565 4.305 94.885 4.565 ;
      RECT 91.125 4.305 91.445 4.565 ;
      RECT 79.885 4.865 80.205 5.125 ;
      RECT 79.285 3.185 79.965 3.445 ;
      RECT 79.405 4.865 79.725 5.125 ;
      RECT 77.925 4.865 78.245 5.125 ;
      RECT 77.445 3.185 77.765 3.445 ;
      RECT 76.725 4.305 77.045 4.565 ;
      RECT 76.005 4.305 76.325 4.565 ;
      RECT 72.565 4.305 72.885 4.565 ;
      RECT 61.325 4.865 61.645 5.125 ;
      RECT 60.725 3.185 61.405 3.445 ;
      RECT 60.845 4.865 61.165 5.125 ;
      RECT 59.365 4.865 59.685 5.125 ;
      RECT 58.885 3.185 59.205 3.445 ;
      RECT 58.165 4.305 58.485 4.565 ;
      RECT 57.445 4.305 57.765 4.565 ;
      RECT 54.005 4.305 54.325 4.565 ;
      RECT 42.765 4.865 43.085 5.125 ;
      RECT 42.165 3.185 42.845 3.445 ;
      RECT 42.285 4.865 42.605 5.125 ;
      RECT 40.805 4.865 41.125 5.125 ;
      RECT 40.325 3.185 40.645 3.445 ;
      RECT 39.605 4.305 39.925 4.565 ;
      RECT 38.885 4.305 39.205 4.565 ;
      RECT 35.445 4.305 35.765 4.565 ;
      RECT 24.205 4.865 24.525 5.125 ;
      RECT 23.605 3.185 24.285 3.445 ;
      RECT 23.725 4.865 24.045 5.125 ;
      RECT 22.245 4.865 22.565 5.125 ;
      RECT 21.765 3.185 22.085 3.445 ;
      RECT 21.045 4.305 21.365 4.565 ;
      RECT 20.325 4.305 20.645 4.565 ;
      RECT 16.885 4.305 17.205 4.565 ;
    LAYER mcon ;
      RECT 107.18 8.61 107.35 8.78 ;
      RECT 107.185 8.605 107.355 8.775 ;
      RECT 88.62 8.61 88.79 8.78 ;
      RECT 88.625 8.605 88.795 8.775 ;
      RECT 70.06 8.61 70.23 8.78 ;
      RECT 70.065 8.605 70.235 8.775 ;
      RECT 51.5 8.61 51.67 8.78 ;
      RECT 51.505 8.605 51.675 8.775 ;
      RECT 32.94 8.61 33.11 8.78 ;
      RECT 32.945 8.605 33.115 8.775 ;
      RECT 107.18 10.09 107.35 10.26 ;
      RECT 106.83 5.455 107 5.625 ;
      RECT 106.83 6.84 107 7.01 ;
      RECT 106.81 4.055 106.98 4.225 ;
      RECT 106.81 8.24 106.98 8.41 ;
      RECT 106.19 2.205 106.36 2.375 ;
      RECT 106.19 3.685 106.36 3.855 ;
      RECT 106.19 8.61 106.36 8.78 ;
      RECT 106.19 10.09 106.36 10.26 ;
      RECT 105.84 5.455 106.01 5.625 ;
      RECT 105.84 6.84 106.01 7.01 ;
      RECT 105.82 4.055 105.99 4.225 ;
      RECT 105.82 8.24 105.99 8.41 ;
      RECT 105.14 5.46 105.31 5.63 ;
      RECT 105.14 6.835 105.31 7.005 ;
      RECT 104.83 3.32 105 3.49 ;
      RECT 104.83 8.975 105 9.145 ;
      RECT 104.4 2.21 104.57 2.38 ;
      RECT 104.4 2.95 104.57 3.12 ;
      RECT 104.4 9.345 104.57 9.515 ;
      RECT 104.4 10.085 104.57 10.255 ;
      RECT 104.025 3.69 104.195 3.86 ;
      RECT 104.025 8.605 104.195 8.775 ;
      RECT 101.555 5.43 101.725 5.6 ;
      RECT 101.095 5.43 101.265 5.6 ;
      RECT 100.72 4.07 100.89 4.24 ;
      RECT 100.635 5.43 100.805 5.6 ;
      RECT 100.48 3.23 100.65 3.4 ;
      RECT 100.24 4.35 100.41 4.52 ;
      RECT 100.175 5.43 100.345 5.6 ;
      RECT 99.76 3.79 99.93 3.96 ;
      RECT 99.715 5.43 99.885 5.6 ;
      RECT 99.525 6.835 99.695 7.005 ;
      RECT 99.52 3.23 99.69 3.4 ;
      RECT 99.52 4.35 99.69 4.52 ;
      RECT 99.52 4.91 99.69 5.08 ;
      RECT 99.255 5.43 99.425 5.6 ;
      RECT 99.215 8.975 99.385 9.145 ;
      RECT 99.04 4.35 99.21 4.52 ;
      RECT 98.795 5.43 98.965 5.6 ;
      RECT 98.785 9.345 98.955 9.515 ;
      RECT 98.785 10.085 98.955 10.255 ;
      RECT 98.52 4.07 98.69 4.24 ;
      RECT 98.52 4.91 98.69 5.08 ;
      RECT 98.335 5.43 98.505 5.6 ;
      RECT 98.04 3.23 98.21 3.4 ;
      RECT 98.04 4.91 98.21 5.08 ;
      RECT 97.875 5.43 98.045 5.6 ;
      RECT 97.415 5.43 97.585 5.6 ;
      RECT 97.08 3.23 97.25 3.4 ;
      RECT 97.08 3.79 97.25 3.96 ;
      RECT 97.08 4.35 97.25 4.52 ;
      RECT 97.08 4.91 97.25 5.08 ;
      RECT 96.955 5.43 97.125 5.6 ;
      RECT 96.56 4.91 96.73 5.08 ;
      RECT 96.495 5.43 96.665 5.6 ;
      RECT 96.08 3.23 96.25 3.4 ;
      RECT 96.035 5.43 96.205 5.6 ;
      RECT 95.84 3.79 96.01 3.96 ;
      RECT 95.575 5.43 95.745 5.6 ;
      RECT 95.36 3.79 95.53 3.96 ;
      RECT 95.36 4.35 95.53 4.52 ;
      RECT 95.12 3.23 95.29 3.4 ;
      RECT 95.115 5.43 95.285 5.6 ;
      RECT 94.655 5.43 94.825 5.6 ;
      RECT 94.64 4.35 94.81 4.52 ;
      RECT 94.195 5.43 94.365 5.6 ;
      RECT 94.12 3.79 94.29 3.96 ;
      RECT 94.12 4.63 94.29 4.8 ;
      RECT 93.735 5.43 93.905 5.6 ;
      RECT 93.64 3.23 93.81 3.4 ;
      RECT 93.64 4.35 93.81 4.52 ;
      RECT 93.275 5.43 93.445 5.6 ;
      RECT 93.16 4.63 93.33 4.8 ;
      RECT 92.92 4.07 93.09 4.24 ;
      RECT 92.815 5.43 92.985 5.6 ;
      RECT 92.355 5.43 92.525 5.6 ;
      RECT 92.115 3.79 92.285 3.96 ;
      RECT 91.895 5.43 92.065 5.6 ;
      RECT 91.435 5.43 91.605 5.6 ;
      RECT 91.2 3.23 91.37 3.4 ;
      RECT 91.2 4.35 91.37 4.52 ;
      RECT 90.975 5.43 91.145 5.6 ;
      RECT 90.96 3.79 91.13 3.96 ;
      RECT 90.515 5.43 90.685 5.6 ;
      RECT 90.24 3.23 90.41 3.4 ;
      RECT 90.24 4.77 90.41 4.94 ;
      RECT 90.055 5.43 90.225 5.6 ;
      RECT 88.62 10.09 88.79 10.26 ;
      RECT 88.27 5.455 88.44 5.625 ;
      RECT 88.27 6.84 88.44 7.01 ;
      RECT 88.25 4.055 88.42 4.225 ;
      RECT 88.25 8.24 88.42 8.41 ;
      RECT 87.63 2.205 87.8 2.375 ;
      RECT 87.63 3.685 87.8 3.855 ;
      RECT 87.63 8.61 87.8 8.78 ;
      RECT 87.63 10.09 87.8 10.26 ;
      RECT 87.28 5.455 87.45 5.625 ;
      RECT 87.28 6.84 87.45 7.01 ;
      RECT 87.26 4.055 87.43 4.225 ;
      RECT 87.26 8.24 87.43 8.41 ;
      RECT 86.58 5.46 86.75 5.63 ;
      RECT 86.58 6.835 86.75 7.005 ;
      RECT 86.27 3.32 86.44 3.49 ;
      RECT 86.27 8.975 86.44 9.145 ;
      RECT 85.84 2.21 86.01 2.38 ;
      RECT 85.84 2.95 86.01 3.12 ;
      RECT 85.84 9.345 86.01 9.515 ;
      RECT 85.84 10.085 86.01 10.255 ;
      RECT 85.465 3.69 85.635 3.86 ;
      RECT 85.465 8.605 85.635 8.775 ;
      RECT 82.995 5.43 83.165 5.6 ;
      RECT 82.535 5.43 82.705 5.6 ;
      RECT 82.16 4.07 82.33 4.24 ;
      RECT 82.075 5.43 82.245 5.6 ;
      RECT 81.92 3.23 82.09 3.4 ;
      RECT 81.68 4.35 81.85 4.52 ;
      RECT 81.615 5.43 81.785 5.6 ;
      RECT 81.2 3.79 81.37 3.96 ;
      RECT 81.155 5.43 81.325 5.6 ;
      RECT 80.965 6.835 81.135 7.005 ;
      RECT 80.96 3.23 81.13 3.4 ;
      RECT 80.96 4.35 81.13 4.52 ;
      RECT 80.96 4.91 81.13 5.08 ;
      RECT 80.695 5.43 80.865 5.6 ;
      RECT 80.655 8.975 80.825 9.145 ;
      RECT 80.48 4.35 80.65 4.52 ;
      RECT 80.235 5.43 80.405 5.6 ;
      RECT 80.225 9.345 80.395 9.515 ;
      RECT 80.225 10.085 80.395 10.255 ;
      RECT 79.96 4.07 80.13 4.24 ;
      RECT 79.96 4.91 80.13 5.08 ;
      RECT 79.775 5.43 79.945 5.6 ;
      RECT 79.48 3.23 79.65 3.4 ;
      RECT 79.48 4.91 79.65 5.08 ;
      RECT 79.315 5.43 79.485 5.6 ;
      RECT 78.855 5.43 79.025 5.6 ;
      RECT 78.52 3.23 78.69 3.4 ;
      RECT 78.52 3.79 78.69 3.96 ;
      RECT 78.52 4.35 78.69 4.52 ;
      RECT 78.52 4.91 78.69 5.08 ;
      RECT 78.395 5.43 78.565 5.6 ;
      RECT 78 4.91 78.17 5.08 ;
      RECT 77.935 5.43 78.105 5.6 ;
      RECT 77.52 3.23 77.69 3.4 ;
      RECT 77.475 5.43 77.645 5.6 ;
      RECT 77.28 3.79 77.45 3.96 ;
      RECT 77.015 5.43 77.185 5.6 ;
      RECT 76.8 3.79 76.97 3.96 ;
      RECT 76.8 4.35 76.97 4.52 ;
      RECT 76.56 3.23 76.73 3.4 ;
      RECT 76.555 5.43 76.725 5.6 ;
      RECT 76.095 5.43 76.265 5.6 ;
      RECT 76.08 4.35 76.25 4.52 ;
      RECT 75.635 5.43 75.805 5.6 ;
      RECT 75.56 3.79 75.73 3.96 ;
      RECT 75.56 4.63 75.73 4.8 ;
      RECT 75.175 5.43 75.345 5.6 ;
      RECT 75.08 3.23 75.25 3.4 ;
      RECT 75.08 4.35 75.25 4.52 ;
      RECT 74.715 5.43 74.885 5.6 ;
      RECT 74.6 4.63 74.77 4.8 ;
      RECT 74.36 4.07 74.53 4.24 ;
      RECT 74.255 5.43 74.425 5.6 ;
      RECT 73.795 5.43 73.965 5.6 ;
      RECT 73.555 3.79 73.725 3.96 ;
      RECT 73.335 5.43 73.505 5.6 ;
      RECT 72.875 5.43 73.045 5.6 ;
      RECT 72.64 3.23 72.81 3.4 ;
      RECT 72.64 4.35 72.81 4.52 ;
      RECT 72.415 5.43 72.585 5.6 ;
      RECT 72.4 3.79 72.57 3.96 ;
      RECT 71.955 5.43 72.125 5.6 ;
      RECT 71.68 3.23 71.85 3.4 ;
      RECT 71.68 4.77 71.85 4.94 ;
      RECT 71.495 5.43 71.665 5.6 ;
      RECT 70.06 10.09 70.23 10.26 ;
      RECT 69.71 5.455 69.88 5.625 ;
      RECT 69.71 6.84 69.88 7.01 ;
      RECT 69.69 4.055 69.86 4.225 ;
      RECT 69.69 8.24 69.86 8.41 ;
      RECT 69.07 2.205 69.24 2.375 ;
      RECT 69.07 3.685 69.24 3.855 ;
      RECT 69.07 8.61 69.24 8.78 ;
      RECT 69.07 10.09 69.24 10.26 ;
      RECT 68.72 5.455 68.89 5.625 ;
      RECT 68.72 6.84 68.89 7.01 ;
      RECT 68.7 4.055 68.87 4.225 ;
      RECT 68.7 8.24 68.87 8.41 ;
      RECT 68.02 5.46 68.19 5.63 ;
      RECT 68.02 6.835 68.19 7.005 ;
      RECT 67.71 3.32 67.88 3.49 ;
      RECT 67.71 8.975 67.88 9.145 ;
      RECT 67.28 2.21 67.45 2.38 ;
      RECT 67.28 2.95 67.45 3.12 ;
      RECT 67.28 9.345 67.45 9.515 ;
      RECT 67.28 10.085 67.45 10.255 ;
      RECT 66.905 3.69 67.075 3.86 ;
      RECT 66.905 8.605 67.075 8.775 ;
      RECT 64.435 5.43 64.605 5.6 ;
      RECT 63.975 5.43 64.145 5.6 ;
      RECT 63.6 4.07 63.77 4.24 ;
      RECT 63.515 5.43 63.685 5.6 ;
      RECT 63.36 3.23 63.53 3.4 ;
      RECT 63.12 4.35 63.29 4.52 ;
      RECT 63.055 5.43 63.225 5.6 ;
      RECT 62.64 3.79 62.81 3.96 ;
      RECT 62.595 5.43 62.765 5.6 ;
      RECT 62.405 6.835 62.575 7.005 ;
      RECT 62.4 3.23 62.57 3.4 ;
      RECT 62.4 4.35 62.57 4.52 ;
      RECT 62.4 4.91 62.57 5.08 ;
      RECT 62.135 5.43 62.305 5.6 ;
      RECT 62.095 8.975 62.265 9.145 ;
      RECT 61.92 4.35 62.09 4.52 ;
      RECT 61.675 5.43 61.845 5.6 ;
      RECT 61.665 9.345 61.835 9.515 ;
      RECT 61.665 10.085 61.835 10.255 ;
      RECT 61.4 4.07 61.57 4.24 ;
      RECT 61.4 4.91 61.57 5.08 ;
      RECT 61.215 5.43 61.385 5.6 ;
      RECT 60.92 3.23 61.09 3.4 ;
      RECT 60.92 4.91 61.09 5.08 ;
      RECT 60.755 5.43 60.925 5.6 ;
      RECT 60.295 5.43 60.465 5.6 ;
      RECT 59.96 3.23 60.13 3.4 ;
      RECT 59.96 3.79 60.13 3.96 ;
      RECT 59.96 4.35 60.13 4.52 ;
      RECT 59.96 4.91 60.13 5.08 ;
      RECT 59.835 5.43 60.005 5.6 ;
      RECT 59.44 4.91 59.61 5.08 ;
      RECT 59.375 5.43 59.545 5.6 ;
      RECT 58.96 3.23 59.13 3.4 ;
      RECT 58.915 5.43 59.085 5.6 ;
      RECT 58.72 3.79 58.89 3.96 ;
      RECT 58.455 5.43 58.625 5.6 ;
      RECT 58.24 3.79 58.41 3.96 ;
      RECT 58.24 4.35 58.41 4.52 ;
      RECT 58 3.23 58.17 3.4 ;
      RECT 57.995 5.43 58.165 5.6 ;
      RECT 57.535 5.43 57.705 5.6 ;
      RECT 57.52 4.35 57.69 4.52 ;
      RECT 57.075 5.43 57.245 5.6 ;
      RECT 57 3.79 57.17 3.96 ;
      RECT 57 4.63 57.17 4.8 ;
      RECT 56.615 5.43 56.785 5.6 ;
      RECT 56.52 3.23 56.69 3.4 ;
      RECT 56.52 4.35 56.69 4.52 ;
      RECT 56.155 5.43 56.325 5.6 ;
      RECT 56.04 4.63 56.21 4.8 ;
      RECT 55.8 4.07 55.97 4.24 ;
      RECT 55.695 5.43 55.865 5.6 ;
      RECT 55.235 5.43 55.405 5.6 ;
      RECT 54.995 3.79 55.165 3.96 ;
      RECT 54.775 5.43 54.945 5.6 ;
      RECT 54.315 5.43 54.485 5.6 ;
      RECT 54.08 3.23 54.25 3.4 ;
      RECT 54.08 4.35 54.25 4.52 ;
      RECT 53.855 5.43 54.025 5.6 ;
      RECT 53.84 3.79 54.01 3.96 ;
      RECT 53.395 5.43 53.565 5.6 ;
      RECT 53.12 3.23 53.29 3.4 ;
      RECT 53.12 4.77 53.29 4.94 ;
      RECT 52.935 5.43 53.105 5.6 ;
      RECT 51.5 10.09 51.67 10.26 ;
      RECT 51.15 5.455 51.32 5.625 ;
      RECT 51.15 6.84 51.32 7.01 ;
      RECT 51.13 4.055 51.3 4.225 ;
      RECT 51.13 8.24 51.3 8.41 ;
      RECT 50.51 2.205 50.68 2.375 ;
      RECT 50.51 3.685 50.68 3.855 ;
      RECT 50.51 8.61 50.68 8.78 ;
      RECT 50.51 10.09 50.68 10.26 ;
      RECT 50.16 5.455 50.33 5.625 ;
      RECT 50.16 6.84 50.33 7.01 ;
      RECT 50.14 4.055 50.31 4.225 ;
      RECT 50.14 8.24 50.31 8.41 ;
      RECT 49.46 5.46 49.63 5.63 ;
      RECT 49.46 6.835 49.63 7.005 ;
      RECT 49.15 3.32 49.32 3.49 ;
      RECT 49.15 8.975 49.32 9.145 ;
      RECT 48.72 2.21 48.89 2.38 ;
      RECT 48.72 2.95 48.89 3.12 ;
      RECT 48.72 9.345 48.89 9.515 ;
      RECT 48.72 10.085 48.89 10.255 ;
      RECT 48.345 3.69 48.515 3.86 ;
      RECT 48.345 8.605 48.515 8.775 ;
      RECT 45.875 5.43 46.045 5.6 ;
      RECT 45.415 5.43 45.585 5.6 ;
      RECT 45.04 4.07 45.21 4.24 ;
      RECT 44.955 5.43 45.125 5.6 ;
      RECT 44.8 3.23 44.97 3.4 ;
      RECT 44.56 4.35 44.73 4.52 ;
      RECT 44.495 5.43 44.665 5.6 ;
      RECT 44.08 3.79 44.25 3.96 ;
      RECT 44.035 5.43 44.205 5.6 ;
      RECT 43.845 6.835 44.015 7.005 ;
      RECT 43.84 3.23 44.01 3.4 ;
      RECT 43.84 4.35 44.01 4.52 ;
      RECT 43.84 4.91 44.01 5.08 ;
      RECT 43.575 5.43 43.745 5.6 ;
      RECT 43.535 8.975 43.705 9.145 ;
      RECT 43.36 4.35 43.53 4.52 ;
      RECT 43.115 5.43 43.285 5.6 ;
      RECT 43.105 9.345 43.275 9.515 ;
      RECT 43.105 10.085 43.275 10.255 ;
      RECT 42.84 4.07 43.01 4.24 ;
      RECT 42.84 4.91 43.01 5.08 ;
      RECT 42.655 5.43 42.825 5.6 ;
      RECT 42.36 3.23 42.53 3.4 ;
      RECT 42.36 4.91 42.53 5.08 ;
      RECT 42.195 5.43 42.365 5.6 ;
      RECT 41.735 5.43 41.905 5.6 ;
      RECT 41.4 3.23 41.57 3.4 ;
      RECT 41.4 3.79 41.57 3.96 ;
      RECT 41.4 4.35 41.57 4.52 ;
      RECT 41.4 4.91 41.57 5.08 ;
      RECT 41.275 5.43 41.445 5.6 ;
      RECT 40.88 4.91 41.05 5.08 ;
      RECT 40.815 5.43 40.985 5.6 ;
      RECT 40.4 3.23 40.57 3.4 ;
      RECT 40.355 5.43 40.525 5.6 ;
      RECT 40.16 3.79 40.33 3.96 ;
      RECT 39.895 5.43 40.065 5.6 ;
      RECT 39.68 3.79 39.85 3.96 ;
      RECT 39.68 4.35 39.85 4.52 ;
      RECT 39.44 3.23 39.61 3.4 ;
      RECT 39.435 5.43 39.605 5.6 ;
      RECT 38.975 5.43 39.145 5.6 ;
      RECT 38.96 4.35 39.13 4.52 ;
      RECT 38.515 5.43 38.685 5.6 ;
      RECT 38.44 3.79 38.61 3.96 ;
      RECT 38.44 4.63 38.61 4.8 ;
      RECT 38.055 5.43 38.225 5.6 ;
      RECT 37.96 3.23 38.13 3.4 ;
      RECT 37.96 4.35 38.13 4.52 ;
      RECT 37.595 5.43 37.765 5.6 ;
      RECT 37.48 4.63 37.65 4.8 ;
      RECT 37.24 4.07 37.41 4.24 ;
      RECT 37.135 5.43 37.305 5.6 ;
      RECT 36.675 5.43 36.845 5.6 ;
      RECT 36.435 3.79 36.605 3.96 ;
      RECT 36.215 5.43 36.385 5.6 ;
      RECT 35.755 5.43 35.925 5.6 ;
      RECT 35.52 3.23 35.69 3.4 ;
      RECT 35.52 4.35 35.69 4.52 ;
      RECT 35.295 5.43 35.465 5.6 ;
      RECT 35.28 3.79 35.45 3.96 ;
      RECT 34.835 5.43 35.005 5.6 ;
      RECT 34.56 3.23 34.73 3.4 ;
      RECT 34.56 4.77 34.73 4.94 ;
      RECT 34.375 5.43 34.545 5.6 ;
      RECT 32.94 10.09 33.11 10.26 ;
      RECT 32.59 5.455 32.76 5.625 ;
      RECT 32.59 6.84 32.76 7.01 ;
      RECT 32.57 4.055 32.74 4.225 ;
      RECT 32.57 8.24 32.74 8.41 ;
      RECT 31.95 2.205 32.12 2.375 ;
      RECT 31.95 3.685 32.12 3.855 ;
      RECT 31.95 8.61 32.12 8.78 ;
      RECT 31.95 10.09 32.12 10.26 ;
      RECT 31.6 5.455 31.77 5.625 ;
      RECT 31.6 6.84 31.77 7.01 ;
      RECT 31.58 4.055 31.75 4.225 ;
      RECT 31.58 8.24 31.75 8.41 ;
      RECT 30.9 5.46 31.07 5.63 ;
      RECT 30.9 6.835 31.07 7.005 ;
      RECT 30.59 3.32 30.76 3.49 ;
      RECT 30.59 8.975 30.76 9.145 ;
      RECT 30.16 2.21 30.33 2.38 ;
      RECT 30.16 2.95 30.33 3.12 ;
      RECT 30.16 9.345 30.33 9.515 ;
      RECT 30.16 10.085 30.33 10.255 ;
      RECT 29.785 3.69 29.955 3.86 ;
      RECT 29.785 8.605 29.955 8.775 ;
      RECT 27.315 5.43 27.485 5.6 ;
      RECT 26.855 5.43 27.025 5.6 ;
      RECT 26.48 4.07 26.65 4.24 ;
      RECT 26.395 5.43 26.565 5.6 ;
      RECT 26.24 3.23 26.41 3.4 ;
      RECT 26 4.35 26.17 4.52 ;
      RECT 25.935 5.43 26.105 5.6 ;
      RECT 25.52 3.79 25.69 3.96 ;
      RECT 25.475 5.43 25.645 5.6 ;
      RECT 25.285 6.835 25.455 7.005 ;
      RECT 25.28 3.23 25.45 3.4 ;
      RECT 25.28 4.35 25.45 4.52 ;
      RECT 25.28 4.91 25.45 5.08 ;
      RECT 25.015 5.43 25.185 5.6 ;
      RECT 24.975 8.975 25.145 9.145 ;
      RECT 24.8 4.35 24.97 4.52 ;
      RECT 24.555 5.43 24.725 5.6 ;
      RECT 24.545 9.345 24.715 9.515 ;
      RECT 24.545 10.085 24.715 10.255 ;
      RECT 24.28 4.07 24.45 4.24 ;
      RECT 24.28 4.91 24.45 5.08 ;
      RECT 24.095 5.43 24.265 5.6 ;
      RECT 23.8 3.23 23.97 3.4 ;
      RECT 23.8 4.91 23.97 5.08 ;
      RECT 23.635 5.43 23.805 5.6 ;
      RECT 23.175 5.43 23.345 5.6 ;
      RECT 22.84 3.23 23.01 3.4 ;
      RECT 22.84 3.79 23.01 3.96 ;
      RECT 22.84 4.35 23.01 4.52 ;
      RECT 22.84 4.91 23.01 5.08 ;
      RECT 22.715 5.43 22.885 5.6 ;
      RECT 22.32 4.91 22.49 5.08 ;
      RECT 22.255 5.43 22.425 5.6 ;
      RECT 21.84 3.23 22.01 3.4 ;
      RECT 21.795 5.43 21.965 5.6 ;
      RECT 21.6 3.79 21.77 3.96 ;
      RECT 21.335 5.43 21.505 5.6 ;
      RECT 21.12 3.79 21.29 3.96 ;
      RECT 21.12 4.35 21.29 4.52 ;
      RECT 20.88 3.23 21.05 3.4 ;
      RECT 20.875 5.43 21.045 5.6 ;
      RECT 20.415 5.43 20.585 5.6 ;
      RECT 20.4 4.35 20.57 4.52 ;
      RECT 19.955 5.43 20.125 5.6 ;
      RECT 19.88 3.79 20.05 3.96 ;
      RECT 19.88 4.63 20.05 4.8 ;
      RECT 19.495 5.43 19.665 5.6 ;
      RECT 19.4 3.23 19.57 3.4 ;
      RECT 19.4 4.35 19.57 4.52 ;
      RECT 19.035 5.43 19.205 5.6 ;
      RECT 18.92 4.63 19.09 4.8 ;
      RECT 18.68 4.07 18.85 4.24 ;
      RECT 18.575 5.43 18.745 5.6 ;
      RECT 18.115 5.43 18.285 5.6 ;
      RECT 17.875 3.79 18.045 3.96 ;
      RECT 17.655 5.43 17.825 5.6 ;
      RECT 17.195 5.43 17.365 5.6 ;
      RECT 16.96 3.23 17.13 3.4 ;
      RECT 16.96 4.35 17.13 4.52 ;
      RECT 16.735 5.43 16.905 5.6 ;
      RECT 16.72 3.79 16.89 3.96 ;
      RECT 16.275 5.43 16.445 5.6 ;
      RECT 16 3.23 16.17 3.4 ;
      RECT 16 4.77 16.17 4.94 ;
      RECT 15.815 5.43 15.985 5.6 ;
      RECT 14.47 6.835 14.64 7.005 ;
      RECT 14.16 8.975 14.33 9.145 ;
      RECT 13.73 9.345 13.9 9.515 ;
      RECT 13.73 10.085 13.9 10.255 ;
      RECT 13.355 8.605 13.525 8.775 ;
    LAYER li1 ;
      RECT 14.16 5.44 14.33 10.595 ;
      RECT 106.75 4.695 106.92 7.77 ;
      RECT 105.76 4.695 105.93 7.77 ;
      RECT 88.19 4.695 88.36 7.77 ;
      RECT 87.2 4.695 87.37 7.77 ;
      RECT 69.63 4.695 69.8 7.77 ;
      RECT 68.64 4.695 68.81 7.77 ;
      RECT 51.07 4.695 51.24 7.77 ;
      RECT 50.08 4.695 50.25 7.77 ;
      RECT 32.51 4.695 32.68 7.77 ;
      RECT 31.52 4.695 31.69 7.77 ;
      RECT 103.02 4.7 103.19 7.765 ;
      RECT 97.405 5.43 97.575 7.765 ;
      RECT 84.46 4.7 84.63 7.765 ;
      RECT 78.845 5.43 79.015 7.765 ;
      RECT 65.9 4.7 66.07 7.765 ;
      RECT 60.285 5.43 60.455 7.765 ;
      RECT 47.34 4.7 47.51 7.765 ;
      RECT 41.725 5.43 41.895 7.765 ;
      RECT 28.78 4.7 28.95 7.765 ;
      RECT 23.165 5.43 23.335 7.765 ;
      RECT 12.35 5.44 12.52 7.765 ;
      RECT 12.13 5.44 107.625 7.04 ;
      RECT 89.91 5.43 107.725 7.035 ;
      RECT 71.35 5.43 89.165 7.04 ;
      RECT 52.79 5.43 70.605 7.04 ;
      RECT 34.23 5.43 52.045 7.04 ;
      RECT 15.67 5.43 33.485 7.04 ;
      RECT 105.59 5.425 107.57 7.04 ;
      RECT 100 4.93 100.17 7.04 ;
      RECT 97.56 4.93 97.73 7.04 ;
      RECT 95.6 4.93 95.77 7.04 ;
      RECT 94.64 4.93 94.81 7.04 ;
      RECT 92.68 4.93 92.85 7.04 ;
      RECT 91.68 4.93 91.85 7.04 ;
      RECT 90.72 4.93 90.89 7.04 ;
      RECT 87.03 5.425 89.01 7.04 ;
      RECT 81.44 4.93 81.61 7.04 ;
      RECT 79 4.93 79.17 7.04 ;
      RECT 77.04 4.93 77.21 7.04 ;
      RECT 76.08 4.93 76.25 7.04 ;
      RECT 74.12 4.93 74.29 7.04 ;
      RECT 73.12 4.93 73.29 7.04 ;
      RECT 72.16 4.93 72.33 7.04 ;
      RECT 68.47 5.425 70.45 7.04 ;
      RECT 62.88 4.93 63.05 7.04 ;
      RECT 60.44 4.93 60.61 7.04 ;
      RECT 58.48 4.93 58.65 7.04 ;
      RECT 57.52 4.93 57.69 7.04 ;
      RECT 55.56 4.93 55.73 7.04 ;
      RECT 54.56 4.93 54.73 7.04 ;
      RECT 53.6 4.93 53.77 7.04 ;
      RECT 49.91 5.425 51.89 7.04 ;
      RECT 44.32 4.93 44.49 7.04 ;
      RECT 41.88 4.93 42.05 7.04 ;
      RECT 39.92 4.93 40.09 7.04 ;
      RECT 38.96 4.93 39.13 7.04 ;
      RECT 37 4.93 37.17 7.04 ;
      RECT 36 4.93 36.17 7.04 ;
      RECT 35.04 4.93 35.21 7.04 ;
      RECT 31.35 5.425 33.33 7.04 ;
      RECT 25.76 4.93 25.93 7.04 ;
      RECT 23.32 4.93 23.49 7.04 ;
      RECT 21.36 4.93 21.53 7.04 ;
      RECT 20.4 4.93 20.57 7.04 ;
      RECT 18.44 4.93 18.61 7.04 ;
      RECT 17.44 4.93 17.61 7.04 ;
      RECT 16.48 4.93 16.65 7.04 ;
      RECT 107.18 7.31 107.35 8.78 ;
      RECT 107.18 8.605 107.355 8.775 ;
      RECT 106.81 3.035 106.98 4.225 ;
      RECT 106.81 3.035 107.28 3.205 ;
      RECT 106.81 9.26 107.28 9.43 ;
      RECT 106.81 8.24 106.98 9.43 ;
      RECT 105.82 3.035 105.99 4.225 ;
      RECT 105.82 3.035 106.29 3.205 ;
      RECT 105.82 9.26 106.29 9.43 ;
      RECT 105.82 8.24 105.99 9.43 ;
      RECT 103.97 3.93 104.14 5.16 ;
      RECT 104.025 2.15 104.195 4.1 ;
      RECT 103.97 1.87 104.14 2.32 ;
      RECT 103.97 10.145 104.14 10.595 ;
      RECT 104.025 8.365 104.195 10.315 ;
      RECT 103.97 7.305 104.14 8.535 ;
      RECT 103.45 1.87 103.62 5.16 ;
      RECT 103.45 3.37 103.855 3.7 ;
      RECT 103.45 2.53 103.855 2.86 ;
      RECT 103.45 7.305 103.62 10.595 ;
      RECT 103.45 9.605 103.855 9.935 ;
      RECT 103.45 8.765 103.855 9.095 ;
      RECT 100.24 4.52 101.21 4.69 ;
      RECT 100.24 4.35 100.41 4.69 ;
      RECT 99.76 3.79 99.93 4.12 ;
      RECT 99.76 3.87 100.49 4.04 ;
      RECT 99.4 4.91 99.69 5.08 ;
      RECT 99.4 3.87 99.57 5.08 ;
      RECT 99.4 4.35 99.69 4.52 ;
      RECT 99.2 3.87 99.57 4.04 ;
      RECT 98.52 3.97 98.69 4.24 ;
      RECT 98.28 3.97 98.69 4.14 ;
      RECT 98.2 3.87 98.53 4.04 ;
      RECT 98.04 4.91 98.69 5.08 ;
      RECT 98.52 4.44 98.69 5.08 ;
      RECT 98.4 4.52 98.69 5.08 ;
      RECT 97.835 7.305 98.005 10.595 ;
      RECT 97.835 9.605 98.24 9.935 ;
      RECT 97.835 8.765 98.24 9.095 ;
      RECT 97.08 4.21 97.25 4.52 ;
      RECT 97.08 4.21 97.97 4.38 ;
      RECT 97.8 3.79 97.97 4.38 ;
      RECT 97.08 3.87 97.57 4.04 ;
      RECT 97.08 3.79 97.25 4.04 ;
      RECT 95.04 4.52 95.53 4.69 ;
      RECT 96.2 3.87 96.37 4.52 ;
      RECT 95.36 4.35 96.37 4.52 ;
      RECT 96.32 3.79 96.49 4.12 ;
      RECT 95.12 3.13 95.29 3.4 ;
      RECT 94.56 3.13 95.29 3.3 ;
      RECT 94.64 3.87 94.81 4.52 ;
      RECT 94.64 3.87 95.13 4.04 ;
      RECT 93.8 3.87 94.29 4.04 ;
      RECT 94.12 3.79 94.29 4.04 ;
      RECT 93.64 3.13 93.81 3.4 ;
      RECT 93.08 3.13 93.81 3.3 ;
      RECT 93.16 4.52 93.33 4.8 ;
      RECT 92.12 4.52 93.41 4.69 ;
      RECT 92.115 3.87 92.69 4.04 ;
      RECT 92.115 3.79 92.285 4.04 ;
      RECT 91.2 3.13 91.37 3.4 ;
      RECT 91.2 3.13 91.93 3.3 ;
      RECT 91.2 4.35 91.37 4.77 ;
      RECT 90.58 4.435 91.37 4.605 ;
      RECT 90.58 4.21 90.75 4.605 ;
      RECT 90.48 3.79 90.65 4.38 ;
      RECT 90.24 3.87 90.65 4.14 ;
      RECT 88.62 7.31 88.79 8.78 ;
      RECT 88.62 8.605 88.795 8.775 ;
      RECT 88.25 3.035 88.42 4.225 ;
      RECT 88.25 3.035 88.72 3.205 ;
      RECT 88.25 9.26 88.72 9.43 ;
      RECT 88.25 8.24 88.42 9.43 ;
      RECT 87.26 3.035 87.43 4.225 ;
      RECT 87.26 3.035 87.73 3.205 ;
      RECT 87.26 9.26 87.73 9.43 ;
      RECT 87.26 8.24 87.43 9.43 ;
      RECT 85.41 3.93 85.58 5.16 ;
      RECT 85.465 2.15 85.635 4.1 ;
      RECT 85.41 1.87 85.58 2.32 ;
      RECT 85.41 10.145 85.58 10.595 ;
      RECT 85.465 8.365 85.635 10.315 ;
      RECT 85.41 7.305 85.58 8.535 ;
      RECT 84.89 1.87 85.06 5.16 ;
      RECT 84.89 3.37 85.295 3.7 ;
      RECT 84.89 2.53 85.295 2.86 ;
      RECT 84.89 7.305 85.06 10.595 ;
      RECT 84.89 9.605 85.295 9.935 ;
      RECT 84.89 8.765 85.295 9.095 ;
      RECT 81.68 4.52 82.65 4.69 ;
      RECT 81.68 4.35 81.85 4.69 ;
      RECT 81.2 3.79 81.37 4.12 ;
      RECT 81.2 3.87 81.93 4.04 ;
      RECT 80.84 4.91 81.13 5.08 ;
      RECT 80.84 3.87 81.01 5.08 ;
      RECT 80.84 4.35 81.13 4.52 ;
      RECT 80.64 3.87 81.01 4.04 ;
      RECT 79.96 3.97 80.13 4.24 ;
      RECT 79.72 3.97 80.13 4.14 ;
      RECT 79.64 3.87 79.97 4.04 ;
      RECT 79.48 4.91 80.13 5.08 ;
      RECT 79.96 4.44 80.13 5.08 ;
      RECT 79.84 4.52 80.13 5.08 ;
      RECT 79.275 7.305 79.445 10.595 ;
      RECT 79.275 9.605 79.68 9.935 ;
      RECT 79.275 8.765 79.68 9.095 ;
      RECT 78.52 4.21 78.69 4.52 ;
      RECT 78.52 4.21 79.41 4.38 ;
      RECT 79.24 3.79 79.41 4.38 ;
      RECT 78.52 3.87 79.01 4.04 ;
      RECT 78.52 3.79 78.69 4.04 ;
      RECT 76.48 4.52 76.97 4.69 ;
      RECT 77.64 3.87 77.81 4.52 ;
      RECT 76.8 4.35 77.81 4.52 ;
      RECT 77.76 3.79 77.93 4.12 ;
      RECT 76.56 3.13 76.73 3.4 ;
      RECT 76 3.13 76.73 3.3 ;
      RECT 76.08 3.87 76.25 4.52 ;
      RECT 76.08 3.87 76.57 4.04 ;
      RECT 75.24 3.87 75.73 4.04 ;
      RECT 75.56 3.79 75.73 4.04 ;
      RECT 75.08 3.13 75.25 3.4 ;
      RECT 74.52 3.13 75.25 3.3 ;
      RECT 74.6 4.52 74.77 4.8 ;
      RECT 73.56 4.52 74.85 4.69 ;
      RECT 73.555 3.87 74.13 4.04 ;
      RECT 73.555 3.79 73.725 4.04 ;
      RECT 72.64 3.13 72.81 3.4 ;
      RECT 72.64 3.13 73.37 3.3 ;
      RECT 72.64 4.35 72.81 4.77 ;
      RECT 72.02 4.435 72.81 4.605 ;
      RECT 72.02 4.21 72.19 4.605 ;
      RECT 71.92 3.79 72.09 4.38 ;
      RECT 71.68 3.87 72.09 4.14 ;
      RECT 70.06 7.31 70.23 8.78 ;
      RECT 70.06 8.605 70.235 8.775 ;
      RECT 69.69 3.035 69.86 4.225 ;
      RECT 69.69 3.035 70.16 3.205 ;
      RECT 69.69 9.26 70.16 9.43 ;
      RECT 69.69 8.24 69.86 9.43 ;
      RECT 68.7 3.035 68.87 4.225 ;
      RECT 68.7 3.035 69.17 3.205 ;
      RECT 68.7 9.26 69.17 9.43 ;
      RECT 68.7 8.24 68.87 9.43 ;
      RECT 66.85 3.93 67.02 5.16 ;
      RECT 66.905 2.15 67.075 4.1 ;
      RECT 66.85 1.87 67.02 2.32 ;
      RECT 66.85 10.145 67.02 10.595 ;
      RECT 66.905 8.365 67.075 10.315 ;
      RECT 66.85 7.305 67.02 8.535 ;
      RECT 66.33 1.87 66.5 5.16 ;
      RECT 66.33 3.37 66.735 3.7 ;
      RECT 66.33 2.53 66.735 2.86 ;
      RECT 66.33 7.305 66.5 10.595 ;
      RECT 66.33 9.605 66.735 9.935 ;
      RECT 66.33 8.765 66.735 9.095 ;
      RECT 63.12 4.52 64.09 4.69 ;
      RECT 63.12 4.35 63.29 4.69 ;
      RECT 62.64 3.79 62.81 4.12 ;
      RECT 62.64 3.87 63.37 4.04 ;
      RECT 62.28 4.91 62.57 5.08 ;
      RECT 62.28 3.87 62.45 5.08 ;
      RECT 62.28 4.35 62.57 4.52 ;
      RECT 62.08 3.87 62.45 4.04 ;
      RECT 61.4 3.97 61.57 4.24 ;
      RECT 61.16 3.97 61.57 4.14 ;
      RECT 61.08 3.87 61.41 4.04 ;
      RECT 60.92 4.91 61.57 5.08 ;
      RECT 61.4 4.44 61.57 5.08 ;
      RECT 61.28 4.52 61.57 5.08 ;
      RECT 60.715 7.305 60.885 10.595 ;
      RECT 60.715 9.605 61.12 9.935 ;
      RECT 60.715 8.765 61.12 9.095 ;
      RECT 59.96 4.21 60.13 4.52 ;
      RECT 59.96 4.21 60.85 4.38 ;
      RECT 60.68 3.79 60.85 4.38 ;
      RECT 59.96 3.87 60.45 4.04 ;
      RECT 59.96 3.79 60.13 4.04 ;
      RECT 57.92 4.52 58.41 4.69 ;
      RECT 59.08 3.87 59.25 4.52 ;
      RECT 58.24 4.35 59.25 4.52 ;
      RECT 59.2 3.79 59.37 4.12 ;
      RECT 58 3.13 58.17 3.4 ;
      RECT 57.44 3.13 58.17 3.3 ;
      RECT 57.52 3.87 57.69 4.52 ;
      RECT 57.52 3.87 58.01 4.04 ;
      RECT 56.68 3.87 57.17 4.04 ;
      RECT 57 3.79 57.17 4.04 ;
      RECT 56.52 3.13 56.69 3.4 ;
      RECT 55.96 3.13 56.69 3.3 ;
      RECT 56.04 4.52 56.21 4.8 ;
      RECT 55 4.52 56.29 4.69 ;
      RECT 54.995 3.87 55.57 4.04 ;
      RECT 54.995 3.79 55.165 4.04 ;
      RECT 54.08 3.13 54.25 3.4 ;
      RECT 54.08 3.13 54.81 3.3 ;
      RECT 54.08 4.35 54.25 4.77 ;
      RECT 53.46 4.435 54.25 4.605 ;
      RECT 53.46 4.21 53.63 4.605 ;
      RECT 53.36 3.79 53.53 4.38 ;
      RECT 53.12 3.87 53.53 4.14 ;
      RECT 51.5 7.31 51.67 8.78 ;
      RECT 51.5 8.605 51.675 8.775 ;
      RECT 51.13 3.035 51.3 4.225 ;
      RECT 51.13 3.035 51.6 3.205 ;
      RECT 51.13 9.26 51.6 9.43 ;
      RECT 51.13 8.24 51.3 9.43 ;
      RECT 50.14 3.035 50.31 4.225 ;
      RECT 50.14 3.035 50.61 3.205 ;
      RECT 50.14 9.26 50.61 9.43 ;
      RECT 50.14 8.24 50.31 9.43 ;
      RECT 48.29 3.93 48.46 5.16 ;
      RECT 48.345 2.15 48.515 4.1 ;
      RECT 48.29 1.87 48.46 2.32 ;
      RECT 48.29 10.145 48.46 10.595 ;
      RECT 48.345 8.365 48.515 10.315 ;
      RECT 48.29 7.305 48.46 8.535 ;
      RECT 47.77 1.87 47.94 5.16 ;
      RECT 47.77 3.37 48.175 3.7 ;
      RECT 47.77 2.53 48.175 2.86 ;
      RECT 47.77 7.305 47.94 10.595 ;
      RECT 47.77 9.605 48.175 9.935 ;
      RECT 47.77 8.765 48.175 9.095 ;
      RECT 44.56 4.52 45.53 4.69 ;
      RECT 44.56 4.35 44.73 4.69 ;
      RECT 44.08 3.79 44.25 4.12 ;
      RECT 44.08 3.87 44.81 4.04 ;
      RECT 43.72 4.91 44.01 5.08 ;
      RECT 43.72 3.87 43.89 5.08 ;
      RECT 43.72 4.35 44.01 4.52 ;
      RECT 43.52 3.87 43.89 4.04 ;
      RECT 42.84 3.97 43.01 4.24 ;
      RECT 42.6 3.97 43.01 4.14 ;
      RECT 42.52 3.87 42.85 4.04 ;
      RECT 42.36 4.91 43.01 5.08 ;
      RECT 42.84 4.44 43.01 5.08 ;
      RECT 42.72 4.52 43.01 5.08 ;
      RECT 42.155 7.305 42.325 10.595 ;
      RECT 42.155 9.605 42.56 9.935 ;
      RECT 42.155 8.765 42.56 9.095 ;
      RECT 41.4 4.21 41.57 4.52 ;
      RECT 41.4 4.21 42.29 4.38 ;
      RECT 42.12 3.79 42.29 4.38 ;
      RECT 41.4 3.87 41.89 4.04 ;
      RECT 41.4 3.79 41.57 4.04 ;
      RECT 39.36 4.52 39.85 4.69 ;
      RECT 40.52 3.87 40.69 4.52 ;
      RECT 39.68 4.35 40.69 4.52 ;
      RECT 40.64 3.79 40.81 4.12 ;
      RECT 39.44 3.13 39.61 3.4 ;
      RECT 38.88 3.13 39.61 3.3 ;
      RECT 38.96 3.87 39.13 4.52 ;
      RECT 38.96 3.87 39.45 4.04 ;
      RECT 38.12 3.87 38.61 4.04 ;
      RECT 38.44 3.79 38.61 4.04 ;
      RECT 37.96 3.13 38.13 3.4 ;
      RECT 37.4 3.13 38.13 3.3 ;
      RECT 37.48 4.52 37.65 4.8 ;
      RECT 36.44 4.52 37.73 4.69 ;
      RECT 36.435 3.87 37.01 4.04 ;
      RECT 36.435 3.79 36.605 4.04 ;
      RECT 35.52 3.13 35.69 3.4 ;
      RECT 35.52 3.13 36.25 3.3 ;
      RECT 35.52 4.35 35.69 4.77 ;
      RECT 34.9 4.435 35.69 4.605 ;
      RECT 34.9 4.21 35.07 4.605 ;
      RECT 34.8 3.79 34.97 4.38 ;
      RECT 34.56 3.87 34.97 4.14 ;
      RECT 32.94 7.31 33.11 8.78 ;
      RECT 32.94 8.605 33.115 8.775 ;
      RECT 32.57 3.035 32.74 4.225 ;
      RECT 32.57 3.035 33.04 3.205 ;
      RECT 32.57 9.26 33.04 9.43 ;
      RECT 32.57 8.24 32.74 9.43 ;
      RECT 31.58 3.035 31.75 4.225 ;
      RECT 31.58 3.035 32.05 3.205 ;
      RECT 31.58 9.26 32.05 9.43 ;
      RECT 31.58 8.24 31.75 9.43 ;
      RECT 29.73 3.93 29.9 5.16 ;
      RECT 29.785 2.15 29.955 4.1 ;
      RECT 29.73 1.87 29.9 2.32 ;
      RECT 29.73 10.145 29.9 10.595 ;
      RECT 29.785 8.365 29.955 10.315 ;
      RECT 29.73 7.305 29.9 8.535 ;
      RECT 29.21 1.87 29.38 5.16 ;
      RECT 29.21 3.37 29.615 3.7 ;
      RECT 29.21 2.53 29.615 2.86 ;
      RECT 29.21 7.305 29.38 10.595 ;
      RECT 29.21 9.605 29.615 9.935 ;
      RECT 29.21 8.765 29.615 9.095 ;
      RECT 26 4.52 26.97 4.69 ;
      RECT 26 4.35 26.17 4.69 ;
      RECT 25.52 3.79 25.69 4.12 ;
      RECT 25.52 3.87 26.25 4.04 ;
      RECT 25.16 4.91 25.45 5.08 ;
      RECT 25.16 3.87 25.33 5.08 ;
      RECT 25.16 4.35 25.45 4.52 ;
      RECT 24.96 3.87 25.33 4.04 ;
      RECT 24.28 3.97 24.45 4.24 ;
      RECT 24.04 3.97 24.45 4.14 ;
      RECT 23.96 3.87 24.29 4.04 ;
      RECT 23.8 4.91 24.45 5.08 ;
      RECT 24.28 4.44 24.45 5.08 ;
      RECT 24.16 4.52 24.45 5.08 ;
      RECT 23.595 7.305 23.765 10.595 ;
      RECT 23.595 9.605 24 9.935 ;
      RECT 23.595 8.765 24 9.095 ;
      RECT 22.84 4.21 23.01 4.52 ;
      RECT 22.84 4.21 23.73 4.38 ;
      RECT 23.56 3.79 23.73 4.38 ;
      RECT 22.84 3.87 23.33 4.04 ;
      RECT 22.84 3.79 23.01 4.04 ;
      RECT 20.8 4.52 21.29 4.69 ;
      RECT 21.96 3.87 22.13 4.52 ;
      RECT 21.12 4.35 22.13 4.52 ;
      RECT 22.08 3.79 22.25 4.12 ;
      RECT 20.88 3.13 21.05 3.4 ;
      RECT 20.32 3.13 21.05 3.3 ;
      RECT 20.4 3.87 20.57 4.52 ;
      RECT 20.4 3.87 20.89 4.04 ;
      RECT 19.56 3.87 20.05 4.04 ;
      RECT 19.88 3.79 20.05 4.04 ;
      RECT 19.4 3.13 19.57 3.4 ;
      RECT 18.84 3.13 19.57 3.3 ;
      RECT 18.92 4.52 19.09 4.8 ;
      RECT 17.88 4.52 19.17 4.69 ;
      RECT 17.875 3.87 18.45 4.04 ;
      RECT 17.875 3.79 18.045 4.04 ;
      RECT 16.96 3.13 17.13 3.4 ;
      RECT 16.96 3.13 17.69 3.3 ;
      RECT 16.96 4.35 17.13 4.77 ;
      RECT 16.34 4.435 17.13 4.605 ;
      RECT 16.34 4.21 16.51 4.605 ;
      RECT 16.24 3.79 16.41 4.38 ;
      RECT 16 3.87 16.41 4.14 ;
      RECT 13.3 10.145 13.47 10.595 ;
      RECT 13.355 8.365 13.525 10.315 ;
      RECT 13.3 7.305 13.47 8.535 ;
      RECT 12.78 7.305 12.95 10.595 ;
      RECT 12.78 9.605 13.185 9.935 ;
      RECT 12.78 8.765 13.185 9.095 ;
      RECT 107.18 10.09 107.35 10.6 ;
      RECT 106.19 1.865 106.36 2.375 ;
      RECT 106.19 3.685 106.36 5.155 ;
      RECT 106.19 7.31 106.36 8.78 ;
      RECT 106.19 10.09 106.36 10.6 ;
      RECT 104.83 1.87 105 5.16 ;
      RECT 104.83 7.305 105 10.595 ;
      RECT 104.4 1.87 104.57 2.38 ;
      RECT 104.4 2.95 104.57 5.16 ;
      RECT 104.4 7.305 104.57 9.515 ;
      RECT 104.4 10.085 104.57 10.595 ;
      RECT 100.72 3.79 100.89 4.24 ;
      RECT 100.48 3.05 100.65 3.4 ;
      RECT 99.52 3.05 99.69 3.4 ;
      RECT 99.215 7.305 99.385 10.595 ;
      RECT 99.04 4.35 99.21 4.77 ;
      RECT 98.785 7.305 98.955 9.515 ;
      RECT 98.785 10.085 98.955 10.595 ;
      RECT 98.04 3.05 98.21 3.4 ;
      RECT 97.08 3.05 97.25 3.4 ;
      RECT 97.08 4.78 97.25 5.11 ;
      RECT 96.56 4.44 96.73 5.08 ;
      RECT 96.08 3.05 96.25 3.4 ;
      RECT 95.84 3.79 96.01 4.12 ;
      RECT 95.36 3.79 95.53 4.12 ;
      RECT 94.12 4.44 94.29 4.8 ;
      RECT 93.64 4.35 93.81 4.77 ;
      RECT 92.92 3.79 93.09 4.24 ;
      RECT 90.96 3.79 91.13 4.12 ;
      RECT 90.24 3.05 90.41 3.4 ;
      RECT 90.24 4.58 90.41 4.94 ;
      RECT 88.62 10.09 88.79 10.6 ;
      RECT 87.63 1.865 87.8 2.375 ;
      RECT 87.63 3.685 87.8 5.155 ;
      RECT 87.63 7.31 87.8 8.78 ;
      RECT 87.63 10.09 87.8 10.6 ;
      RECT 86.27 1.87 86.44 5.16 ;
      RECT 86.27 7.305 86.44 10.595 ;
      RECT 85.84 1.87 86.01 2.38 ;
      RECT 85.84 2.95 86.01 5.16 ;
      RECT 85.84 7.305 86.01 9.515 ;
      RECT 85.84 10.085 86.01 10.595 ;
      RECT 82.16 3.79 82.33 4.24 ;
      RECT 81.92 3.05 82.09 3.4 ;
      RECT 80.96 3.05 81.13 3.4 ;
      RECT 80.655 7.305 80.825 10.595 ;
      RECT 80.48 4.35 80.65 4.77 ;
      RECT 80.225 7.305 80.395 9.515 ;
      RECT 80.225 10.085 80.395 10.595 ;
      RECT 79.48 3.05 79.65 3.4 ;
      RECT 78.52 3.05 78.69 3.4 ;
      RECT 78.52 4.78 78.69 5.11 ;
      RECT 78 4.44 78.17 5.08 ;
      RECT 77.52 3.05 77.69 3.4 ;
      RECT 77.28 3.79 77.45 4.12 ;
      RECT 76.8 3.79 76.97 4.12 ;
      RECT 75.56 4.44 75.73 4.8 ;
      RECT 75.08 4.35 75.25 4.77 ;
      RECT 74.36 3.79 74.53 4.24 ;
      RECT 72.4 3.79 72.57 4.12 ;
      RECT 71.68 3.05 71.85 3.4 ;
      RECT 71.68 4.58 71.85 4.94 ;
      RECT 70.06 10.09 70.23 10.6 ;
      RECT 69.07 1.865 69.24 2.375 ;
      RECT 69.07 3.685 69.24 5.155 ;
      RECT 69.07 7.31 69.24 8.78 ;
      RECT 69.07 10.09 69.24 10.6 ;
      RECT 67.71 1.87 67.88 5.16 ;
      RECT 67.71 7.305 67.88 10.595 ;
      RECT 67.28 1.87 67.45 2.38 ;
      RECT 67.28 2.95 67.45 5.16 ;
      RECT 67.28 7.305 67.45 9.515 ;
      RECT 67.28 10.085 67.45 10.595 ;
      RECT 63.6 3.79 63.77 4.24 ;
      RECT 63.36 3.05 63.53 3.4 ;
      RECT 62.4 3.05 62.57 3.4 ;
      RECT 62.095 7.305 62.265 10.595 ;
      RECT 61.92 4.35 62.09 4.77 ;
      RECT 61.665 7.305 61.835 9.515 ;
      RECT 61.665 10.085 61.835 10.595 ;
      RECT 60.92 3.05 61.09 3.4 ;
      RECT 59.96 3.05 60.13 3.4 ;
      RECT 59.96 4.78 60.13 5.11 ;
      RECT 59.44 4.44 59.61 5.08 ;
      RECT 58.96 3.05 59.13 3.4 ;
      RECT 58.72 3.79 58.89 4.12 ;
      RECT 58.24 3.79 58.41 4.12 ;
      RECT 57 4.44 57.17 4.8 ;
      RECT 56.52 4.35 56.69 4.77 ;
      RECT 55.8 3.79 55.97 4.24 ;
      RECT 53.84 3.79 54.01 4.12 ;
      RECT 53.12 3.05 53.29 3.4 ;
      RECT 53.12 4.58 53.29 4.94 ;
      RECT 51.5 10.09 51.67 10.6 ;
      RECT 50.51 1.865 50.68 2.375 ;
      RECT 50.51 3.685 50.68 5.155 ;
      RECT 50.51 7.31 50.68 8.78 ;
      RECT 50.51 10.09 50.68 10.6 ;
      RECT 49.15 1.87 49.32 5.16 ;
      RECT 49.15 7.305 49.32 10.595 ;
      RECT 48.72 1.87 48.89 2.38 ;
      RECT 48.72 2.95 48.89 5.16 ;
      RECT 48.72 7.305 48.89 9.515 ;
      RECT 48.72 10.085 48.89 10.595 ;
      RECT 45.04 3.79 45.21 4.24 ;
      RECT 44.8 3.05 44.97 3.4 ;
      RECT 43.84 3.05 44.01 3.4 ;
      RECT 43.535 7.305 43.705 10.595 ;
      RECT 43.36 4.35 43.53 4.77 ;
      RECT 43.105 7.305 43.275 9.515 ;
      RECT 43.105 10.085 43.275 10.595 ;
      RECT 42.36 3.05 42.53 3.4 ;
      RECT 41.4 3.05 41.57 3.4 ;
      RECT 41.4 4.78 41.57 5.11 ;
      RECT 40.88 4.44 41.05 5.08 ;
      RECT 40.4 3.05 40.57 3.4 ;
      RECT 40.16 3.79 40.33 4.12 ;
      RECT 39.68 3.79 39.85 4.12 ;
      RECT 38.44 4.44 38.61 4.8 ;
      RECT 37.96 4.35 38.13 4.77 ;
      RECT 37.24 3.79 37.41 4.24 ;
      RECT 35.28 3.79 35.45 4.12 ;
      RECT 34.56 3.05 34.73 3.4 ;
      RECT 34.56 4.58 34.73 4.94 ;
      RECT 32.94 10.09 33.11 10.6 ;
      RECT 31.95 1.865 32.12 2.375 ;
      RECT 31.95 3.685 32.12 5.155 ;
      RECT 31.95 7.31 32.12 8.78 ;
      RECT 31.95 10.09 32.12 10.6 ;
      RECT 30.59 1.87 30.76 5.16 ;
      RECT 30.59 7.305 30.76 10.595 ;
      RECT 30.16 1.87 30.33 2.38 ;
      RECT 30.16 2.95 30.33 5.16 ;
      RECT 30.16 7.305 30.33 9.515 ;
      RECT 30.16 10.085 30.33 10.595 ;
      RECT 26.48 3.79 26.65 4.24 ;
      RECT 26.24 3.05 26.41 3.4 ;
      RECT 25.28 3.05 25.45 3.4 ;
      RECT 24.975 7.305 25.145 10.595 ;
      RECT 24.8 4.35 24.97 4.77 ;
      RECT 24.545 7.305 24.715 9.515 ;
      RECT 24.545 10.085 24.715 10.595 ;
      RECT 23.8 3.05 23.97 3.4 ;
      RECT 22.84 3.05 23.01 3.4 ;
      RECT 22.84 4.78 23.01 5.11 ;
      RECT 22.32 4.44 22.49 5.08 ;
      RECT 21.84 3.05 22.01 3.4 ;
      RECT 21.6 3.79 21.77 4.12 ;
      RECT 21.12 3.79 21.29 4.12 ;
      RECT 19.88 4.44 20.05 4.8 ;
      RECT 19.4 4.35 19.57 4.77 ;
      RECT 18.68 3.79 18.85 4.24 ;
      RECT 16.72 3.79 16.89 4.12 ;
      RECT 16 3.05 16.17 3.4 ;
      RECT 16 4.58 16.17 4.94 ;
      RECT 13.73 7.305 13.9 9.515 ;
      RECT 13.73 10.085 13.9 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  ORIGIN -8.83 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r1 ;
  SIZE 79.095 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 26.34 1.865 26.51 2.375 ;
        RECT 26.34 3.685 26.51 5.155 ;
      LAYER met1 ;
        RECT 26.28 3.655 26.57 3.885 ;
        RECT 26.28 2.175 26.57 2.405 ;
        RECT 26.34 2.175 26.51 3.885 ;
      LAYER mcon ;
        RECT 26.34 3.685 26.51 3.855 ;
        RECT 26.34 2.205 26.51 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 41.6 1.865 41.77 2.375 ;
        RECT 41.6 3.685 41.77 5.155 ;
      LAYER met1 ;
        RECT 41.54 3.655 41.83 3.885 ;
        RECT 41.54 2.175 41.83 2.405 ;
        RECT 41.6 2.175 41.77 3.885 ;
      LAYER mcon ;
        RECT 41.6 3.685 41.77 3.855 ;
        RECT 41.6 2.205 41.77 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 56.86 1.865 57.03 2.375 ;
        RECT 56.86 3.685 57.03 5.155 ;
      LAYER met1 ;
        RECT 56.8 3.655 57.09 3.885 ;
        RECT 56.8 2.175 57.09 2.405 ;
        RECT 56.86 2.175 57.03 3.885 ;
      LAYER mcon ;
        RECT 56.86 3.685 57.03 3.855 ;
        RECT 56.86 2.205 57.03 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 72.12 1.865 72.29 2.375 ;
        RECT 72.12 3.685 72.29 5.155 ;
      LAYER met1 ;
        RECT 72.06 3.655 72.35 3.885 ;
        RECT 72.06 2.175 72.35 2.405 ;
        RECT 72.12 2.175 72.29 3.885 ;
      LAYER mcon ;
        RECT 72.12 3.685 72.29 3.855 ;
        RECT 72.12 2.205 72.29 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 87.38 1.865 87.55 2.375 ;
        RECT 87.38 3.685 87.55 5.155 ;
      LAYER met1 ;
        RECT 87.32 3.655 87.61 3.885 ;
        RECT 87.32 2.175 87.61 2.405 ;
        RECT 87.38 2.175 87.55 3.885 ;
      LAYER mcon ;
        RECT 87.38 3.685 87.55 3.855 ;
        RECT 87.38 2.205 87.55 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 22.11 8.15 22.45 8.5 ;
        RECT 22.11 4 22.45 4.35 ;
        RECT 22.19 4 22.36 8.5 ;
      LAYER li1 ;
        RECT 22.19 2.955 22.36 4.23 ;
        RECT 22.19 8.235 22.36 9.51 ;
        RECT 16.575 8.235 16.745 9.51 ;
      LAYER met1 ;
        RECT 22.11 4.06 22.59 4.23 ;
        RECT 22.11 4 22.45 4.35 ;
        RECT 16.515 8.235 22.59 8.405 ;
        RECT 22.11 8.15 22.45 8.5 ;
        RECT 16.515 8.205 16.805 8.435 ;
      LAYER via1 ;
        RECT 22.21 8.25 22.36 8.4 ;
        RECT 22.21 4.1 22.36 4.25 ;
      LAYER mcon ;
        RECT 16.575 8.235 16.745 8.405 ;
        RECT 22.19 8.235 22.36 8.405 ;
        RECT 22.19 4.06 22.36 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 37.37 8.15 37.71 8.5 ;
        RECT 37.37 4 37.71 4.35 ;
        RECT 37.45 4 37.62 8.5 ;
      LAYER li1 ;
        RECT 37.45 2.955 37.62 4.23 ;
        RECT 37.45 8.235 37.62 9.51 ;
        RECT 31.835 8.235 32.005 9.51 ;
      LAYER met1 ;
        RECT 37.37 4.06 37.85 4.23 ;
        RECT 37.37 4 37.71 4.35 ;
        RECT 31.775 8.235 37.85 8.405 ;
        RECT 37.37 8.15 37.71 8.5 ;
        RECT 31.775 8.205 32.065 8.435 ;
      LAYER via1 ;
        RECT 37.47 8.25 37.62 8.4 ;
        RECT 37.47 4.1 37.62 4.25 ;
      LAYER mcon ;
        RECT 31.835 8.235 32.005 8.405 ;
        RECT 37.45 8.235 37.62 8.405 ;
        RECT 37.45 4.06 37.62 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 52.63 8.15 52.97 8.5 ;
        RECT 52.63 4 52.97 4.35 ;
        RECT 52.71 4 52.88 8.5 ;
      LAYER li1 ;
        RECT 52.71 2.955 52.88 4.23 ;
        RECT 52.71 8.235 52.88 9.51 ;
        RECT 47.095 8.235 47.265 9.51 ;
      LAYER met1 ;
        RECT 52.63 4.06 53.11 4.23 ;
        RECT 52.63 4 52.97 4.35 ;
        RECT 47.035 8.235 53.11 8.405 ;
        RECT 52.63 8.15 52.97 8.5 ;
        RECT 47.035 8.205 47.325 8.435 ;
      LAYER via1 ;
        RECT 52.73 8.25 52.88 8.4 ;
        RECT 52.73 4.1 52.88 4.25 ;
      LAYER mcon ;
        RECT 47.095 8.235 47.265 8.405 ;
        RECT 52.71 8.235 52.88 8.405 ;
        RECT 52.71 4.06 52.88 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 67.89 8.15 68.23 8.5 ;
        RECT 67.89 4 68.23 4.35 ;
        RECT 67.97 4 68.14 8.5 ;
      LAYER li1 ;
        RECT 67.97 2.955 68.14 4.23 ;
        RECT 67.97 8.235 68.14 9.51 ;
        RECT 62.355 8.235 62.525 9.51 ;
      LAYER met1 ;
        RECT 67.89 4.06 68.37 4.23 ;
        RECT 67.89 4 68.23 4.35 ;
        RECT 62.295 8.235 68.37 8.405 ;
        RECT 67.89 8.15 68.23 8.5 ;
        RECT 62.295 8.205 62.585 8.435 ;
      LAYER via1 ;
        RECT 67.99 8.25 68.14 8.4 ;
        RECT 67.99 4.1 68.14 4.25 ;
      LAYER mcon ;
        RECT 62.355 8.235 62.525 8.405 ;
        RECT 67.97 8.235 68.14 8.405 ;
        RECT 67.97 4.06 68.14 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 83.15 8.15 83.49 8.5 ;
        RECT 83.15 4 83.49 4.35 ;
        RECT 83.23 4 83.4 8.5 ;
      LAYER li1 ;
        RECT 83.23 2.955 83.4 4.23 ;
        RECT 83.23 8.235 83.4 9.51 ;
        RECT 77.615 8.235 77.785 9.51 ;
      LAYER met1 ;
        RECT 83.15 4.06 83.63 4.23 ;
        RECT 83.15 4 83.49 4.35 ;
        RECT 77.555 8.235 83.63 8.405 ;
        RECT 83.15 8.15 83.49 8.5 ;
        RECT 77.555 8.205 77.845 8.435 ;
      LAYER via1 ;
        RECT 83.25 8.25 83.4 8.4 ;
        RECT 83.25 4.1 83.4 4.25 ;
      LAYER mcon ;
        RECT 77.615 8.235 77.785 8.405 ;
        RECT 83.23 8.235 83.4 8.405 ;
        RECT 83.23 4.06 83.4 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 9.06 8.235 9.23 9.51 ;
      LAYER met1 ;
        RECT 9 8.235 9.46 8.405 ;
        RECT 9 8.205 9.29 8.435 ;
      LAYER mcon ;
        RECT 9.06 8.235 9.23 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 10.495 6.555 11.3 6.935 ;
      LAYER met2 ;
        RECT 10.685 6.555 11.065 6.935 ;
      LAYER li1 ;
        RECT 8.875 5.435 87.925 7.035 ;
        RECT 73.415 5.43 87.925 7.035 ;
        RECT 85.79 5.425 87.77 7.04 ;
        RECT 86.95 4.695 87.12 7.77 ;
        RECT 85.96 4.695 86.13 7.77 ;
        RECT 83.22 4.7 83.39 7.765 ;
        RECT 80.445 4.93 80.615 7.035 ;
        RECT 78.525 4.93 78.695 7.035 ;
        RECT 77.605 5.43 77.775 7.765 ;
        RECT 77.585 4.93 77.755 7.035 ;
        RECT 76.125 4.93 76.295 7.035 ;
        RECT 74.205 4.93 74.375 7.035 ;
        RECT 58.155 5.43 72.665 7.035 ;
        RECT 70.53 5.425 72.51 7.04 ;
        RECT 71.69 4.695 71.86 7.77 ;
        RECT 70.7 4.695 70.87 7.77 ;
        RECT 67.96 4.7 68.13 7.765 ;
        RECT 65.185 4.93 65.355 7.035 ;
        RECT 63.265 4.93 63.435 7.035 ;
        RECT 62.345 5.43 62.515 7.765 ;
        RECT 62.325 4.93 62.495 7.035 ;
        RECT 60.865 4.93 61.035 7.035 ;
        RECT 58.945 4.93 59.115 7.035 ;
        RECT 42.895 5.43 57.405 7.035 ;
        RECT 55.27 5.425 57.25 7.04 ;
        RECT 56.43 4.695 56.6 7.77 ;
        RECT 55.44 4.695 55.61 7.77 ;
        RECT 52.7 4.7 52.87 7.765 ;
        RECT 49.925 4.93 50.095 7.035 ;
        RECT 48.005 4.93 48.175 7.035 ;
        RECT 47.085 5.43 47.255 7.765 ;
        RECT 47.065 4.93 47.235 7.035 ;
        RECT 45.605 4.93 45.775 7.035 ;
        RECT 43.685 4.93 43.855 7.035 ;
        RECT 27.635 5.43 42.145 7.035 ;
        RECT 40.01 5.425 41.99 7.04 ;
        RECT 41.17 4.695 41.34 7.77 ;
        RECT 40.18 4.695 40.35 7.77 ;
        RECT 37.44 4.7 37.61 7.765 ;
        RECT 34.665 4.93 34.835 7.035 ;
        RECT 32.745 4.93 32.915 7.035 ;
        RECT 31.825 5.43 31.995 7.765 ;
        RECT 31.805 4.93 31.975 7.035 ;
        RECT 30.345 4.93 30.515 7.035 ;
        RECT 28.425 4.93 28.595 7.035 ;
        RECT 12.375 5.43 26.885 7.035 ;
        RECT 24.75 5.425 26.73 7.04 ;
        RECT 25.91 4.695 26.08 7.77 ;
        RECT 24.92 4.695 25.09 7.77 ;
        RECT 22.18 4.7 22.35 7.765 ;
        RECT 19.405 4.93 19.575 7.035 ;
        RECT 17.485 4.93 17.655 7.035 ;
        RECT 16.565 5.43 16.735 7.765 ;
        RECT 16.545 4.93 16.715 7.035 ;
        RECT 15.085 4.93 15.255 7.035 ;
        RECT 13.165 4.93 13.335 7.035 ;
        RECT 10.86 5.435 11.03 10.595 ;
        RECT 9.05 5.435 9.22 7.765 ;
      LAYER met1 ;
        RECT 8.875 5.435 87.925 7.035 ;
        RECT 73.415 5.43 87.925 7.035 ;
        RECT 85.79 5.425 87.77 7.04 ;
        RECT 73.415 5.275 82.155 7.035 ;
        RECT 58.155 5.43 72.665 7.035 ;
        RECT 70.53 5.425 72.51 7.04 ;
        RECT 58.155 5.275 66.895 7.035 ;
        RECT 42.895 5.43 57.405 7.035 ;
        RECT 55.27 5.425 57.25 7.04 ;
        RECT 42.895 5.275 51.635 7.035 ;
        RECT 27.635 5.43 42.145 7.035 ;
        RECT 40.01 5.425 41.99 7.04 ;
        RECT 27.635 5.275 36.375 7.035 ;
        RECT 12.375 5.43 26.885 7.035 ;
        RECT 24.75 5.425 26.73 7.04 ;
        RECT 12.375 5.275 21.115 7.035 ;
        RECT 10.8 8.945 11.09 9.175 ;
        RECT 10.63 8.975 11.09 9.145 ;
      LAYER via2 ;
        RECT 10.775 6.645 10.975 6.845 ;
      LAYER via1 ;
        RECT 10.8 6.67 10.95 6.82 ;
      LAYER mcon ;
        RECT 10.86 8.975 11.03 9.145 ;
        RECT 11.17 6.835 11.34 7.005 ;
        RECT 12.52 5.43 12.69 5.6 ;
        RECT 12.98 5.43 13.15 5.6 ;
        RECT 13.44 5.43 13.61 5.6 ;
        RECT 13.9 5.43 14.07 5.6 ;
        RECT 14.36 5.43 14.53 5.6 ;
        RECT 14.82 5.43 14.99 5.6 ;
        RECT 15.28 5.43 15.45 5.6 ;
        RECT 15.74 5.43 15.91 5.6 ;
        RECT 16.2 5.43 16.37 5.6 ;
        RECT 16.66 5.43 16.83 5.6 ;
        RECT 17.12 5.43 17.29 5.6 ;
        RECT 17.58 5.43 17.75 5.6 ;
        RECT 18.04 5.43 18.21 5.6 ;
        RECT 18.5 5.43 18.67 5.6 ;
        RECT 18.685 6.835 18.855 7.005 ;
        RECT 18.96 5.43 19.13 5.6 ;
        RECT 19.42 5.43 19.59 5.6 ;
        RECT 19.88 5.43 20.05 5.6 ;
        RECT 20.34 5.43 20.51 5.6 ;
        RECT 20.8 5.43 20.97 5.6 ;
        RECT 24.3 6.835 24.47 7.005 ;
        RECT 24.3 5.46 24.47 5.63 ;
        RECT 25 6.84 25.17 7.01 ;
        RECT 25 5.455 25.17 5.625 ;
        RECT 25.99 6.84 26.16 7.01 ;
        RECT 25.99 5.455 26.16 5.625 ;
        RECT 27.78 5.43 27.95 5.6 ;
        RECT 28.24 5.43 28.41 5.6 ;
        RECT 28.7 5.43 28.87 5.6 ;
        RECT 29.16 5.43 29.33 5.6 ;
        RECT 29.62 5.43 29.79 5.6 ;
        RECT 30.08 5.43 30.25 5.6 ;
        RECT 30.54 5.43 30.71 5.6 ;
        RECT 31 5.43 31.17 5.6 ;
        RECT 31.46 5.43 31.63 5.6 ;
        RECT 31.92 5.43 32.09 5.6 ;
        RECT 32.38 5.43 32.55 5.6 ;
        RECT 32.84 5.43 33.01 5.6 ;
        RECT 33.3 5.43 33.47 5.6 ;
        RECT 33.76 5.43 33.93 5.6 ;
        RECT 33.945 6.835 34.115 7.005 ;
        RECT 34.22 5.43 34.39 5.6 ;
        RECT 34.68 5.43 34.85 5.6 ;
        RECT 35.14 5.43 35.31 5.6 ;
        RECT 35.6 5.43 35.77 5.6 ;
        RECT 36.06 5.43 36.23 5.6 ;
        RECT 39.56 6.835 39.73 7.005 ;
        RECT 39.56 5.46 39.73 5.63 ;
        RECT 40.26 6.84 40.43 7.01 ;
        RECT 40.26 5.455 40.43 5.625 ;
        RECT 41.25 6.84 41.42 7.01 ;
        RECT 41.25 5.455 41.42 5.625 ;
        RECT 43.04 5.43 43.21 5.6 ;
        RECT 43.5 5.43 43.67 5.6 ;
        RECT 43.96 5.43 44.13 5.6 ;
        RECT 44.42 5.43 44.59 5.6 ;
        RECT 44.88 5.43 45.05 5.6 ;
        RECT 45.34 5.43 45.51 5.6 ;
        RECT 45.8 5.43 45.97 5.6 ;
        RECT 46.26 5.43 46.43 5.6 ;
        RECT 46.72 5.43 46.89 5.6 ;
        RECT 47.18 5.43 47.35 5.6 ;
        RECT 47.64 5.43 47.81 5.6 ;
        RECT 48.1 5.43 48.27 5.6 ;
        RECT 48.56 5.43 48.73 5.6 ;
        RECT 49.02 5.43 49.19 5.6 ;
        RECT 49.205 6.835 49.375 7.005 ;
        RECT 49.48 5.43 49.65 5.6 ;
        RECT 49.94 5.43 50.11 5.6 ;
        RECT 50.4 5.43 50.57 5.6 ;
        RECT 50.86 5.43 51.03 5.6 ;
        RECT 51.32 5.43 51.49 5.6 ;
        RECT 54.82 6.835 54.99 7.005 ;
        RECT 54.82 5.46 54.99 5.63 ;
        RECT 55.52 6.84 55.69 7.01 ;
        RECT 55.52 5.455 55.69 5.625 ;
        RECT 56.51 6.84 56.68 7.01 ;
        RECT 56.51 5.455 56.68 5.625 ;
        RECT 58.3 5.43 58.47 5.6 ;
        RECT 58.76 5.43 58.93 5.6 ;
        RECT 59.22 5.43 59.39 5.6 ;
        RECT 59.68 5.43 59.85 5.6 ;
        RECT 60.14 5.43 60.31 5.6 ;
        RECT 60.6 5.43 60.77 5.6 ;
        RECT 61.06 5.43 61.23 5.6 ;
        RECT 61.52 5.43 61.69 5.6 ;
        RECT 61.98 5.43 62.15 5.6 ;
        RECT 62.44 5.43 62.61 5.6 ;
        RECT 62.9 5.43 63.07 5.6 ;
        RECT 63.36 5.43 63.53 5.6 ;
        RECT 63.82 5.43 63.99 5.6 ;
        RECT 64.28 5.43 64.45 5.6 ;
        RECT 64.465 6.835 64.635 7.005 ;
        RECT 64.74 5.43 64.91 5.6 ;
        RECT 65.2 5.43 65.37 5.6 ;
        RECT 65.66 5.43 65.83 5.6 ;
        RECT 66.12 5.43 66.29 5.6 ;
        RECT 66.58 5.43 66.75 5.6 ;
        RECT 70.08 6.835 70.25 7.005 ;
        RECT 70.08 5.46 70.25 5.63 ;
        RECT 70.78 6.84 70.95 7.01 ;
        RECT 70.78 5.455 70.95 5.625 ;
        RECT 71.77 6.84 71.94 7.01 ;
        RECT 71.77 5.455 71.94 5.625 ;
        RECT 73.56 5.43 73.73 5.6 ;
        RECT 74.02 5.43 74.19 5.6 ;
        RECT 74.48 5.43 74.65 5.6 ;
        RECT 74.94 5.43 75.11 5.6 ;
        RECT 75.4 5.43 75.57 5.6 ;
        RECT 75.86 5.43 76.03 5.6 ;
        RECT 76.32 5.43 76.49 5.6 ;
        RECT 76.78 5.43 76.95 5.6 ;
        RECT 77.24 5.43 77.41 5.6 ;
        RECT 77.7 5.43 77.87 5.6 ;
        RECT 78.16 5.43 78.33 5.6 ;
        RECT 78.62 5.43 78.79 5.6 ;
        RECT 79.08 5.43 79.25 5.6 ;
        RECT 79.54 5.43 79.71 5.6 ;
        RECT 79.725 6.835 79.895 7.005 ;
        RECT 80 5.43 80.17 5.6 ;
        RECT 80.46 5.43 80.63 5.6 ;
        RECT 80.92 5.43 81.09 5.6 ;
        RECT 81.38 5.43 81.55 5.6 ;
        RECT 81.84 5.43 82.01 5.6 ;
        RECT 85.34 6.835 85.51 7.005 ;
        RECT 85.34 5.46 85.51 5.63 ;
        RECT 86.04 6.84 86.21 7.01 ;
        RECT 86.04 5.455 86.21 5.625 ;
        RECT 87.03 6.84 87.2 7.01 ;
        RECT 87.03 5.455 87.2 5.625 ;
    END
  END vccd1
  OBS
    LAYER met4 ;
      RECT 75.565 4.27 75.895 4.6 ;
      RECT 75.58 3.795 75.895 4.6 ;
      RECT 77.725 3.78 78.055 4.135 ;
      RECT 75.58 3.795 78.055 4.095 ;
      RECT 60.305 4.27 60.635 4.6 ;
      RECT 60.32 3.795 60.635 4.6 ;
      RECT 62.465 3.78 62.795 4.135 ;
      RECT 60.32 3.795 62.795 4.095 ;
      RECT 45.045 4.27 45.375 4.6 ;
      RECT 45.06 3.795 45.375 4.6 ;
      RECT 47.205 3.78 47.535 4.135 ;
      RECT 45.06 3.795 47.535 4.095 ;
      RECT 29.785 4.27 30.115 4.6 ;
      RECT 29.8 3.795 30.115 4.6 ;
      RECT 31.945 3.78 32.275 4.135 ;
      RECT 29.8 3.795 32.275 4.095 ;
      RECT 14.525 4.27 14.855 4.6 ;
      RECT 14.54 3.795 14.855 4.6 ;
      RECT 16.685 3.78 17.015 4.135 ;
      RECT 14.54 3.795 17.015 4.095 ;
    LAYER via3 ;
      RECT 77.79 3.87 77.99 4.07 ;
      RECT 75.63 4.335 75.83 4.535 ;
      RECT 62.53 3.87 62.73 4.07 ;
      RECT 60.37 4.335 60.57 4.535 ;
      RECT 47.27 3.87 47.47 4.07 ;
      RECT 45.11 4.335 45.31 4.535 ;
      RECT 32.01 3.87 32.21 4.07 ;
      RECT 29.85 4.335 30.05 4.535 ;
      RECT 16.75 3.87 16.95 4.07 ;
      RECT 14.59 4.335 14.79 4.535 ;
    LAYER met3 ;
      RECT 78.885 9.345 79.255 9.715 ;
      RECT 78.92 5.77 79.22 9.715 ;
      RECT 77.48 5.77 79.22 7.065 ;
      RECT 74.685 5.55 77.78 6.845 ;
      RECT 77.48 3.81 77.78 7.065 ;
      RECT 74.685 4.27 74.985 6.845 ;
      RECT 78.205 4.805 78.535 5.16 ;
      RECT 76.3 4.845 78.535 5.145 ;
      RECT 76.3 3.71 76.6 5.145 ;
      RECT 74.38 4.27 75.11 4.6 ;
      RECT 77.275 3.815 78.055 4.16 ;
      RECT 77.75 3.78 78.055 4.16 ;
      RECT 76.285 3.71 76.615 4.04 ;
      RECT 75.57 3.71 75.89 4.625 ;
      RECT 75.57 3.71 75.9 4.245 ;
      RECT 63.625 9.345 63.995 9.715 ;
      RECT 63.66 5.77 63.96 9.715 ;
      RECT 62.22 5.77 63.96 7.065 ;
      RECT 59.425 5.55 62.52 6.845 ;
      RECT 62.22 3.81 62.52 7.065 ;
      RECT 59.425 4.27 59.725 6.845 ;
      RECT 62.945 4.805 63.275 5.16 ;
      RECT 61.04 4.845 63.275 5.145 ;
      RECT 61.04 3.71 61.34 5.145 ;
      RECT 59.12 4.27 59.85 4.6 ;
      RECT 62.015 3.815 62.795 4.16 ;
      RECT 62.49 3.78 62.795 4.16 ;
      RECT 61.025 3.71 61.355 4.04 ;
      RECT 60.31 3.71 60.63 4.625 ;
      RECT 60.31 3.71 60.64 4.245 ;
      RECT 48.365 9.345 48.735 9.715 ;
      RECT 48.4 5.77 48.7 9.715 ;
      RECT 46.96 5.77 48.7 7.065 ;
      RECT 44.165 5.55 47.26 6.845 ;
      RECT 46.96 3.81 47.26 7.065 ;
      RECT 44.165 4.27 44.465 6.845 ;
      RECT 47.685 4.805 48.015 5.16 ;
      RECT 45.78 4.845 48.015 5.145 ;
      RECT 45.78 3.71 46.08 5.145 ;
      RECT 43.86 4.27 44.59 4.6 ;
      RECT 46.755 3.815 47.535 4.16 ;
      RECT 47.23 3.78 47.535 4.16 ;
      RECT 45.765 3.71 46.095 4.04 ;
      RECT 45.05 3.71 45.37 4.625 ;
      RECT 45.05 3.71 45.38 4.245 ;
      RECT 33.105 9.345 33.475 9.715 ;
      RECT 33.14 5.77 33.44 9.715 ;
      RECT 31.7 5.77 33.44 7.065 ;
      RECT 28.905 5.55 32 6.845 ;
      RECT 31.7 3.81 32 7.065 ;
      RECT 28.905 4.27 29.205 6.845 ;
      RECT 32.425 4.805 32.755 5.16 ;
      RECT 30.52 4.845 32.755 5.145 ;
      RECT 30.52 3.71 30.82 5.145 ;
      RECT 28.6 4.27 29.33 4.6 ;
      RECT 31.495 3.815 32.275 4.16 ;
      RECT 31.97 3.78 32.275 4.16 ;
      RECT 30.505 3.71 30.835 4.04 ;
      RECT 29.79 3.71 30.11 4.625 ;
      RECT 29.79 3.71 30.12 4.245 ;
      RECT 17.845 9.345 18.215 9.715 ;
      RECT 17.88 5.77 18.18 9.715 ;
      RECT 16.44 5.77 18.18 7.065 ;
      RECT 13.645 5.55 16.74 6.845 ;
      RECT 16.44 3.81 16.74 7.065 ;
      RECT 13.645 4.27 13.945 6.845 ;
      RECT 17.165 4.805 17.495 5.16 ;
      RECT 15.26 4.845 17.495 5.145 ;
      RECT 15.26 3.71 15.56 5.145 ;
      RECT 13.34 4.27 14.07 4.6 ;
      RECT 16.235 3.815 17.015 4.16 ;
      RECT 16.71 3.78 17.015 4.16 ;
      RECT 15.245 3.71 15.575 4.04 ;
      RECT 14.53 3.71 14.85 4.625 ;
      RECT 14.53 3.71 14.86 4.245 ;
      RECT 81.125 3.15 81.855 3.48 ;
      RECT 79.435 3.165 80.165 3.495 ;
      RECT 78.4 3.15 79.13 3.5 ;
      RECT 76.85 3.175 77.58 3.505 ;
      RECT 74.245 3.15 74.975 3.48 ;
      RECT 65.865 3.15 66.595 3.48 ;
      RECT 64.175 3.165 64.905 3.495 ;
      RECT 63.14 3.15 63.87 3.5 ;
      RECT 61.59 3.175 62.32 3.505 ;
      RECT 58.985 3.15 59.715 3.48 ;
      RECT 50.605 3.15 51.335 3.48 ;
      RECT 48.915 3.165 49.645 3.495 ;
      RECT 47.88 3.15 48.61 3.5 ;
      RECT 46.33 3.175 47.06 3.505 ;
      RECT 43.725 3.15 44.455 3.48 ;
      RECT 35.345 3.15 36.075 3.48 ;
      RECT 33.655 3.165 34.385 3.495 ;
      RECT 32.62 3.15 33.35 3.5 ;
      RECT 31.07 3.175 31.8 3.505 ;
      RECT 28.465 3.15 29.195 3.48 ;
      RECT 20.085 3.15 20.815 3.48 ;
      RECT 18.395 3.165 19.125 3.495 ;
      RECT 17.36 3.15 18.09 3.5 ;
      RECT 15.81 3.175 16.54 3.505 ;
      RECT 13.205 3.15 13.935 3.48 ;
    LAYER via2 ;
      RECT 81.36 3.215 81.56 3.415 ;
      RECT 79.5 3.23 79.7 3.43 ;
      RECT 78.97 9.43 79.17 9.63 ;
      RECT 78.48 3.235 78.68 3.435 ;
      RECT 78.27 4.87 78.47 5.07 ;
      RECT 77.79 3.87 77.99 4.07 ;
      RECT 77.04 3.24 77.24 3.44 ;
      RECT 76.35 3.775 76.55 3.975 ;
      RECT 75.635 3.775 75.835 3.975 ;
      RECT 74.67 4.335 74.87 4.535 ;
      RECT 74.43 3.215 74.63 3.415 ;
      RECT 66.1 3.215 66.3 3.415 ;
      RECT 64.24 3.23 64.44 3.43 ;
      RECT 63.71 9.43 63.91 9.63 ;
      RECT 63.22 3.235 63.42 3.435 ;
      RECT 63.01 4.87 63.21 5.07 ;
      RECT 62.53 3.87 62.73 4.07 ;
      RECT 61.78 3.24 61.98 3.44 ;
      RECT 61.09 3.775 61.29 3.975 ;
      RECT 60.375 3.775 60.575 3.975 ;
      RECT 59.41 4.335 59.61 4.535 ;
      RECT 59.17 3.215 59.37 3.415 ;
      RECT 50.84 3.215 51.04 3.415 ;
      RECT 48.98 3.23 49.18 3.43 ;
      RECT 48.45 9.43 48.65 9.63 ;
      RECT 47.96 3.235 48.16 3.435 ;
      RECT 47.75 4.87 47.95 5.07 ;
      RECT 47.27 3.87 47.47 4.07 ;
      RECT 46.52 3.24 46.72 3.44 ;
      RECT 45.83 3.775 46.03 3.975 ;
      RECT 45.115 3.775 45.315 3.975 ;
      RECT 44.15 4.335 44.35 4.535 ;
      RECT 43.91 3.215 44.11 3.415 ;
      RECT 35.58 3.215 35.78 3.415 ;
      RECT 33.72 3.23 33.92 3.43 ;
      RECT 33.19 9.43 33.39 9.63 ;
      RECT 32.7 3.235 32.9 3.435 ;
      RECT 32.49 4.87 32.69 5.07 ;
      RECT 32.01 3.87 32.21 4.07 ;
      RECT 31.26 3.24 31.46 3.44 ;
      RECT 30.57 3.775 30.77 3.975 ;
      RECT 29.855 3.775 30.055 3.975 ;
      RECT 28.89 4.335 29.09 4.535 ;
      RECT 28.65 3.215 28.85 3.415 ;
      RECT 20.32 3.215 20.52 3.415 ;
      RECT 18.46 3.23 18.66 3.43 ;
      RECT 17.93 9.43 18.13 9.63 ;
      RECT 17.44 3.235 17.64 3.435 ;
      RECT 17.23 4.87 17.43 5.07 ;
      RECT 16.75 3.87 16.95 4.07 ;
      RECT 16 3.24 16.2 3.44 ;
      RECT 15.31 3.775 15.51 3.975 ;
      RECT 14.595 3.775 14.795 3.975 ;
      RECT 13.63 4.335 13.83 4.535 ;
      RECT 13.39 3.215 13.59 3.415 ;
    LAYER met2 ;
      RECT 10.055 10.69 87.555 10.86 ;
      RECT 87.385 9.565 87.555 10.86 ;
      RECT 10.055 8.545 10.225 10.86 ;
      RECT 87.355 9.565 87.705 9.915 ;
      RECT 9.995 8.545 10.285 8.895 ;
      RECT 84.195 8.51 84.515 8.835 ;
      RECT 84.225 7.985 84.395 8.835 ;
      RECT 84.225 7.985 84.4 8.335 ;
      RECT 84.225 7.985 85.2 8.16 ;
      RECT 85.025 3.26 85.2 8.16 ;
      RECT 84.97 3.26 85.32 3.61 ;
      RECT 84.995 8.945 85.32 9.27 ;
      RECT 83.88 9.035 85.32 9.205 ;
      RECT 83.88 3.69 84.04 9.205 ;
      RECT 84.195 3.66 84.515 3.98 ;
      RECT 83.88 3.69 84.515 3.86 ;
      RECT 81.33 4.835 81.59 5.155 ;
      RECT 81.39 3.13 81.53 5.155 ;
      RECT 82.59 3.995 82.93 4.345 ;
      RECT 81.965 4.065 82.93 4.265 ;
      RECT 81.965 3.235 82.165 4.265 ;
      RECT 81.215 3.69 81.53 4.06 ;
      RECT 82.68 3.99 82.85 4.345 ;
      RECT 81.285 3.245 81.53 4.06 ;
      RECT 81.32 3.13 81.6 3.5 ;
      RECT 81.32 3.235 82.165 3.435 ;
      RECT 80.64 3.715 80.9 4.035 ;
      RECT 79.98 3.805 80.9 3.945 ;
      RECT 79.98 2.865 80.12 3.945 ;
      RECT 76.44 3.155 76.7 3.475 ;
      RECT 76.62 2.865 76.76 3.385 ;
      RECT 76.62 2.865 80.12 3.005 ;
      RECT 72.07 8.945 72.42 9.295 ;
      RECT 79.555 8.9 79.905 9.25 ;
      RECT 72.07 8.975 79.905 9.175 ;
      RECT 79.47 4.555 79.73 4.875 ;
      RECT 79.53 3.145 79.67 4.875 ;
      RECT 79.46 3.145 79.74 3.515 ;
      RECT 76.86 5.305 79.295 5.445 ;
      RECT 79.155 3.995 79.295 5.445 ;
      RECT 76.86 4.925 77 5.445 ;
      RECT 76.56 4.925 77 5.155 ;
      RECT 74.22 4.925 77 5.065 ;
      RECT 76.56 4.835 76.82 5.155 ;
      RECT 74.22 4.645 74.36 5.065 ;
      RECT 73.71 4.555 73.97 4.875 ;
      RECT 73.71 4.645 74.36 4.785 ;
      RECT 73.77 3.155 73.91 4.875 ;
      RECT 79.095 3.995 79.355 4.315 ;
      RECT 73.71 3.155 73.97 3.475 ;
      RECT 78.72 4.835 78.98 5.155 ;
      RECT 78.78 3.245 78.92 5.155 ;
      RECT 78.44 3.245 78.92 3.52 ;
      RECT 78.24 3.15 78.72 3.495 ;
      RECT 78.23 4.785 78.51 5.155 ;
      RECT 78.3 3.69 78.44 5.155 ;
      RECT 78.24 3.69 78.5 4.315 ;
      RECT 78.23 3.69 78.51 4.06 ;
      RECT 77.16 4.835 77.42 5.155 ;
      RECT 77.16 4.645 77.36 5.155 ;
      RECT 76.965 4.645 77.36 4.785 ;
      RECT 76.965 3.155 77.105 4.785 ;
      RECT 76.965 3.155 77.28 3.525 ;
      RECT 76.905 3.155 77.28 3.475 ;
      RECT 74.63 4.25 74.91 4.62 ;
      RECT 76.08 4.275 76.34 4.595 ;
      RECT 74.46 4.365 76.34 4.505 ;
      RECT 74.46 4.25 74.91 4.505 ;
      RECT 74.4 3.69 74.66 4.315 ;
      RECT 74.39 3.69 74.67 4.06 ;
      RECT 75.47 3.69 75.88 4.06 ;
      RECT 74.88 3.715 75.14 4.035 ;
      RECT 74.88 3.805 75.88 3.945 ;
      RECT 74.39 3.13 74.67 3.5 ;
      RECT 74.39 3.155 74.78 3.475 ;
      RECT 68.935 8.51 69.255 8.835 ;
      RECT 68.965 7.985 69.135 8.835 ;
      RECT 68.965 7.985 69.14 8.335 ;
      RECT 68.965 7.985 69.94 8.16 ;
      RECT 69.765 3.26 69.94 8.16 ;
      RECT 69.71 3.26 70.06 3.61 ;
      RECT 69.735 8.945 70.06 9.27 ;
      RECT 68.62 9.035 70.06 9.205 ;
      RECT 68.62 3.69 68.78 9.205 ;
      RECT 68.935 3.66 69.255 3.98 ;
      RECT 68.62 3.69 69.255 3.86 ;
      RECT 66.07 4.835 66.33 5.155 ;
      RECT 66.13 3.13 66.27 5.155 ;
      RECT 67.33 3.995 67.67 4.345 ;
      RECT 66.705 4.065 67.67 4.265 ;
      RECT 66.705 3.235 66.905 4.265 ;
      RECT 65.955 3.69 66.27 4.06 ;
      RECT 67.42 3.99 67.59 4.345 ;
      RECT 66.025 3.245 66.27 4.06 ;
      RECT 66.06 3.13 66.34 3.5 ;
      RECT 66.06 3.235 66.905 3.435 ;
      RECT 65.38 3.715 65.64 4.035 ;
      RECT 64.72 3.805 65.64 3.945 ;
      RECT 64.72 2.865 64.86 3.945 ;
      RECT 61.18 3.155 61.44 3.475 ;
      RECT 61.36 2.865 61.5 3.385 ;
      RECT 61.36 2.865 64.86 3.005 ;
      RECT 56.81 8.945 57.16 9.295 ;
      RECT 64.3 8.9 64.65 9.25 ;
      RECT 56.81 8.975 64.65 9.175 ;
      RECT 64.21 4.555 64.47 4.875 ;
      RECT 64.27 3.145 64.41 4.875 ;
      RECT 64.2 3.145 64.48 3.515 ;
      RECT 61.6 5.305 64.035 5.445 ;
      RECT 63.895 3.995 64.035 5.445 ;
      RECT 61.6 4.925 61.74 5.445 ;
      RECT 61.3 4.925 61.74 5.155 ;
      RECT 58.96 4.925 61.74 5.065 ;
      RECT 61.3 4.835 61.56 5.155 ;
      RECT 58.96 4.645 59.1 5.065 ;
      RECT 58.45 4.555 58.71 4.875 ;
      RECT 58.45 4.645 59.1 4.785 ;
      RECT 58.51 3.155 58.65 4.875 ;
      RECT 63.835 3.995 64.095 4.315 ;
      RECT 58.45 3.155 58.71 3.475 ;
      RECT 63.46 4.835 63.72 5.155 ;
      RECT 63.52 3.245 63.66 5.155 ;
      RECT 63.18 3.245 63.66 3.52 ;
      RECT 62.98 3.15 63.46 3.495 ;
      RECT 62.97 4.785 63.25 5.155 ;
      RECT 63.04 3.69 63.18 5.155 ;
      RECT 62.98 3.69 63.24 4.315 ;
      RECT 62.97 3.69 63.25 4.06 ;
      RECT 61.9 4.835 62.16 5.155 ;
      RECT 61.9 4.645 62.1 5.155 ;
      RECT 61.705 4.645 62.1 4.785 ;
      RECT 61.705 3.155 61.845 4.785 ;
      RECT 61.705 3.155 62.02 3.525 ;
      RECT 61.645 3.155 62.02 3.475 ;
      RECT 59.37 4.25 59.65 4.62 ;
      RECT 60.82 4.275 61.08 4.595 ;
      RECT 59.2 4.365 61.08 4.505 ;
      RECT 59.2 4.25 59.65 4.505 ;
      RECT 59.14 3.69 59.4 4.315 ;
      RECT 59.13 3.69 59.41 4.06 ;
      RECT 60.21 3.69 60.62 4.06 ;
      RECT 59.62 3.715 59.88 4.035 ;
      RECT 59.62 3.805 60.62 3.945 ;
      RECT 59.13 3.13 59.41 3.5 ;
      RECT 59.13 3.155 59.52 3.475 ;
      RECT 53.675 8.51 53.995 8.835 ;
      RECT 53.705 7.985 53.875 8.835 ;
      RECT 53.705 7.985 53.88 8.335 ;
      RECT 53.705 7.985 54.68 8.16 ;
      RECT 54.505 3.26 54.68 8.16 ;
      RECT 54.45 3.26 54.8 3.61 ;
      RECT 54.475 8.945 54.8 9.27 ;
      RECT 53.36 9.035 54.8 9.205 ;
      RECT 53.36 3.69 53.52 9.205 ;
      RECT 53.675 3.66 53.995 3.98 ;
      RECT 53.36 3.69 53.995 3.86 ;
      RECT 50.81 4.835 51.07 5.155 ;
      RECT 50.87 3.13 51.01 5.155 ;
      RECT 52.07 3.995 52.41 4.345 ;
      RECT 51.445 4.065 52.41 4.265 ;
      RECT 51.445 3.235 51.645 4.265 ;
      RECT 50.695 3.69 51.01 4.06 ;
      RECT 52.16 3.99 52.33 4.345 ;
      RECT 50.765 3.245 51.01 4.06 ;
      RECT 50.8 3.13 51.08 3.5 ;
      RECT 50.8 3.235 51.645 3.435 ;
      RECT 50.12 3.715 50.38 4.035 ;
      RECT 49.46 3.805 50.38 3.945 ;
      RECT 49.46 2.865 49.6 3.945 ;
      RECT 45.92 3.155 46.18 3.475 ;
      RECT 46.1 2.865 46.24 3.385 ;
      RECT 46.1 2.865 49.6 3.005 ;
      RECT 41.595 8.95 41.945 9.3 ;
      RECT 49.035 8.905 49.385 9.255 ;
      RECT 41.595 8.98 49.385 9.18 ;
      RECT 48.95 4.555 49.21 4.875 ;
      RECT 49.01 3.145 49.15 4.875 ;
      RECT 48.94 3.145 49.22 3.515 ;
      RECT 46.34 5.305 48.775 5.445 ;
      RECT 48.635 3.995 48.775 5.445 ;
      RECT 46.34 4.925 46.48 5.445 ;
      RECT 46.04 4.925 46.48 5.155 ;
      RECT 43.7 4.925 46.48 5.065 ;
      RECT 46.04 4.835 46.3 5.155 ;
      RECT 43.7 4.645 43.84 5.065 ;
      RECT 43.19 4.555 43.45 4.875 ;
      RECT 43.19 4.645 43.84 4.785 ;
      RECT 43.25 3.155 43.39 4.875 ;
      RECT 48.575 3.995 48.835 4.315 ;
      RECT 43.19 3.155 43.45 3.475 ;
      RECT 48.2 4.835 48.46 5.155 ;
      RECT 48.26 3.245 48.4 5.155 ;
      RECT 47.92 3.245 48.4 3.52 ;
      RECT 47.72 3.15 48.2 3.495 ;
      RECT 47.71 4.785 47.99 5.155 ;
      RECT 47.78 3.69 47.92 5.155 ;
      RECT 47.72 3.69 47.98 4.315 ;
      RECT 47.71 3.69 47.99 4.06 ;
      RECT 46.64 4.835 46.9 5.155 ;
      RECT 46.64 4.645 46.84 5.155 ;
      RECT 46.445 4.645 46.84 4.785 ;
      RECT 46.445 3.155 46.585 4.785 ;
      RECT 46.445 3.155 46.76 3.525 ;
      RECT 46.385 3.155 46.76 3.475 ;
      RECT 44.11 4.25 44.39 4.62 ;
      RECT 45.56 4.275 45.82 4.595 ;
      RECT 43.94 4.365 45.82 4.505 ;
      RECT 43.94 4.25 44.39 4.505 ;
      RECT 43.88 3.69 44.14 4.315 ;
      RECT 43.87 3.69 44.15 4.06 ;
      RECT 44.95 3.69 45.36 4.06 ;
      RECT 44.36 3.715 44.62 4.035 ;
      RECT 44.36 3.805 45.36 3.945 ;
      RECT 43.87 3.13 44.15 3.5 ;
      RECT 43.87 3.155 44.26 3.475 ;
      RECT 38.415 8.51 38.735 8.835 ;
      RECT 38.445 7.985 38.615 8.835 ;
      RECT 38.445 7.985 38.62 8.335 ;
      RECT 38.445 7.985 39.42 8.16 ;
      RECT 39.245 3.26 39.42 8.16 ;
      RECT 39.19 3.26 39.54 3.61 ;
      RECT 39.215 8.945 39.54 9.27 ;
      RECT 38.1 9.035 39.54 9.205 ;
      RECT 38.1 3.69 38.26 9.205 ;
      RECT 38.415 3.66 38.735 3.98 ;
      RECT 38.1 3.69 38.735 3.86 ;
      RECT 35.55 4.835 35.81 5.155 ;
      RECT 35.61 3.13 35.75 5.155 ;
      RECT 36.81 3.995 37.15 4.345 ;
      RECT 36.185 4.065 37.15 4.265 ;
      RECT 36.185 3.235 36.385 4.265 ;
      RECT 35.435 3.69 35.75 4.06 ;
      RECT 36.9 3.99 37.07 4.345 ;
      RECT 35.505 3.245 35.75 4.06 ;
      RECT 35.54 3.13 35.82 3.5 ;
      RECT 35.54 3.235 36.385 3.435 ;
      RECT 34.86 3.715 35.12 4.035 ;
      RECT 34.2 3.805 35.12 3.945 ;
      RECT 34.2 2.865 34.34 3.945 ;
      RECT 30.66 3.155 30.92 3.475 ;
      RECT 30.84 2.865 30.98 3.385 ;
      RECT 30.84 2.865 34.34 3.005 ;
      RECT 26.335 8.945 26.685 9.295 ;
      RECT 33.775 8.9 34.125 9.25 ;
      RECT 26.335 8.975 34.125 9.175 ;
      RECT 33.69 4.555 33.95 4.875 ;
      RECT 33.75 3.145 33.89 4.875 ;
      RECT 33.68 3.145 33.96 3.515 ;
      RECT 31.08 5.305 33.515 5.445 ;
      RECT 33.375 3.995 33.515 5.445 ;
      RECT 31.08 4.925 31.22 5.445 ;
      RECT 30.78 4.925 31.22 5.155 ;
      RECT 28.44 4.925 31.22 5.065 ;
      RECT 30.78 4.835 31.04 5.155 ;
      RECT 28.44 4.645 28.58 5.065 ;
      RECT 27.93 4.555 28.19 4.875 ;
      RECT 27.93 4.645 28.58 4.785 ;
      RECT 27.99 3.155 28.13 4.875 ;
      RECT 33.315 3.995 33.575 4.315 ;
      RECT 27.93 3.155 28.19 3.475 ;
      RECT 32.94 4.835 33.2 5.155 ;
      RECT 33 3.245 33.14 5.155 ;
      RECT 32.66 3.245 33.14 3.52 ;
      RECT 32.46 3.15 32.94 3.495 ;
      RECT 32.45 4.785 32.73 5.155 ;
      RECT 32.52 3.69 32.66 5.155 ;
      RECT 32.46 3.69 32.72 4.315 ;
      RECT 32.45 3.69 32.73 4.06 ;
      RECT 31.38 4.835 31.64 5.155 ;
      RECT 31.38 4.645 31.58 5.155 ;
      RECT 31.185 4.645 31.58 4.785 ;
      RECT 31.185 3.155 31.325 4.785 ;
      RECT 31.185 3.155 31.5 3.525 ;
      RECT 31.125 3.155 31.5 3.475 ;
      RECT 28.85 4.25 29.13 4.62 ;
      RECT 30.3 4.275 30.56 4.595 ;
      RECT 28.68 4.365 30.56 4.505 ;
      RECT 28.68 4.25 29.13 4.505 ;
      RECT 28.62 3.69 28.88 4.315 ;
      RECT 28.61 3.69 28.89 4.06 ;
      RECT 29.69 3.69 30.1 4.06 ;
      RECT 29.1 3.715 29.36 4.035 ;
      RECT 29.1 3.805 30.1 3.945 ;
      RECT 28.61 3.13 28.89 3.5 ;
      RECT 28.61 3.155 29 3.475 ;
      RECT 23.155 8.51 23.475 8.835 ;
      RECT 23.185 7.985 23.355 8.835 ;
      RECT 23.185 7.985 23.36 8.335 ;
      RECT 23.185 7.985 24.16 8.16 ;
      RECT 23.985 3.26 24.16 8.16 ;
      RECT 23.93 3.26 24.28 3.61 ;
      RECT 23.955 8.945 24.28 9.27 ;
      RECT 22.84 9.035 24.28 9.205 ;
      RECT 22.84 3.69 23 9.205 ;
      RECT 23.155 3.66 23.475 3.98 ;
      RECT 22.84 3.69 23.475 3.86 ;
      RECT 20.29 4.835 20.55 5.155 ;
      RECT 20.35 3.13 20.49 5.155 ;
      RECT 21.55 3.995 21.89 4.345 ;
      RECT 20.925 4.065 21.89 4.265 ;
      RECT 20.925 3.235 21.125 4.265 ;
      RECT 20.175 3.69 20.49 4.06 ;
      RECT 21.64 3.99 21.81 4.345 ;
      RECT 20.245 3.245 20.49 4.06 ;
      RECT 20.28 3.13 20.56 3.5 ;
      RECT 20.28 3.235 21.125 3.435 ;
      RECT 19.6 3.715 19.86 4.035 ;
      RECT 18.94 3.805 19.86 3.945 ;
      RECT 18.94 2.865 19.08 3.945 ;
      RECT 15.4 3.155 15.66 3.475 ;
      RECT 15.58 2.865 15.72 3.385 ;
      RECT 15.58 2.865 19.08 3.005 ;
      RECT 10.37 9.285 10.66 9.635 ;
      RECT 10.37 9.355 11.59 9.525 ;
      RECT 11.42 8.975 11.59 9.525 ;
      RECT 18.515 8.895 18.865 9.245 ;
      RECT 11.42 8.975 18.865 9.145 ;
      RECT 18.43 4.555 18.69 4.875 ;
      RECT 18.49 3.145 18.63 4.875 ;
      RECT 18.42 3.145 18.7 3.515 ;
      RECT 15.82 5.305 18.255 5.445 ;
      RECT 18.115 3.995 18.255 5.445 ;
      RECT 15.82 4.925 15.96 5.445 ;
      RECT 15.52 4.925 15.96 5.155 ;
      RECT 13.18 4.925 15.96 5.065 ;
      RECT 15.52 4.835 15.78 5.155 ;
      RECT 13.18 4.645 13.32 5.065 ;
      RECT 12.67 4.555 12.93 4.875 ;
      RECT 12.67 4.645 13.32 4.785 ;
      RECT 12.73 3.155 12.87 4.875 ;
      RECT 18.055 3.995 18.315 4.315 ;
      RECT 12.67 3.155 12.93 3.475 ;
      RECT 17.68 4.835 17.94 5.155 ;
      RECT 17.74 3.245 17.88 5.155 ;
      RECT 17.4 3.245 17.88 3.52 ;
      RECT 17.2 3.15 17.68 3.495 ;
      RECT 17.19 4.785 17.47 5.155 ;
      RECT 17.26 3.69 17.4 5.155 ;
      RECT 17.2 3.69 17.46 4.315 ;
      RECT 17.19 3.69 17.47 4.06 ;
      RECT 16.12 4.835 16.38 5.155 ;
      RECT 16.12 4.645 16.32 5.155 ;
      RECT 15.925 4.645 16.32 4.785 ;
      RECT 15.925 3.155 16.065 4.785 ;
      RECT 15.925 3.155 16.24 3.525 ;
      RECT 15.865 3.155 16.24 3.475 ;
      RECT 13.59 4.25 13.87 4.62 ;
      RECT 15.04 4.275 15.3 4.595 ;
      RECT 13.42 4.365 15.3 4.505 ;
      RECT 13.42 4.25 13.87 4.505 ;
      RECT 13.36 3.69 13.62 4.315 ;
      RECT 13.35 3.69 13.63 4.06 ;
      RECT 14.43 3.69 14.84 4.06 ;
      RECT 13.84 3.715 14.1 4.035 ;
      RECT 13.84 3.805 14.84 3.945 ;
      RECT 13.35 3.13 13.63 3.5 ;
      RECT 13.35 3.155 13.74 3.475 ;
      RECT 78.885 9.345 79.255 9.715 ;
      RECT 77.75 3.69 78.03 4.155 ;
      RECT 77.51 3.155 77.79 3.5 ;
      RECT 76.31 3.69 76.59 4.06 ;
      RECT 63.625 9.345 63.995 9.715 ;
      RECT 62.49 3.69 62.77 4.155 ;
      RECT 62.25 3.155 62.53 3.5 ;
      RECT 61.05 3.69 61.33 4.06 ;
      RECT 48.365 9.345 48.735 9.715 ;
      RECT 47.23 3.69 47.51 4.155 ;
      RECT 46.99 3.155 47.27 3.5 ;
      RECT 45.79 3.69 46.07 4.06 ;
      RECT 33.105 9.345 33.475 9.715 ;
      RECT 31.97 3.69 32.25 4.155 ;
      RECT 31.73 3.155 32.01 3.5 ;
      RECT 30.53 3.69 30.81 4.06 ;
      RECT 17.845 9.345 18.215 9.715 ;
      RECT 16.71 3.69 16.99 4.155 ;
      RECT 16.47 3.155 16.75 3.5 ;
      RECT 15.27 3.69 15.55 4.06 ;
    LAYER via1 ;
      RECT 87.455 9.665 87.605 9.815 ;
      RECT 85.085 9.03 85.235 9.18 ;
      RECT 85.07 3.36 85.22 3.51 ;
      RECT 84.28 3.745 84.43 3.895 ;
      RECT 84.28 8.615 84.43 8.765 ;
      RECT 82.69 4.095 82.84 4.245 ;
      RECT 81.385 3.24 81.535 3.39 ;
      RECT 81.385 4.92 81.535 5.07 ;
      RECT 80.695 3.8 80.845 3.95 ;
      RECT 79.655 9 79.805 9.15 ;
      RECT 79.525 3.24 79.675 3.39 ;
      RECT 79.525 4.64 79.675 4.79 ;
      RECT 79.15 4.08 79.3 4.23 ;
      RECT 78.995 9.455 79.145 9.605 ;
      RECT 78.775 4.92 78.925 5.07 ;
      RECT 78.295 3.24 78.445 3.39 ;
      RECT 78.295 4.08 78.445 4.23 ;
      RECT 77.815 3.8 77.965 3.95 ;
      RECT 77.575 3.24 77.725 3.39 ;
      RECT 77.215 4.92 77.365 5.07 ;
      RECT 76.96 3.24 77.11 3.39 ;
      RECT 76.615 4.92 76.765 5.07 ;
      RECT 76.495 3.24 76.645 3.39 ;
      RECT 76.375 3.8 76.525 3.95 ;
      RECT 76.135 4.36 76.285 4.51 ;
      RECT 74.935 3.8 75.085 3.95 ;
      RECT 74.575 3.24 74.725 3.39 ;
      RECT 74.455 4.08 74.605 4.23 ;
      RECT 73.765 3.24 73.915 3.39 ;
      RECT 73.765 4.64 73.915 4.79 ;
      RECT 72.17 9.045 72.32 9.195 ;
      RECT 69.825 9.03 69.975 9.18 ;
      RECT 69.81 3.36 69.96 3.51 ;
      RECT 69.02 3.745 69.17 3.895 ;
      RECT 69.02 8.615 69.17 8.765 ;
      RECT 67.43 4.095 67.58 4.245 ;
      RECT 66.125 3.24 66.275 3.39 ;
      RECT 66.125 4.92 66.275 5.07 ;
      RECT 65.435 3.8 65.585 3.95 ;
      RECT 64.4 9 64.55 9.15 ;
      RECT 64.265 3.24 64.415 3.39 ;
      RECT 64.265 4.64 64.415 4.79 ;
      RECT 63.89 4.08 64.04 4.23 ;
      RECT 63.735 9.455 63.885 9.605 ;
      RECT 63.515 4.92 63.665 5.07 ;
      RECT 63.035 3.24 63.185 3.39 ;
      RECT 63.035 4.08 63.185 4.23 ;
      RECT 62.555 3.8 62.705 3.95 ;
      RECT 62.315 3.24 62.465 3.39 ;
      RECT 61.955 4.92 62.105 5.07 ;
      RECT 61.7 3.24 61.85 3.39 ;
      RECT 61.355 4.92 61.505 5.07 ;
      RECT 61.235 3.24 61.385 3.39 ;
      RECT 61.115 3.8 61.265 3.95 ;
      RECT 60.875 4.36 61.025 4.51 ;
      RECT 59.675 3.8 59.825 3.95 ;
      RECT 59.315 3.24 59.465 3.39 ;
      RECT 59.195 4.08 59.345 4.23 ;
      RECT 58.505 3.24 58.655 3.39 ;
      RECT 58.505 4.64 58.655 4.79 ;
      RECT 56.91 9.045 57.06 9.195 ;
      RECT 54.565 9.03 54.715 9.18 ;
      RECT 54.55 3.36 54.7 3.51 ;
      RECT 53.76 3.745 53.91 3.895 ;
      RECT 53.76 8.615 53.91 8.765 ;
      RECT 52.17 4.095 52.32 4.245 ;
      RECT 50.865 3.24 51.015 3.39 ;
      RECT 50.865 4.92 51.015 5.07 ;
      RECT 50.175 3.8 50.325 3.95 ;
      RECT 49.135 9.005 49.285 9.155 ;
      RECT 49.005 3.24 49.155 3.39 ;
      RECT 49.005 4.64 49.155 4.79 ;
      RECT 48.63 4.08 48.78 4.23 ;
      RECT 48.475 9.455 48.625 9.605 ;
      RECT 48.255 4.92 48.405 5.07 ;
      RECT 47.775 3.24 47.925 3.39 ;
      RECT 47.775 4.08 47.925 4.23 ;
      RECT 47.295 3.8 47.445 3.95 ;
      RECT 47.055 3.24 47.205 3.39 ;
      RECT 46.695 4.92 46.845 5.07 ;
      RECT 46.44 3.24 46.59 3.39 ;
      RECT 46.095 4.92 46.245 5.07 ;
      RECT 45.975 3.24 46.125 3.39 ;
      RECT 45.855 3.8 46.005 3.95 ;
      RECT 45.615 4.36 45.765 4.51 ;
      RECT 44.415 3.8 44.565 3.95 ;
      RECT 44.055 3.24 44.205 3.39 ;
      RECT 43.935 4.08 44.085 4.23 ;
      RECT 43.245 3.24 43.395 3.39 ;
      RECT 43.245 4.64 43.395 4.79 ;
      RECT 41.695 9.05 41.845 9.2 ;
      RECT 39.305 9.03 39.455 9.18 ;
      RECT 39.29 3.36 39.44 3.51 ;
      RECT 38.5 3.745 38.65 3.895 ;
      RECT 38.5 8.615 38.65 8.765 ;
      RECT 36.91 4.095 37.06 4.245 ;
      RECT 35.605 3.24 35.755 3.39 ;
      RECT 35.605 4.92 35.755 5.07 ;
      RECT 34.915 3.8 35.065 3.95 ;
      RECT 33.875 9 34.025 9.15 ;
      RECT 33.745 3.24 33.895 3.39 ;
      RECT 33.745 4.64 33.895 4.79 ;
      RECT 33.37 4.08 33.52 4.23 ;
      RECT 33.215 9.455 33.365 9.605 ;
      RECT 32.995 4.92 33.145 5.07 ;
      RECT 32.515 3.24 32.665 3.39 ;
      RECT 32.515 4.08 32.665 4.23 ;
      RECT 32.035 3.8 32.185 3.95 ;
      RECT 31.795 3.24 31.945 3.39 ;
      RECT 31.435 4.92 31.585 5.07 ;
      RECT 31.18 3.24 31.33 3.39 ;
      RECT 30.835 4.92 30.985 5.07 ;
      RECT 30.715 3.24 30.865 3.39 ;
      RECT 30.595 3.8 30.745 3.95 ;
      RECT 30.355 4.36 30.505 4.51 ;
      RECT 29.155 3.8 29.305 3.95 ;
      RECT 28.795 3.24 28.945 3.39 ;
      RECT 28.675 4.08 28.825 4.23 ;
      RECT 27.985 3.24 28.135 3.39 ;
      RECT 27.985 4.64 28.135 4.79 ;
      RECT 26.435 9.045 26.585 9.195 ;
      RECT 24.045 9.03 24.195 9.18 ;
      RECT 24.03 3.36 24.18 3.51 ;
      RECT 23.24 3.745 23.39 3.895 ;
      RECT 23.24 8.615 23.39 8.765 ;
      RECT 21.65 4.095 21.8 4.245 ;
      RECT 20.345 3.24 20.495 3.39 ;
      RECT 20.345 4.92 20.495 5.07 ;
      RECT 19.655 3.8 19.805 3.95 ;
      RECT 18.615 8.995 18.765 9.145 ;
      RECT 18.485 3.24 18.635 3.39 ;
      RECT 18.485 4.64 18.635 4.79 ;
      RECT 18.11 4.08 18.26 4.23 ;
      RECT 17.955 9.455 18.105 9.605 ;
      RECT 17.735 4.92 17.885 5.07 ;
      RECT 17.255 3.24 17.405 3.39 ;
      RECT 17.255 4.08 17.405 4.23 ;
      RECT 16.775 3.8 16.925 3.95 ;
      RECT 16.535 3.24 16.685 3.39 ;
      RECT 16.175 4.92 16.325 5.07 ;
      RECT 15.92 3.24 16.07 3.39 ;
      RECT 15.575 4.92 15.725 5.07 ;
      RECT 15.455 3.24 15.605 3.39 ;
      RECT 15.335 3.8 15.485 3.95 ;
      RECT 15.095 4.36 15.245 4.51 ;
      RECT 13.895 3.8 14.045 3.95 ;
      RECT 13.535 3.24 13.685 3.39 ;
      RECT 13.415 4.08 13.565 4.23 ;
      RECT 12.725 3.24 12.875 3.39 ;
      RECT 12.725 4.64 12.875 4.79 ;
      RECT 10.44 9.385 10.59 9.535 ;
      RECT 10.065 8.645 10.215 8.795 ;
    LAYER met1 ;
      RECT 73.905 4.04 74.195 4.27 ;
      RECT 58.645 4.04 58.935 4.27 ;
      RECT 43.385 4.04 43.675 4.27 ;
      RECT 28.125 4.04 28.415 4.27 ;
      RECT 12.865 4.04 13.155 4.27 ;
      RECT 73.98 3.225 74.12 4.27 ;
      RECT 58.72 3.665 58.86 4.27 ;
      RECT 43.46 3.665 43.6 4.27 ;
      RECT 28.2 3.665 28.34 4.27 ;
      RECT 12.94 3.665 13.08 4.27 ;
      RECT 73.98 3.665 74.6 3.805 ;
      RECT 74.46 0 74.6 3.805 ;
      RECT 58.72 3.665 59.34 3.805 ;
      RECT 59.2 0 59.34 3.805 ;
      RECT 43.46 3.665 44.08 3.805 ;
      RECT 43.94 0 44.08 3.805 ;
      RECT 28.2 3.665 28.82 3.805 ;
      RECT 28.68 0 28.82 3.805 ;
      RECT 12.94 3.665 13.56 3.805 ;
      RECT 13.42 0 13.56 3.805 ;
      RECT 73.68 3.185 74 3.685 ;
      RECT 73.595 3.225 74.165 3.685 ;
      RECT 74.22 3.245 74.6 3.505 ;
      RECT 58.96 3.245 59.34 3.505 ;
      RECT 43.7 3.245 44.08 3.505 ;
      RECT 28.44 3.245 28.82 3.505 ;
      RECT 13.18 3.245 13.56 3.505 ;
      RECT 74.4 3.185 74.81 3.445 ;
      RECT 59.14 3.185 59.55 3.445 ;
      RECT 43.88 3.185 44.29 3.445 ;
      RECT 28.62 3.185 29.03 3.445 ;
      RECT 13.36 3.185 13.77 3.445 ;
      RECT 75.105 3.2 75.395 3.43 ;
      RECT 59.845 3.2 60.135 3.43 ;
      RECT 44.585 3.2 44.875 3.43 ;
      RECT 29.325 3.2 29.615 3.43 ;
      RECT 14.065 3.2 14.355 3.43 ;
      RECT 74.22 3.245 75.395 3.385 ;
      RECT 58.96 3.245 60.135 3.385 ;
      RECT 43.7 3.245 44.875 3.385 ;
      RECT 28.44 3.245 29.615 3.385 ;
      RECT 13.18 3.245 14.355 3.385 ;
      RECT 74.4 0 74.69 3.445 ;
      RECT 59.14 0 59.43 3.445 ;
      RECT 43.88 0 44.17 3.445 ;
      RECT 28.62 0 28.91 3.445 ;
      RECT 13.36 0 13.65 3.445 ;
      RECT 73.415 0 82.155 3.035 ;
      RECT 58.155 0 66.895 3.035 ;
      RECT 42.895 0 51.635 3.035 ;
      RECT 27.635 0 36.375 3.035 ;
      RECT 12.375 0 21.115 3.035 ;
      RECT 8.875 0 87.925 1.6 ;
      RECT 8.83 10.865 87.925 12.465 ;
      RECT 78.385 8.605 78.555 12.465 ;
      RECT 63.125 8.605 63.295 12.465 ;
      RECT 47.865 8.605 48.035 12.465 ;
      RECT 32.605 8.605 32.775 12.465 ;
      RECT 17.345 8.605 17.515 12.465 ;
      RECT 78.55 8.575 78.84 8.805 ;
      RECT 63.29 8.575 63.58 8.805 ;
      RECT 48.03 8.575 48.32 8.805 ;
      RECT 32.77 8.575 33.06 8.805 ;
      RECT 17.51 8.575 17.8 8.805 ;
      RECT 78.38 8.605 78.84 8.775 ;
      RECT 63.12 8.605 63.58 8.775 ;
      RECT 47.86 8.605 48.32 8.775 ;
      RECT 32.6 8.605 33.06 8.775 ;
      RECT 17.34 8.605 17.8 8.775 ;
      RECT 87.32 10.06 87.61 10.29 ;
      RECT 87.38 8.58 87.55 10.29 ;
      RECT 87.355 9.565 87.705 9.915 ;
      RECT 87.32 8.58 87.61 8.81 ;
      RECT 86.915 3.69 87.02 4.26 ;
      RECT 86.915 4.025 87.24 4.255 ;
      RECT 86.915 4.055 87.41 4.225 ;
      RECT 86.915 3.69 87.105 4.255 ;
      RECT 86.33 3.655 86.62 3.885 ;
      RECT 86.33 3.69 87.105 3.86 ;
      RECT 86.39 2.175 86.56 3.885 ;
      RECT 86.33 2.175 86.62 2.405 ;
      RECT 86.33 10.06 86.62 10.29 ;
      RECT 86.39 8.58 86.56 10.29 ;
      RECT 86.33 8.58 86.62 8.81 ;
      RECT 86.33 8.615 87.18 8.775 ;
      RECT 87.015 8.21 87.18 8.775 ;
      RECT 86.33 8.61 86.725 8.775 ;
      RECT 86.95 8.21 87.24 8.44 ;
      RECT 86.95 8.24 87.41 8.41 ;
      RECT 85.96 4.025 86.25 4.255 ;
      RECT 85.96 4.055 86.42 4.225 ;
      RECT 86.025 2.95 86.19 4.255 ;
      RECT 84.54 2.92 84.83 3.15 ;
      RECT 84.54 2.95 86.19 3.12 ;
      RECT 84.6 2.18 84.77 3.15 ;
      RECT 84.54 2.18 84.83 2.41 ;
      RECT 84.54 10.055 84.83 10.285 ;
      RECT 84.6 9.315 84.77 10.285 ;
      RECT 84.6 9.41 86.19 9.58 ;
      RECT 86.02 8.21 86.19 9.58 ;
      RECT 84.54 9.315 84.83 9.545 ;
      RECT 85.96 8.21 86.25 8.44 ;
      RECT 85.96 8.24 86.42 8.41 ;
      RECT 82.59 3.995 82.93 4.345 ;
      RECT 82.68 3.32 82.85 4.345 ;
      RECT 84.97 3.26 85.32 3.61 ;
      RECT 82.68 3.32 85.32 3.49 ;
      RECT 84.995 8.945 85.32 9.27 ;
      RECT 79.555 8.9 79.905 9.25 ;
      RECT 84.97 8.945 85.32 9.175 ;
      RECT 79.355 8.945 79.905 9.175 ;
      RECT 79.185 8.975 85.32 9.145 ;
      RECT 84.195 3.66 84.515 3.98 ;
      RECT 84.165 3.66 84.515 3.89 ;
      RECT 83.995 3.69 84.515 3.86 ;
      RECT 84.195 8.545 84.515 8.835 ;
      RECT 84.165 8.575 84.515 8.805 ;
      RECT 83.995 8.605 84.515 8.775 ;
      RECT 81.3 3.185 81.62 3.445 ;
      RECT 80.865 3.2 81.155 3.43 ;
      RECT 80.865 3.245 81.62 3.385 ;
      RECT 81.3 4.865 81.62 5.125 ;
      RECT 80.865 4.88 81.155 5.11 ;
      RECT 80.865 4.925 81.62 5.065 ;
      RECT 80.625 4.32 80.915 4.55 ;
      RECT 80.625 4.365 81.2 4.505 ;
      RECT 81.06 4.225 81.32 4.365 ;
      RECT 81.105 4.04 81.395 4.27 ;
      RECT 79.26 4.225 80.36 4.365 ;
      RECT 79.065 4.025 79.385 4.285 ;
      RECT 80.145 4.04 80.435 4.27 ;
      RECT 79.065 4.04 79.475 4.285 ;
      RECT 79.44 3.185 79.76 3.445 ;
      RECT 79.905 3.2 80.195 3.43 ;
      RECT 79.44 3.245 80.195 3.385 ;
      RECT 76.74 4.45 78.92 4.59 ;
      RECT 78.78 3.46 78.92 4.59 ;
      RECT 76.74 4.365 78.035 4.59 ;
      RECT 77.745 4.32 78.035 4.59 ;
      RECT 76.74 4.085 77.075 4.59 ;
      RECT 76.785 4.04 77.075 4.59 ;
      RECT 79.665 3.76 79.955 3.99 ;
      RECT 78.78 3.665 79.88 3.805 ;
      RECT 78.705 3.46 78.995 3.71 ;
      RECT 78.925 10.055 79.215 10.285 ;
      RECT 78.985 9.315 79.155 10.285 ;
      RECT 78.885 9.345 79.255 9.715 ;
      RECT 78.925 9.315 79.215 9.715 ;
      RECT 78.69 4.865 79.01 5.125 ;
      RECT 78.69 4.88 79.205 5.11 ;
      RECT 77.265 3.76 77.555 3.99 ;
      RECT 77.415 3.365 77.555 3.99 ;
      RECT 77.415 3.365 77.72 3.505 ;
      RECT 78.21 3.185 78.53 3.445 ;
      RECT 77.49 3.185 77.81 3.445 ;
      RECT 77.985 3.2 78.53 3.43 ;
      RECT 77.49 3.245 78.53 3.385 ;
      RECT 77.13 4.865 77.45 5.125 ;
      RECT 77.025 4.88 77.45 5.11 ;
      RECT 75.105 4.32 75.395 4.55 ;
      RECT 75.105 4.32 75.56 4.505 ;
      RECT 75.42 3.845 75.56 4.505 ;
      RECT 75.54 3.245 75.68 3.985 ;
      RECT 76.41 3.185 76.73 3.445 ;
      RECT 75.585 3.2 75.875 3.43 ;
      RECT 75.54 3.245 76.73 3.385 ;
      RECT 76.29 3.745 76.61 4.005 ;
      RECT 75.825 3.76 76.115 3.99 ;
      RECT 75.825 3.805 76.61 3.945 ;
      RECT 76.05 4.305 76.37 4.565 ;
      RECT 76.05 4.32 76.595 4.55 ;
      RECT 75.585 4.88 75.875 5.11 ;
      RECT 74.7 4.76 75.8 4.9 ;
      RECT 74.625 4.6 74.915 4.83 ;
      RECT 72.06 10.06 72.35 10.29 ;
      RECT 72.12 8.58 72.29 10.29 ;
      RECT 72.07 8.945 72.42 9.295 ;
      RECT 72.06 8.58 72.35 8.81 ;
      RECT 71.655 3.69 71.76 4.26 ;
      RECT 71.655 4.025 71.98 4.255 ;
      RECT 71.655 4.055 72.15 4.225 ;
      RECT 71.655 3.69 71.845 4.255 ;
      RECT 71.07 3.655 71.36 3.885 ;
      RECT 71.07 3.69 71.845 3.86 ;
      RECT 71.13 2.175 71.3 3.885 ;
      RECT 71.07 2.175 71.36 2.405 ;
      RECT 71.07 10.06 71.36 10.29 ;
      RECT 71.13 8.58 71.3 10.29 ;
      RECT 71.07 8.58 71.36 8.81 ;
      RECT 71.07 8.615 71.92 8.775 ;
      RECT 71.755 8.21 71.92 8.775 ;
      RECT 71.07 8.61 71.465 8.775 ;
      RECT 71.69 8.21 71.98 8.44 ;
      RECT 71.69 8.24 72.15 8.41 ;
      RECT 70.7 4.025 70.99 4.255 ;
      RECT 70.7 4.055 71.16 4.225 ;
      RECT 70.765 2.95 70.93 4.255 ;
      RECT 69.28 2.92 69.57 3.15 ;
      RECT 69.28 2.95 70.93 3.12 ;
      RECT 69.34 2.18 69.51 3.15 ;
      RECT 69.28 2.18 69.57 2.41 ;
      RECT 69.28 10.055 69.57 10.285 ;
      RECT 69.34 9.315 69.51 10.285 ;
      RECT 69.34 9.41 70.93 9.58 ;
      RECT 70.76 8.21 70.93 9.58 ;
      RECT 69.28 9.315 69.57 9.545 ;
      RECT 70.7 8.21 70.99 8.44 ;
      RECT 70.7 8.24 71.16 8.41 ;
      RECT 67.33 3.995 67.67 4.345 ;
      RECT 67.42 3.32 67.59 4.345 ;
      RECT 69.71 3.26 70.06 3.61 ;
      RECT 67.42 3.32 70.06 3.49 ;
      RECT 69.735 8.945 70.06 9.27 ;
      RECT 64.3 8.9 64.65 9.25 ;
      RECT 69.71 8.945 70.06 9.175 ;
      RECT 64.095 8.945 64.65 9.175 ;
      RECT 63.925 8.975 70.06 9.145 ;
      RECT 68.935 3.66 69.255 3.98 ;
      RECT 68.905 3.66 69.255 3.89 ;
      RECT 68.735 3.69 69.255 3.86 ;
      RECT 68.935 8.545 69.255 8.835 ;
      RECT 68.905 8.575 69.255 8.805 ;
      RECT 68.735 8.605 69.255 8.775 ;
      RECT 66.04 3.185 66.36 3.445 ;
      RECT 65.605 3.2 65.895 3.43 ;
      RECT 65.605 3.245 66.36 3.385 ;
      RECT 66.04 4.865 66.36 5.125 ;
      RECT 65.605 4.88 65.895 5.11 ;
      RECT 65.605 4.925 66.36 5.065 ;
      RECT 65.365 4.32 65.655 4.55 ;
      RECT 65.365 4.365 65.94 4.505 ;
      RECT 65.8 4.225 66.06 4.365 ;
      RECT 65.845 4.04 66.135 4.27 ;
      RECT 64 4.225 65.1 4.365 ;
      RECT 63.805 4.025 64.125 4.285 ;
      RECT 64.885 4.04 65.175 4.27 ;
      RECT 63.805 4.04 64.215 4.285 ;
      RECT 64.18 3.185 64.5 3.445 ;
      RECT 64.645 3.2 64.935 3.43 ;
      RECT 64.18 3.245 64.935 3.385 ;
      RECT 61.48 4.45 63.66 4.59 ;
      RECT 63.52 3.46 63.66 4.59 ;
      RECT 61.48 4.365 62.775 4.59 ;
      RECT 62.485 4.32 62.775 4.59 ;
      RECT 61.48 4.085 61.815 4.59 ;
      RECT 61.525 4.04 61.815 4.59 ;
      RECT 64.405 3.76 64.695 3.99 ;
      RECT 63.52 3.665 64.62 3.805 ;
      RECT 63.445 3.46 63.735 3.71 ;
      RECT 63.665 10.055 63.955 10.285 ;
      RECT 63.725 9.315 63.895 10.285 ;
      RECT 63.625 9.345 63.995 9.715 ;
      RECT 63.665 9.315 63.955 9.715 ;
      RECT 63.43 4.865 63.75 5.125 ;
      RECT 63.43 4.88 63.945 5.11 ;
      RECT 62.005 3.76 62.295 3.99 ;
      RECT 62.155 3.365 62.295 3.99 ;
      RECT 62.155 3.365 62.46 3.505 ;
      RECT 62.95 3.185 63.27 3.445 ;
      RECT 62.23 3.185 62.55 3.445 ;
      RECT 62.725 3.2 63.27 3.43 ;
      RECT 62.23 3.245 63.27 3.385 ;
      RECT 61.87 4.865 62.19 5.125 ;
      RECT 61.765 4.88 62.19 5.11 ;
      RECT 59.845 4.32 60.135 4.55 ;
      RECT 59.845 4.32 60.3 4.505 ;
      RECT 60.16 3.845 60.3 4.505 ;
      RECT 60.28 3.245 60.42 3.985 ;
      RECT 61.15 3.185 61.47 3.445 ;
      RECT 60.325 3.2 60.615 3.43 ;
      RECT 60.28 3.245 61.47 3.385 ;
      RECT 61.03 3.745 61.35 4.005 ;
      RECT 60.565 3.76 60.855 3.99 ;
      RECT 60.565 3.805 61.35 3.945 ;
      RECT 60.79 4.305 61.11 4.565 ;
      RECT 60.79 4.32 61.335 4.55 ;
      RECT 60.325 4.88 60.615 5.11 ;
      RECT 59.44 4.76 60.54 4.9 ;
      RECT 59.365 4.6 59.655 4.83 ;
      RECT 56.8 10.06 57.09 10.29 ;
      RECT 56.86 8.58 57.03 10.29 ;
      RECT 56.81 8.945 57.16 9.295 ;
      RECT 56.8 8.58 57.09 8.81 ;
      RECT 56.395 3.69 56.5 4.26 ;
      RECT 56.395 4.025 56.72 4.255 ;
      RECT 56.395 4.055 56.89 4.225 ;
      RECT 56.395 3.69 56.585 4.255 ;
      RECT 55.81 3.655 56.1 3.885 ;
      RECT 55.81 3.69 56.585 3.86 ;
      RECT 55.87 2.175 56.04 3.885 ;
      RECT 55.81 2.175 56.1 2.405 ;
      RECT 55.81 10.06 56.1 10.29 ;
      RECT 55.87 8.58 56.04 10.29 ;
      RECT 55.81 8.58 56.1 8.81 ;
      RECT 55.81 8.615 56.66 8.775 ;
      RECT 56.495 8.21 56.66 8.775 ;
      RECT 55.81 8.61 56.205 8.775 ;
      RECT 56.43 8.21 56.72 8.44 ;
      RECT 56.43 8.24 56.89 8.41 ;
      RECT 55.44 4.025 55.73 4.255 ;
      RECT 55.44 4.055 55.9 4.225 ;
      RECT 55.505 2.95 55.67 4.255 ;
      RECT 54.02 2.92 54.31 3.15 ;
      RECT 54.02 2.95 55.67 3.12 ;
      RECT 54.08 2.18 54.25 3.15 ;
      RECT 54.02 2.18 54.31 2.41 ;
      RECT 54.02 10.055 54.31 10.285 ;
      RECT 54.08 9.315 54.25 10.285 ;
      RECT 54.08 9.41 55.67 9.58 ;
      RECT 55.5 8.21 55.67 9.58 ;
      RECT 54.02 9.315 54.31 9.545 ;
      RECT 55.44 8.21 55.73 8.44 ;
      RECT 55.44 8.24 55.9 8.41 ;
      RECT 52.07 3.995 52.41 4.345 ;
      RECT 52.16 3.32 52.33 4.345 ;
      RECT 54.45 3.26 54.8 3.61 ;
      RECT 52.16 3.32 54.8 3.49 ;
      RECT 54.475 8.945 54.8 9.27 ;
      RECT 49.035 8.905 49.385 9.255 ;
      RECT 54.45 8.945 54.8 9.175 ;
      RECT 48.835 8.945 49.385 9.175 ;
      RECT 48.665 8.975 54.8 9.145 ;
      RECT 53.675 3.66 53.995 3.98 ;
      RECT 53.645 3.66 53.995 3.89 ;
      RECT 53.475 3.69 53.995 3.86 ;
      RECT 53.675 8.545 53.995 8.835 ;
      RECT 53.645 8.575 53.995 8.805 ;
      RECT 53.475 8.605 53.995 8.775 ;
      RECT 50.78 3.185 51.1 3.445 ;
      RECT 50.345 3.2 50.635 3.43 ;
      RECT 50.345 3.245 51.1 3.385 ;
      RECT 50.78 4.865 51.1 5.125 ;
      RECT 50.345 4.88 50.635 5.11 ;
      RECT 50.345 4.925 51.1 5.065 ;
      RECT 50.105 4.32 50.395 4.55 ;
      RECT 50.105 4.365 50.68 4.505 ;
      RECT 50.54 4.225 50.8 4.365 ;
      RECT 50.585 4.04 50.875 4.27 ;
      RECT 48.74 4.225 49.84 4.365 ;
      RECT 48.545 4.025 48.865 4.285 ;
      RECT 49.625 4.04 49.915 4.27 ;
      RECT 48.545 4.04 48.955 4.285 ;
      RECT 48.92 3.185 49.24 3.445 ;
      RECT 49.385 3.2 49.675 3.43 ;
      RECT 48.92 3.245 49.675 3.385 ;
      RECT 46.22 4.45 48.4 4.59 ;
      RECT 48.26 3.46 48.4 4.59 ;
      RECT 46.22 4.365 47.515 4.59 ;
      RECT 47.225 4.32 47.515 4.59 ;
      RECT 46.22 4.085 46.555 4.59 ;
      RECT 46.265 4.04 46.555 4.59 ;
      RECT 49.145 3.76 49.435 3.99 ;
      RECT 48.26 3.665 49.36 3.805 ;
      RECT 48.185 3.46 48.475 3.71 ;
      RECT 48.405 10.055 48.695 10.285 ;
      RECT 48.465 9.315 48.635 10.285 ;
      RECT 48.365 9.345 48.735 9.715 ;
      RECT 48.405 9.315 48.695 9.715 ;
      RECT 48.17 4.865 48.49 5.125 ;
      RECT 48.17 4.88 48.685 5.11 ;
      RECT 46.745 3.76 47.035 3.99 ;
      RECT 46.895 3.365 47.035 3.99 ;
      RECT 46.895 3.365 47.2 3.505 ;
      RECT 47.69 3.185 48.01 3.445 ;
      RECT 46.97 3.185 47.29 3.445 ;
      RECT 47.465 3.2 48.01 3.43 ;
      RECT 46.97 3.245 48.01 3.385 ;
      RECT 46.61 4.865 46.93 5.125 ;
      RECT 46.505 4.88 46.93 5.11 ;
      RECT 44.585 4.32 44.875 4.55 ;
      RECT 44.585 4.32 45.04 4.505 ;
      RECT 44.9 3.845 45.04 4.505 ;
      RECT 45.02 3.245 45.16 3.985 ;
      RECT 45.89 3.185 46.21 3.445 ;
      RECT 45.065 3.2 45.355 3.43 ;
      RECT 45.02 3.245 46.21 3.385 ;
      RECT 45.77 3.745 46.09 4.005 ;
      RECT 45.305 3.76 45.595 3.99 ;
      RECT 45.305 3.805 46.09 3.945 ;
      RECT 45.53 4.305 45.85 4.565 ;
      RECT 45.53 4.32 46.075 4.55 ;
      RECT 45.065 4.88 45.355 5.11 ;
      RECT 44.18 4.76 45.28 4.9 ;
      RECT 44.105 4.6 44.395 4.83 ;
      RECT 41.54 10.06 41.83 10.29 ;
      RECT 41.6 8.58 41.77 10.29 ;
      RECT 41.59 8.95 41.945 9.305 ;
      RECT 41.54 8.58 41.83 8.81 ;
      RECT 41.135 3.69 41.24 4.26 ;
      RECT 41.135 4.025 41.46 4.255 ;
      RECT 41.135 4.055 41.63 4.225 ;
      RECT 41.135 3.69 41.325 4.255 ;
      RECT 40.55 3.655 40.84 3.885 ;
      RECT 40.55 3.69 41.325 3.86 ;
      RECT 40.61 2.175 40.78 3.885 ;
      RECT 40.55 2.175 40.84 2.405 ;
      RECT 40.55 10.06 40.84 10.29 ;
      RECT 40.61 8.58 40.78 10.29 ;
      RECT 40.55 8.58 40.84 8.81 ;
      RECT 40.55 8.615 41.4 8.775 ;
      RECT 41.235 8.21 41.4 8.775 ;
      RECT 40.55 8.61 40.945 8.775 ;
      RECT 41.17 8.21 41.46 8.44 ;
      RECT 41.17 8.24 41.63 8.41 ;
      RECT 40.18 4.025 40.47 4.255 ;
      RECT 40.18 4.055 40.64 4.225 ;
      RECT 40.245 2.95 40.41 4.255 ;
      RECT 38.76 2.92 39.05 3.15 ;
      RECT 38.76 2.95 40.41 3.12 ;
      RECT 38.82 2.18 38.99 3.15 ;
      RECT 38.76 2.18 39.05 2.41 ;
      RECT 38.76 10.055 39.05 10.285 ;
      RECT 38.82 9.315 38.99 10.285 ;
      RECT 38.82 9.41 40.41 9.58 ;
      RECT 40.24 8.21 40.41 9.58 ;
      RECT 38.76 9.315 39.05 9.545 ;
      RECT 40.18 8.21 40.47 8.44 ;
      RECT 40.18 8.24 40.64 8.41 ;
      RECT 36.81 3.995 37.15 4.345 ;
      RECT 36.9 3.32 37.07 4.345 ;
      RECT 39.19 3.26 39.54 3.61 ;
      RECT 36.9 3.32 39.54 3.49 ;
      RECT 39.215 8.945 39.54 9.27 ;
      RECT 33.775 8.9 34.125 9.25 ;
      RECT 39.19 8.945 39.54 9.175 ;
      RECT 33.575 8.945 34.125 9.175 ;
      RECT 33.405 8.975 39.54 9.145 ;
      RECT 38.415 3.66 38.735 3.98 ;
      RECT 38.385 3.66 38.735 3.89 ;
      RECT 38.215 3.69 38.735 3.86 ;
      RECT 38.415 8.545 38.735 8.835 ;
      RECT 38.385 8.575 38.735 8.805 ;
      RECT 38.215 8.605 38.735 8.775 ;
      RECT 35.52 3.185 35.84 3.445 ;
      RECT 35.085 3.2 35.375 3.43 ;
      RECT 35.085 3.245 35.84 3.385 ;
      RECT 35.52 4.865 35.84 5.125 ;
      RECT 35.085 4.88 35.375 5.11 ;
      RECT 35.085 4.925 35.84 5.065 ;
      RECT 34.845 4.32 35.135 4.55 ;
      RECT 34.845 4.365 35.42 4.505 ;
      RECT 35.28 4.225 35.54 4.365 ;
      RECT 35.325 4.04 35.615 4.27 ;
      RECT 33.48 4.225 34.58 4.365 ;
      RECT 33.285 4.025 33.605 4.285 ;
      RECT 34.365 4.04 34.655 4.27 ;
      RECT 33.285 4.04 33.695 4.285 ;
      RECT 33.66 3.185 33.98 3.445 ;
      RECT 34.125 3.2 34.415 3.43 ;
      RECT 33.66 3.245 34.415 3.385 ;
      RECT 30.96 4.45 33.14 4.59 ;
      RECT 33 3.46 33.14 4.59 ;
      RECT 30.96 4.365 32.255 4.59 ;
      RECT 31.965 4.32 32.255 4.59 ;
      RECT 30.96 4.085 31.295 4.59 ;
      RECT 31.005 4.04 31.295 4.59 ;
      RECT 33.885 3.76 34.175 3.99 ;
      RECT 33 3.665 34.1 3.805 ;
      RECT 32.925 3.46 33.215 3.71 ;
      RECT 33.145 10.055 33.435 10.285 ;
      RECT 33.205 9.315 33.375 10.285 ;
      RECT 33.105 9.345 33.475 9.715 ;
      RECT 33.145 9.315 33.435 9.715 ;
      RECT 32.91 4.865 33.23 5.125 ;
      RECT 32.91 4.88 33.425 5.11 ;
      RECT 31.485 3.76 31.775 3.99 ;
      RECT 31.635 3.365 31.775 3.99 ;
      RECT 31.635 3.365 31.94 3.505 ;
      RECT 32.43 3.185 32.75 3.445 ;
      RECT 31.71 3.185 32.03 3.445 ;
      RECT 32.205 3.2 32.75 3.43 ;
      RECT 31.71 3.245 32.75 3.385 ;
      RECT 31.35 4.865 31.67 5.125 ;
      RECT 31.245 4.88 31.67 5.11 ;
      RECT 29.325 4.32 29.615 4.55 ;
      RECT 29.325 4.32 29.78 4.505 ;
      RECT 29.64 3.845 29.78 4.505 ;
      RECT 29.76 3.245 29.9 3.985 ;
      RECT 30.63 3.185 30.95 3.445 ;
      RECT 29.805 3.2 30.095 3.43 ;
      RECT 29.76 3.245 30.95 3.385 ;
      RECT 30.51 3.745 30.83 4.005 ;
      RECT 30.045 3.76 30.335 3.99 ;
      RECT 30.045 3.805 30.83 3.945 ;
      RECT 30.27 4.305 30.59 4.565 ;
      RECT 30.27 4.32 30.815 4.55 ;
      RECT 29.805 4.88 30.095 5.11 ;
      RECT 28.92 4.76 30.02 4.9 ;
      RECT 28.845 4.6 29.135 4.83 ;
      RECT 26.28 10.06 26.57 10.29 ;
      RECT 26.34 8.58 26.51 10.29 ;
      RECT 26.335 8.945 26.685 9.295 ;
      RECT 26.28 8.58 26.57 8.81 ;
      RECT 25.875 3.69 25.98 4.26 ;
      RECT 25.875 4.025 26.2 4.255 ;
      RECT 25.875 4.055 26.37 4.225 ;
      RECT 25.875 3.69 26.065 4.255 ;
      RECT 25.29 3.655 25.58 3.885 ;
      RECT 25.29 3.69 26.065 3.86 ;
      RECT 25.35 2.175 25.52 3.885 ;
      RECT 25.29 2.175 25.58 2.405 ;
      RECT 25.29 10.06 25.58 10.29 ;
      RECT 25.35 8.58 25.52 10.29 ;
      RECT 25.29 8.58 25.58 8.81 ;
      RECT 25.29 8.615 26.14 8.775 ;
      RECT 25.975 8.21 26.14 8.775 ;
      RECT 25.29 8.61 25.685 8.775 ;
      RECT 25.91 8.21 26.2 8.44 ;
      RECT 25.91 8.24 26.37 8.41 ;
      RECT 24.92 4.025 25.21 4.255 ;
      RECT 24.92 4.055 25.38 4.225 ;
      RECT 24.985 2.95 25.15 4.255 ;
      RECT 23.5 2.92 23.79 3.15 ;
      RECT 23.5 2.95 25.15 3.12 ;
      RECT 23.56 2.18 23.73 3.15 ;
      RECT 23.5 2.18 23.79 2.41 ;
      RECT 23.5 10.055 23.79 10.285 ;
      RECT 23.56 9.315 23.73 10.285 ;
      RECT 23.56 9.41 25.15 9.58 ;
      RECT 24.98 8.21 25.15 9.58 ;
      RECT 23.5 9.315 23.79 9.545 ;
      RECT 24.92 8.21 25.21 8.44 ;
      RECT 24.92 8.24 25.38 8.41 ;
      RECT 21.55 3.995 21.89 4.345 ;
      RECT 21.64 3.32 21.81 4.345 ;
      RECT 23.93 3.26 24.28 3.61 ;
      RECT 21.64 3.32 24.28 3.49 ;
      RECT 23.955 8.945 24.28 9.27 ;
      RECT 18.515 8.895 18.865 9.245 ;
      RECT 23.93 8.945 24.28 9.175 ;
      RECT 18.315 8.945 18.865 9.175 ;
      RECT 18.145 8.975 24.28 9.145 ;
      RECT 23.155 3.66 23.475 3.98 ;
      RECT 23.125 3.66 23.475 3.89 ;
      RECT 22.955 3.69 23.475 3.86 ;
      RECT 23.155 8.545 23.475 8.835 ;
      RECT 23.125 8.575 23.475 8.805 ;
      RECT 22.955 8.605 23.475 8.775 ;
      RECT 20.26 3.185 20.58 3.445 ;
      RECT 19.825 3.2 20.115 3.43 ;
      RECT 19.825 3.245 20.58 3.385 ;
      RECT 20.26 4.865 20.58 5.125 ;
      RECT 19.825 4.88 20.115 5.11 ;
      RECT 19.825 4.925 20.58 5.065 ;
      RECT 19.585 4.32 19.875 4.55 ;
      RECT 19.585 4.365 20.16 4.505 ;
      RECT 20.02 4.225 20.28 4.365 ;
      RECT 20.065 4.04 20.355 4.27 ;
      RECT 18.22 4.225 19.32 4.365 ;
      RECT 18.025 4.025 18.345 4.285 ;
      RECT 19.105 4.04 19.395 4.27 ;
      RECT 18.025 4.04 18.435 4.285 ;
      RECT 18.4 3.185 18.72 3.445 ;
      RECT 18.865 3.2 19.155 3.43 ;
      RECT 18.4 3.245 19.155 3.385 ;
      RECT 15.7 4.45 17.88 4.59 ;
      RECT 17.74 3.46 17.88 4.59 ;
      RECT 15.7 4.365 16.995 4.59 ;
      RECT 16.705 4.32 16.995 4.59 ;
      RECT 15.7 4.085 16.035 4.59 ;
      RECT 15.745 4.04 16.035 4.59 ;
      RECT 18.625 3.76 18.915 3.99 ;
      RECT 17.74 3.665 18.84 3.805 ;
      RECT 17.665 3.46 17.955 3.71 ;
      RECT 17.885 10.055 18.175 10.285 ;
      RECT 17.945 9.315 18.115 10.285 ;
      RECT 17.845 9.345 18.215 9.715 ;
      RECT 17.885 9.315 18.175 9.715 ;
      RECT 17.65 4.865 17.97 5.125 ;
      RECT 17.65 4.88 18.165 5.11 ;
      RECT 16.225 3.76 16.515 3.99 ;
      RECT 16.375 3.365 16.515 3.99 ;
      RECT 16.375 3.365 16.68 3.505 ;
      RECT 17.17 3.185 17.49 3.445 ;
      RECT 16.45 3.185 16.77 3.445 ;
      RECT 16.945 3.2 17.49 3.43 ;
      RECT 16.45 3.245 17.49 3.385 ;
      RECT 16.09 4.865 16.41 5.125 ;
      RECT 15.985 4.88 16.41 5.11 ;
      RECT 14.065 4.32 14.355 4.55 ;
      RECT 14.065 4.32 14.52 4.505 ;
      RECT 14.38 3.845 14.52 4.505 ;
      RECT 14.5 3.245 14.64 3.985 ;
      RECT 15.37 3.185 15.69 3.445 ;
      RECT 14.545 3.2 14.835 3.43 ;
      RECT 14.5 3.245 15.69 3.385 ;
      RECT 15.25 3.745 15.57 4.005 ;
      RECT 14.785 3.76 15.075 3.99 ;
      RECT 14.785 3.805 15.57 3.945 ;
      RECT 15.01 4.305 15.33 4.565 ;
      RECT 15.01 4.32 15.555 4.55 ;
      RECT 14.545 4.88 14.835 5.11 ;
      RECT 13.66 4.76 14.76 4.9 ;
      RECT 13.585 4.6 13.875 4.83 ;
      RECT 10.37 10.055 10.66 10.285 ;
      RECT 10.43 9.315 10.6 10.285 ;
      RECT 10.34 9.315 10.69 9.605 ;
      RECT 9.965 8.575 10.315 8.865 ;
      RECT 9.825 8.605 10.315 8.775 ;
      RECT 80.61 3.745 80.93 4.005 ;
      RECT 79.44 4.585 79.76 4.845 ;
      RECT 78.21 4.025 78.53 4.285 ;
      RECT 77.73 3.745 78.05 4.005 ;
      RECT 76.875 3.185 77.275 3.445 ;
      RECT 76.53 4.865 76.85 5.125 ;
      RECT 74.85 3.745 75.17 4.005 ;
      RECT 74.37 4.025 74.69 4.285 ;
      RECT 73.68 4.585 74 4.845 ;
      RECT 65.35 3.745 65.67 4.005 ;
      RECT 64.18 4.585 64.5 4.845 ;
      RECT 62.95 4.025 63.27 4.285 ;
      RECT 62.47 3.745 62.79 4.005 ;
      RECT 61.615 3.185 62.015 3.445 ;
      RECT 61.27 4.865 61.59 5.125 ;
      RECT 59.59 3.745 59.91 4.005 ;
      RECT 59.11 4.025 59.43 4.285 ;
      RECT 58.42 3.185 58.74 3.445 ;
      RECT 58.42 4.585 58.74 4.845 ;
      RECT 50.09 3.745 50.41 4.005 ;
      RECT 48.92 4.585 49.24 4.845 ;
      RECT 47.69 4.025 48.01 4.285 ;
      RECT 47.21 3.745 47.53 4.005 ;
      RECT 46.355 3.185 46.755 3.445 ;
      RECT 46.01 4.865 46.33 5.125 ;
      RECT 44.33 3.745 44.65 4.005 ;
      RECT 43.85 4.025 44.17 4.285 ;
      RECT 43.16 3.185 43.48 3.445 ;
      RECT 43.16 4.585 43.48 4.845 ;
      RECT 34.83 3.745 35.15 4.005 ;
      RECT 33.66 4.585 33.98 4.845 ;
      RECT 32.43 4.025 32.75 4.285 ;
      RECT 31.95 3.745 32.27 4.005 ;
      RECT 31.095 3.185 31.495 3.445 ;
      RECT 30.75 4.865 31.07 5.125 ;
      RECT 29.07 3.745 29.39 4.005 ;
      RECT 28.59 4.025 28.91 4.285 ;
      RECT 27.9 3.185 28.22 3.445 ;
      RECT 27.9 4.585 28.22 4.845 ;
      RECT 19.57 3.745 19.89 4.005 ;
      RECT 18.4 4.585 18.72 4.845 ;
      RECT 17.17 4.025 17.49 4.285 ;
      RECT 16.69 3.745 17.01 4.005 ;
      RECT 15.835 3.185 16.235 3.445 ;
      RECT 15.49 4.865 15.81 5.125 ;
      RECT 13.81 3.745 14.13 4.005 ;
      RECT 13.33 4.025 13.65 4.285 ;
      RECT 12.64 3.185 12.96 3.445 ;
      RECT 12.64 4.585 12.96 4.845 ;
    LAYER mcon ;
      RECT 87.38 8.61 87.55 8.78 ;
      RECT 87.38 10.09 87.55 10.26 ;
      RECT 87.03 1.395 87.2 1.565 ;
      RECT 87.03 10.9 87.2 11.07 ;
      RECT 87.01 4.055 87.18 4.225 ;
      RECT 87.01 8.24 87.18 8.41 ;
      RECT 86.39 2.205 86.56 2.375 ;
      RECT 86.39 3.685 86.56 3.855 ;
      RECT 86.39 8.61 86.56 8.78 ;
      RECT 86.39 10.09 86.56 10.26 ;
      RECT 86.04 1.395 86.21 1.565 ;
      RECT 86.04 10.9 86.21 11.07 ;
      RECT 86.02 4.055 86.19 4.225 ;
      RECT 86.02 8.24 86.19 8.41 ;
      RECT 85.34 1.4 85.51 1.57 ;
      RECT 85.34 10.895 85.51 11.065 ;
      RECT 85.03 3.32 85.2 3.49 ;
      RECT 85.03 8.975 85.2 9.145 ;
      RECT 84.66 1.4 84.83 1.57 ;
      RECT 84.66 10.895 84.83 11.065 ;
      RECT 84.6 2.21 84.77 2.38 ;
      RECT 84.6 2.95 84.77 3.12 ;
      RECT 84.6 9.345 84.77 9.515 ;
      RECT 84.6 10.085 84.77 10.255 ;
      RECT 84.225 3.69 84.395 3.86 ;
      RECT 84.225 8.605 84.395 8.775 ;
      RECT 83.98 1.4 84.15 1.57 ;
      RECT 83.98 10.895 84.15 11.065 ;
      RECT 83.3 1.4 83.47 1.57 ;
      RECT 83.3 10.895 83.47 11.065 ;
      RECT 81.84 2.71 82.01 2.88 ;
      RECT 81.38 2.71 81.55 2.88 ;
      RECT 81.165 4.07 81.335 4.24 ;
      RECT 80.925 3.23 81.095 3.4 ;
      RECT 80.925 4.91 81.095 5.08 ;
      RECT 80.92 2.71 81.09 2.88 ;
      RECT 80.685 3.79 80.855 3.96 ;
      RECT 80.685 4.35 80.855 4.52 ;
      RECT 80.46 2.71 80.63 2.88 ;
      RECT 80.205 4.07 80.375 4.24 ;
      RECT 80 2.71 80.17 2.88 ;
      RECT 79.965 3.23 80.135 3.4 ;
      RECT 79.725 3.79 79.895 3.96 ;
      RECT 79.725 10.895 79.895 11.065 ;
      RECT 79.54 2.71 79.71 2.88 ;
      RECT 79.515 4.63 79.685 4.8 ;
      RECT 79.415 8.975 79.585 9.145 ;
      RECT 79.245 4.07 79.415 4.24 ;
      RECT 79.08 2.71 79.25 2.88 ;
      RECT 79.045 10.895 79.215 11.065 ;
      RECT 78.985 9.345 79.155 9.515 ;
      RECT 78.985 10.085 79.155 10.255 ;
      RECT 78.975 4.91 79.145 5.08 ;
      RECT 78.765 3.49 78.935 3.66 ;
      RECT 78.62 2.71 78.79 2.88 ;
      RECT 78.61 8.605 78.78 8.775 ;
      RECT 78.365 10.895 78.535 11.065 ;
      RECT 78.285 4.07 78.455 4.24 ;
      RECT 78.16 2.71 78.33 2.88 ;
      RECT 78.045 3.23 78.215 3.4 ;
      RECT 77.805 3.79 77.975 3.96 ;
      RECT 77.805 4.35 77.975 4.52 ;
      RECT 77.7 2.71 77.87 2.88 ;
      RECT 77.685 10.895 77.855 11.065 ;
      RECT 77.325 3.79 77.495 3.96 ;
      RECT 77.24 2.71 77.41 2.88 ;
      RECT 77.085 4.91 77.255 5.08 ;
      RECT 77.045 3.23 77.215 3.4 ;
      RECT 76.845 4.07 77.015 4.24 ;
      RECT 76.78 2.71 76.95 2.88 ;
      RECT 76.605 4.91 76.775 5.08 ;
      RECT 76.365 4.35 76.535 4.52 ;
      RECT 76.32 2.71 76.49 2.88 ;
      RECT 75.885 3.79 76.055 3.96 ;
      RECT 75.86 2.71 76.03 2.88 ;
      RECT 75.645 3.23 75.815 3.4 ;
      RECT 75.645 4.91 75.815 5.08 ;
      RECT 75.4 2.71 75.57 2.88 ;
      RECT 75.165 3.23 75.335 3.4 ;
      RECT 75.165 4.35 75.335 4.52 ;
      RECT 74.94 2.71 75.11 2.88 ;
      RECT 74.925 3.79 75.095 3.96 ;
      RECT 74.685 4.63 74.855 4.8 ;
      RECT 74.48 2.71 74.65 2.88 ;
      RECT 74.445 4.07 74.615 4.24 ;
      RECT 74.02 2.71 74.19 2.88 ;
      RECT 73.965 4.07 74.135 4.24 ;
      RECT 73.755 3.23 73.925 3.4 ;
      RECT 73.755 4.63 73.925 4.8 ;
      RECT 73.56 2.71 73.73 2.88 ;
      RECT 72.12 8.61 72.29 8.78 ;
      RECT 72.12 10.09 72.29 10.26 ;
      RECT 71.77 1.395 71.94 1.565 ;
      RECT 71.77 10.9 71.94 11.07 ;
      RECT 71.75 4.055 71.92 4.225 ;
      RECT 71.75 8.24 71.92 8.41 ;
      RECT 71.13 2.205 71.3 2.375 ;
      RECT 71.13 3.685 71.3 3.855 ;
      RECT 71.13 8.61 71.3 8.78 ;
      RECT 71.13 10.09 71.3 10.26 ;
      RECT 70.78 1.395 70.95 1.565 ;
      RECT 70.78 10.9 70.95 11.07 ;
      RECT 70.76 4.055 70.93 4.225 ;
      RECT 70.76 8.24 70.93 8.41 ;
      RECT 70.08 1.4 70.25 1.57 ;
      RECT 70.08 10.895 70.25 11.065 ;
      RECT 69.77 3.32 69.94 3.49 ;
      RECT 69.77 8.975 69.94 9.145 ;
      RECT 69.4 1.4 69.57 1.57 ;
      RECT 69.4 10.895 69.57 11.065 ;
      RECT 69.34 2.21 69.51 2.38 ;
      RECT 69.34 2.95 69.51 3.12 ;
      RECT 69.34 9.345 69.51 9.515 ;
      RECT 69.34 10.085 69.51 10.255 ;
      RECT 68.965 3.69 69.135 3.86 ;
      RECT 68.965 8.605 69.135 8.775 ;
      RECT 68.72 1.4 68.89 1.57 ;
      RECT 68.72 10.895 68.89 11.065 ;
      RECT 68.04 1.4 68.21 1.57 ;
      RECT 68.04 10.895 68.21 11.065 ;
      RECT 66.58 2.71 66.75 2.88 ;
      RECT 66.12 2.71 66.29 2.88 ;
      RECT 65.905 4.07 66.075 4.24 ;
      RECT 65.665 3.23 65.835 3.4 ;
      RECT 65.665 4.91 65.835 5.08 ;
      RECT 65.66 2.71 65.83 2.88 ;
      RECT 65.425 3.79 65.595 3.96 ;
      RECT 65.425 4.35 65.595 4.52 ;
      RECT 65.2 2.71 65.37 2.88 ;
      RECT 64.945 4.07 65.115 4.24 ;
      RECT 64.74 2.71 64.91 2.88 ;
      RECT 64.705 3.23 64.875 3.4 ;
      RECT 64.465 3.79 64.635 3.96 ;
      RECT 64.465 10.895 64.635 11.065 ;
      RECT 64.28 2.71 64.45 2.88 ;
      RECT 64.255 4.63 64.425 4.8 ;
      RECT 64.155 8.975 64.325 9.145 ;
      RECT 63.985 4.07 64.155 4.24 ;
      RECT 63.82 2.71 63.99 2.88 ;
      RECT 63.785 10.895 63.955 11.065 ;
      RECT 63.725 9.345 63.895 9.515 ;
      RECT 63.725 10.085 63.895 10.255 ;
      RECT 63.715 4.91 63.885 5.08 ;
      RECT 63.505 3.49 63.675 3.66 ;
      RECT 63.36 2.71 63.53 2.88 ;
      RECT 63.35 8.605 63.52 8.775 ;
      RECT 63.105 10.895 63.275 11.065 ;
      RECT 63.025 4.07 63.195 4.24 ;
      RECT 62.9 2.71 63.07 2.88 ;
      RECT 62.785 3.23 62.955 3.4 ;
      RECT 62.545 3.79 62.715 3.96 ;
      RECT 62.545 4.35 62.715 4.52 ;
      RECT 62.44 2.71 62.61 2.88 ;
      RECT 62.425 10.895 62.595 11.065 ;
      RECT 62.065 3.79 62.235 3.96 ;
      RECT 61.98 2.71 62.15 2.88 ;
      RECT 61.825 4.91 61.995 5.08 ;
      RECT 61.785 3.23 61.955 3.4 ;
      RECT 61.585 4.07 61.755 4.24 ;
      RECT 61.52 2.71 61.69 2.88 ;
      RECT 61.345 4.91 61.515 5.08 ;
      RECT 61.105 4.35 61.275 4.52 ;
      RECT 61.06 2.71 61.23 2.88 ;
      RECT 60.625 3.79 60.795 3.96 ;
      RECT 60.6 2.71 60.77 2.88 ;
      RECT 60.385 3.23 60.555 3.4 ;
      RECT 60.385 4.91 60.555 5.08 ;
      RECT 60.14 2.71 60.31 2.88 ;
      RECT 59.905 3.23 60.075 3.4 ;
      RECT 59.905 4.35 60.075 4.52 ;
      RECT 59.68 2.71 59.85 2.88 ;
      RECT 59.665 3.79 59.835 3.96 ;
      RECT 59.425 4.63 59.595 4.8 ;
      RECT 59.22 2.71 59.39 2.88 ;
      RECT 59.185 4.07 59.355 4.24 ;
      RECT 58.76 2.71 58.93 2.88 ;
      RECT 58.705 4.07 58.875 4.24 ;
      RECT 58.495 3.23 58.665 3.4 ;
      RECT 58.495 4.63 58.665 4.8 ;
      RECT 58.3 2.71 58.47 2.88 ;
      RECT 56.86 8.61 57.03 8.78 ;
      RECT 56.86 10.09 57.03 10.26 ;
      RECT 56.51 1.395 56.68 1.565 ;
      RECT 56.51 10.9 56.68 11.07 ;
      RECT 56.49 4.055 56.66 4.225 ;
      RECT 56.49 8.24 56.66 8.41 ;
      RECT 55.87 2.205 56.04 2.375 ;
      RECT 55.87 3.685 56.04 3.855 ;
      RECT 55.87 8.61 56.04 8.78 ;
      RECT 55.87 10.09 56.04 10.26 ;
      RECT 55.52 1.395 55.69 1.565 ;
      RECT 55.52 10.9 55.69 11.07 ;
      RECT 55.5 4.055 55.67 4.225 ;
      RECT 55.5 8.24 55.67 8.41 ;
      RECT 54.82 1.4 54.99 1.57 ;
      RECT 54.82 10.895 54.99 11.065 ;
      RECT 54.51 3.32 54.68 3.49 ;
      RECT 54.51 8.975 54.68 9.145 ;
      RECT 54.14 1.4 54.31 1.57 ;
      RECT 54.14 10.895 54.31 11.065 ;
      RECT 54.08 2.21 54.25 2.38 ;
      RECT 54.08 2.95 54.25 3.12 ;
      RECT 54.08 9.345 54.25 9.515 ;
      RECT 54.08 10.085 54.25 10.255 ;
      RECT 53.705 3.69 53.875 3.86 ;
      RECT 53.705 8.605 53.875 8.775 ;
      RECT 53.46 1.4 53.63 1.57 ;
      RECT 53.46 10.895 53.63 11.065 ;
      RECT 52.78 1.4 52.95 1.57 ;
      RECT 52.78 10.895 52.95 11.065 ;
      RECT 51.32 2.71 51.49 2.88 ;
      RECT 50.86 2.71 51.03 2.88 ;
      RECT 50.645 4.07 50.815 4.24 ;
      RECT 50.405 3.23 50.575 3.4 ;
      RECT 50.405 4.91 50.575 5.08 ;
      RECT 50.4 2.71 50.57 2.88 ;
      RECT 50.165 3.79 50.335 3.96 ;
      RECT 50.165 4.35 50.335 4.52 ;
      RECT 49.94 2.71 50.11 2.88 ;
      RECT 49.685 4.07 49.855 4.24 ;
      RECT 49.48 2.71 49.65 2.88 ;
      RECT 49.445 3.23 49.615 3.4 ;
      RECT 49.205 3.79 49.375 3.96 ;
      RECT 49.205 10.895 49.375 11.065 ;
      RECT 49.02 2.71 49.19 2.88 ;
      RECT 48.995 4.63 49.165 4.8 ;
      RECT 48.895 8.975 49.065 9.145 ;
      RECT 48.725 4.07 48.895 4.24 ;
      RECT 48.56 2.71 48.73 2.88 ;
      RECT 48.525 10.895 48.695 11.065 ;
      RECT 48.465 9.345 48.635 9.515 ;
      RECT 48.465 10.085 48.635 10.255 ;
      RECT 48.455 4.91 48.625 5.08 ;
      RECT 48.245 3.49 48.415 3.66 ;
      RECT 48.1 2.71 48.27 2.88 ;
      RECT 48.09 8.605 48.26 8.775 ;
      RECT 47.845 10.895 48.015 11.065 ;
      RECT 47.765 4.07 47.935 4.24 ;
      RECT 47.64 2.71 47.81 2.88 ;
      RECT 47.525 3.23 47.695 3.4 ;
      RECT 47.285 3.79 47.455 3.96 ;
      RECT 47.285 4.35 47.455 4.52 ;
      RECT 47.18 2.71 47.35 2.88 ;
      RECT 47.165 10.895 47.335 11.065 ;
      RECT 46.805 3.79 46.975 3.96 ;
      RECT 46.72 2.71 46.89 2.88 ;
      RECT 46.565 4.91 46.735 5.08 ;
      RECT 46.525 3.23 46.695 3.4 ;
      RECT 46.325 4.07 46.495 4.24 ;
      RECT 46.26 2.71 46.43 2.88 ;
      RECT 46.085 4.91 46.255 5.08 ;
      RECT 45.845 4.35 46.015 4.52 ;
      RECT 45.8 2.71 45.97 2.88 ;
      RECT 45.365 3.79 45.535 3.96 ;
      RECT 45.34 2.71 45.51 2.88 ;
      RECT 45.125 3.23 45.295 3.4 ;
      RECT 45.125 4.91 45.295 5.08 ;
      RECT 44.88 2.71 45.05 2.88 ;
      RECT 44.645 3.23 44.815 3.4 ;
      RECT 44.645 4.35 44.815 4.52 ;
      RECT 44.42 2.71 44.59 2.88 ;
      RECT 44.405 3.79 44.575 3.96 ;
      RECT 44.165 4.63 44.335 4.8 ;
      RECT 43.96 2.71 44.13 2.88 ;
      RECT 43.925 4.07 44.095 4.24 ;
      RECT 43.5 2.71 43.67 2.88 ;
      RECT 43.445 4.07 43.615 4.24 ;
      RECT 43.235 3.23 43.405 3.4 ;
      RECT 43.235 4.63 43.405 4.8 ;
      RECT 43.04 2.71 43.21 2.88 ;
      RECT 41.6 8.61 41.77 8.78 ;
      RECT 41.6 10.09 41.77 10.26 ;
      RECT 41.25 1.395 41.42 1.565 ;
      RECT 41.25 10.9 41.42 11.07 ;
      RECT 41.23 4.055 41.4 4.225 ;
      RECT 41.23 8.24 41.4 8.41 ;
      RECT 40.61 2.205 40.78 2.375 ;
      RECT 40.61 3.685 40.78 3.855 ;
      RECT 40.61 8.61 40.78 8.78 ;
      RECT 40.61 10.09 40.78 10.26 ;
      RECT 40.26 1.395 40.43 1.565 ;
      RECT 40.26 10.9 40.43 11.07 ;
      RECT 40.24 4.055 40.41 4.225 ;
      RECT 40.24 8.24 40.41 8.41 ;
      RECT 39.56 1.4 39.73 1.57 ;
      RECT 39.56 10.895 39.73 11.065 ;
      RECT 39.25 3.32 39.42 3.49 ;
      RECT 39.25 8.975 39.42 9.145 ;
      RECT 38.88 1.4 39.05 1.57 ;
      RECT 38.88 10.895 39.05 11.065 ;
      RECT 38.82 2.21 38.99 2.38 ;
      RECT 38.82 2.95 38.99 3.12 ;
      RECT 38.82 9.345 38.99 9.515 ;
      RECT 38.82 10.085 38.99 10.255 ;
      RECT 38.445 3.69 38.615 3.86 ;
      RECT 38.445 8.605 38.615 8.775 ;
      RECT 38.2 1.4 38.37 1.57 ;
      RECT 38.2 10.895 38.37 11.065 ;
      RECT 37.52 1.4 37.69 1.57 ;
      RECT 37.52 10.895 37.69 11.065 ;
      RECT 36.06 2.71 36.23 2.88 ;
      RECT 35.6 2.71 35.77 2.88 ;
      RECT 35.385 4.07 35.555 4.24 ;
      RECT 35.145 3.23 35.315 3.4 ;
      RECT 35.145 4.91 35.315 5.08 ;
      RECT 35.14 2.71 35.31 2.88 ;
      RECT 34.905 3.79 35.075 3.96 ;
      RECT 34.905 4.35 35.075 4.52 ;
      RECT 34.68 2.71 34.85 2.88 ;
      RECT 34.425 4.07 34.595 4.24 ;
      RECT 34.22 2.71 34.39 2.88 ;
      RECT 34.185 3.23 34.355 3.4 ;
      RECT 33.945 3.79 34.115 3.96 ;
      RECT 33.945 10.895 34.115 11.065 ;
      RECT 33.76 2.71 33.93 2.88 ;
      RECT 33.735 4.63 33.905 4.8 ;
      RECT 33.635 8.975 33.805 9.145 ;
      RECT 33.465 4.07 33.635 4.24 ;
      RECT 33.3 2.71 33.47 2.88 ;
      RECT 33.265 10.895 33.435 11.065 ;
      RECT 33.205 9.345 33.375 9.515 ;
      RECT 33.205 10.085 33.375 10.255 ;
      RECT 33.195 4.91 33.365 5.08 ;
      RECT 32.985 3.49 33.155 3.66 ;
      RECT 32.84 2.71 33.01 2.88 ;
      RECT 32.83 8.605 33 8.775 ;
      RECT 32.585 10.895 32.755 11.065 ;
      RECT 32.505 4.07 32.675 4.24 ;
      RECT 32.38 2.71 32.55 2.88 ;
      RECT 32.265 3.23 32.435 3.4 ;
      RECT 32.025 3.79 32.195 3.96 ;
      RECT 32.025 4.35 32.195 4.52 ;
      RECT 31.92 2.71 32.09 2.88 ;
      RECT 31.905 10.895 32.075 11.065 ;
      RECT 31.545 3.79 31.715 3.96 ;
      RECT 31.46 2.71 31.63 2.88 ;
      RECT 31.305 4.91 31.475 5.08 ;
      RECT 31.265 3.23 31.435 3.4 ;
      RECT 31.065 4.07 31.235 4.24 ;
      RECT 31 2.71 31.17 2.88 ;
      RECT 30.825 4.91 30.995 5.08 ;
      RECT 30.585 4.35 30.755 4.52 ;
      RECT 30.54 2.71 30.71 2.88 ;
      RECT 30.105 3.79 30.275 3.96 ;
      RECT 30.08 2.71 30.25 2.88 ;
      RECT 29.865 3.23 30.035 3.4 ;
      RECT 29.865 4.91 30.035 5.08 ;
      RECT 29.62 2.71 29.79 2.88 ;
      RECT 29.385 3.23 29.555 3.4 ;
      RECT 29.385 4.35 29.555 4.52 ;
      RECT 29.16 2.71 29.33 2.88 ;
      RECT 29.145 3.79 29.315 3.96 ;
      RECT 28.905 4.63 29.075 4.8 ;
      RECT 28.7 2.71 28.87 2.88 ;
      RECT 28.665 4.07 28.835 4.24 ;
      RECT 28.24 2.71 28.41 2.88 ;
      RECT 28.185 4.07 28.355 4.24 ;
      RECT 27.975 3.23 28.145 3.4 ;
      RECT 27.975 4.63 28.145 4.8 ;
      RECT 27.78 2.71 27.95 2.88 ;
      RECT 26.34 8.61 26.51 8.78 ;
      RECT 26.34 10.09 26.51 10.26 ;
      RECT 25.99 1.395 26.16 1.565 ;
      RECT 25.99 10.9 26.16 11.07 ;
      RECT 25.97 4.055 26.14 4.225 ;
      RECT 25.97 8.24 26.14 8.41 ;
      RECT 25.35 2.205 25.52 2.375 ;
      RECT 25.35 3.685 25.52 3.855 ;
      RECT 25.35 8.61 25.52 8.78 ;
      RECT 25.35 10.09 25.52 10.26 ;
      RECT 25 1.395 25.17 1.565 ;
      RECT 25 10.9 25.17 11.07 ;
      RECT 24.98 4.055 25.15 4.225 ;
      RECT 24.98 8.24 25.15 8.41 ;
      RECT 24.3 1.4 24.47 1.57 ;
      RECT 24.3 10.895 24.47 11.065 ;
      RECT 23.99 3.32 24.16 3.49 ;
      RECT 23.99 8.975 24.16 9.145 ;
      RECT 23.62 1.4 23.79 1.57 ;
      RECT 23.62 10.895 23.79 11.065 ;
      RECT 23.56 2.21 23.73 2.38 ;
      RECT 23.56 2.95 23.73 3.12 ;
      RECT 23.56 9.345 23.73 9.515 ;
      RECT 23.56 10.085 23.73 10.255 ;
      RECT 23.185 3.69 23.355 3.86 ;
      RECT 23.185 8.605 23.355 8.775 ;
      RECT 22.94 1.4 23.11 1.57 ;
      RECT 22.94 10.895 23.11 11.065 ;
      RECT 22.26 1.4 22.43 1.57 ;
      RECT 22.26 10.895 22.43 11.065 ;
      RECT 20.8 2.71 20.97 2.88 ;
      RECT 20.34 2.71 20.51 2.88 ;
      RECT 20.125 4.07 20.295 4.24 ;
      RECT 19.885 3.23 20.055 3.4 ;
      RECT 19.885 4.91 20.055 5.08 ;
      RECT 19.88 2.71 20.05 2.88 ;
      RECT 19.645 3.79 19.815 3.96 ;
      RECT 19.645 4.35 19.815 4.52 ;
      RECT 19.42 2.71 19.59 2.88 ;
      RECT 19.165 4.07 19.335 4.24 ;
      RECT 18.96 2.71 19.13 2.88 ;
      RECT 18.925 3.23 19.095 3.4 ;
      RECT 18.685 3.79 18.855 3.96 ;
      RECT 18.685 10.895 18.855 11.065 ;
      RECT 18.5 2.71 18.67 2.88 ;
      RECT 18.475 4.63 18.645 4.8 ;
      RECT 18.375 8.975 18.545 9.145 ;
      RECT 18.205 4.07 18.375 4.24 ;
      RECT 18.04 2.71 18.21 2.88 ;
      RECT 18.005 10.895 18.175 11.065 ;
      RECT 17.945 9.345 18.115 9.515 ;
      RECT 17.945 10.085 18.115 10.255 ;
      RECT 17.935 4.91 18.105 5.08 ;
      RECT 17.725 3.49 17.895 3.66 ;
      RECT 17.58 2.71 17.75 2.88 ;
      RECT 17.57 8.605 17.74 8.775 ;
      RECT 17.325 10.895 17.495 11.065 ;
      RECT 17.245 4.07 17.415 4.24 ;
      RECT 17.12 2.71 17.29 2.88 ;
      RECT 17.005 3.23 17.175 3.4 ;
      RECT 16.765 3.79 16.935 3.96 ;
      RECT 16.765 4.35 16.935 4.52 ;
      RECT 16.66 2.71 16.83 2.88 ;
      RECT 16.645 10.895 16.815 11.065 ;
      RECT 16.285 3.79 16.455 3.96 ;
      RECT 16.2 2.71 16.37 2.88 ;
      RECT 16.045 4.91 16.215 5.08 ;
      RECT 16.005 3.23 16.175 3.4 ;
      RECT 15.805 4.07 15.975 4.24 ;
      RECT 15.74 2.71 15.91 2.88 ;
      RECT 15.565 4.91 15.735 5.08 ;
      RECT 15.325 4.35 15.495 4.52 ;
      RECT 15.28 2.71 15.45 2.88 ;
      RECT 14.845 3.79 15.015 3.96 ;
      RECT 14.82 2.71 14.99 2.88 ;
      RECT 14.605 3.23 14.775 3.4 ;
      RECT 14.605 4.91 14.775 5.08 ;
      RECT 14.36 2.71 14.53 2.88 ;
      RECT 14.125 3.23 14.295 3.4 ;
      RECT 14.125 4.35 14.295 4.52 ;
      RECT 13.9 2.71 14.07 2.88 ;
      RECT 13.885 3.79 14.055 3.96 ;
      RECT 13.645 4.63 13.815 4.8 ;
      RECT 13.44 2.71 13.61 2.88 ;
      RECT 13.405 4.07 13.575 4.24 ;
      RECT 12.98 2.71 13.15 2.88 ;
      RECT 12.925 4.07 13.095 4.24 ;
      RECT 12.715 3.23 12.885 3.4 ;
      RECT 12.715 4.63 12.885 4.8 ;
      RECT 12.52 2.71 12.69 2.88 ;
      RECT 11.17 10.895 11.34 11.065 ;
      RECT 10.49 10.895 10.66 11.065 ;
      RECT 10.43 9.345 10.6 9.515 ;
      RECT 10.43 10.085 10.6 10.255 ;
      RECT 10.055 8.605 10.225 8.775 ;
      RECT 9.81 10.895 9.98 11.065 ;
      RECT 9.13 10.895 9.3 11.065 ;
    LAYER li1 ;
      RECT 81.385 0 81.555 3.38 ;
      RECT 80.445 0 80.615 3.38 ;
      RECT 79.485 0 79.655 3.38 ;
      RECT 77.565 0 77.735 3.38 ;
      RECT 76.605 0 76.775 3.38 ;
      RECT 74.685 0 74.855 3.38 ;
      RECT 66.125 0 66.295 3.38 ;
      RECT 65.185 0 65.355 3.38 ;
      RECT 64.225 0 64.395 3.38 ;
      RECT 62.305 0 62.475 3.38 ;
      RECT 61.345 0 61.515 3.38 ;
      RECT 59.425 0 59.595 3.38 ;
      RECT 50.865 0 51.035 3.38 ;
      RECT 49.925 0 50.095 3.38 ;
      RECT 48.965 0 49.135 3.38 ;
      RECT 47.045 0 47.215 3.38 ;
      RECT 46.085 0 46.255 3.38 ;
      RECT 44.165 0 44.335 3.38 ;
      RECT 35.605 0 35.775 3.38 ;
      RECT 34.665 0 34.835 3.38 ;
      RECT 33.705 0 33.875 3.38 ;
      RECT 31.785 0 31.955 3.38 ;
      RECT 30.825 0 30.995 3.38 ;
      RECT 28.905 0 29.075 3.38 ;
      RECT 20.345 0 20.515 3.38 ;
      RECT 19.405 0 19.575 3.38 ;
      RECT 18.445 0 18.615 3.38 ;
      RECT 16.525 0 16.695 3.38 ;
      RECT 15.565 0 15.735 3.38 ;
      RECT 13.645 0 13.815 3.38 ;
      RECT 78.44 0 78.635 2.89 ;
      RECT 74.685 0 74.96 2.89 ;
      RECT 63.18 0 63.375 2.89 ;
      RECT 59.425 0 59.7 2.89 ;
      RECT 47.92 0 48.115 2.89 ;
      RECT 44.165 0 44.44 2.89 ;
      RECT 32.66 0 32.855 2.89 ;
      RECT 28.905 0 29.18 2.89 ;
      RECT 17.4 0 17.595 2.89 ;
      RECT 13.645 0 13.92 2.89 ;
      RECT 73.415 0 82.155 2.88 ;
      RECT 58.155 0 66.895 2.88 ;
      RECT 42.895 0 51.635 2.88 ;
      RECT 27.635 0 36.375 2.88 ;
      RECT 12.375 0 21.115 2.88 ;
      RECT 83.22 0 83.39 2.23 ;
      RECT 67.96 0 68.13 2.23 ;
      RECT 52.7 0 52.87 2.23 ;
      RECT 37.44 0 37.61 2.23 ;
      RECT 22.18 0 22.35 2.23 ;
      RECT 86.95 0 87.12 2.225 ;
      RECT 85.96 0 86.13 2.225 ;
      RECT 71.69 0 71.86 2.225 ;
      RECT 70.7 0 70.87 2.225 ;
      RECT 56.43 0 56.6 2.225 ;
      RECT 55.44 0 55.61 2.225 ;
      RECT 41.17 0 41.34 2.225 ;
      RECT 40.18 0 40.35 2.225 ;
      RECT 25.91 0 26.08 2.225 ;
      RECT 24.92 0 25.09 2.225 ;
      RECT 8.88 0 87.925 1.6 ;
      RECT 8.83 10.865 87.925 12.465 ;
      RECT 86.95 10.24 87.12 12.465 ;
      RECT 85.96 10.24 86.13 12.465 ;
      RECT 83.22 10.235 83.39 12.465 ;
      RECT 77.605 10.235 77.775 12.465 ;
      RECT 71.69 10.24 71.86 12.465 ;
      RECT 70.7 10.24 70.87 12.465 ;
      RECT 67.96 10.235 68.13 12.465 ;
      RECT 62.345 10.235 62.515 12.465 ;
      RECT 56.43 10.24 56.6 12.465 ;
      RECT 55.44 10.24 55.61 12.465 ;
      RECT 52.7 10.235 52.87 12.465 ;
      RECT 47.085 10.235 47.255 12.465 ;
      RECT 41.17 10.24 41.34 12.465 ;
      RECT 40.18 10.24 40.35 12.465 ;
      RECT 37.44 10.235 37.61 12.465 ;
      RECT 31.825 10.235 31.995 12.465 ;
      RECT 25.91 10.24 26.08 12.465 ;
      RECT 24.92 10.24 25.09 12.465 ;
      RECT 22.18 10.235 22.35 12.465 ;
      RECT 16.565 10.235 16.735 12.465 ;
      RECT 9.05 10.235 9.22 12.465 ;
      RECT 87.01 3.035 87.18 4.225 ;
      RECT 87.01 3.035 87.48 3.205 ;
      RECT 87.01 9.26 87.48 9.43 ;
      RECT 87.01 8.24 87.18 9.43 ;
      RECT 86.02 3.035 86.19 4.225 ;
      RECT 86.02 3.035 86.49 3.205 ;
      RECT 86.02 9.26 86.49 9.43 ;
      RECT 86.02 8.24 86.19 9.43 ;
      RECT 84.17 3.93 84.34 5.16 ;
      RECT 84.225 2.15 84.395 4.1 ;
      RECT 84.17 1.87 84.34 2.32 ;
      RECT 84.17 10.145 84.34 10.595 ;
      RECT 84.225 8.365 84.395 10.315 ;
      RECT 84.17 7.305 84.34 8.535 ;
      RECT 83.65 1.87 83.82 5.16 ;
      RECT 83.65 3.37 84.055 3.7 ;
      RECT 83.65 2.53 84.055 2.86 ;
      RECT 83.65 7.305 83.82 10.595 ;
      RECT 83.65 9.605 84.055 9.935 ;
      RECT 83.65 8.765 84.055 9.095 ;
      RECT 80.925 4.91 81.44 5.08 ;
      RECT 81.27 4.52 81.44 5.08 ;
      RECT 81.375 4.44 81.545 4.77 ;
      RECT 81.165 3.83 81.44 4.24 ;
      RECT 81.045 3.83 81.44 4.04 ;
      RECT 79.515 4.44 79.685 4.8 ;
      RECT 79.515 4.52 80.855 4.69 ;
      RECT 80.685 4.35 80.855 4.69 ;
      RECT 79.245 3.87 79.415 4.24 ;
      RECT 78.765 3.87 79.415 4.14 ;
      RECT 78.685 3.87 79.495 4.04 ;
      RECT 78.045 3.11 78.215 3.4 ;
      RECT 78.045 3.11 79.285 3.28 ;
      RECT 78.765 3.45 78.935 3.66 ;
      RECT 78.405 3.45 78.935 3.62 ;
      RECT 78.555 10.145 78.725 10.595 ;
      RECT 78.61 8.365 78.78 10.315 ;
      RECT 78.555 7.305 78.725 8.535 ;
      RECT 78.035 7.305 78.205 10.595 ;
      RECT 78.035 9.605 78.44 9.935 ;
      RECT 78.035 8.765 78.44 9.095 ;
      RECT 77.805 4.52 78.295 4.69 ;
      RECT 77.805 4.35 77.975 4.69 ;
      RECT 77.085 4.52 77.255 5.08 ;
      RECT 76.975 4.52 77.305 4.69 ;
      RECT 77.045 3.13 77.215 3.4 ;
      RECT 77.085 3.05 77.255 3.38 ;
      RECT 76.95 3.13 77.255 3.35 ;
      RECT 75.525 4.52 75.815 5.08 ;
      RECT 75.645 4.44 75.815 5.08 ;
      RECT 75.285 3.87 75.655 4.04 ;
      RECT 75.285 3.23 75.455 4.04 ;
      RECT 75.165 3.23 75.455 3.4 ;
      RECT 73.595 3.225 74.165 3.685 ;
      RECT 73.755 3.05 73.925 3.685 ;
      RECT 71.75 3.035 71.92 4.225 ;
      RECT 71.75 3.035 72.22 3.205 ;
      RECT 71.75 9.26 72.22 9.43 ;
      RECT 71.75 8.24 71.92 9.43 ;
      RECT 70.76 3.035 70.93 4.225 ;
      RECT 70.76 3.035 71.23 3.205 ;
      RECT 70.76 9.26 71.23 9.43 ;
      RECT 70.76 8.24 70.93 9.43 ;
      RECT 68.91 3.93 69.08 5.16 ;
      RECT 68.965 2.15 69.135 4.1 ;
      RECT 68.91 1.87 69.08 2.32 ;
      RECT 68.91 10.145 69.08 10.595 ;
      RECT 68.965 8.365 69.135 10.315 ;
      RECT 68.91 7.305 69.08 8.535 ;
      RECT 68.39 1.87 68.56 5.16 ;
      RECT 68.39 3.37 68.795 3.7 ;
      RECT 68.39 2.53 68.795 2.86 ;
      RECT 68.39 7.305 68.56 10.595 ;
      RECT 68.39 9.605 68.795 9.935 ;
      RECT 68.39 8.765 68.795 9.095 ;
      RECT 65.665 4.91 66.18 5.08 ;
      RECT 66.01 4.52 66.18 5.08 ;
      RECT 66.115 4.44 66.285 4.77 ;
      RECT 65.905 3.83 66.18 4.24 ;
      RECT 65.785 3.83 66.18 4.04 ;
      RECT 64.255 4.44 64.425 4.8 ;
      RECT 64.255 4.52 65.595 4.69 ;
      RECT 65.425 4.35 65.595 4.69 ;
      RECT 63.985 3.87 64.155 4.24 ;
      RECT 63.505 3.87 64.155 4.14 ;
      RECT 63.425 3.87 64.235 4.04 ;
      RECT 62.785 3.11 62.955 3.4 ;
      RECT 62.785 3.11 64.025 3.28 ;
      RECT 63.505 3.45 63.675 3.66 ;
      RECT 63.145 3.45 63.675 3.62 ;
      RECT 63.295 10.145 63.465 10.595 ;
      RECT 63.35 8.365 63.52 10.315 ;
      RECT 63.295 7.305 63.465 8.535 ;
      RECT 62.775 7.305 62.945 10.595 ;
      RECT 62.775 9.605 63.18 9.935 ;
      RECT 62.775 8.765 63.18 9.095 ;
      RECT 62.545 4.52 63.035 4.69 ;
      RECT 62.545 4.35 62.715 4.69 ;
      RECT 61.825 4.52 61.995 5.08 ;
      RECT 61.715 4.52 62.045 4.69 ;
      RECT 61.785 3.13 61.955 3.4 ;
      RECT 61.825 3.05 61.995 3.38 ;
      RECT 61.69 3.13 61.995 3.35 ;
      RECT 60.265 4.52 60.555 5.08 ;
      RECT 60.385 4.44 60.555 5.08 ;
      RECT 60.025 3.87 60.395 4.04 ;
      RECT 60.025 3.23 60.195 4.04 ;
      RECT 59.905 3.23 60.195 3.4 ;
      RECT 56.49 3.035 56.66 4.225 ;
      RECT 56.49 3.035 56.96 3.205 ;
      RECT 56.49 9.26 56.96 9.43 ;
      RECT 56.49 8.24 56.66 9.43 ;
      RECT 55.5 3.035 55.67 4.225 ;
      RECT 55.5 3.035 55.97 3.205 ;
      RECT 55.5 9.26 55.97 9.43 ;
      RECT 55.5 8.24 55.67 9.43 ;
      RECT 53.65 3.93 53.82 5.16 ;
      RECT 53.705 2.15 53.875 4.1 ;
      RECT 53.65 1.87 53.82 2.32 ;
      RECT 53.65 10.145 53.82 10.595 ;
      RECT 53.705 8.365 53.875 10.315 ;
      RECT 53.65 7.305 53.82 8.535 ;
      RECT 53.13 1.87 53.3 5.16 ;
      RECT 53.13 3.37 53.535 3.7 ;
      RECT 53.13 2.53 53.535 2.86 ;
      RECT 53.13 7.305 53.3 10.595 ;
      RECT 53.13 9.605 53.535 9.935 ;
      RECT 53.13 8.765 53.535 9.095 ;
      RECT 50.405 4.91 50.92 5.08 ;
      RECT 50.75 4.52 50.92 5.08 ;
      RECT 50.855 4.44 51.025 4.77 ;
      RECT 50.645 3.83 50.92 4.24 ;
      RECT 50.525 3.83 50.92 4.04 ;
      RECT 48.995 4.44 49.165 4.8 ;
      RECT 48.995 4.52 50.335 4.69 ;
      RECT 50.165 4.35 50.335 4.69 ;
      RECT 48.725 3.87 48.895 4.24 ;
      RECT 48.245 3.87 48.895 4.14 ;
      RECT 48.165 3.87 48.975 4.04 ;
      RECT 47.525 3.11 47.695 3.4 ;
      RECT 47.525 3.11 48.765 3.28 ;
      RECT 48.245 3.45 48.415 3.66 ;
      RECT 47.885 3.45 48.415 3.62 ;
      RECT 48.035 10.145 48.205 10.595 ;
      RECT 48.09 8.365 48.26 10.315 ;
      RECT 48.035 7.305 48.205 8.535 ;
      RECT 47.515 7.305 47.685 10.595 ;
      RECT 47.515 9.605 47.92 9.935 ;
      RECT 47.515 8.765 47.92 9.095 ;
      RECT 47.285 4.52 47.775 4.69 ;
      RECT 47.285 4.35 47.455 4.69 ;
      RECT 46.565 4.52 46.735 5.08 ;
      RECT 46.455 4.52 46.785 4.69 ;
      RECT 46.525 3.13 46.695 3.4 ;
      RECT 46.565 3.05 46.735 3.38 ;
      RECT 46.43 3.13 46.735 3.35 ;
      RECT 45.005 4.52 45.295 5.08 ;
      RECT 45.125 4.44 45.295 5.08 ;
      RECT 44.765 3.87 45.135 4.04 ;
      RECT 44.765 3.23 44.935 4.04 ;
      RECT 44.645 3.23 44.935 3.4 ;
      RECT 41.23 3.035 41.4 4.225 ;
      RECT 41.23 3.035 41.7 3.205 ;
      RECT 41.23 9.26 41.7 9.43 ;
      RECT 41.23 8.24 41.4 9.43 ;
      RECT 40.24 3.035 40.41 4.225 ;
      RECT 40.24 3.035 40.71 3.205 ;
      RECT 40.24 9.26 40.71 9.43 ;
      RECT 40.24 8.24 40.41 9.43 ;
      RECT 38.39 3.93 38.56 5.16 ;
      RECT 38.445 2.15 38.615 4.1 ;
      RECT 38.39 1.87 38.56 2.32 ;
      RECT 38.39 10.145 38.56 10.595 ;
      RECT 38.445 8.365 38.615 10.315 ;
      RECT 38.39 7.305 38.56 8.535 ;
      RECT 37.87 1.87 38.04 5.16 ;
      RECT 37.87 3.37 38.275 3.7 ;
      RECT 37.87 2.53 38.275 2.86 ;
      RECT 37.87 7.305 38.04 10.595 ;
      RECT 37.87 9.605 38.275 9.935 ;
      RECT 37.87 8.765 38.275 9.095 ;
      RECT 35.145 4.91 35.66 5.08 ;
      RECT 35.49 4.52 35.66 5.08 ;
      RECT 35.595 4.44 35.765 4.77 ;
      RECT 35.385 3.83 35.66 4.24 ;
      RECT 35.265 3.83 35.66 4.04 ;
      RECT 33.735 4.44 33.905 4.8 ;
      RECT 33.735 4.52 35.075 4.69 ;
      RECT 34.905 4.35 35.075 4.69 ;
      RECT 33.465 3.87 33.635 4.24 ;
      RECT 32.985 3.87 33.635 4.14 ;
      RECT 32.905 3.87 33.715 4.04 ;
      RECT 32.265 3.11 32.435 3.4 ;
      RECT 32.265 3.11 33.505 3.28 ;
      RECT 32.985 3.45 33.155 3.66 ;
      RECT 32.625 3.45 33.155 3.62 ;
      RECT 32.775 10.145 32.945 10.595 ;
      RECT 32.83 8.365 33 10.315 ;
      RECT 32.775 7.305 32.945 8.535 ;
      RECT 32.255 7.305 32.425 10.595 ;
      RECT 32.255 9.605 32.66 9.935 ;
      RECT 32.255 8.765 32.66 9.095 ;
      RECT 32.025 4.52 32.515 4.69 ;
      RECT 32.025 4.35 32.195 4.69 ;
      RECT 31.305 4.52 31.475 5.08 ;
      RECT 31.195 4.52 31.525 4.69 ;
      RECT 31.265 3.13 31.435 3.4 ;
      RECT 31.305 3.05 31.475 3.38 ;
      RECT 31.17 3.13 31.475 3.35 ;
      RECT 29.745 4.52 30.035 5.08 ;
      RECT 29.865 4.44 30.035 5.08 ;
      RECT 29.505 3.87 29.875 4.04 ;
      RECT 29.505 3.23 29.675 4.04 ;
      RECT 29.385 3.23 29.675 3.4 ;
      RECT 25.97 3.035 26.14 4.225 ;
      RECT 25.97 3.035 26.44 3.205 ;
      RECT 25.97 9.26 26.44 9.43 ;
      RECT 25.97 8.24 26.14 9.43 ;
      RECT 24.98 3.035 25.15 4.225 ;
      RECT 24.98 3.035 25.45 3.205 ;
      RECT 24.98 9.26 25.45 9.43 ;
      RECT 24.98 8.24 25.15 9.43 ;
      RECT 23.13 3.93 23.3 5.16 ;
      RECT 23.185 2.15 23.355 4.1 ;
      RECT 23.13 1.87 23.3 2.32 ;
      RECT 23.13 10.145 23.3 10.595 ;
      RECT 23.185 8.365 23.355 10.315 ;
      RECT 23.13 7.305 23.3 8.535 ;
      RECT 22.61 1.87 22.78 5.16 ;
      RECT 22.61 3.37 23.015 3.7 ;
      RECT 22.61 2.53 23.015 2.86 ;
      RECT 22.61 7.305 22.78 10.595 ;
      RECT 22.61 9.605 23.015 9.935 ;
      RECT 22.61 8.765 23.015 9.095 ;
      RECT 19.885 4.91 20.4 5.08 ;
      RECT 20.23 4.52 20.4 5.08 ;
      RECT 20.335 4.44 20.505 4.77 ;
      RECT 20.125 3.83 20.4 4.24 ;
      RECT 20.005 3.83 20.4 4.04 ;
      RECT 18.475 4.44 18.645 4.8 ;
      RECT 18.475 4.52 19.815 4.69 ;
      RECT 19.645 4.35 19.815 4.69 ;
      RECT 18.205 3.87 18.375 4.24 ;
      RECT 17.725 3.87 18.375 4.14 ;
      RECT 17.645 3.87 18.455 4.04 ;
      RECT 17.005 3.11 17.175 3.4 ;
      RECT 17.005 3.11 18.245 3.28 ;
      RECT 17.725 3.45 17.895 3.66 ;
      RECT 17.365 3.45 17.895 3.62 ;
      RECT 17.515 10.145 17.685 10.595 ;
      RECT 17.57 8.365 17.74 10.315 ;
      RECT 17.515 7.305 17.685 8.535 ;
      RECT 16.995 7.305 17.165 10.595 ;
      RECT 16.995 9.605 17.4 9.935 ;
      RECT 16.995 8.765 17.4 9.095 ;
      RECT 16.765 4.52 17.255 4.69 ;
      RECT 16.765 4.35 16.935 4.69 ;
      RECT 16.045 4.52 16.215 5.08 ;
      RECT 15.935 4.52 16.265 4.69 ;
      RECT 16.005 3.13 16.175 3.4 ;
      RECT 16.045 3.05 16.215 3.38 ;
      RECT 15.91 3.13 16.215 3.35 ;
      RECT 14.485 4.52 14.775 5.08 ;
      RECT 14.605 4.44 14.775 5.08 ;
      RECT 14.245 3.87 14.615 4.04 ;
      RECT 14.245 3.23 14.415 4.04 ;
      RECT 14.125 3.23 14.415 3.4 ;
      RECT 10 10.145 10.17 10.595 ;
      RECT 10.055 8.365 10.225 10.315 ;
      RECT 10 7.305 10.17 8.535 ;
      RECT 9.48 7.305 9.65 10.595 ;
      RECT 9.48 9.605 9.885 9.935 ;
      RECT 9.48 8.765 9.885 9.095 ;
      RECT 87.38 7.31 87.55 8.78 ;
      RECT 87.38 10.09 87.55 10.6 ;
      RECT 86.39 1.865 86.56 2.375 ;
      RECT 86.39 3.685 86.56 5.155 ;
      RECT 86.39 7.31 86.56 8.78 ;
      RECT 86.39 10.09 86.56 10.6 ;
      RECT 85.03 1.87 85.2 5.16 ;
      RECT 85.03 7.305 85.2 10.595 ;
      RECT 84.6 1.87 84.77 2.38 ;
      RECT 84.6 2.95 84.77 5.16 ;
      RECT 84.6 7.305 84.77 9.515 ;
      RECT 84.6 10.085 84.77 10.595 ;
      RECT 80.925 3.05 81.095 3.4 ;
      RECT 80.685 3.79 80.855 4.12 ;
      RECT 80.205 3.79 80.375 4.24 ;
      RECT 79.965 3.05 80.135 3.4 ;
      RECT 79.725 3.79 79.895 4.12 ;
      RECT 79.415 7.305 79.585 10.595 ;
      RECT 78.985 7.305 79.155 9.515 ;
      RECT 78.985 10.085 79.155 10.595 ;
      RECT 78.975 4.78 79.145 5.11 ;
      RECT 78.285 3.79 78.455 4.24 ;
      RECT 77.805 3.79 77.975 4.12 ;
      RECT 77.325 3.79 77.495 4.12 ;
      RECT 76.845 3.79 77.015 4.24 ;
      RECT 76.605 4.78 76.775 5.11 ;
      RECT 76.365 3.79 76.535 4.52 ;
      RECT 75.885 3.79 76.055 4.12 ;
      RECT 75.645 3.05 75.815 3.4 ;
      RECT 75.165 4.35 75.335 4.77 ;
      RECT 74.925 3.79 75.095 4.12 ;
      RECT 74.685 4.44 74.855 4.8 ;
      RECT 74.445 3.79 74.615 4.24 ;
      RECT 73.965 3.79 74.135 4.24 ;
      RECT 73.755 4.44 73.925 4.8 ;
      RECT 72.12 7.31 72.29 8.78 ;
      RECT 72.12 10.09 72.29 10.6 ;
      RECT 71.13 1.865 71.3 2.375 ;
      RECT 71.13 3.685 71.3 5.155 ;
      RECT 71.13 7.31 71.3 8.78 ;
      RECT 71.13 10.09 71.3 10.6 ;
      RECT 69.77 1.87 69.94 5.16 ;
      RECT 69.77 7.305 69.94 10.595 ;
      RECT 69.34 1.87 69.51 2.38 ;
      RECT 69.34 2.95 69.51 5.16 ;
      RECT 69.34 7.305 69.51 9.515 ;
      RECT 69.34 10.085 69.51 10.595 ;
      RECT 65.665 3.05 65.835 3.4 ;
      RECT 65.425 3.79 65.595 4.12 ;
      RECT 64.945 3.79 65.115 4.24 ;
      RECT 64.705 3.05 64.875 3.4 ;
      RECT 64.465 3.79 64.635 4.12 ;
      RECT 64.155 7.305 64.325 10.595 ;
      RECT 63.725 7.305 63.895 9.515 ;
      RECT 63.725 10.085 63.895 10.595 ;
      RECT 63.715 4.78 63.885 5.11 ;
      RECT 63.025 3.79 63.195 4.24 ;
      RECT 62.545 3.79 62.715 4.12 ;
      RECT 62.065 3.79 62.235 4.12 ;
      RECT 61.585 3.79 61.755 4.24 ;
      RECT 61.345 4.78 61.515 5.11 ;
      RECT 61.105 3.79 61.275 4.52 ;
      RECT 60.625 3.79 60.795 4.12 ;
      RECT 60.385 3.05 60.555 3.4 ;
      RECT 59.905 4.35 60.075 4.77 ;
      RECT 59.665 3.79 59.835 4.12 ;
      RECT 59.425 4.44 59.595 4.8 ;
      RECT 59.185 3.79 59.355 4.24 ;
      RECT 58.705 3.79 58.875 4.24 ;
      RECT 58.495 3.05 58.665 3.4 ;
      RECT 58.495 4.44 58.665 4.8 ;
      RECT 56.86 7.31 57.03 8.78 ;
      RECT 56.86 10.09 57.03 10.6 ;
      RECT 55.87 1.865 56.04 2.375 ;
      RECT 55.87 3.685 56.04 5.155 ;
      RECT 55.87 7.31 56.04 8.78 ;
      RECT 55.87 10.09 56.04 10.6 ;
      RECT 54.51 1.87 54.68 5.16 ;
      RECT 54.51 7.305 54.68 10.595 ;
      RECT 54.08 1.87 54.25 2.38 ;
      RECT 54.08 2.95 54.25 5.16 ;
      RECT 54.08 7.305 54.25 9.515 ;
      RECT 54.08 10.085 54.25 10.595 ;
      RECT 50.405 3.05 50.575 3.4 ;
      RECT 50.165 3.79 50.335 4.12 ;
      RECT 49.685 3.79 49.855 4.24 ;
      RECT 49.445 3.05 49.615 3.4 ;
      RECT 49.205 3.79 49.375 4.12 ;
      RECT 48.895 7.305 49.065 10.595 ;
      RECT 48.465 7.305 48.635 9.515 ;
      RECT 48.465 10.085 48.635 10.595 ;
      RECT 48.455 4.78 48.625 5.11 ;
      RECT 47.765 3.79 47.935 4.24 ;
      RECT 47.285 3.79 47.455 4.12 ;
      RECT 46.805 3.79 46.975 4.12 ;
      RECT 46.325 3.79 46.495 4.24 ;
      RECT 46.085 4.78 46.255 5.11 ;
      RECT 45.845 3.79 46.015 4.52 ;
      RECT 45.365 3.79 45.535 4.12 ;
      RECT 45.125 3.05 45.295 3.4 ;
      RECT 44.645 4.35 44.815 4.77 ;
      RECT 44.405 3.79 44.575 4.12 ;
      RECT 44.165 4.44 44.335 4.8 ;
      RECT 43.925 3.79 44.095 4.24 ;
      RECT 43.445 3.79 43.615 4.24 ;
      RECT 43.235 3.05 43.405 3.4 ;
      RECT 43.235 4.44 43.405 4.8 ;
      RECT 41.6 7.31 41.77 8.78 ;
      RECT 41.6 10.09 41.77 10.6 ;
      RECT 40.61 1.865 40.78 2.375 ;
      RECT 40.61 3.685 40.78 5.155 ;
      RECT 40.61 7.31 40.78 8.78 ;
      RECT 40.61 10.09 40.78 10.6 ;
      RECT 39.25 1.87 39.42 5.16 ;
      RECT 39.25 7.305 39.42 10.595 ;
      RECT 38.82 1.87 38.99 2.38 ;
      RECT 38.82 2.95 38.99 5.16 ;
      RECT 38.82 7.305 38.99 9.515 ;
      RECT 38.82 10.085 38.99 10.595 ;
      RECT 35.145 3.05 35.315 3.4 ;
      RECT 34.905 3.79 35.075 4.12 ;
      RECT 34.425 3.79 34.595 4.24 ;
      RECT 34.185 3.05 34.355 3.4 ;
      RECT 33.945 3.79 34.115 4.12 ;
      RECT 33.635 7.305 33.805 10.595 ;
      RECT 33.205 7.305 33.375 9.515 ;
      RECT 33.205 10.085 33.375 10.595 ;
      RECT 33.195 4.78 33.365 5.11 ;
      RECT 32.505 3.79 32.675 4.24 ;
      RECT 32.025 3.79 32.195 4.12 ;
      RECT 31.545 3.79 31.715 4.12 ;
      RECT 31.065 3.79 31.235 4.24 ;
      RECT 30.825 4.78 30.995 5.11 ;
      RECT 30.585 3.79 30.755 4.52 ;
      RECT 30.105 3.79 30.275 4.12 ;
      RECT 29.865 3.05 30.035 3.4 ;
      RECT 29.385 4.35 29.555 4.77 ;
      RECT 29.145 3.79 29.315 4.12 ;
      RECT 28.905 4.44 29.075 4.8 ;
      RECT 28.665 3.79 28.835 4.24 ;
      RECT 28.185 3.79 28.355 4.24 ;
      RECT 27.975 3.05 28.145 3.4 ;
      RECT 27.975 4.44 28.145 4.8 ;
      RECT 26.34 7.31 26.51 8.78 ;
      RECT 26.34 10.09 26.51 10.6 ;
      RECT 25.35 1.865 25.52 2.375 ;
      RECT 25.35 3.685 25.52 5.155 ;
      RECT 25.35 7.31 25.52 8.78 ;
      RECT 25.35 10.09 25.52 10.6 ;
      RECT 23.99 1.87 24.16 5.16 ;
      RECT 23.99 7.305 24.16 10.595 ;
      RECT 23.56 1.87 23.73 2.38 ;
      RECT 23.56 2.95 23.73 5.16 ;
      RECT 23.56 7.305 23.73 9.515 ;
      RECT 23.56 10.085 23.73 10.595 ;
      RECT 19.885 3.05 20.055 3.4 ;
      RECT 19.645 3.79 19.815 4.12 ;
      RECT 19.165 3.79 19.335 4.24 ;
      RECT 18.925 3.05 19.095 3.4 ;
      RECT 18.685 3.79 18.855 4.12 ;
      RECT 18.375 7.305 18.545 10.595 ;
      RECT 17.945 7.305 18.115 9.515 ;
      RECT 17.945 10.085 18.115 10.595 ;
      RECT 17.935 4.78 18.105 5.11 ;
      RECT 17.245 3.79 17.415 4.24 ;
      RECT 16.765 3.79 16.935 4.12 ;
      RECT 16.285 3.79 16.455 4.12 ;
      RECT 15.805 3.79 15.975 4.24 ;
      RECT 15.565 4.78 15.735 5.11 ;
      RECT 15.325 3.79 15.495 4.52 ;
      RECT 14.845 3.79 15.015 4.12 ;
      RECT 14.605 3.05 14.775 3.4 ;
      RECT 14.125 4.35 14.295 4.77 ;
      RECT 13.885 3.79 14.055 4.12 ;
      RECT 13.645 4.44 13.815 4.8 ;
      RECT 13.405 3.79 13.575 4.24 ;
      RECT 12.925 3.79 13.095 4.24 ;
      RECT 12.715 3.05 12.885 3.4 ;
      RECT 12.715 4.44 12.885 4.8 ;
      RECT 10.43 7.305 10.6 9.515 ;
      RECT 10.43 10.085 10.6 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r2 ;
  SIZE 79.1 BY 12.47 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 17.515 1.87 17.685 2.38 ;
        RECT 17.515 3.69 17.685 5.16 ;
      LAYER met1 ;
        RECT 17.455 3.66 17.745 3.89 ;
        RECT 17.455 2.18 17.745 2.41 ;
        RECT 17.515 2.18 17.685 3.89 ;
      LAYER mcon ;
        RECT 17.515 3.69 17.685 3.86 ;
        RECT 17.515 2.21 17.685 2.38 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 32.775 1.87 32.945 2.38 ;
        RECT 32.775 3.69 32.945 5.16 ;
      LAYER met1 ;
        RECT 32.715 3.66 33.005 3.89 ;
        RECT 32.715 2.18 33.005 2.41 ;
        RECT 32.775 2.18 32.945 3.89 ;
      LAYER mcon ;
        RECT 32.775 3.69 32.945 3.86 ;
        RECT 32.775 2.21 32.945 2.38 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 48.035 1.87 48.205 2.38 ;
        RECT 48.035 3.69 48.205 5.16 ;
      LAYER met1 ;
        RECT 47.975 3.66 48.265 3.89 ;
        RECT 47.975 2.18 48.265 2.41 ;
        RECT 48.035 2.18 48.205 3.89 ;
      LAYER mcon ;
        RECT 48.035 3.69 48.205 3.86 ;
        RECT 48.035 2.21 48.205 2.38 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 63.295 1.87 63.465 2.38 ;
        RECT 63.295 3.69 63.465 5.16 ;
      LAYER met1 ;
        RECT 63.235 3.66 63.525 3.89 ;
        RECT 63.235 2.18 63.525 2.41 ;
        RECT 63.295 2.18 63.465 3.89 ;
      LAYER mcon ;
        RECT 63.295 3.69 63.465 3.86 ;
        RECT 63.295 2.21 63.465 2.38 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 78.555 1.87 78.725 2.38 ;
        RECT 78.555 3.69 78.725 5.16 ;
      LAYER met1 ;
        RECT 78.495 3.66 78.785 3.89 ;
        RECT 78.495 2.18 78.785 2.41 ;
        RECT 78.555 2.18 78.725 3.89 ;
      LAYER mcon ;
        RECT 78.555 3.69 78.725 3.86 ;
        RECT 78.555 2.21 78.725 2.38 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 13.285 8.155 13.625 8.505 ;
        RECT 13.285 4.005 13.625 4.355 ;
        RECT 13.365 4.005 13.535 8.505 ;
      LAYER li1 ;
        RECT 13.365 2.96 13.535 4.235 ;
        RECT 13.365 8.24 13.535 9.515 ;
        RECT 7.75 8.24 7.92 9.515 ;
      LAYER met1 ;
        RECT 13.285 4.065 13.765 4.235 ;
        RECT 13.285 4.005 13.625 4.355 ;
        RECT 7.69 8.24 13.765 8.41 ;
        RECT 13.285 8.155 13.625 8.505 ;
        RECT 7.69 8.21 7.98 8.44 ;
      LAYER via1 ;
        RECT 13.385 8.255 13.535 8.405 ;
        RECT 13.385 4.105 13.535 4.255 ;
      LAYER mcon ;
        RECT 7.75 8.24 7.92 8.41 ;
        RECT 13.365 8.24 13.535 8.41 ;
        RECT 13.365 4.065 13.535 4.235 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 28.545 8.155 28.885 8.505 ;
        RECT 28.545 4.005 28.885 4.355 ;
        RECT 28.625 4.005 28.795 8.505 ;
      LAYER li1 ;
        RECT 28.625 2.96 28.795 4.235 ;
        RECT 28.625 8.24 28.795 9.515 ;
        RECT 23.01 8.24 23.18 9.515 ;
      LAYER met1 ;
        RECT 28.545 4.065 29.025 4.235 ;
        RECT 28.545 4.005 28.885 4.355 ;
        RECT 22.95 8.24 29.025 8.41 ;
        RECT 28.545 8.155 28.885 8.505 ;
        RECT 22.95 8.21 23.24 8.44 ;
      LAYER via1 ;
        RECT 28.645 8.255 28.795 8.405 ;
        RECT 28.645 4.105 28.795 4.255 ;
      LAYER mcon ;
        RECT 23.01 8.24 23.18 8.41 ;
        RECT 28.625 8.24 28.795 8.41 ;
        RECT 28.625 4.065 28.795 4.235 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 43.805 8.155 44.145 8.505 ;
        RECT 43.805 4.005 44.145 4.355 ;
        RECT 43.885 4.005 44.055 8.505 ;
      LAYER li1 ;
        RECT 43.885 2.96 44.055 4.235 ;
        RECT 43.885 8.24 44.055 9.515 ;
        RECT 38.27 8.24 38.44 9.515 ;
      LAYER met1 ;
        RECT 43.805 4.065 44.285 4.235 ;
        RECT 43.805 4.005 44.145 4.355 ;
        RECT 38.21 8.24 44.285 8.41 ;
        RECT 43.805 8.155 44.145 8.505 ;
        RECT 38.21 8.21 38.5 8.44 ;
      LAYER via1 ;
        RECT 43.905 8.255 44.055 8.405 ;
        RECT 43.905 4.105 44.055 4.255 ;
      LAYER mcon ;
        RECT 38.27 8.24 38.44 8.41 ;
        RECT 43.885 8.24 44.055 8.41 ;
        RECT 43.885 4.065 44.055 4.235 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 59.065 8.155 59.405 8.505 ;
        RECT 59.065 4.005 59.405 4.355 ;
        RECT 59.145 4.005 59.315 8.505 ;
      LAYER li1 ;
        RECT 59.145 2.96 59.315 4.235 ;
        RECT 59.145 8.24 59.315 9.515 ;
        RECT 53.53 8.24 53.7 9.515 ;
      LAYER met1 ;
        RECT 59.065 4.065 59.545 4.235 ;
        RECT 59.065 4.005 59.405 4.355 ;
        RECT 53.47 8.24 59.545 8.41 ;
        RECT 59.065 8.155 59.405 8.505 ;
        RECT 53.47 8.21 53.76 8.44 ;
      LAYER via1 ;
        RECT 59.165 8.255 59.315 8.405 ;
        RECT 59.165 4.105 59.315 4.255 ;
      LAYER mcon ;
        RECT 53.53 8.24 53.7 8.41 ;
        RECT 59.145 8.24 59.315 8.41 ;
        RECT 59.145 4.065 59.315 4.235 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 74.325 8.155 74.665 8.505 ;
        RECT 74.325 4.005 74.665 4.355 ;
        RECT 74.405 4.005 74.575 8.505 ;
      LAYER li1 ;
        RECT 74.405 2.96 74.575 4.235 ;
        RECT 74.405 8.24 74.575 9.515 ;
        RECT 68.79 8.24 68.96 9.515 ;
      LAYER met1 ;
        RECT 74.325 4.065 74.805 4.235 ;
        RECT 74.325 4.005 74.665 4.355 ;
        RECT 68.73 8.24 74.805 8.41 ;
        RECT 74.325 8.155 74.665 8.505 ;
        RECT 68.73 8.21 69.02 8.44 ;
      LAYER via1 ;
        RECT 74.425 8.255 74.575 8.405 ;
        RECT 74.425 4.105 74.575 4.255 ;
      LAYER mcon ;
        RECT 68.79 8.24 68.96 8.41 ;
        RECT 74.405 8.24 74.575 8.41 ;
        RECT 74.405 4.065 74.575 4.235 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.235 8.24 0.405 9.515 ;
      LAYER met1 ;
        RECT 0.175 8.24 0.635 8.41 ;
        RECT 0.175 8.21 0.465 8.44 ;
      LAYER mcon ;
        RECT 0.235 8.24 0.405 8.41 ;
    END
  END start
  OBS
    LAYER met4 ;
      RECT 66.74 4.275 67.07 4.605 ;
      RECT 66.755 3.8 67.07 4.605 ;
      RECT 68.9 3.785 69.23 4.14 ;
      RECT 66.755 3.8 69.23 4.1 ;
      RECT 51.48 4.275 51.81 4.605 ;
      RECT 51.495 3.8 51.81 4.605 ;
      RECT 53.64 3.785 53.97 4.14 ;
      RECT 51.495 3.8 53.97 4.1 ;
      RECT 36.22 4.275 36.55 4.605 ;
      RECT 36.235 3.8 36.55 4.605 ;
      RECT 38.38 3.785 38.71 4.14 ;
      RECT 36.235 3.8 38.71 4.1 ;
      RECT 20.96 4.275 21.29 4.605 ;
      RECT 20.975 3.8 21.29 4.605 ;
      RECT 23.12 3.785 23.45 4.14 ;
      RECT 20.975 3.8 23.45 4.1 ;
      RECT 5.7 4.275 6.03 4.605 ;
      RECT 5.715 3.8 6.03 4.605 ;
      RECT 7.86 3.785 8.19 4.14 ;
      RECT 5.715 3.8 8.19 4.1 ;
    LAYER via3 ;
      RECT 68.965 3.875 69.165 4.075 ;
      RECT 66.805 4.34 67.005 4.54 ;
      RECT 53.705 3.875 53.905 4.075 ;
      RECT 51.545 4.34 51.745 4.54 ;
      RECT 38.445 3.875 38.645 4.075 ;
      RECT 36.285 4.34 36.485 4.54 ;
      RECT 23.185 3.875 23.385 4.075 ;
      RECT 21.025 4.34 21.225 4.54 ;
      RECT 7.925 3.875 8.125 4.075 ;
      RECT 5.765 4.34 5.965 4.54 ;
    LAYER met3 ;
      RECT 73.765 2.405 74.105 4.365 ;
      RECT 68.025 3.18 68.755 3.51 ;
      RECT 68.175 2.405 68.475 3.51 ;
      RECT 68.175 2.405 74.105 2.705 ;
      RECT 70.06 9.35 70.43 9.72 ;
      RECT 70.095 5.775 70.395 9.72 ;
      RECT 68.655 5.775 70.395 7.07 ;
      RECT 65.86 5.555 68.955 6.85 ;
      RECT 68.655 3.815 68.955 7.07 ;
      RECT 65.86 4.275 66.16 6.85 ;
      RECT 69.38 4.81 69.71 5.165 ;
      RECT 67.475 4.85 69.71 5.15 ;
      RECT 67.475 3.715 67.775 5.15 ;
      RECT 65.555 4.275 66.285 4.605 ;
      RECT 68.45 3.82 69.23 4.165 ;
      RECT 68.925 3.785 69.23 4.165 ;
      RECT 67.46 3.715 67.79 4.045 ;
      RECT 66.745 3.715 67.065 4.63 ;
      RECT 66.745 3.715 67.075 4.25 ;
      RECT 58.505 2.405 58.845 4.365 ;
      RECT 52.765 3.18 53.495 3.51 ;
      RECT 52.915 2.405 53.215 3.51 ;
      RECT 52.915 2.405 58.845 2.705 ;
      RECT 54.8 9.35 55.17 9.72 ;
      RECT 54.835 5.775 55.135 9.72 ;
      RECT 53.395 5.775 55.135 7.07 ;
      RECT 50.6 5.555 53.695 6.85 ;
      RECT 53.395 3.815 53.695 7.07 ;
      RECT 50.6 4.275 50.9 6.85 ;
      RECT 54.12 4.81 54.45 5.165 ;
      RECT 52.215 4.85 54.45 5.15 ;
      RECT 52.215 3.715 52.515 5.15 ;
      RECT 50.295 4.275 51.025 4.605 ;
      RECT 53.19 3.82 53.97 4.165 ;
      RECT 53.665 3.785 53.97 4.165 ;
      RECT 52.2 3.715 52.53 4.045 ;
      RECT 51.485 3.715 51.805 4.63 ;
      RECT 51.485 3.715 51.815 4.25 ;
      RECT 43.245 2.405 43.585 4.365 ;
      RECT 37.505 3.18 38.235 3.51 ;
      RECT 37.655 2.405 37.955 3.51 ;
      RECT 37.655 2.405 43.585 2.705 ;
      RECT 39.54 9.35 39.91 9.72 ;
      RECT 39.575 5.775 39.875 9.72 ;
      RECT 38.135 5.775 39.875 7.07 ;
      RECT 35.34 5.555 38.435 6.85 ;
      RECT 38.135 3.815 38.435 7.07 ;
      RECT 35.34 4.275 35.64 6.85 ;
      RECT 38.86 4.81 39.19 5.165 ;
      RECT 36.955 4.85 39.19 5.15 ;
      RECT 36.955 3.715 37.255 5.15 ;
      RECT 35.035 4.275 35.765 4.605 ;
      RECT 37.93 3.82 38.71 4.165 ;
      RECT 38.405 3.785 38.71 4.165 ;
      RECT 36.94 3.715 37.27 4.045 ;
      RECT 36.225 3.715 36.545 4.63 ;
      RECT 36.225 3.715 36.555 4.25 ;
      RECT 27.985 2.405 28.325 4.365 ;
      RECT 22.245 3.18 22.975 3.51 ;
      RECT 22.395 2.405 22.695 3.51 ;
      RECT 22.395 2.405 28.325 2.705 ;
      RECT 24.28 9.35 24.65 9.72 ;
      RECT 24.315 5.775 24.615 9.72 ;
      RECT 22.875 5.775 24.615 7.07 ;
      RECT 20.08 5.555 23.175 6.85 ;
      RECT 22.875 3.815 23.175 7.07 ;
      RECT 20.08 4.275 20.38 6.85 ;
      RECT 23.6 4.81 23.93 5.165 ;
      RECT 21.695 4.85 23.93 5.15 ;
      RECT 21.695 3.715 21.995 5.15 ;
      RECT 19.775 4.275 20.505 4.605 ;
      RECT 22.67 3.82 23.45 4.165 ;
      RECT 23.145 3.785 23.45 4.165 ;
      RECT 21.68 3.715 22.01 4.045 ;
      RECT 20.965 3.715 21.285 4.63 ;
      RECT 20.965 3.715 21.295 4.25 ;
      RECT 12.725 2.405 13.065 4.365 ;
      RECT 6.985 3.18 7.715 3.51 ;
      RECT 7.135 2.405 7.435 3.51 ;
      RECT 7.135 2.405 13.065 2.705 ;
      RECT 9.02 9.35 9.39 9.72 ;
      RECT 9.055 5.775 9.355 9.72 ;
      RECT 7.615 5.775 9.355 7.07 ;
      RECT 4.82 5.555 7.915 6.85 ;
      RECT 7.615 3.815 7.915 7.07 ;
      RECT 4.82 4.275 5.12 6.85 ;
      RECT 8.34 4.81 8.67 5.165 ;
      RECT 6.435 4.85 8.67 5.15 ;
      RECT 6.435 3.715 6.735 5.15 ;
      RECT 4.515 4.275 5.245 4.605 ;
      RECT 7.41 3.82 8.19 4.165 ;
      RECT 7.885 3.785 8.19 4.165 ;
      RECT 6.42 3.715 6.75 4.045 ;
      RECT 5.705 3.715 6.025 4.63 ;
      RECT 5.705 3.715 6.035 4.25 ;
      RECT 72.3 3.155 73.03 3.485 ;
      RECT 70.61 3.17 71.34 3.5 ;
      RECT 69.575 3.155 70.305 3.505 ;
      RECT 65.42 3.155 66.15 3.485 ;
      RECT 57.04 3.155 57.77 3.485 ;
      RECT 55.35 3.17 56.08 3.5 ;
      RECT 54.315 3.155 55.045 3.505 ;
      RECT 50.16 3.155 50.89 3.485 ;
      RECT 41.78 3.155 42.51 3.485 ;
      RECT 40.09 3.17 40.82 3.5 ;
      RECT 39.055 3.155 39.785 3.505 ;
      RECT 34.9 3.155 35.63 3.485 ;
      RECT 26.52 3.155 27.25 3.485 ;
      RECT 24.83 3.17 25.56 3.5 ;
      RECT 23.795 3.155 24.525 3.505 ;
      RECT 19.64 3.155 20.37 3.485 ;
      RECT 11.26 3.155 11.99 3.485 ;
      RECT 9.57 3.17 10.3 3.5 ;
      RECT 8.535 3.155 9.265 3.505 ;
      RECT 4.38 3.155 5.11 3.485 ;
      RECT 0.01 10.795 0.815 11.175 ;
      RECT 0.005 0.005 0.81 0.385 ;
    LAYER via2 ;
      RECT 73.84 4.075 74.04 4.275 ;
      RECT 72.535 3.22 72.735 3.42 ;
      RECT 70.675 3.235 70.875 3.435 ;
      RECT 70.145 9.435 70.345 9.635 ;
      RECT 69.655 3.24 69.855 3.44 ;
      RECT 69.445 4.875 69.645 5.075 ;
      RECT 68.965 3.875 69.165 4.075 ;
      RECT 68.215 3.245 68.415 3.445 ;
      RECT 67.525 3.78 67.725 3.98 ;
      RECT 66.81 3.78 67.01 3.98 ;
      RECT 65.845 4.34 66.045 4.54 ;
      RECT 65.605 3.22 65.805 3.42 ;
      RECT 58.58 4.075 58.78 4.275 ;
      RECT 57.275 3.22 57.475 3.42 ;
      RECT 55.415 3.235 55.615 3.435 ;
      RECT 54.885 9.435 55.085 9.635 ;
      RECT 54.395 3.24 54.595 3.44 ;
      RECT 54.185 4.875 54.385 5.075 ;
      RECT 53.705 3.875 53.905 4.075 ;
      RECT 52.955 3.245 53.155 3.445 ;
      RECT 52.265 3.78 52.465 3.98 ;
      RECT 51.55 3.78 51.75 3.98 ;
      RECT 50.585 4.34 50.785 4.54 ;
      RECT 50.345 3.22 50.545 3.42 ;
      RECT 43.32 4.075 43.52 4.275 ;
      RECT 42.015 3.22 42.215 3.42 ;
      RECT 40.155 3.235 40.355 3.435 ;
      RECT 39.625 9.435 39.825 9.635 ;
      RECT 39.135 3.24 39.335 3.44 ;
      RECT 38.925 4.875 39.125 5.075 ;
      RECT 38.445 3.875 38.645 4.075 ;
      RECT 37.695 3.245 37.895 3.445 ;
      RECT 37.005 3.78 37.205 3.98 ;
      RECT 36.29 3.78 36.49 3.98 ;
      RECT 35.325 4.34 35.525 4.54 ;
      RECT 35.085 3.22 35.285 3.42 ;
      RECT 28.06 4.075 28.26 4.275 ;
      RECT 26.755 3.22 26.955 3.42 ;
      RECT 24.895 3.235 25.095 3.435 ;
      RECT 24.365 9.435 24.565 9.635 ;
      RECT 23.875 3.24 24.075 3.44 ;
      RECT 23.665 4.875 23.865 5.075 ;
      RECT 23.185 3.875 23.385 4.075 ;
      RECT 22.435 3.245 22.635 3.445 ;
      RECT 21.745 3.78 21.945 3.98 ;
      RECT 21.03 3.78 21.23 3.98 ;
      RECT 20.065 4.34 20.265 4.54 ;
      RECT 19.825 3.22 20.025 3.42 ;
      RECT 12.8 4.075 13 4.275 ;
      RECT 11.495 3.22 11.695 3.42 ;
      RECT 9.635 3.235 9.835 3.435 ;
      RECT 9.105 9.435 9.305 9.635 ;
      RECT 8.615 3.24 8.815 3.44 ;
      RECT 8.405 4.875 8.605 5.075 ;
      RECT 7.925 3.875 8.125 4.075 ;
      RECT 7.175 3.245 7.375 3.445 ;
      RECT 6.485 3.78 6.685 3.98 ;
      RECT 5.77 3.78 5.97 3.98 ;
      RECT 4.805 4.34 5.005 4.54 ;
      RECT 4.565 3.22 4.765 3.42 ;
      RECT 0.29 10.885 0.49 11.085 ;
      RECT 0.285 0.095 0.485 0.295 ;
    LAYER met2 ;
      RECT 1.235 10.695 78.73 10.865 ;
      RECT 78.56 9.57 78.73 10.865 ;
      RECT 1.235 8.55 1.405 10.865 ;
      RECT 78.53 9.57 78.88 9.92 ;
      RECT 1.17 8.55 1.46 8.9 ;
      RECT 75.37 8.515 75.69 8.84 ;
      RECT 75.4 7.99 75.57 8.84 ;
      RECT 75.4 7.99 75.575 8.34 ;
      RECT 75.4 7.99 76.375 8.165 ;
      RECT 76.2 3.265 76.375 8.165 ;
      RECT 76.145 3.265 76.495 3.615 ;
      RECT 76.17 8.95 76.495 9.275 ;
      RECT 75.055 9.04 76.495 9.21 ;
      RECT 75.055 3.695 75.215 9.21 ;
      RECT 75.37 3.665 75.69 3.985 ;
      RECT 75.055 3.695 75.69 3.865 ;
      RECT 73.795 3.985 74.085 4.365 ;
      RECT 73.765 4 74.105 4.35 ;
      RECT 72.505 4.84 72.765 5.16 ;
      RECT 72.565 3.135 72.705 5.16 ;
      RECT 72.39 3.695 72.705 4.065 ;
      RECT 72.46 3.25 72.705 4.065 ;
      RECT 72.495 3.135 72.775 3.505 ;
      RECT 71.815 3.72 72.075 4.04 ;
      RECT 71.155 3.81 72.075 3.95 ;
      RECT 71.155 2.87 71.295 3.95 ;
      RECT 67.615 3.16 67.875 3.48 ;
      RECT 67.795 2.87 67.935 3.39 ;
      RECT 67.795 2.87 71.295 3.01 ;
      RECT 63.245 8.95 63.595 9.3 ;
      RECT 70.73 8.905 71.08 9.255 ;
      RECT 63.245 8.98 71.08 9.18 ;
      RECT 70.645 4.56 70.905 4.88 ;
      RECT 70.705 3.15 70.845 4.88 ;
      RECT 70.635 3.15 70.915 3.52 ;
      RECT 68.035 5.31 70.47 5.45 ;
      RECT 70.33 4 70.47 5.45 ;
      RECT 68.035 4.93 68.175 5.45 ;
      RECT 67.735 4.93 68.175 5.16 ;
      RECT 65.395 4.93 68.175 5.07 ;
      RECT 67.735 4.84 67.995 5.16 ;
      RECT 65.395 4.65 65.535 5.07 ;
      RECT 64.885 4.56 65.145 4.88 ;
      RECT 64.885 4.65 65.535 4.79 ;
      RECT 64.945 3.16 65.085 4.88 ;
      RECT 70.27 4 70.53 4.32 ;
      RECT 64.885 3.16 65.145 3.48 ;
      RECT 69.895 4.84 70.155 5.16 ;
      RECT 69.955 3.25 70.095 5.16 ;
      RECT 69.615 3.25 70.095 3.525 ;
      RECT 69.415 3.155 69.895 3.5 ;
      RECT 69.405 4.79 69.685 5.16 ;
      RECT 69.475 3.695 69.615 5.16 ;
      RECT 69.415 3.695 69.675 4.32 ;
      RECT 69.405 3.695 69.685 4.065 ;
      RECT 68.335 4.84 68.595 5.16 ;
      RECT 68.335 4.65 68.535 5.16 ;
      RECT 68.14 4.65 68.535 4.79 ;
      RECT 68.14 3.16 68.28 4.79 ;
      RECT 68.14 3.16 68.455 3.53 ;
      RECT 68.08 3.16 68.455 3.48 ;
      RECT 65.805 4.255 66.085 4.625 ;
      RECT 67.255 4.28 67.515 4.6 ;
      RECT 65.635 4.37 67.515 4.51 ;
      RECT 65.635 4.255 66.085 4.51 ;
      RECT 65.575 3.695 65.835 4.32 ;
      RECT 65.565 3.695 65.845 4.065 ;
      RECT 66.645 3.695 67.055 4.065 ;
      RECT 66.055 3.72 66.315 4.04 ;
      RECT 66.055 3.81 67.055 3.95 ;
      RECT 65.565 3.135 65.845 3.505 ;
      RECT 65.565 3.16 65.955 3.48 ;
      RECT 60.11 8.515 60.43 8.84 ;
      RECT 60.14 7.99 60.31 8.84 ;
      RECT 60.14 7.99 60.315 8.34 ;
      RECT 60.14 7.99 61.115 8.165 ;
      RECT 60.94 3.265 61.115 8.165 ;
      RECT 60.885 3.265 61.235 3.615 ;
      RECT 60.91 8.95 61.235 9.275 ;
      RECT 59.795 9.04 61.235 9.21 ;
      RECT 59.795 3.695 59.955 9.21 ;
      RECT 60.11 3.665 60.43 3.985 ;
      RECT 59.795 3.695 60.43 3.865 ;
      RECT 58.535 3.985 58.825 4.365 ;
      RECT 58.505 4 58.845 4.35 ;
      RECT 57.245 4.84 57.505 5.16 ;
      RECT 57.305 3.135 57.445 5.16 ;
      RECT 57.13 3.695 57.445 4.065 ;
      RECT 57.2 3.25 57.445 4.065 ;
      RECT 57.235 3.135 57.515 3.505 ;
      RECT 56.555 3.72 56.815 4.04 ;
      RECT 55.895 3.81 56.815 3.95 ;
      RECT 55.895 2.87 56.035 3.95 ;
      RECT 52.355 3.16 52.615 3.48 ;
      RECT 52.535 2.87 52.675 3.39 ;
      RECT 52.535 2.87 56.035 3.01 ;
      RECT 47.985 8.95 48.335 9.3 ;
      RECT 55.475 8.905 55.825 9.255 ;
      RECT 47.985 8.98 55.825 9.18 ;
      RECT 55.385 4.56 55.645 4.88 ;
      RECT 55.445 3.15 55.585 4.88 ;
      RECT 55.375 3.15 55.655 3.52 ;
      RECT 52.775 5.31 55.21 5.45 ;
      RECT 55.07 4 55.21 5.45 ;
      RECT 52.775 4.93 52.915 5.45 ;
      RECT 52.475 4.93 52.915 5.16 ;
      RECT 50.135 4.93 52.915 5.07 ;
      RECT 52.475 4.84 52.735 5.16 ;
      RECT 50.135 4.65 50.275 5.07 ;
      RECT 49.625 4.56 49.885 4.88 ;
      RECT 49.625 4.65 50.275 4.79 ;
      RECT 49.685 3.16 49.825 4.88 ;
      RECT 55.01 4 55.27 4.32 ;
      RECT 49.625 3.16 49.885 3.48 ;
      RECT 54.635 4.84 54.895 5.16 ;
      RECT 54.695 3.25 54.835 5.16 ;
      RECT 54.355 3.25 54.835 3.525 ;
      RECT 54.155 3.155 54.635 3.5 ;
      RECT 54.145 4.79 54.425 5.16 ;
      RECT 54.215 3.695 54.355 5.16 ;
      RECT 54.155 3.695 54.415 4.32 ;
      RECT 54.145 3.695 54.425 4.065 ;
      RECT 53.075 4.84 53.335 5.16 ;
      RECT 53.075 4.65 53.275 5.16 ;
      RECT 52.88 4.65 53.275 4.79 ;
      RECT 52.88 3.16 53.02 4.79 ;
      RECT 52.88 3.16 53.195 3.53 ;
      RECT 52.82 3.16 53.195 3.48 ;
      RECT 50.545 4.255 50.825 4.625 ;
      RECT 51.995 4.28 52.255 4.6 ;
      RECT 50.375 4.37 52.255 4.51 ;
      RECT 50.375 4.255 50.825 4.51 ;
      RECT 50.315 3.695 50.575 4.32 ;
      RECT 50.305 3.695 50.585 4.065 ;
      RECT 51.385 3.695 51.795 4.065 ;
      RECT 50.795 3.72 51.055 4.04 ;
      RECT 50.795 3.81 51.795 3.95 ;
      RECT 50.305 3.135 50.585 3.505 ;
      RECT 50.305 3.16 50.695 3.48 ;
      RECT 44.85 8.515 45.17 8.84 ;
      RECT 44.88 7.99 45.05 8.84 ;
      RECT 44.88 7.99 45.055 8.34 ;
      RECT 44.88 7.99 45.855 8.165 ;
      RECT 45.68 3.265 45.855 8.165 ;
      RECT 45.625 3.265 45.975 3.615 ;
      RECT 45.65 8.95 45.975 9.275 ;
      RECT 44.535 9.04 45.975 9.21 ;
      RECT 44.535 3.695 44.695 9.21 ;
      RECT 44.85 3.665 45.17 3.985 ;
      RECT 44.535 3.695 45.17 3.865 ;
      RECT 43.275 3.985 43.565 4.365 ;
      RECT 43.245 4 43.585 4.35 ;
      RECT 41.985 4.84 42.245 5.16 ;
      RECT 42.045 3.135 42.185 5.16 ;
      RECT 41.87 3.695 42.185 4.065 ;
      RECT 41.94 3.25 42.185 4.065 ;
      RECT 41.975 3.135 42.255 3.505 ;
      RECT 41.295 3.72 41.555 4.04 ;
      RECT 40.635 3.81 41.555 3.95 ;
      RECT 40.635 2.87 40.775 3.95 ;
      RECT 37.095 3.16 37.355 3.48 ;
      RECT 37.275 2.87 37.415 3.39 ;
      RECT 37.275 2.87 40.775 3.01 ;
      RECT 32.77 8.955 33.12 9.305 ;
      RECT 40.21 8.91 40.56 9.26 ;
      RECT 32.77 8.985 40.56 9.185 ;
      RECT 40.125 4.56 40.385 4.88 ;
      RECT 40.185 3.15 40.325 4.88 ;
      RECT 40.115 3.15 40.395 3.52 ;
      RECT 37.515 5.31 39.95 5.45 ;
      RECT 39.81 4 39.95 5.45 ;
      RECT 37.515 4.93 37.655 5.45 ;
      RECT 37.215 4.93 37.655 5.16 ;
      RECT 34.875 4.93 37.655 5.07 ;
      RECT 37.215 4.84 37.475 5.16 ;
      RECT 34.875 4.65 35.015 5.07 ;
      RECT 34.365 4.56 34.625 4.88 ;
      RECT 34.365 4.65 35.015 4.79 ;
      RECT 34.425 3.16 34.565 4.88 ;
      RECT 39.75 4 40.01 4.32 ;
      RECT 34.365 3.16 34.625 3.48 ;
      RECT 39.375 4.84 39.635 5.16 ;
      RECT 39.435 3.25 39.575 5.16 ;
      RECT 39.095 3.25 39.575 3.525 ;
      RECT 38.895 3.155 39.375 3.5 ;
      RECT 38.885 4.79 39.165 5.16 ;
      RECT 38.955 3.695 39.095 5.16 ;
      RECT 38.895 3.695 39.155 4.32 ;
      RECT 38.885 3.695 39.165 4.065 ;
      RECT 37.815 4.84 38.075 5.16 ;
      RECT 37.815 4.65 38.015 5.16 ;
      RECT 37.62 4.65 38.015 4.79 ;
      RECT 37.62 3.16 37.76 4.79 ;
      RECT 37.62 3.16 37.935 3.53 ;
      RECT 37.56 3.16 37.935 3.48 ;
      RECT 35.285 4.255 35.565 4.625 ;
      RECT 36.735 4.28 36.995 4.6 ;
      RECT 35.115 4.37 36.995 4.51 ;
      RECT 35.115 4.255 35.565 4.51 ;
      RECT 35.055 3.695 35.315 4.32 ;
      RECT 35.045 3.695 35.325 4.065 ;
      RECT 36.125 3.695 36.535 4.065 ;
      RECT 35.535 3.72 35.795 4.04 ;
      RECT 35.535 3.81 36.535 3.95 ;
      RECT 35.045 3.135 35.325 3.505 ;
      RECT 35.045 3.16 35.435 3.48 ;
      RECT 29.59 8.515 29.91 8.84 ;
      RECT 29.62 7.99 29.79 8.84 ;
      RECT 29.62 7.99 29.795 8.34 ;
      RECT 29.62 7.99 30.595 8.165 ;
      RECT 30.42 3.265 30.595 8.165 ;
      RECT 30.365 3.265 30.715 3.615 ;
      RECT 30.39 8.95 30.715 9.275 ;
      RECT 29.275 9.04 30.715 9.21 ;
      RECT 29.275 3.695 29.435 9.21 ;
      RECT 29.59 3.665 29.91 3.985 ;
      RECT 29.275 3.695 29.91 3.865 ;
      RECT 28.015 3.985 28.305 4.365 ;
      RECT 27.985 4 28.325 4.35 ;
      RECT 26.725 4.84 26.985 5.16 ;
      RECT 26.785 3.135 26.925 5.16 ;
      RECT 26.61 3.695 26.925 4.065 ;
      RECT 26.68 3.25 26.925 4.065 ;
      RECT 26.715 3.135 26.995 3.505 ;
      RECT 26.035 3.72 26.295 4.04 ;
      RECT 25.375 3.81 26.295 3.95 ;
      RECT 25.375 2.87 25.515 3.95 ;
      RECT 21.835 3.16 22.095 3.48 ;
      RECT 22.015 2.87 22.155 3.39 ;
      RECT 22.015 2.87 25.515 3.01 ;
      RECT 17.51 8.95 17.86 9.3 ;
      RECT 24.95 8.905 25.3 9.255 ;
      RECT 17.51 8.98 25.3 9.18 ;
      RECT 24.865 4.56 25.125 4.88 ;
      RECT 24.925 3.15 25.065 4.88 ;
      RECT 24.855 3.15 25.135 3.52 ;
      RECT 22.255 5.31 24.69 5.45 ;
      RECT 24.55 4 24.69 5.45 ;
      RECT 22.255 4.93 22.395 5.45 ;
      RECT 21.955 4.93 22.395 5.16 ;
      RECT 19.615 4.93 22.395 5.07 ;
      RECT 21.955 4.84 22.215 5.16 ;
      RECT 19.615 4.65 19.755 5.07 ;
      RECT 19.105 4.56 19.365 4.88 ;
      RECT 19.105 4.65 19.755 4.79 ;
      RECT 19.165 3.16 19.305 4.88 ;
      RECT 24.49 4 24.75 4.32 ;
      RECT 19.105 3.16 19.365 3.48 ;
      RECT 24.115 4.84 24.375 5.16 ;
      RECT 24.175 3.25 24.315 5.16 ;
      RECT 23.835 3.25 24.315 3.525 ;
      RECT 23.635 3.155 24.115 3.5 ;
      RECT 23.625 4.79 23.905 5.16 ;
      RECT 23.695 3.695 23.835 5.16 ;
      RECT 23.635 3.695 23.895 4.32 ;
      RECT 23.625 3.695 23.905 4.065 ;
      RECT 22.555 4.84 22.815 5.16 ;
      RECT 22.555 4.65 22.755 5.16 ;
      RECT 22.36 4.65 22.755 4.79 ;
      RECT 22.36 3.16 22.5 4.79 ;
      RECT 22.36 3.16 22.675 3.53 ;
      RECT 22.3 3.16 22.675 3.48 ;
      RECT 20.025 4.255 20.305 4.625 ;
      RECT 21.475 4.28 21.735 4.6 ;
      RECT 19.855 4.37 21.735 4.51 ;
      RECT 19.855 4.255 20.305 4.51 ;
      RECT 19.795 3.695 20.055 4.32 ;
      RECT 19.785 3.695 20.065 4.065 ;
      RECT 20.865 3.695 21.275 4.065 ;
      RECT 20.275 3.72 20.535 4.04 ;
      RECT 20.275 3.81 21.275 3.95 ;
      RECT 19.785 3.135 20.065 3.505 ;
      RECT 19.785 3.16 20.175 3.48 ;
      RECT 14.33 8.515 14.65 8.84 ;
      RECT 14.36 7.99 14.53 8.84 ;
      RECT 14.36 7.99 14.535 8.34 ;
      RECT 14.36 7.99 15.335 8.165 ;
      RECT 15.16 3.265 15.335 8.165 ;
      RECT 15.105 3.265 15.455 3.615 ;
      RECT 15.13 8.95 15.455 9.275 ;
      RECT 14.015 9.04 15.455 9.21 ;
      RECT 14.015 3.695 14.175 9.21 ;
      RECT 14.33 3.665 14.65 3.985 ;
      RECT 14.015 3.695 14.65 3.865 ;
      RECT 12.755 3.985 13.045 4.365 ;
      RECT 12.725 4 13.065 4.35 ;
      RECT 11.465 4.84 11.725 5.16 ;
      RECT 11.525 3.135 11.665 5.16 ;
      RECT 11.35 3.695 11.665 4.065 ;
      RECT 11.42 3.25 11.665 4.065 ;
      RECT 11.455 3.135 11.735 3.505 ;
      RECT 10.775 3.72 11.035 4.04 ;
      RECT 10.115 3.81 11.035 3.95 ;
      RECT 10.115 2.87 10.255 3.95 ;
      RECT 6.575 3.16 6.835 3.48 ;
      RECT 6.755 2.87 6.895 3.39 ;
      RECT 6.755 2.87 10.255 3.01 ;
      RECT 1.545 9.29 1.835 9.64 ;
      RECT 1.545 9.345 2.8 9.515 ;
      RECT 2.63 8.98 2.8 9.515 ;
      RECT 9.69 8.9 10.04 9.25 ;
      RECT 2.63 8.98 10.04 9.15 ;
      RECT 9.605 4.56 9.865 4.88 ;
      RECT 9.665 3.15 9.805 4.88 ;
      RECT 9.595 3.15 9.875 3.52 ;
      RECT 6.995 5.31 9.43 5.45 ;
      RECT 9.29 4 9.43 5.45 ;
      RECT 6.995 4.93 7.135 5.45 ;
      RECT 6.695 4.93 7.135 5.16 ;
      RECT 4.355 4.93 7.135 5.07 ;
      RECT 6.695 4.84 6.955 5.16 ;
      RECT 4.355 4.65 4.495 5.07 ;
      RECT 3.845 4.56 4.105 4.88 ;
      RECT 3.845 4.65 4.495 4.79 ;
      RECT 3.905 3.16 4.045 4.88 ;
      RECT 9.23 4 9.49 4.32 ;
      RECT 3.845 3.16 4.105 3.48 ;
      RECT 8.855 4.84 9.115 5.16 ;
      RECT 8.915 3.25 9.055 5.16 ;
      RECT 8.575 3.25 9.055 3.525 ;
      RECT 8.375 3.155 8.855 3.5 ;
      RECT 8.365 4.79 8.645 5.16 ;
      RECT 8.435 3.695 8.575 5.16 ;
      RECT 8.375 3.695 8.635 4.32 ;
      RECT 8.365 3.695 8.645 4.065 ;
      RECT 7.295 4.84 7.555 5.16 ;
      RECT 7.295 4.65 7.495 5.16 ;
      RECT 7.1 4.65 7.495 4.79 ;
      RECT 7.1 3.16 7.24 4.79 ;
      RECT 7.1 3.16 7.415 3.53 ;
      RECT 7.04 3.16 7.415 3.48 ;
      RECT 4.765 4.255 5.045 4.625 ;
      RECT 6.215 4.28 6.475 4.6 ;
      RECT 4.595 4.37 6.475 4.51 ;
      RECT 4.595 4.255 5.045 4.51 ;
      RECT 4.535 3.695 4.795 4.32 ;
      RECT 4.525 3.695 4.805 4.065 ;
      RECT 5.605 3.695 6.015 4.065 ;
      RECT 5.015 3.72 5.275 4.04 ;
      RECT 5.015 3.81 6.015 3.95 ;
      RECT 4.525 3.135 4.805 3.505 ;
      RECT 4.525 3.16 4.915 3.48 ;
      RECT 0.2 10.795 0.58 11.175 ;
      RECT 0.24 0.005 0.405 11.175 ;
      RECT 0.195 0.005 0.575 0.385 ;
      RECT 70.06 9.35 70.43 9.72 ;
      RECT 68.925 3.695 69.205 4.16 ;
      RECT 68.685 3.16 68.965 3.505 ;
      RECT 67.485 3.695 67.765 4.065 ;
      RECT 64.925 2.515 65.295 2.52 ;
      RECT 54.8 9.35 55.17 9.72 ;
      RECT 53.665 3.695 53.945 4.16 ;
      RECT 53.425 3.16 53.705 3.505 ;
      RECT 52.225 3.695 52.505 4.065 ;
      RECT 49.665 2.515 50.035 2.52 ;
      RECT 39.54 9.35 39.91 9.72 ;
      RECT 38.405 3.695 38.685 4.16 ;
      RECT 38.165 3.16 38.445 3.505 ;
      RECT 36.965 3.695 37.245 4.065 ;
      RECT 34.405 2.515 34.775 2.52 ;
      RECT 24.28 9.35 24.65 9.72 ;
      RECT 23.145 3.695 23.425 4.16 ;
      RECT 22.905 3.16 23.185 3.505 ;
      RECT 21.705 3.695 21.985 4.065 ;
      RECT 19.145 2.515 19.515 2.52 ;
      RECT 9.02 9.35 9.39 9.72 ;
      RECT 7.885 3.695 8.165 4.16 ;
      RECT 7.645 3.16 7.925 3.505 ;
      RECT 6.445 3.695 6.725 4.065 ;
      RECT 3.885 2.515 4.255 2.52 ;
    LAYER via1 ;
      RECT 78.63 9.67 78.78 9.82 ;
      RECT 76.26 9.035 76.41 9.185 ;
      RECT 76.245 3.365 76.395 3.515 ;
      RECT 75.455 3.75 75.605 3.9 ;
      RECT 75.455 8.62 75.605 8.77 ;
      RECT 73.865 4.1 74.015 4.25 ;
      RECT 72.56 3.245 72.71 3.395 ;
      RECT 72.56 4.925 72.71 5.075 ;
      RECT 71.87 3.805 72.02 3.955 ;
      RECT 70.83 9.005 70.98 9.155 ;
      RECT 70.7 3.245 70.85 3.395 ;
      RECT 70.7 4.645 70.85 4.795 ;
      RECT 70.325 4.085 70.475 4.235 ;
      RECT 70.17 9.46 70.32 9.61 ;
      RECT 69.95 4.925 70.1 5.075 ;
      RECT 69.47 3.245 69.62 3.395 ;
      RECT 69.47 4.085 69.62 4.235 ;
      RECT 68.99 3.805 69.14 3.955 ;
      RECT 68.75 3.245 68.9 3.395 ;
      RECT 68.39 4.925 68.54 5.075 ;
      RECT 68.135 3.245 68.285 3.395 ;
      RECT 67.79 4.925 67.94 5.075 ;
      RECT 67.67 3.245 67.82 3.395 ;
      RECT 67.55 3.805 67.7 3.955 ;
      RECT 67.31 4.365 67.46 4.515 ;
      RECT 66.11 3.805 66.26 3.955 ;
      RECT 65.75 3.245 65.9 3.395 ;
      RECT 65.63 4.085 65.78 4.235 ;
      RECT 64.94 3.245 65.09 3.395 ;
      RECT 64.94 4.645 65.09 4.795 ;
      RECT 63.345 9.05 63.495 9.2 ;
      RECT 61 9.035 61.15 9.185 ;
      RECT 60.985 3.365 61.135 3.515 ;
      RECT 60.195 3.75 60.345 3.9 ;
      RECT 60.195 8.62 60.345 8.77 ;
      RECT 58.605 4.1 58.755 4.25 ;
      RECT 57.3 3.245 57.45 3.395 ;
      RECT 57.3 4.925 57.45 5.075 ;
      RECT 56.61 3.805 56.76 3.955 ;
      RECT 55.575 9.005 55.725 9.155 ;
      RECT 55.44 3.245 55.59 3.395 ;
      RECT 55.44 4.645 55.59 4.795 ;
      RECT 55.065 4.085 55.215 4.235 ;
      RECT 54.91 9.46 55.06 9.61 ;
      RECT 54.69 4.925 54.84 5.075 ;
      RECT 54.21 3.245 54.36 3.395 ;
      RECT 54.21 4.085 54.36 4.235 ;
      RECT 53.73 3.805 53.88 3.955 ;
      RECT 53.49 3.245 53.64 3.395 ;
      RECT 53.13 4.925 53.28 5.075 ;
      RECT 52.875 3.245 53.025 3.395 ;
      RECT 52.53 4.925 52.68 5.075 ;
      RECT 52.41 3.245 52.56 3.395 ;
      RECT 52.29 3.805 52.44 3.955 ;
      RECT 52.05 4.365 52.2 4.515 ;
      RECT 50.85 3.805 51 3.955 ;
      RECT 50.49 3.245 50.64 3.395 ;
      RECT 50.37 4.085 50.52 4.235 ;
      RECT 49.68 3.245 49.83 3.395 ;
      RECT 49.68 4.645 49.83 4.795 ;
      RECT 48.085 9.05 48.235 9.2 ;
      RECT 45.74 9.035 45.89 9.185 ;
      RECT 45.725 3.365 45.875 3.515 ;
      RECT 44.935 3.75 45.085 3.9 ;
      RECT 44.935 8.62 45.085 8.77 ;
      RECT 43.345 4.1 43.495 4.25 ;
      RECT 42.04 3.245 42.19 3.395 ;
      RECT 42.04 4.925 42.19 5.075 ;
      RECT 41.35 3.805 41.5 3.955 ;
      RECT 40.31 9.01 40.46 9.16 ;
      RECT 40.18 3.245 40.33 3.395 ;
      RECT 40.18 4.645 40.33 4.795 ;
      RECT 39.805 4.085 39.955 4.235 ;
      RECT 39.65 9.46 39.8 9.61 ;
      RECT 39.43 4.925 39.58 5.075 ;
      RECT 38.95 3.245 39.1 3.395 ;
      RECT 38.95 4.085 39.1 4.235 ;
      RECT 38.47 3.805 38.62 3.955 ;
      RECT 38.23 3.245 38.38 3.395 ;
      RECT 37.87 4.925 38.02 5.075 ;
      RECT 37.615 3.245 37.765 3.395 ;
      RECT 37.27 4.925 37.42 5.075 ;
      RECT 37.15 3.245 37.3 3.395 ;
      RECT 37.03 3.805 37.18 3.955 ;
      RECT 36.79 4.365 36.94 4.515 ;
      RECT 35.59 3.805 35.74 3.955 ;
      RECT 35.23 3.245 35.38 3.395 ;
      RECT 35.11 4.085 35.26 4.235 ;
      RECT 34.42 3.245 34.57 3.395 ;
      RECT 34.42 4.645 34.57 4.795 ;
      RECT 32.87 9.055 33.02 9.205 ;
      RECT 30.48 9.035 30.63 9.185 ;
      RECT 30.465 3.365 30.615 3.515 ;
      RECT 29.675 3.75 29.825 3.9 ;
      RECT 29.675 8.62 29.825 8.77 ;
      RECT 28.085 4.1 28.235 4.25 ;
      RECT 26.78 3.245 26.93 3.395 ;
      RECT 26.78 4.925 26.93 5.075 ;
      RECT 26.09 3.805 26.24 3.955 ;
      RECT 25.05 9.005 25.2 9.155 ;
      RECT 24.92 3.245 25.07 3.395 ;
      RECT 24.92 4.645 25.07 4.795 ;
      RECT 24.545 4.085 24.695 4.235 ;
      RECT 24.39 9.46 24.54 9.61 ;
      RECT 24.17 4.925 24.32 5.075 ;
      RECT 23.69 3.245 23.84 3.395 ;
      RECT 23.69 4.085 23.84 4.235 ;
      RECT 23.21 3.805 23.36 3.955 ;
      RECT 22.97 3.245 23.12 3.395 ;
      RECT 22.61 4.925 22.76 5.075 ;
      RECT 22.355 3.245 22.505 3.395 ;
      RECT 22.01 4.925 22.16 5.075 ;
      RECT 21.89 3.245 22.04 3.395 ;
      RECT 21.77 3.805 21.92 3.955 ;
      RECT 21.53 4.365 21.68 4.515 ;
      RECT 20.33 3.805 20.48 3.955 ;
      RECT 19.97 3.245 20.12 3.395 ;
      RECT 19.85 4.085 20 4.235 ;
      RECT 19.16 3.245 19.31 3.395 ;
      RECT 19.16 4.645 19.31 4.795 ;
      RECT 17.61 9.05 17.76 9.2 ;
      RECT 15.22 9.035 15.37 9.185 ;
      RECT 15.205 3.365 15.355 3.515 ;
      RECT 14.415 3.75 14.565 3.9 ;
      RECT 14.415 8.62 14.565 8.77 ;
      RECT 12.825 4.1 12.975 4.25 ;
      RECT 11.52 3.245 11.67 3.395 ;
      RECT 11.52 4.925 11.67 5.075 ;
      RECT 10.83 3.805 10.98 3.955 ;
      RECT 9.79 9 9.94 9.15 ;
      RECT 9.66 3.245 9.81 3.395 ;
      RECT 9.66 4.645 9.81 4.795 ;
      RECT 9.285 4.085 9.435 4.235 ;
      RECT 9.13 9.46 9.28 9.61 ;
      RECT 8.91 4.925 9.06 5.075 ;
      RECT 8.43 3.245 8.58 3.395 ;
      RECT 8.43 4.085 8.58 4.235 ;
      RECT 7.95 3.805 8.1 3.955 ;
      RECT 7.71 3.245 7.86 3.395 ;
      RECT 7.35 4.925 7.5 5.075 ;
      RECT 7.095 3.245 7.245 3.395 ;
      RECT 6.75 4.925 6.9 5.075 ;
      RECT 6.63 3.245 6.78 3.395 ;
      RECT 6.51 3.805 6.66 3.955 ;
      RECT 6.27 4.365 6.42 4.515 ;
      RECT 5.07 3.805 5.22 3.955 ;
      RECT 4.71 3.245 4.86 3.395 ;
      RECT 4.59 4.085 4.74 4.235 ;
      RECT 3.9 3.245 4.05 3.395 ;
      RECT 3.9 4.645 4.05 4.795 ;
      RECT 1.615 9.39 1.765 9.54 ;
      RECT 1.24 8.65 1.39 8.8 ;
      RECT 0.315 10.91 0.465 11.06 ;
      RECT 0.31 0.12 0.46 0.27 ;
    LAYER met1 ;
      RECT 65.08 4.045 65.37 4.275 ;
      RECT 49.82 4.045 50.11 4.275 ;
      RECT 34.56 4.045 34.85 4.275 ;
      RECT 19.3 4.045 19.59 4.275 ;
      RECT 4.04 4.045 4.33 4.275 ;
      RECT 65.155 3.23 65.295 4.275 ;
      RECT 49.895 3.67 50.035 4.275 ;
      RECT 34.635 3.67 34.775 4.275 ;
      RECT 19.375 3.67 19.515 4.275 ;
      RECT 4.115 3.67 4.255 4.275 ;
      RECT 65.155 3.67 65.775 3.81 ;
      RECT 65.635 0.005 65.775 3.81 ;
      RECT 49.895 3.67 50.515 3.81 ;
      RECT 50.375 0.005 50.515 3.81 ;
      RECT 34.635 3.67 35.255 3.81 ;
      RECT 35.115 0.005 35.255 3.81 ;
      RECT 19.375 3.67 19.995 3.81 ;
      RECT 19.855 0.005 19.995 3.81 ;
      RECT 4.115 3.67 4.735 3.81 ;
      RECT 4.595 0.005 4.735 3.81 ;
      RECT 64.855 3.19 65.175 3.69 ;
      RECT 64.77 3.23 65.34 3.69 ;
      RECT 65.395 3.25 65.775 3.51 ;
      RECT 50.135 3.25 50.515 3.51 ;
      RECT 34.875 3.25 35.255 3.51 ;
      RECT 19.615 3.25 19.995 3.51 ;
      RECT 4.355 3.25 4.735 3.51 ;
      RECT 65.575 3.19 65.985 3.45 ;
      RECT 50.315 3.19 50.725 3.45 ;
      RECT 35.055 3.19 35.465 3.45 ;
      RECT 19.795 3.19 20.205 3.45 ;
      RECT 4.535 3.19 4.945 3.45 ;
      RECT 66.28 3.205 66.57 3.435 ;
      RECT 51.02 3.205 51.31 3.435 ;
      RECT 35.76 3.205 36.05 3.435 ;
      RECT 20.5 3.205 20.79 3.435 ;
      RECT 5.24 3.205 5.53 3.435 ;
      RECT 65.395 3.25 66.57 3.39 ;
      RECT 50.135 3.25 51.31 3.39 ;
      RECT 34.875 3.25 36.05 3.39 ;
      RECT 19.615 3.25 20.79 3.39 ;
      RECT 4.355 3.25 5.53 3.39 ;
      RECT 65.575 0.005 65.865 3.45 ;
      RECT 50.315 0.005 50.605 3.45 ;
      RECT 35.055 0.005 35.345 3.45 ;
      RECT 19.795 0.005 20.085 3.45 ;
      RECT 4.535 0.005 4.825 3.45 ;
      RECT 64.59 0.005 73.33 3.04 ;
      RECT 49.33 0.005 58.07 3.04 ;
      RECT 34.07 0.005 42.81 3.04 ;
      RECT 18.81 0.005 27.55 3.04 ;
      RECT 3.55 0.005 12.29 3.04 ;
      RECT 0.005 0.005 79.1 1.605 ;
      RECT 76.965 5.43 78.945 7.045 ;
      RECT 61.705 5.43 63.685 7.045 ;
      RECT 46.445 5.43 48.425 7.045 ;
      RECT 31.185 5.43 33.165 7.045 ;
      RECT 15.925 5.43 17.905 7.045 ;
      RECT 0.005 5.44 79.1 7.04 ;
      RECT 64.59 5.435 79.1 7.04 ;
      RECT 49.33 5.435 63.84 7.04 ;
      RECT 34.07 5.435 48.58 7.04 ;
      RECT 18.81 5.435 33.32 7.04 ;
      RECT 3.55 5.435 18.06 7.04 ;
      RECT 64.59 5.28 73.33 7.04 ;
      RECT 49.33 5.28 58.07 7.04 ;
      RECT 34.07 5.28 42.81 7.04 ;
      RECT 18.81 5.28 27.55 7.04 ;
      RECT 3.55 5.28 12.29 7.04 ;
      RECT 0.005 10.87 79.1 12.47 ;
      RECT 69.56 8.61 69.73 12.47 ;
      RECT 54.3 8.61 54.47 12.47 ;
      RECT 39.04 8.61 39.21 12.47 ;
      RECT 23.78 8.61 23.95 12.47 ;
      RECT 8.52 8.61 8.69 12.47 ;
      RECT 0.01 10.86 0.815 12.47 ;
      RECT 0.215 10.84 0.565 12.47 ;
      RECT 69.725 8.58 70.015 8.81 ;
      RECT 54.465 8.58 54.755 8.81 ;
      RECT 39.205 8.58 39.495 8.81 ;
      RECT 23.945 8.58 24.235 8.81 ;
      RECT 8.685 8.58 8.975 8.81 ;
      RECT 69.555 8.61 70.015 8.78 ;
      RECT 54.295 8.61 54.755 8.78 ;
      RECT 39.035 8.61 39.495 8.78 ;
      RECT 23.775 8.61 24.235 8.78 ;
      RECT 8.515 8.61 8.975 8.78 ;
      RECT 78.495 10.065 78.785 10.295 ;
      RECT 78.555 8.585 78.725 10.295 ;
      RECT 78.53 9.57 78.88 9.92 ;
      RECT 78.495 8.585 78.785 8.815 ;
      RECT 78.09 3.695 78.195 4.265 ;
      RECT 78.09 4.03 78.415 4.26 ;
      RECT 78.09 4.06 78.585 4.23 ;
      RECT 78.09 3.695 78.28 4.26 ;
      RECT 77.505 3.66 77.795 3.89 ;
      RECT 77.505 3.695 78.28 3.865 ;
      RECT 77.565 2.18 77.735 3.89 ;
      RECT 77.505 2.18 77.795 2.41 ;
      RECT 77.505 10.065 77.795 10.295 ;
      RECT 77.565 8.585 77.735 10.295 ;
      RECT 77.505 8.585 77.795 8.815 ;
      RECT 77.505 8.62 78.36 8.78 ;
      RECT 78.19 8.215 78.36 8.78 ;
      RECT 77.505 8.615 77.9 8.78 ;
      RECT 78.125 8.215 78.415 8.445 ;
      RECT 78.125 8.245 78.585 8.415 ;
      RECT 77.135 4.03 77.425 4.26 ;
      RECT 77.135 4.06 77.595 4.23 ;
      RECT 77.2 2.955 77.365 4.26 ;
      RECT 75.715 2.925 76.005 3.155 ;
      RECT 75.715 2.955 77.365 3.125 ;
      RECT 75.775 2.185 75.945 3.155 ;
      RECT 75.715 2.185 76.005 2.415 ;
      RECT 75.715 10.06 76.005 10.29 ;
      RECT 75.775 9.32 75.945 10.29 ;
      RECT 75.775 9.415 77.365 9.585 ;
      RECT 77.195 8.215 77.365 9.585 ;
      RECT 75.715 9.32 76.005 9.55 ;
      RECT 77.135 8.215 77.425 8.445 ;
      RECT 77.135 8.245 77.595 8.415 ;
      RECT 73.765 4 74.105 4.35 ;
      RECT 73.855 3.325 74.025 4.35 ;
      RECT 76.145 3.265 76.495 3.615 ;
      RECT 73.855 3.325 76.495 3.495 ;
      RECT 76.17 8.95 76.495 9.275 ;
      RECT 70.73 8.905 71.08 9.255 ;
      RECT 76.145 8.95 76.495 9.18 ;
      RECT 70.53 8.95 71.08 9.18 ;
      RECT 70.36 8.98 76.495 9.15 ;
      RECT 75.37 3.665 75.69 3.985 ;
      RECT 75.34 3.665 75.69 3.895 ;
      RECT 75.17 3.695 75.69 3.865 ;
      RECT 75.37 8.55 75.69 8.84 ;
      RECT 75.34 8.58 75.69 8.81 ;
      RECT 75.17 8.61 75.69 8.78 ;
      RECT 72.475 3.19 72.795 3.45 ;
      RECT 72.04 3.205 72.33 3.435 ;
      RECT 72.04 3.25 72.795 3.39 ;
      RECT 72.475 4.87 72.795 5.13 ;
      RECT 72.04 4.885 72.33 5.115 ;
      RECT 72.04 4.93 72.795 5.07 ;
      RECT 71.8 4.325 72.09 4.555 ;
      RECT 71.8 4.37 72.375 4.51 ;
      RECT 72.235 4.23 72.495 4.37 ;
      RECT 72.28 4.045 72.57 4.275 ;
      RECT 70.435 4.23 71.535 4.37 ;
      RECT 70.24 4.03 70.56 4.29 ;
      RECT 71.32 4.045 71.61 4.275 ;
      RECT 70.24 4.045 70.65 4.29 ;
      RECT 70.615 3.19 70.935 3.45 ;
      RECT 71.08 3.205 71.37 3.435 ;
      RECT 70.615 3.25 71.37 3.39 ;
      RECT 67.915 4.455 70.095 4.595 ;
      RECT 69.955 3.465 70.095 4.595 ;
      RECT 67.915 4.37 69.21 4.595 ;
      RECT 68.92 4.325 69.21 4.595 ;
      RECT 67.915 4.09 68.25 4.595 ;
      RECT 67.96 4.045 68.25 4.595 ;
      RECT 70.84 3.765 71.13 3.995 ;
      RECT 69.955 3.67 71.055 3.81 ;
      RECT 69.88 3.465 70.17 3.715 ;
      RECT 70.1 10.06 70.39 10.29 ;
      RECT 70.16 9.32 70.33 10.29 ;
      RECT 70.06 9.35 70.43 9.72 ;
      RECT 70.1 9.32 70.39 9.72 ;
      RECT 69.865 4.87 70.185 5.13 ;
      RECT 69.865 4.885 70.38 5.115 ;
      RECT 68.44 3.765 68.73 3.995 ;
      RECT 68.59 3.37 68.73 3.995 ;
      RECT 68.59 3.37 68.895 3.51 ;
      RECT 69.385 3.19 69.705 3.45 ;
      RECT 68.665 3.19 68.985 3.45 ;
      RECT 69.16 3.205 69.705 3.435 ;
      RECT 68.665 3.25 69.705 3.39 ;
      RECT 68.305 4.87 68.625 5.13 ;
      RECT 68.2 4.885 68.625 5.115 ;
      RECT 66.28 4.325 66.57 4.555 ;
      RECT 66.28 4.325 66.735 4.51 ;
      RECT 66.595 3.85 66.735 4.51 ;
      RECT 66.715 3.25 66.855 3.99 ;
      RECT 67.585 3.19 67.905 3.45 ;
      RECT 66.76 3.205 67.05 3.435 ;
      RECT 66.715 3.25 67.905 3.39 ;
      RECT 67.465 3.75 67.785 4.01 ;
      RECT 67 3.765 67.29 3.995 ;
      RECT 67 3.81 67.785 3.95 ;
      RECT 67.225 4.31 67.545 4.57 ;
      RECT 67.225 4.325 67.77 4.555 ;
      RECT 66.76 4.885 67.05 5.115 ;
      RECT 65.875 4.765 66.975 4.905 ;
      RECT 65.8 4.605 66.09 4.835 ;
      RECT 63.235 10.065 63.525 10.295 ;
      RECT 63.295 8.585 63.465 10.295 ;
      RECT 63.245 8.95 63.595 9.3 ;
      RECT 63.235 8.585 63.525 8.815 ;
      RECT 62.83 3.695 62.935 4.265 ;
      RECT 62.83 4.03 63.155 4.26 ;
      RECT 62.83 4.06 63.325 4.23 ;
      RECT 62.83 3.695 63.02 4.26 ;
      RECT 62.245 3.66 62.535 3.89 ;
      RECT 62.245 3.695 63.02 3.865 ;
      RECT 62.305 2.18 62.475 3.89 ;
      RECT 62.245 2.18 62.535 2.41 ;
      RECT 62.245 10.065 62.535 10.295 ;
      RECT 62.305 8.585 62.475 10.295 ;
      RECT 62.245 8.585 62.535 8.815 ;
      RECT 62.245 8.62 63.1 8.78 ;
      RECT 62.93 8.215 63.1 8.78 ;
      RECT 62.245 8.615 62.64 8.78 ;
      RECT 62.865 8.215 63.155 8.445 ;
      RECT 62.865 8.245 63.325 8.415 ;
      RECT 61.875 4.03 62.165 4.26 ;
      RECT 61.875 4.06 62.335 4.23 ;
      RECT 61.94 2.955 62.105 4.26 ;
      RECT 60.455 2.925 60.745 3.155 ;
      RECT 60.455 2.955 62.105 3.125 ;
      RECT 60.515 2.185 60.685 3.155 ;
      RECT 60.455 2.185 60.745 2.415 ;
      RECT 60.455 10.06 60.745 10.29 ;
      RECT 60.515 9.32 60.685 10.29 ;
      RECT 60.515 9.415 62.105 9.585 ;
      RECT 61.935 8.215 62.105 9.585 ;
      RECT 60.455 9.32 60.745 9.55 ;
      RECT 61.875 8.215 62.165 8.445 ;
      RECT 61.875 8.245 62.335 8.415 ;
      RECT 58.505 4 58.845 4.35 ;
      RECT 58.595 3.325 58.765 4.35 ;
      RECT 60.885 3.265 61.235 3.615 ;
      RECT 58.595 3.325 61.235 3.495 ;
      RECT 60.91 8.95 61.235 9.275 ;
      RECT 55.475 8.905 55.825 9.255 ;
      RECT 60.885 8.95 61.235 9.18 ;
      RECT 55.27 8.95 55.825 9.18 ;
      RECT 55.1 8.98 61.235 9.15 ;
      RECT 60.11 3.665 60.43 3.985 ;
      RECT 60.08 3.665 60.43 3.895 ;
      RECT 59.91 3.695 60.43 3.865 ;
      RECT 60.11 8.55 60.43 8.84 ;
      RECT 60.08 8.58 60.43 8.81 ;
      RECT 59.91 8.61 60.43 8.78 ;
      RECT 57.215 3.19 57.535 3.45 ;
      RECT 56.78 3.205 57.07 3.435 ;
      RECT 56.78 3.25 57.535 3.39 ;
      RECT 57.215 4.87 57.535 5.13 ;
      RECT 56.78 4.885 57.07 5.115 ;
      RECT 56.78 4.93 57.535 5.07 ;
      RECT 56.54 4.325 56.83 4.555 ;
      RECT 56.54 4.37 57.115 4.51 ;
      RECT 56.975 4.23 57.235 4.37 ;
      RECT 57.02 4.045 57.31 4.275 ;
      RECT 55.175 4.23 56.275 4.37 ;
      RECT 54.98 4.03 55.3 4.29 ;
      RECT 56.06 4.045 56.35 4.275 ;
      RECT 54.98 4.045 55.39 4.29 ;
      RECT 55.355 3.19 55.675 3.45 ;
      RECT 55.82 3.205 56.11 3.435 ;
      RECT 55.355 3.25 56.11 3.39 ;
      RECT 52.655 4.455 54.835 4.595 ;
      RECT 54.695 3.465 54.835 4.595 ;
      RECT 52.655 4.37 53.95 4.595 ;
      RECT 53.66 4.325 53.95 4.595 ;
      RECT 52.655 4.09 52.99 4.595 ;
      RECT 52.7 4.045 52.99 4.595 ;
      RECT 55.58 3.765 55.87 3.995 ;
      RECT 54.695 3.67 55.795 3.81 ;
      RECT 54.62 3.465 54.91 3.715 ;
      RECT 54.84 10.06 55.13 10.29 ;
      RECT 54.9 9.32 55.07 10.29 ;
      RECT 54.8 9.35 55.17 9.72 ;
      RECT 54.84 9.32 55.13 9.72 ;
      RECT 54.605 4.87 54.925 5.13 ;
      RECT 54.605 4.885 55.12 5.115 ;
      RECT 53.18 3.765 53.47 3.995 ;
      RECT 53.33 3.37 53.47 3.995 ;
      RECT 53.33 3.37 53.635 3.51 ;
      RECT 54.125 3.19 54.445 3.45 ;
      RECT 53.405 3.19 53.725 3.45 ;
      RECT 53.9 3.205 54.445 3.435 ;
      RECT 53.405 3.25 54.445 3.39 ;
      RECT 53.045 4.87 53.365 5.13 ;
      RECT 52.94 4.885 53.365 5.115 ;
      RECT 51.02 4.325 51.31 4.555 ;
      RECT 51.02 4.325 51.475 4.51 ;
      RECT 51.335 3.85 51.475 4.51 ;
      RECT 51.455 3.25 51.595 3.99 ;
      RECT 52.325 3.19 52.645 3.45 ;
      RECT 51.5 3.205 51.79 3.435 ;
      RECT 51.455 3.25 52.645 3.39 ;
      RECT 52.205 3.75 52.525 4.01 ;
      RECT 51.74 3.765 52.03 3.995 ;
      RECT 51.74 3.81 52.525 3.95 ;
      RECT 51.965 4.31 52.285 4.57 ;
      RECT 51.965 4.325 52.51 4.555 ;
      RECT 51.5 4.885 51.79 5.115 ;
      RECT 50.615 4.765 51.715 4.905 ;
      RECT 50.54 4.605 50.83 4.835 ;
      RECT 47.975 10.065 48.265 10.295 ;
      RECT 48.035 8.585 48.205 10.295 ;
      RECT 47.985 8.95 48.335 9.3 ;
      RECT 47.975 8.585 48.265 8.815 ;
      RECT 47.57 3.695 47.675 4.265 ;
      RECT 47.57 4.03 47.895 4.26 ;
      RECT 47.57 4.06 48.065 4.23 ;
      RECT 47.57 3.695 47.76 4.26 ;
      RECT 46.985 3.66 47.275 3.89 ;
      RECT 46.985 3.695 47.76 3.865 ;
      RECT 47.045 2.18 47.215 3.89 ;
      RECT 46.985 2.18 47.275 2.41 ;
      RECT 46.985 10.065 47.275 10.295 ;
      RECT 47.045 8.585 47.215 10.295 ;
      RECT 46.985 8.585 47.275 8.815 ;
      RECT 46.985 8.62 47.84 8.78 ;
      RECT 47.67 8.215 47.84 8.78 ;
      RECT 46.985 8.615 47.38 8.78 ;
      RECT 47.605 8.215 47.895 8.445 ;
      RECT 47.605 8.245 48.065 8.415 ;
      RECT 46.615 4.03 46.905 4.26 ;
      RECT 46.615 4.06 47.075 4.23 ;
      RECT 46.68 2.955 46.845 4.26 ;
      RECT 45.195 2.925 45.485 3.155 ;
      RECT 45.195 2.955 46.845 3.125 ;
      RECT 45.255 2.185 45.425 3.155 ;
      RECT 45.195 2.185 45.485 2.415 ;
      RECT 45.195 10.06 45.485 10.29 ;
      RECT 45.255 9.32 45.425 10.29 ;
      RECT 45.255 9.415 46.845 9.585 ;
      RECT 46.675 8.215 46.845 9.585 ;
      RECT 45.195 9.32 45.485 9.55 ;
      RECT 46.615 8.215 46.905 8.445 ;
      RECT 46.615 8.245 47.075 8.415 ;
      RECT 43.245 4 43.585 4.35 ;
      RECT 43.335 3.325 43.505 4.35 ;
      RECT 45.625 3.265 45.975 3.615 ;
      RECT 43.335 3.325 45.975 3.495 ;
      RECT 45.65 8.95 45.975 9.275 ;
      RECT 40.21 8.91 40.56 9.26 ;
      RECT 45.625 8.95 45.975 9.18 ;
      RECT 40.01 8.95 40.56 9.18 ;
      RECT 39.84 8.98 45.975 9.15 ;
      RECT 44.85 3.665 45.17 3.985 ;
      RECT 44.82 3.665 45.17 3.895 ;
      RECT 44.65 3.695 45.17 3.865 ;
      RECT 44.85 8.55 45.17 8.84 ;
      RECT 44.82 8.58 45.17 8.81 ;
      RECT 44.65 8.61 45.17 8.78 ;
      RECT 41.955 3.19 42.275 3.45 ;
      RECT 41.52 3.205 41.81 3.435 ;
      RECT 41.52 3.25 42.275 3.39 ;
      RECT 41.955 4.87 42.275 5.13 ;
      RECT 41.52 4.885 41.81 5.115 ;
      RECT 41.52 4.93 42.275 5.07 ;
      RECT 41.28 4.325 41.57 4.555 ;
      RECT 41.28 4.37 41.855 4.51 ;
      RECT 41.715 4.23 41.975 4.37 ;
      RECT 41.76 4.045 42.05 4.275 ;
      RECT 39.915 4.23 41.015 4.37 ;
      RECT 39.72 4.03 40.04 4.29 ;
      RECT 40.8 4.045 41.09 4.275 ;
      RECT 39.72 4.045 40.13 4.29 ;
      RECT 40.095 3.19 40.415 3.45 ;
      RECT 40.56 3.205 40.85 3.435 ;
      RECT 40.095 3.25 40.85 3.39 ;
      RECT 37.395 4.455 39.575 4.595 ;
      RECT 39.435 3.465 39.575 4.595 ;
      RECT 37.395 4.37 38.69 4.595 ;
      RECT 38.4 4.325 38.69 4.595 ;
      RECT 37.395 4.09 37.73 4.595 ;
      RECT 37.44 4.045 37.73 4.595 ;
      RECT 40.32 3.765 40.61 3.995 ;
      RECT 39.435 3.67 40.535 3.81 ;
      RECT 39.36 3.465 39.65 3.715 ;
      RECT 39.58 10.06 39.87 10.29 ;
      RECT 39.64 9.32 39.81 10.29 ;
      RECT 39.54 9.35 39.91 9.72 ;
      RECT 39.58 9.32 39.87 9.72 ;
      RECT 39.345 4.87 39.665 5.13 ;
      RECT 39.345 4.885 39.86 5.115 ;
      RECT 37.92 3.765 38.21 3.995 ;
      RECT 38.07 3.37 38.21 3.995 ;
      RECT 38.07 3.37 38.375 3.51 ;
      RECT 38.865 3.19 39.185 3.45 ;
      RECT 38.145 3.19 38.465 3.45 ;
      RECT 38.64 3.205 39.185 3.435 ;
      RECT 38.145 3.25 39.185 3.39 ;
      RECT 37.785 4.87 38.105 5.13 ;
      RECT 37.68 4.885 38.105 5.115 ;
      RECT 35.76 4.325 36.05 4.555 ;
      RECT 35.76 4.325 36.215 4.51 ;
      RECT 36.075 3.85 36.215 4.51 ;
      RECT 36.195 3.25 36.335 3.99 ;
      RECT 37.065 3.19 37.385 3.45 ;
      RECT 36.24 3.205 36.53 3.435 ;
      RECT 36.195 3.25 37.385 3.39 ;
      RECT 36.945 3.75 37.265 4.01 ;
      RECT 36.48 3.765 36.77 3.995 ;
      RECT 36.48 3.81 37.265 3.95 ;
      RECT 36.705 4.31 37.025 4.57 ;
      RECT 36.705 4.325 37.25 4.555 ;
      RECT 36.24 4.885 36.53 5.115 ;
      RECT 35.355 4.765 36.455 4.905 ;
      RECT 35.28 4.605 35.57 4.835 ;
      RECT 32.715 10.065 33.005 10.295 ;
      RECT 32.775 8.585 32.945 10.295 ;
      RECT 32.765 8.955 33.12 9.31 ;
      RECT 32.715 8.585 33.005 8.815 ;
      RECT 32.31 3.695 32.415 4.265 ;
      RECT 32.31 4.03 32.635 4.26 ;
      RECT 32.31 4.06 32.805 4.23 ;
      RECT 32.31 3.695 32.5 4.26 ;
      RECT 31.725 3.66 32.015 3.89 ;
      RECT 31.725 3.695 32.5 3.865 ;
      RECT 31.785 2.18 31.955 3.89 ;
      RECT 31.725 2.18 32.015 2.41 ;
      RECT 31.725 10.065 32.015 10.295 ;
      RECT 31.785 8.585 31.955 10.295 ;
      RECT 31.725 8.585 32.015 8.815 ;
      RECT 31.725 8.62 32.58 8.78 ;
      RECT 32.41 8.215 32.58 8.78 ;
      RECT 31.725 8.615 32.12 8.78 ;
      RECT 32.345 8.215 32.635 8.445 ;
      RECT 32.345 8.245 32.805 8.415 ;
      RECT 31.355 4.03 31.645 4.26 ;
      RECT 31.355 4.06 31.815 4.23 ;
      RECT 31.42 2.955 31.585 4.26 ;
      RECT 29.935 2.925 30.225 3.155 ;
      RECT 29.935 2.955 31.585 3.125 ;
      RECT 29.995 2.185 30.165 3.155 ;
      RECT 29.935 2.185 30.225 2.415 ;
      RECT 29.935 10.06 30.225 10.29 ;
      RECT 29.995 9.32 30.165 10.29 ;
      RECT 29.995 9.415 31.585 9.585 ;
      RECT 31.415 8.215 31.585 9.585 ;
      RECT 29.935 9.32 30.225 9.55 ;
      RECT 31.355 8.215 31.645 8.445 ;
      RECT 31.355 8.245 31.815 8.415 ;
      RECT 27.985 4 28.325 4.35 ;
      RECT 28.075 3.325 28.245 4.35 ;
      RECT 30.365 3.265 30.715 3.615 ;
      RECT 28.075 3.325 30.715 3.495 ;
      RECT 30.39 8.95 30.715 9.275 ;
      RECT 24.95 8.905 25.3 9.255 ;
      RECT 30.365 8.95 30.715 9.18 ;
      RECT 24.75 8.95 25.3 9.18 ;
      RECT 24.58 8.98 30.715 9.15 ;
      RECT 29.59 3.665 29.91 3.985 ;
      RECT 29.56 3.665 29.91 3.895 ;
      RECT 29.39 3.695 29.91 3.865 ;
      RECT 29.59 8.55 29.91 8.84 ;
      RECT 29.56 8.58 29.91 8.81 ;
      RECT 29.39 8.61 29.91 8.78 ;
      RECT 26.695 3.19 27.015 3.45 ;
      RECT 26.26 3.205 26.55 3.435 ;
      RECT 26.26 3.25 27.015 3.39 ;
      RECT 26.695 4.87 27.015 5.13 ;
      RECT 26.26 4.885 26.55 5.115 ;
      RECT 26.26 4.93 27.015 5.07 ;
      RECT 26.02 4.325 26.31 4.555 ;
      RECT 26.02 4.37 26.595 4.51 ;
      RECT 26.455 4.23 26.715 4.37 ;
      RECT 26.5 4.045 26.79 4.275 ;
      RECT 24.655 4.23 25.755 4.37 ;
      RECT 24.46 4.03 24.78 4.29 ;
      RECT 25.54 4.045 25.83 4.275 ;
      RECT 24.46 4.045 24.87 4.29 ;
      RECT 24.835 3.19 25.155 3.45 ;
      RECT 25.3 3.205 25.59 3.435 ;
      RECT 24.835 3.25 25.59 3.39 ;
      RECT 22.135 4.455 24.315 4.595 ;
      RECT 24.175 3.465 24.315 4.595 ;
      RECT 22.135 4.37 23.43 4.595 ;
      RECT 23.14 4.325 23.43 4.595 ;
      RECT 22.135 4.09 22.47 4.595 ;
      RECT 22.18 4.045 22.47 4.595 ;
      RECT 25.06 3.765 25.35 3.995 ;
      RECT 24.175 3.67 25.275 3.81 ;
      RECT 24.1 3.465 24.39 3.715 ;
      RECT 24.32 10.06 24.61 10.29 ;
      RECT 24.38 9.32 24.55 10.29 ;
      RECT 24.28 9.35 24.65 9.72 ;
      RECT 24.32 9.32 24.61 9.72 ;
      RECT 24.085 4.87 24.405 5.13 ;
      RECT 24.085 4.885 24.6 5.115 ;
      RECT 22.66 3.765 22.95 3.995 ;
      RECT 22.81 3.37 22.95 3.995 ;
      RECT 22.81 3.37 23.115 3.51 ;
      RECT 23.605 3.19 23.925 3.45 ;
      RECT 22.885 3.19 23.205 3.45 ;
      RECT 23.38 3.205 23.925 3.435 ;
      RECT 22.885 3.25 23.925 3.39 ;
      RECT 22.525 4.87 22.845 5.13 ;
      RECT 22.42 4.885 22.845 5.115 ;
      RECT 20.5 4.325 20.79 4.555 ;
      RECT 20.5 4.325 20.955 4.51 ;
      RECT 20.815 3.85 20.955 4.51 ;
      RECT 20.935 3.25 21.075 3.99 ;
      RECT 21.805 3.19 22.125 3.45 ;
      RECT 20.98 3.205 21.27 3.435 ;
      RECT 20.935 3.25 22.125 3.39 ;
      RECT 21.685 3.75 22.005 4.01 ;
      RECT 21.22 3.765 21.51 3.995 ;
      RECT 21.22 3.81 22.005 3.95 ;
      RECT 21.445 4.31 21.765 4.57 ;
      RECT 21.445 4.325 21.99 4.555 ;
      RECT 20.98 4.885 21.27 5.115 ;
      RECT 20.095 4.765 21.195 4.905 ;
      RECT 20.02 4.605 20.31 4.835 ;
      RECT 17.455 10.065 17.745 10.295 ;
      RECT 17.515 8.585 17.685 10.295 ;
      RECT 17.51 8.95 17.86 9.3 ;
      RECT 17.455 8.585 17.745 8.815 ;
      RECT 17.05 3.695 17.155 4.265 ;
      RECT 17.05 4.03 17.375 4.26 ;
      RECT 17.05 4.06 17.545 4.23 ;
      RECT 17.05 3.695 17.24 4.26 ;
      RECT 16.465 3.66 16.755 3.89 ;
      RECT 16.465 3.695 17.24 3.865 ;
      RECT 16.525 2.18 16.695 3.89 ;
      RECT 16.465 2.18 16.755 2.41 ;
      RECT 16.465 10.065 16.755 10.295 ;
      RECT 16.525 8.585 16.695 10.295 ;
      RECT 16.465 8.585 16.755 8.815 ;
      RECT 16.465 8.62 17.32 8.78 ;
      RECT 17.15 8.215 17.32 8.78 ;
      RECT 16.465 8.615 16.86 8.78 ;
      RECT 17.085 8.215 17.375 8.445 ;
      RECT 17.085 8.245 17.545 8.415 ;
      RECT 16.095 4.03 16.385 4.26 ;
      RECT 16.095 4.06 16.555 4.23 ;
      RECT 16.16 2.955 16.325 4.26 ;
      RECT 14.675 2.925 14.965 3.155 ;
      RECT 14.675 2.955 16.325 3.125 ;
      RECT 14.735 2.185 14.905 3.155 ;
      RECT 14.675 2.185 14.965 2.415 ;
      RECT 14.675 10.06 14.965 10.29 ;
      RECT 14.735 9.32 14.905 10.29 ;
      RECT 14.735 9.415 16.325 9.585 ;
      RECT 16.155 8.215 16.325 9.585 ;
      RECT 14.675 9.32 14.965 9.55 ;
      RECT 16.095 8.215 16.385 8.445 ;
      RECT 16.095 8.245 16.555 8.415 ;
      RECT 12.725 4 13.065 4.35 ;
      RECT 12.815 3.325 12.985 4.35 ;
      RECT 15.105 3.265 15.455 3.615 ;
      RECT 12.815 3.325 15.455 3.495 ;
      RECT 15.13 8.95 15.455 9.275 ;
      RECT 9.69 8.9 10.04 9.25 ;
      RECT 15.105 8.95 15.455 9.18 ;
      RECT 9.49 8.95 10.04 9.18 ;
      RECT 9.32 8.98 15.455 9.15 ;
      RECT 14.33 3.665 14.65 3.985 ;
      RECT 14.3 3.665 14.65 3.895 ;
      RECT 14.13 3.695 14.65 3.865 ;
      RECT 14.33 8.55 14.65 8.84 ;
      RECT 14.3 8.58 14.65 8.81 ;
      RECT 14.13 8.61 14.65 8.78 ;
      RECT 11.435 3.19 11.755 3.45 ;
      RECT 11 3.205 11.29 3.435 ;
      RECT 11 3.25 11.755 3.39 ;
      RECT 11.435 4.87 11.755 5.13 ;
      RECT 11 4.885 11.29 5.115 ;
      RECT 11 4.93 11.755 5.07 ;
      RECT 10.76 4.325 11.05 4.555 ;
      RECT 10.76 4.37 11.335 4.51 ;
      RECT 11.195 4.23 11.455 4.37 ;
      RECT 11.24 4.045 11.53 4.275 ;
      RECT 9.395 4.23 10.495 4.37 ;
      RECT 9.2 4.03 9.52 4.29 ;
      RECT 10.28 4.045 10.57 4.275 ;
      RECT 9.2 4.045 9.61 4.29 ;
      RECT 9.575 3.19 9.895 3.45 ;
      RECT 10.04 3.205 10.33 3.435 ;
      RECT 9.575 3.25 10.33 3.39 ;
      RECT 6.875 4.455 9.055 4.595 ;
      RECT 8.915 3.465 9.055 4.595 ;
      RECT 6.875 4.37 8.17 4.595 ;
      RECT 7.88 4.325 8.17 4.595 ;
      RECT 6.875 4.09 7.21 4.595 ;
      RECT 6.92 4.045 7.21 4.595 ;
      RECT 9.8 3.765 10.09 3.995 ;
      RECT 8.915 3.67 10.015 3.81 ;
      RECT 8.84 3.465 9.13 3.715 ;
      RECT 9.06 10.06 9.35 10.29 ;
      RECT 9.12 9.32 9.29 10.29 ;
      RECT 9.02 9.35 9.39 9.72 ;
      RECT 9.06 9.32 9.35 9.72 ;
      RECT 8.825 4.87 9.145 5.13 ;
      RECT 8.825 4.885 9.34 5.115 ;
      RECT 7.4 3.765 7.69 3.995 ;
      RECT 7.55 3.37 7.69 3.995 ;
      RECT 7.55 3.37 7.855 3.51 ;
      RECT 8.345 3.19 8.665 3.45 ;
      RECT 7.625 3.19 7.945 3.45 ;
      RECT 8.12 3.205 8.665 3.435 ;
      RECT 7.625 3.25 8.665 3.39 ;
      RECT 7.265 4.87 7.585 5.13 ;
      RECT 7.16 4.885 7.585 5.115 ;
      RECT 5.24 4.325 5.53 4.555 ;
      RECT 5.24 4.325 5.695 4.51 ;
      RECT 5.555 3.85 5.695 4.51 ;
      RECT 5.675 3.25 5.815 3.99 ;
      RECT 6.545 3.19 6.865 3.45 ;
      RECT 5.72 3.205 6.01 3.435 ;
      RECT 5.675 3.25 6.865 3.39 ;
      RECT 6.425 3.75 6.745 4.01 ;
      RECT 5.96 3.765 6.25 3.995 ;
      RECT 5.96 3.81 6.745 3.95 ;
      RECT 6.185 4.31 6.505 4.57 ;
      RECT 6.185 4.325 6.73 4.555 ;
      RECT 5.72 4.885 6.01 5.115 ;
      RECT 4.835 4.765 5.935 4.905 ;
      RECT 4.76 4.605 5.05 4.835 ;
      RECT 1.975 8.95 2.265 9.18 ;
      RECT 1.805 8.98 2.265 9.15 ;
      RECT 1.545 10.06 1.835 10.29 ;
      RECT 1.605 9.32 1.775 10.29 ;
      RECT 1.515 9.32 1.865 9.61 ;
      RECT 1.14 8.58 1.49 8.87 ;
      RECT 1 8.61 1.49 8.78 ;
      RECT 71.785 3.75 72.105 4.01 ;
      RECT 70.615 4.59 70.935 4.85 ;
      RECT 69.385 4.03 69.705 4.29 ;
      RECT 68.905 3.75 69.225 4.01 ;
      RECT 68.05 3.19 68.45 3.45 ;
      RECT 67.705 4.87 68.025 5.13 ;
      RECT 66.025 3.75 66.345 4.01 ;
      RECT 65.545 4.03 65.865 4.29 ;
      RECT 64.855 4.59 65.175 4.85 ;
      RECT 56.525 3.75 56.845 4.01 ;
      RECT 55.355 4.59 55.675 4.85 ;
      RECT 54.125 4.03 54.445 4.29 ;
      RECT 53.645 3.75 53.965 4.01 ;
      RECT 52.79 3.19 53.19 3.45 ;
      RECT 52.445 4.87 52.765 5.13 ;
      RECT 50.765 3.75 51.085 4.01 ;
      RECT 50.285 4.03 50.605 4.29 ;
      RECT 49.595 3.19 49.915 3.45 ;
      RECT 49.595 4.59 49.915 4.85 ;
      RECT 41.265 3.75 41.585 4.01 ;
      RECT 40.095 4.59 40.415 4.85 ;
      RECT 38.865 4.03 39.185 4.29 ;
      RECT 38.385 3.75 38.705 4.01 ;
      RECT 37.53 3.19 37.93 3.45 ;
      RECT 37.185 4.87 37.505 5.13 ;
      RECT 35.505 3.75 35.825 4.01 ;
      RECT 35.025 4.03 35.345 4.29 ;
      RECT 34.335 3.19 34.655 3.45 ;
      RECT 34.335 4.59 34.655 4.85 ;
      RECT 26.005 3.75 26.325 4.01 ;
      RECT 24.835 4.59 25.155 4.85 ;
      RECT 23.605 4.03 23.925 4.29 ;
      RECT 23.125 3.75 23.445 4.01 ;
      RECT 22.27 3.19 22.67 3.45 ;
      RECT 21.925 4.87 22.245 5.13 ;
      RECT 20.245 3.75 20.565 4.01 ;
      RECT 19.765 4.03 20.085 4.29 ;
      RECT 19.075 3.19 19.395 3.45 ;
      RECT 19.075 4.59 19.395 4.85 ;
      RECT 10.745 3.75 11.065 4.01 ;
      RECT 9.575 4.59 9.895 4.85 ;
      RECT 8.345 4.03 8.665 4.29 ;
      RECT 7.865 3.75 8.185 4.01 ;
      RECT 7.01 3.19 7.41 3.45 ;
      RECT 6.665 4.87 6.985 5.13 ;
      RECT 4.985 3.75 5.305 4.01 ;
      RECT 4.505 4.03 4.825 4.29 ;
      RECT 3.815 3.19 4.135 3.45 ;
      RECT 3.815 4.59 4.135 4.85 ;
    LAYER mcon ;
      RECT 78.555 8.615 78.725 8.785 ;
      RECT 78.555 10.095 78.725 10.265 ;
      RECT 78.205 1.4 78.375 1.57 ;
      RECT 78.205 5.46 78.375 5.63 ;
      RECT 78.205 6.845 78.375 7.015 ;
      RECT 78.205 10.905 78.375 11.075 ;
      RECT 78.185 4.06 78.355 4.23 ;
      RECT 78.185 8.245 78.355 8.415 ;
      RECT 77.565 2.21 77.735 2.38 ;
      RECT 77.565 3.69 77.735 3.86 ;
      RECT 77.565 8.615 77.735 8.785 ;
      RECT 77.565 10.095 77.735 10.265 ;
      RECT 77.215 1.4 77.385 1.57 ;
      RECT 77.215 5.46 77.385 5.63 ;
      RECT 77.215 6.845 77.385 7.015 ;
      RECT 77.215 10.905 77.385 11.075 ;
      RECT 77.195 4.06 77.365 4.23 ;
      RECT 77.195 8.245 77.365 8.415 ;
      RECT 76.515 1.405 76.685 1.575 ;
      RECT 76.515 5.465 76.685 5.635 ;
      RECT 76.515 6.84 76.685 7.01 ;
      RECT 76.515 10.9 76.685 11.07 ;
      RECT 76.205 3.325 76.375 3.495 ;
      RECT 76.205 8.98 76.375 9.15 ;
      RECT 75.835 1.405 76.005 1.575 ;
      RECT 75.835 10.9 76.005 11.07 ;
      RECT 75.775 2.215 75.945 2.385 ;
      RECT 75.775 2.955 75.945 3.125 ;
      RECT 75.775 9.35 75.945 9.52 ;
      RECT 75.775 10.09 75.945 10.26 ;
      RECT 75.4 3.695 75.57 3.865 ;
      RECT 75.4 8.61 75.57 8.78 ;
      RECT 75.155 1.405 75.325 1.575 ;
      RECT 75.155 10.9 75.325 11.07 ;
      RECT 74.475 1.405 74.645 1.575 ;
      RECT 74.475 10.9 74.645 11.07 ;
      RECT 73.015 2.715 73.185 2.885 ;
      RECT 73.015 5.435 73.185 5.605 ;
      RECT 72.555 2.715 72.725 2.885 ;
      RECT 72.555 5.435 72.725 5.605 ;
      RECT 72.34 4.075 72.51 4.245 ;
      RECT 72.1 3.235 72.27 3.405 ;
      RECT 72.1 4.915 72.27 5.085 ;
      RECT 72.095 2.715 72.265 2.885 ;
      RECT 72.095 5.435 72.265 5.605 ;
      RECT 71.86 3.795 72.03 3.965 ;
      RECT 71.86 4.355 72.03 4.525 ;
      RECT 71.635 2.715 71.805 2.885 ;
      RECT 71.635 5.435 71.805 5.605 ;
      RECT 71.38 4.075 71.55 4.245 ;
      RECT 71.175 2.715 71.345 2.885 ;
      RECT 71.175 5.435 71.345 5.605 ;
      RECT 71.14 3.235 71.31 3.405 ;
      RECT 70.9 3.795 71.07 3.965 ;
      RECT 70.9 6.84 71.07 7.01 ;
      RECT 70.9 10.9 71.07 11.07 ;
      RECT 70.715 2.715 70.885 2.885 ;
      RECT 70.715 5.435 70.885 5.605 ;
      RECT 70.69 4.635 70.86 4.805 ;
      RECT 70.59 8.98 70.76 9.15 ;
      RECT 70.42 4.075 70.59 4.245 ;
      RECT 70.255 2.715 70.425 2.885 ;
      RECT 70.255 5.435 70.425 5.605 ;
      RECT 70.22 10.9 70.39 11.07 ;
      RECT 70.16 9.35 70.33 9.52 ;
      RECT 70.16 10.09 70.33 10.26 ;
      RECT 70.15 4.915 70.32 5.085 ;
      RECT 69.94 3.495 70.11 3.665 ;
      RECT 69.795 2.715 69.965 2.885 ;
      RECT 69.795 5.435 69.965 5.605 ;
      RECT 69.785 8.61 69.955 8.78 ;
      RECT 69.54 10.9 69.71 11.07 ;
      RECT 69.46 4.075 69.63 4.245 ;
      RECT 69.335 2.715 69.505 2.885 ;
      RECT 69.335 5.435 69.505 5.605 ;
      RECT 69.22 3.235 69.39 3.405 ;
      RECT 68.98 3.795 69.15 3.965 ;
      RECT 68.98 4.355 69.15 4.525 ;
      RECT 68.875 2.715 69.045 2.885 ;
      RECT 68.875 5.435 69.045 5.605 ;
      RECT 68.86 10.9 69.03 11.07 ;
      RECT 68.5 3.795 68.67 3.965 ;
      RECT 68.415 2.715 68.585 2.885 ;
      RECT 68.415 5.435 68.585 5.605 ;
      RECT 68.26 4.915 68.43 5.085 ;
      RECT 68.22 3.235 68.39 3.405 ;
      RECT 68.02 4.075 68.19 4.245 ;
      RECT 67.955 2.715 68.125 2.885 ;
      RECT 67.955 5.435 68.125 5.605 ;
      RECT 67.78 4.915 67.95 5.085 ;
      RECT 67.54 4.355 67.71 4.525 ;
      RECT 67.495 2.715 67.665 2.885 ;
      RECT 67.495 5.435 67.665 5.605 ;
      RECT 67.06 3.795 67.23 3.965 ;
      RECT 67.035 2.715 67.205 2.885 ;
      RECT 67.035 5.435 67.205 5.605 ;
      RECT 66.82 3.235 66.99 3.405 ;
      RECT 66.82 4.915 66.99 5.085 ;
      RECT 66.575 2.715 66.745 2.885 ;
      RECT 66.575 5.435 66.745 5.605 ;
      RECT 66.34 3.235 66.51 3.405 ;
      RECT 66.34 4.355 66.51 4.525 ;
      RECT 66.115 2.715 66.285 2.885 ;
      RECT 66.115 5.435 66.285 5.605 ;
      RECT 66.1 3.795 66.27 3.965 ;
      RECT 65.86 4.635 66.03 4.805 ;
      RECT 65.655 2.715 65.825 2.885 ;
      RECT 65.655 5.435 65.825 5.605 ;
      RECT 65.62 4.075 65.79 4.245 ;
      RECT 65.195 2.715 65.365 2.885 ;
      RECT 65.195 5.435 65.365 5.605 ;
      RECT 65.14 4.075 65.31 4.245 ;
      RECT 64.93 3.235 65.1 3.405 ;
      RECT 64.93 4.635 65.1 4.805 ;
      RECT 64.735 2.715 64.905 2.885 ;
      RECT 64.735 5.435 64.905 5.605 ;
      RECT 63.295 8.615 63.465 8.785 ;
      RECT 63.295 10.095 63.465 10.265 ;
      RECT 62.945 1.4 63.115 1.57 ;
      RECT 62.945 5.46 63.115 5.63 ;
      RECT 62.945 6.845 63.115 7.015 ;
      RECT 62.945 10.905 63.115 11.075 ;
      RECT 62.925 4.06 63.095 4.23 ;
      RECT 62.925 8.245 63.095 8.415 ;
      RECT 62.305 2.21 62.475 2.38 ;
      RECT 62.305 3.69 62.475 3.86 ;
      RECT 62.305 8.615 62.475 8.785 ;
      RECT 62.305 10.095 62.475 10.265 ;
      RECT 61.955 1.4 62.125 1.57 ;
      RECT 61.955 5.46 62.125 5.63 ;
      RECT 61.955 6.845 62.125 7.015 ;
      RECT 61.955 10.905 62.125 11.075 ;
      RECT 61.935 4.06 62.105 4.23 ;
      RECT 61.935 8.245 62.105 8.415 ;
      RECT 61.255 1.405 61.425 1.575 ;
      RECT 61.255 5.465 61.425 5.635 ;
      RECT 61.255 6.84 61.425 7.01 ;
      RECT 61.255 10.9 61.425 11.07 ;
      RECT 60.945 3.325 61.115 3.495 ;
      RECT 60.945 8.98 61.115 9.15 ;
      RECT 60.575 1.405 60.745 1.575 ;
      RECT 60.575 10.9 60.745 11.07 ;
      RECT 60.515 2.215 60.685 2.385 ;
      RECT 60.515 2.955 60.685 3.125 ;
      RECT 60.515 9.35 60.685 9.52 ;
      RECT 60.515 10.09 60.685 10.26 ;
      RECT 60.14 3.695 60.31 3.865 ;
      RECT 60.14 8.61 60.31 8.78 ;
      RECT 59.895 1.405 60.065 1.575 ;
      RECT 59.895 10.9 60.065 11.07 ;
      RECT 59.215 1.405 59.385 1.575 ;
      RECT 59.215 10.9 59.385 11.07 ;
      RECT 57.755 2.715 57.925 2.885 ;
      RECT 57.755 5.435 57.925 5.605 ;
      RECT 57.295 2.715 57.465 2.885 ;
      RECT 57.295 5.435 57.465 5.605 ;
      RECT 57.08 4.075 57.25 4.245 ;
      RECT 56.84 3.235 57.01 3.405 ;
      RECT 56.84 4.915 57.01 5.085 ;
      RECT 56.835 2.715 57.005 2.885 ;
      RECT 56.835 5.435 57.005 5.605 ;
      RECT 56.6 3.795 56.77 3.965 ;
      RECT 56.6 4.355 56.77 4.525 ;
      RECT 56.375 2.715 56.545 2.885 ;
      RECT 56.375 5.435 56.545 5.605 ;
      RECT 56.12 4.075 56.29 4.245 ;
      RECT 55.915 2.715 56.085 2.885 ;
      RECT 55.915 5.435 56.085 5.605 ;
      RECT 55.88 3.235 56.05 3.405 ;
      RECT 55.64 3.795 55.81 3.965 ;
      RECT 55.64 6.84 55.81 7.01 ;
      RECT 55.64 10.9 55.81 11.07 ;
      RECT 55.455 2.715 55.625 2.885 ;
      RECT 55.455 5.435 55.625 5.605 ;
      RECT 55.43 4.635 55.6 4.805 ;
      RECT 55.33 8.98 55.5 9.15 ;
      RECT 55.16 4.075 55.33 4.245 ;
      RECT 54.995 2.715 55.165 2.885 ;
      RECT 54.995 5.435 55.165 5.605 ;
      RECT 54.96 10.9 55.13 11.07 ;
      RECT 54.9 9.35 55.07 9.52 ;
      RECT 54.9 10.09 55.07 10.26 ;
      RECT 54.89 4.915 55.06 5.085 ;
      RECT 54.68 3.495 54.85 3.665 ;
      RECT 54.535 2.715 54.705 2.885 ;
      RECT 54.535 5.435 54.705 5.605 ;
      RECT 54.525 8.61 54.695 8.78 ;
      RECT 54.28 10.9 54.45 11.07 ;
      RECT 54.2 4.075 54.37 4.245 ;
      RECT 54.075 2.715 54.245 2.885 ;
      RECT 54.075 5.435 54.245 5.605 ;
      RECT 53.96 3.235 54.13 3.405 ;
      RECT 53.72 3.795 53.89 3.965 ;
      RECT 53.72 4.355 53.89 4.525 ;
      RECT 53.615 2.715 53.785 2.885 ;
      RECT 53.615 5.435 53.785 5.605 ;
      RECT 53.6 10.9 53.77 11.07 ;
      RECT 53.24 3.795 53.41 3.965 ;
      RECT 53.155 2.715 53.325 2.885 ;
      RECT 53.155 5.435 53.325 5.605 ;
      RECT 53 4.915 53.17 5.085 ;
      RECT 52.96 3.235 53.13 3.405 ;
      RECT 52.76 4.075 52.93 4.245 ;
      RECT 52.695 2.715 52.865 2.885 ;
      RECT 52.695 5.435 52.865 5.605 ;
      RECT 52.52 4.915 52.69 5.085 ;
      RECT 52.28 4.355 52.45 4.525 ;
      RECT 52.235 2.715 52.405 2.885 ;
      RECT 52.235 5.435 52.405 5.605 ;
      RECT 51.8 3.795 51.97 3.965 ;
      RECT 51.775 2.715 51.945 2.885 ;
      RECT 51.775 5.435 51.945 5.605 ;
      RECT 51.56 3.235 51.73 3.405 ;
      RECT 51.56 4.915 51.73 5.085 ;
      RECT 51.315 2.715 51.485 2.885 ;
      RECT 51.315 5.435 51.485 5.605 ;
      RECT 51.08 3.235 51.25 3.405 ;
      RECT 51.08 4.355 51.25 4.525 ;
      RECT 50.855 2.715 51.025 2.885 ;
      RECT 50.855 5.435 51.025 5.605 ;
      RECT 50.84 3.795 51.01 3.965 ;
      RECT 50.6 4.635 50.77 4.805 ;
      RECT 50.395 2.715 50.565 2.885 ;
      RECT 50.395 5.435 50.565 5.605 ;
      RECT 50.36 4.075 50.53 4.245 ;
      RECT 49.935 2.715 50.105 2.885 ;
      RECT 49.935 5.435 50.105 5.605 ;
      RECT 49.88 4.075 50.05 4.245 ;
      RECT 49.67 3.235 49.84 3.405 ;
      RECT 49.67 4.635 49.84 4.805 ;
      RECT 49.475 2.715 49.645 2.885 ;
      RECT 49.475 5.435 49.645 5.605 ;
      RECT 48.035 8.615 48.205 8.785 ;
      RECT 48.035 10.095 48.205 10.265 ;
      RECT 47.685 1.4 47.855 1.57 ;
      RECT 47.685 5.46 47.855 5.63 ;
      RECT 47.685 6.845 47.855 7.015 ;
      RECT 47.685 10.905 47.855 11.075 ;
      RECT 47.665 4.06 47.835 4.23 ;
      RECT 47.665 8.245 47.835 8.415 ;
      RECT 47.045 2.21 47.215 2.38 ;
      RECT 47.045 3.69 47.215 3.86 ;
      RECT 47.045 8.615 47.215 8.785 ;
      RECT 47.045 10.095 47.215 10.265 ;
      RECT 46.695 1.4 46.865 1.57 ;
      RECT 46.695 5.46 46.865 5.63 ;
      RECT 46.695 6.845 46.865 7.015 ;
      RECT 46.695 10.905 46.865 11.075 ;
      RECT 46.675 4.06 46.845 4.23 ;
      RECT 46.675 8.245 46.845 8.415 ;
      RECT 45.995 1.405 46.165 1.575 ;
      RECT 45.995 5.465 46.165 5.635 ;
      RECT 45.995 6.84 46.165 7.01 ;
      RECT 45.995 10.9 46.165 11.07 ;
      RECT 45.685 3.325 45.855 3.495 ;
      RECT 45.685 8.98 45.855 9.15 ;
      RECT 45.315 1.405 45.485 1.575 ;
      RECT 45.315 10.9 45.485 11.07 ;
      RECT 45.255 2.215 45.425 2.385 ;
      RECT 45.255 2.955 45.425 3.125 ;
      RECT 45.255 9.35 45.425 9.52 ;
      RECT 45.255 10.09 45.425 10.26 ;
      RECT 44.88 3.695 45.05 3.865 ;
      RECT 44.88 8.61 45.05 8.78 ;
      RECT 44.635 1.405 44.805 1.575 ;
      RECT 44.635 10.9 44.805 11.07 ;
      RECT 43.955 1.405 44.125 1.575 ;
      RECT 43.955 10.9 44.125 11.07 ;
      RECT 42.495 2.715 42.665 2.885 ;
      RECT 42.495 5.435 42.665 5.605 ;
      RECT 42.035 2.715 42.205 2.885 ;
      RECT 42.035 5.435 42.205 5.605 ;
      RECT 41.82 4.075 41.99 4.245 ;
      RECT 41.58 3.235 41.75 3.405 ;
      RECT 41.58 4.915 41.75 5.085 ;
      RECT 41.575 2.715 41.745 2.885 ;
      RECT 41.575 5.435 41.745 5.605 ;
      RECT 41.34 3.795 41.51 3.965 ;
      RECT 41.34 4.355 41.51 4.525 ;
      RECT 41.115 2.715 41.285 2.885 ;
      RECT 41.115 5.435 41.285 5.605 ;
      RECT 40.86 4.075 41.03 4.245 ;
      RECT 40.655 2.715 40.825 2.885 ;
      RECT 40.655 5.435 40.825 5.605 ;
      RECT 40.62 3.235 40.79 3.405 ;
      RECT 40.38 3.795 40.55 3.965 ;
      RECT 40.38 6.84 40.55 7.01 ;
      RECT 40.38 10.9 40.55 11.07 ;
      RECT 40.195 2.715 40.365 2.885 ;
      RECT 40.195 5.435 40.365 5.605 ;
      RECT 40.17 4.635 40.34 4.805 ;
      RECT 40.07 8.98 40.24 9.15 ;
      RECT 39.9 4.075 40.07 4.245 ;
      RECT 39.735 2.715 39.905 2.885 ;
      RECT 39.735 5.435 39.905 5.605 ;
      RECT 39.7 10.9 39.87 11.07 ;
      RECT 39.64 9.35 39.81 9.52 ;
      RECT 39.64 10.09 39.81 10.26 ;
      RECT 39.63 4.915 39.8 5.085 ;
      RECT 39.42 3.495 39.59 3.665 ;
      RECT 39.275 2.715 39.445 2.885 ;
      RECT 39.275 5.435 39.445 5.605 ;
      RECT 39.265 8.61 39.435 8.78 ;
      RECT 39.02 10.9 39.19 11.07 ;
      RECT 38.94 4.075 39.11 4.245 ;
      RECT 38.815 2.715 38.985 2.885 ;
      RECT 38.815 5.435 38.985 5.605 ;
      RECT 38.7 3.235 38.87 3.405 ;
      RECT 38.46 3.795 38.63 3.965 ;
      RECT 38.46 4.355 38.63 4.525 ;
      RECT 38.355 2.715 38.525 2.885 ;
      RECT 38.355 5.435 38.525 5.605 ;
      RECT 38.34 10.9 38.51 11.07 ;
      RECT 37.98 3.795 38.15 3.965 ;
      RECT 37.895 2.715 38.065 2.885 ;
      RECT 37.895 5.435 38.065 5.605 ;
      RECT 37.74 4.915 37.91 5.085 ;
      RECT 37.7 3.235 37.87 3.405 ;
      RECT 37.5 4.075 37.67 4.245 ;
      RECT 37.435 2.715 37.605 2.885 ;
      RECT 37.435 5.435 37.605 5.605 ;
      RECT 37.26 4.915 37.43 5.085 ;
      RECT 37.02 4.355 37.19 4.525 ;
      RECT 36.975 2.715 37.145 2.885 ;
      RECT 36.975 5.435 37.145 5.605 ;
      RECT 36.54 3.795 36.71 3.965 ;
      RECT 36.515 2.715 36.685 2.885 ;
      RECT 36.515 5.435 36.685 5.605 ;
      RECT 36.3 3.235 36.47 3.405 ;
      RECT 36.3 4.915 36.47 5.085 ;
      RECT 36.055 2.715 36.225 2.885 ;
      RECT 36.055 5.435 36.225 5.605 ;
      RECT 35.82 3.235 35.99 3.405 ;
      RECT 35.82 4.355 35.99 4.525 ;
      RECT 35.595 2.715 35.765 2.885 ;
      RECT 35.595 5.435 35.765 5.605 ;
      RECT 35.58 3.795 35.75 3.965 ;
      RECT 35.34 4.635 35.51 4.805 ;
      RECT 35.135 2.715 35.305 2.885 ;
      RECT 35.135 5.435 35.305 5.605 ;
      RECT 35.1 4.075 35.27 4.245 ;
      RECT 34.675 2.715 34.845 2.885 ;
      RECT 34.675 5.435 34.845 5.605 ;
      RECT 34.62 4.075 34.79 4.245 ;
      RECT 34.41 3.235 34.58 3.405 ;
      RECT 34.41 4.635 34.58 4.805 ;
      RECT 34.215 2.715 34.385 2.885 ;
      RECT 34.215 5.435 34.385 5.605 ;
      RECT 32.775 8.615 32.945 8.785 ;
      RECT 32.775 10.095 32.945 10.265 ;
      RECT 32.425 1.4 32.595 1.57 ;
      RECT 32.425 5.46 32.595 5.63 ;
      RECT 32.425 6.845 32.595 7.015 ;
      RECT 32.425 10.905 32.595 11.075 ;
      RECT 32.405 4.06 32.575 4.23 ;
      RECT 32.405 8.245 32.575 8.415 ;
      RECT 31.785 2.21 31.955 2.38 ;
      RECT 31.785 3.69 31.955 3.86 ;
      RECT 31.785 8.615 31.955 8.785 ;
      RECT 31.785 10.095 31.955 10.265 ;
      RECT 31.435 1.4 31.605 1.57 ;
      RECT 31.435 5.46 31.605 5.63 ;
      RECT 31.435 6.845 31.605 7.015 ;
      RECT 31.435 10.905 31.605 11.075 ;
      RECT 31.415 4.06 31.585 4.23 ;
      RECT 31.415 8.245 31.585 8.415 ;
      RECT 30.735 1.405 30.905 1.575 ;
      RECT 30.735 5.465 30.905 5.635 ;
      RECT 30.735 6.84 30.905 7.01 ;
      RECT 30.735 10.9 30.905 11.07 ;
      RECT 30.425 3.325 30.595 3.495 ;
      RECT 30.425 8.98 30.595 9.15 ;
      RECT 30.055 1.405 30.225 1.575 ;
      RECT 30.055 10.9 30.225 11.07 ;
      RECT 29.995 2.215 30.165 2.385 ;
      RECT 29.995 2.955 30.165 3.125 ;
      RECT 29.995 9.35 30.165 9.52 ;
      RECT 29.995 10.09 30.165 10.26 ;
      RECT 29.62 3.695 29.79 3.865 ;
      RECT 29.62 8.61 29.79 8.78 ;
      RECT 29.375 1.405 29.545 1.575 ;
      RECT 29.375 10.9 29.545 11.07 ;
      RECT 28.695 1.405 28.865 1.575 ;
      RECT 28.695 10.9 28.865 11.07 ;
      RECT 27.235 2.715 27.405 2.885 ;
      RECT 27.235 5.435 27.405 5.605 ;
      RECT 26.775 2.715 26.945 2.885 ;
      RECT 26.775 5.435 26.945 5.605 ;
      RECT 26.56 4.075 26.73 4.245 ;
      RECT 26.32 3.235 26.49 3.405 ;
      RECT 26.32 4.915 26.49 5.085 ;
      RECT 26.315 2.715 26.485 2.885 ;
      RECT 26.315 5.435 26.485 5.605 ;
      RECT 26.08 3.795 26.25 3.965 ;
      RECT 26.08 4.355 26.25 4.525 ;
      RECT 25.855 2.715 26.025 2.885 ;
      RECT 25.855 5.435 26.025 5.605 ;
      RECT 25.6 4.075 25.77 4.245 ;
      RECT 25.395 2.715 25.565 2.885 ;
      RECT 25.395 5.435 25.565 5.605 ;
      RECT 25.36 3.235 25.53 3.405 ;
      RECT 25.12 3.795 25.29 3.965 ;
      RECT 25.12 6.84 25.29 7.01 ;
      RECT 25.12 10.9 25.29 11.07 ;
      RECT 24.935 2.715 25.105 2.885 ;
      RECT 24.935 5.435 25.105 5.605 ;
      RECT 24.91 4.635 25.08 4.805 ;
      RECT 24.81 8.98 24.98 9.15 ;
      RECT 24.64 4.075 24.81 4.245 ;
      RECT 24.475 2.715 24.645 2.885 ;
      RECT 24.475 5.435 24.645 5.605 ;
      RECT 24.44 10.9 24.61 11.07 ;
      RECT 24.38 9.35 24.55 9.52 ;
      RECT 24.38 10.09 24.55 10.26 ;
      RECT 24.37 4.915 24.54 5.085 ;
      RECT 24.16 3.495 24.33 3.665 ;
      RECT 24.015 2.715 24.185 2.885 ;
      RECT 24.015 5.435 24.185 5.605 ;
      RECT 24.005 8.61 24.175 8.78 ;
      RECT 23.76 10.9 23.93 11.07 ;
      RECT 23.68 4.075 23.85 4.245 ;
      RECT 23.555 2.715 23.725 2.885 ;
      RECT 23.555 5.435 23.725 5.605 ;
      RECT 23.44 3.235 23.61 3.405 ;
      RECT 23.2 3.795 23.37 3.965 ;
      RECT 23.2 4.355 23.37 4.525 ;
      RECT 23.095 2.715 23.265 2.885 ;
      RECT 23.095 5.435 23.265 5.605 ;
      RECT 23.08 10.9 23.25 11.07 ;
      RECT 22.72 3.795 22.89 3.965 ;
      RECT 22.635 2.715 22.805 2.885 ;
      RECT 22.635 5.435 22.805 5.605 ;
      RECT 22.48 4.915 22.65 5.085 ;
      RECT 22.44 3.235 22.61 3.405 ;
      RECT 22.24 4.075 22.41 4.245 ;
      RECT 22.175 2.715 22.345 2.885 ;
      RECT 22.175 5.435 22.345 5.605 ;
      RECT 22 4.915 22.17 5.085 ;
      RECT 21.76 4.355 21.93 4.525 ;
      RECT 21.715 2.715 21.885 2.885 ;
      RECT 21.715 5.435 21.885 5.605 ;
      RECT 21.28 3.795 21.45 3.965 ;
      RECT 21.255 2.715 21.425 2.885 ;
      RECT 21.255 5.435 21.425 5.605 ;
      RECT 21.04 3.235 21.21 3.405 ;
      RECT 21.04 4.915 21.21 5.085 ;
      RECT 20.795 2.715 20.965 2.885 ;
      RECT 20.795 5.435 20.965 5.605 ;
      RECT 20.56 3.235 20.73 3.405 ;
      RECT 20.56 4.355 20.73 4.525 ;
      RECT 20.335 2.715 20.505 2.885 ;
      RECT 20.335 5.435 20.505 5.605 ;
      RECT 20.32 3.795 20.49 3.965 ;
      RECT 20.08 4.635 20.25 4.805 ;
      RECT 19.875 2.715 20.045 2.885 ;
      RECT 19.875 5.435 20.045 5.605 ;
      RECT 19.84 4.075 20.01 4.245 ;
      RECT 19.415 2.715 19.585 2.885 ;
      RECT 19.415 5.435 19.585 5.605 ;
      RECT 19.36 4.075 19.53 4.245 ;
      RECT 19.15 3.235 19.32 3.405 ;
      RECT 19.15 4.635 19.32 4.805 ;
      RECT 18.955 2.715 19.125 2.885 ;
      RECT 18.955 5.435 19.125 5.605 ;
      RECT 17.515 8.615 17.685 8.785 ;
      RECT 17.515 10.095 17.685 10.265 ;
      RECT 17.165 1.4 17.335 1.57 ;
      RECT 17.165 5.46 17.335 5.63 ;
      RECT 17.165 6.845 17.335 7.015 ;
      RECT 17.165 10.905 17.335 11.075 ;
      RECT 17.145 4.06 17.315 4.23 ;
      RECT 17.145 8.245 17.315 8.415 ;
      RECT 16.525 2.21 16.695 2.38 ;
      RECT 16.525 3.69 16.695 3.86 ;
      RECT 16.525 8.615 16.695 8.785 ;
      RECT 16.525 10.095 16.695 10.265 ;
      RECT 16.175 1.4 16.345 1.57 ;
      RECT 16.175 5.46 16.345 5.63 ;
      RECT 16.175 6.845 16.345 7.015 ;
      RECT 16.175 10.905 16.345 11.075 ;
      RECT 16.155 4.06 16.325 4.23 ;
      RECT 16.155 8.245 16.325 8.415 ;
      RECT 15.475 1.405 15.645 1.575 ;
      RECT 15.475 5.465 15.645 5.635 ;
      RECT 15.475 6.84 15.645 7.01 ;
      RECT 15.475 10.9 15.645 11.07 ;
      RECT 15.165 3.325 15.335 3.495 ;
      RECT 15.165 8.98 15.335 9.15 ;
      RECT 14.795 1.405 14.965 1.575 ;
      RECT 14.795 10.9 14.965 11.07 ;
      RECT 14.735 2.215 14.905 2.385 ;
      RECT 14.735 2.955 14.905 3.125 ;
      RECT 14.735 9.35 14.905 9.52 ;
      RECT 14.735 10.09 14.905 10.26 ;
      RECT 14.36 3.695 14.53 3.865 ;
      RECT 14.36 8.61 14.53 8.78 ;
      RECT 14.115 1.405 14.285 1.575 ;
      RECT 14.115 10.9 14.285 11.07 ;
      RECT 13.435 1.405 13.605 1.575 ;
      RECT 13.435 10.9 13.605 11.07 ;
      RECT 11.975 2.715 12.145 2.885 ;
      RECT 11.975 5.435 12.145 5.605 ;
      RECT 11.515 2.715 11.685 2.885 ;
      RECT 11.515 5.435 11.685 5.605 ;
      RECT 11.3 4.075 11.47 4.245 ;
      RECT 11.06 3.235 11.23 3.405 ;
      RECT 11.06 4.915 11.23 5.085 ;
      RECT 11.055 2.715 11.225 2.885 ;
      RECT 11.055 5.435 11.225 5.605 ;
      RECT 10.82 3.795 10.99 3.965 ;
      RECT 10.82 4.355 10.99 4.525 ;
      RECT 10.595 2.715 10.765 2.885 ;
      RECT 10.595 5.435 10.765 5.605 ;
      RECT 10.34 4.075 10.51 4.245 ;
      RECT 10.135 2.715 10.305 2.885 ;
      RECT 10.135 5.435 10.305 5.605 ;
      RECT 10.1 3.235 10.27 3.405 ;
      RECT 9.86 3.795 10.03 3.965 ;
      RECT 9.86 6.84 10.03 7.01 ;
      RECT 9.86 10.9 10.03 11.07 ;
      RECT 9.675 2.715 9.845 2.885 ;
      RECT 9.675 5.435 9.845 5.605 ;
      RECT 9.65 4.635 9.82 4.805 ;
      RECT 9.55 8.98 9.72 9.15 ;
      RECT 9.38 4.075 9.55 4.245 ;
      RECT 9.215 2.715 9.385 2.885 ;
      RECT 9.215 5.435 9.385 5.605 ;
      RECT 9.18 10.9 9.35 11.07 ;
      RECT 9.12 9.35 9.29 9.52 ;
      RECT 9.12 10.09 9.29 10.26 ;
      RECT 9.11 4.915 9.28 5.085 ;
      RECT 8.9 3.495 9.07 3.665 ;
      RECT 8.755 2.715 8.925 2.885 ;
      RECT 8.755 5.435 8.925 5.605 ;
      RECT 8.745 8.61 8.915 8.78 ;
      RECT 8.5 10.9 8.67 11.07 ;
      RECT 8.42 4.075 8.59 4.245 ;
      RECT 8.295 2.715 8.465 2.885 ;
      RECT 8.295 5.435 8.465 5.605 ;
      RECT 8.18 3.235 8.35 3.405 ;
      RECT 7.94 3.795 8.11 3.965 ;
      RECT 7.94 4.355 8.11 4.525 ;
      RECT 7.835 2.715 8.005 2.885 ;
      RECT 7.835 5.435 8.005 5.605 ;
      RECT 7.82 10.9 7.99 11.07 ;
      RECT 7.46 3.795 7.63 3.965 ;
      RECT 7.375 2.715 7.545 2.885 ;
      RECT 7.375 5.435 7.545 5.605 ;
      RECT 7.22 4.915 7.39 5.085 ;
      RECT 7.18 3.235 7.35 3.405 ;
      RECT 6.98 4.075 7.15 4.245 ;
      RECT 6.915 2.715 7.085 2.885 ;
      RECT 6.915 5.435 7.085 5.605 ;
      RECT 6.74 4.915 6.91 5.085 ;
      RECT 6.5 4.355 6.67 4.525 ;
      RECT 6.455 2.715 6.625 2.885 ;
      RECT 6.455 5.435 6.625 5.605 ;
      RECT 6.02 3.795 6.19 3.965 ;
      RECT 5.995 2.715 6.165 2.885 ;
      RECT 5.995 5.435 6.165 5.605 ;
      RECT 5.78 3.235 5.95 3.405 ;
      RECT 5.78 4.915 5.95 5.085 ;
      RECT 5.535 2.715 5.705 2.885 ;
      RECT 5.535 5.435 5.705 5.605 ;
      RECT 5.3 3.235 5.47 3.405 ;
      RECT 5.3 4.355 5.47 4.525 ;
      RECT 5.075 2.715 5.245 2.885 ;
      RECT 5.075 5.435 5.245 5.605 ;
      RECT 5.06 3.795 5.23 3.965 ;
      RECT 4.82 4.635 4.99 4.805 ;
      RECT 4.615 2.715 4.785 2.885 ;
      RECT 4.615 5.435 4.785 5.605 ;
      RECT 4.58 4.075 4.75 4.245 ;
      RECT 4.155 2.715 4.325 2.885 ;
      RECT 4.155 5.435 4.325 5.605 ;
      RECT 4.1 4.075 4.27 4.245 ;
      RECT 3.89 3.235 4.06 3.405 ;
      RECT 3.89 4.635 4.06 4.805 ;
      RECT 3.695 2.715 3.865 2.885 ;
      RECT 3.695 5.435 3.865 5.605 ;
      RECT 2.345 6.84 2.515 7.01 ;
      RECT 2.345 10.9 2.515 11.07 ;
      RECT 2.035 8.98 2.205 9.15 ;
      RECT 1.665 10.9 1.835 11.07 ;
      RECT 1.605 9.35 1.775 9.52 ;
      RECT 1.605 10.09 1.775 10.26 ;
      RECT 1.23 8.61 1.4 8.78 ;
      RECT 0.985 10.9 1.155 11.07 ;
      RECT 0.305 10.9 0.475 11.07 ;
    LAYER li1 ;
      RECT 72.56 0.005 72.73 3.385 ;
      RECT 71.62 0.005 71.79 3.385 ;
      RECT 70.66 0.005 70.83 3.385 ;
      RECT 68.74 0.005 68.91 3.385 ;
      RECT 67.78 0.005 67.95 3.385 ;
      RECT 65.86 0.005 66.03 3.385 ;
      RECT 57.3 0.005 57.47 3.385 ;
      RECT 56.36 0.005 56.53 3.385 ;
      RECT 55.4 0.005 55.57 3.385 ;
      RECT 53.48 0.005 53.65 3.385 ;
      RECT 52.52 0.005 52.69 3.385 ;
      RECT 50.6 0.005 50.77 3.385 ;
      RECT 42.04 0.005 42.21 3.385 ;
      RECT 41.1 0.005 41.27 3.385 ;
      RECT 40.14 0.005 40.31 3.385 ;
      RECT 38.22 0.005 38.39 3.385 ;
      RECT 37.26 0.005 37.43 3.385 ;
      RECT 35.34 0.005 35.51 3.385 ;
      RECT 26.78 0.005 26.95 3.385 ;
      RECT 25.84 0.005 26.01 3.385 ;
      RECT 24.88 0.005 25.05 3.385 ;
      RECT 22.96 0.005 23.13 3.385 ;
      RECT 22 0.005 22.17 3.385 ;
      RECT 20.08 0.005 20.25 3.385 ;
      RECT 11.52 0 11.69 3.385 ;
      RECT 10.58 0 10.75 3.385 ;
      RECT 9.62 0 9.79 3.385 ;
      RECT 7.7 0 7.87 3.385 ;
      RECT 6.74 0 6.91 3.385 ;
      RECT 4.82 0 4.99 3.385 ;
      RECT 69.615 0.005 69.81 2.895 ;
      RECT 65.86 0.005 66.135 2.895 ;
      RECT 54.355 0.005 54.55 2.895 ;
      RECT 50.6 0.005 50.875 2.895 ;
      RECT 39.095 0.005 39.29 2.895 ;
      RECT 35.34 0.005 35.615 2.895 ;
      RECT 23.835 0.005 24.03 2.895 ;
      RECT 20.08 0.005 20.355 2.895 ;
      RECT 8.575 0 8.77 2.895 ;
      RECT 4.82 0 5.095 2.895 ;
      RECT 64.59 0.005 73.33 2.885 ;
      RECT 49.33 0.005 58.07 2.885 ;
      RECT 34.07 0.005 42.81 2.885 ;
      RECT 18.81 0.005 27.55 2.885 ;
      RECT 3.55 0 12.29 2.885 ;
      RECT 74.395 0.005 74.565 2.235 ;
      RECT 59.135 0.005 59.305 2.235 ;
      RECT 43.875 0.005 44.045 2.235 ;
      RECT 28.615 0.005 28.785 2.235 ;
      RECT 13.355 0.005 13.525 2.235 ;
      RECT 78.125 0.005 78.295 2.23 ;
      RECT 77.135 0.005 77.305 2.23 ;
      RECT 62.865 0.005 63.035 2.23 ;
      RECT 61.875 0.005 62.045 2.23 ;
      RECT 47.605 0.005 47.775 2.23 ;
      RECT 46.615 0.005 46.785 2.23 ;
      RECT 32.345 0.005 32.515 2.23 ;
      RECT 31.355 0.005 31.525 2.23 ;
      RECT 17.085 0.005 17.255 2.23 ;
      RECT 16.095 0.005 16.265 2.23 ;
      RECT 2.8 0.005 79.1 1.605 ;
      RECT 0 0 13.43 1.6 ;
      RECT 2.035 5.44 2.205 10.6 ;
      RECT 78.125 4.7 78.295 7.775 ;
      RECT 77.135 4.7 77.305 7.775 ;
      RECT 62.865 4.7 63.035 7.775 ;
      RECT 61.875 4.7 62.045 7.775 ;
      RECT 47.605 4.7 47.775 7.775 ;
      RECT 46.615 4.7 46.785 7.775 ;
      RECT 32.345 4.7 32.515 7.775 ;
      RECT 31.355 4.7 31.525 7.775 ;
      RECT 17.085 4.7 17.255 7.775 ;
      RECT 16.095 4.7 16.265 7.775 ;
      RECT 74.395 4.705 74.565 7.77 ;
      RECT 68.78 5.435 68.95 7.77 ;
      RECT 59.135 4.705 59.305 7.77 ;
      RECT 53.52 5.435 53.69 7.77 ;
      RECT 43.875 4.705 44.045 7.77 ;
      RECT 38.26 5.435 38.43 7.77 ;
      RECT 28.615 4.705 28.785 7.77 ;
      RECT 23 5.435 23.17 7.77 ;
      RECT 13.355 4.705 13.525 7.77 ;
      RECT 7.74 5.435 7.91 7.77 ;
      RECT 0.225 5.44 0.395 7.77 ;
      RECT 76.965 5.43 78.945 7.045 ;
      RECT 61.705 5.43 63.685 7.045 ;
      RECT 46.445 5.43 48.425 7.045 ;
      RECT 31.185 5.43 33.165 7.045 ;
      RECT 15.925 5.43 17.905 7.045 ;
      RECT 0.005 5.44 79.1 7.04 ;
      RECT 64.59 5.435 79.1 7.04 ;
      RECT 49.33 5.435 63.84 7.04 ;
      RECT 34.07 5.435 48.58 7.04 ;
      RECT 18.81 5.435 33.32 7.04 ;
      RECT 3.55 5.435 18.06 7.04 ;
      RECT 71.62 4.935 71.79 7.04 ;
      RECT 69.7 4.935 69.87 7.04 ;
      RECT 68.76 4.935 68.93 7.04 ;
      RECT 67.3 4.935 67.47 7.04 ;
      RECT 65.38 4.935 65.55 7.04 ;
      RECT 56.36 4.935 56.53 7.04 ;
      RECT 54.44 4.935 54.61 7.04 ;
      RECT 53.5 4.935 53.67 7.04 ;
      RECT 52.04 4.935 52.21 7.04 ;
      RECT 50.12 4.935 50.29 7.04 ;
      RECT 41.1 4.935 41.27 7.04 ;
      RECT 39.18 4.935 39.35 7.04 ;
      RECT 38.24 4.935 38.41 7.04 ;
      RECT 36.78 4.935 36.95 7.04 ;
      RECT 34.86 4.935 35.03 7.04 ;
      RECT 25.84 4.935 26.01 7.04 ;
      RECT 23.92 4.935 24.09 7.04 ;
      RECT 22.98 4.935 23.15 7.04 ;
      RECT 21.52 4.935 21.69 7.04 ;
      RECT 19.6 4.935 19.77 7.04 ;
      RECT 10.58 4.935 10.75 7.04 ;
      RECT 8.66 4.935 8.83 7.04 ;
      RECT 7.72 4.935 7.89 7.04 ;
      RECT 6.26 4.935 6.43 7.04 ;
      RECT 4.34 4.935 4.51 7.04 ;
      RECT 0.005 10.87 79.1 12.47 ;
      RECT 78.125 10.245 78.295 12.47 ;
      RECT 77.135 10.245 77.305 12.47 ;
      RECT 74.395 10.24 74.565 12.47 ;
      RECT 68.78 10.24 68.95 12.47 ;
      RECT 62.865 10.245 63.035 12.47 ;
      RECT 61.875 10.245 62.045 12.47 ;
      RECT 59.135 10.24 59.305 12.47 ;
      RECT 53.52 10.24 53.69 12.47 ;
      RECT 47.605 10.245 47.775 12.47 ;
      RECT 46.615 10.245 46.785 12.47 ;
      RECT 43.875 10.24 44.045 12.47 ;
      RECT 38.26 10.24 38.43 12.47 ;
      RECT 32.345 10.245 32.515 12.47 ;
      RECT 31.355 10.245 31.525 12.47 ;
      RECT 28.615 10.24 28.785 12.47 ;
      RECT 23 10.24 23.17 12.47 ;
      RECT 17.085 10.245 17.255 12.47 ;
      RECT 16.095 10.245 16.265 12.47 ;
      RECT 13.355 10.24 13.525 12.47 ;
      RECT 7.74 10.24 7.91 12.47 ;
      RECT 0.01 10.86 0.815 12.47 ;
      RECT 0.225 10.84 0.475 12.47 ;
      RECT 0.225 10.24 0.395 12.47 ;
      RECT 78.185 3.04 78.355 4.23 ;
      RECT 78.185 3.04 78.655 3.21 ;
      RECT 78.185 9.265 78.655 9.435 ;
      RECT 78.185 8.245 78.355 9.435 ;
      RECT 77.195 3.04 77.365 4.23 ;
      RECT 77.195 3.04 77.665 3.21 ;
      RECT 77.195 9.265 77.665 9.435 ;
      RECT 77.195 8.245 77.365 9.435 ;
      RECT 75.345 3.935 75.515 5.165 ;
      RECT 75.4 2.155 75.57 4.105 ;
      RECT 75.345 1.875 75.515 2.325 ;
      RECT 75.345 10.15 75.515 10.6 ;
      RECT 75.4 8.37 75.57 10.32 ;
      RECT 75.345 7.31 75.515 8.54 ;
      RECT 74.825 1.875 74.995 5.165 ;
      RECT 74.825 3.375 75.23 3.705 ;
      RECT 74.825 2.535 75.23 2.865 ;
      RECT 74.825 7.31 74.995 10.6 ;
      RECT 74.825 9.61 75.23 9.94 ;
      RECT 74.825 8.77 75.23 9.1 ;
      RECT 72.1 4.915 72.615 5.085 ;
      RECT 72.445 4.525 72.615 5.085 ;
      RECT 72.55 4.445 72.72 4.775 ;
      RECT 72.34 3.835 72.615 4.245 ;
      RECT 72.22 3.835 72.615 4.045 ;
      RECT 70.69 4.445 70.86 4.805 ;
      RECT 70.69 4.525 72.03 4.695 ;
      RECT 71.86 4.355 72.03 4.695 ;
      RECT 70.42 3.875 70.59 4.245 ;
      RECT 69.94 3.875 70.59 4.145 ;
      RECT 69.86 3.875 70.67 4.045 ;
      RECT 69.22 3.115 69.39 3.405 ;
      RECT 69.22 3.115 70.46 3.285 ;
      RECT 69.94 3.455 70.11 3.665 ;
      RECT 69.58 3.455 70.11 3.625 ;
      RECT 69.73 10.15 69.9 10.6 ;
      RECT 69.785 8.37 69.955 10.32 ;
      RECT 69.73 7.31 69.9 8.54 ;
      RECT 69.21 7.31 69.38 10.6 ;
      RECT 69.21 9.61 69.615 9.94 ;
      RECT 69.21 8.77 69.615 9.1 ;
      RECT 68.98 4.525 69.47 4.695 ;
      RECT 68.98 4.355 69.15 4.695 ;
      RECT 68.26 4.525 68.43 5.085 ;
      RECT 68.15 4.525 68.48 4.695 ;
      RECT 68.22 3.135 68.39 3.405 ;
      RECT 68.26 3.055 68.43 3.385 ;
      RECT 68.125 3.135 68.43 3.355 ;
      RECT 66.7 4.525 66.99 5.085 ;
      RECT 66.82 4.445 66.99 5.085 ;
      RECT 66.46 3.875 66.83 4.045 ;
      RECT 66.46 3.235 66.63 4.045 ;
      RECT 66.34 3.235 66.63 3.405 ;
      RECT 64.77 3.23 65.34 3.69 ;
      RECT 64.93 3.055 65.1 3.69 ;
      RECT 62.925 3.04 63.095 4.23 ;
      RECT 62.925 3.04 63.395 3.21 ;
      RECT 62.925 9.265 63.395 9.435 ;
      RECT 62.925 8.245 63.095 9.435 ;
      RECT 61.935 3.04 62.105 4.23 ;
      RECT 61.935 3.04 62.405 3.21 ;
      RECT 61.935 9.265 62.405 9.435 ;
      RECT 61.935 8.245 62.105 9.435 ;
      RECT 60.085 3.935 60.255 5.165 ;
      RECT 60.14 2.155 60.31 4.105 ;
      RECT 60.085 1.875 60.255 2.325 ;
      RECT 60.085 10.15 60.255 10.6 ;
      RECT 60.14 8.37 60.31 10.32 ;
      RECT 60.085 7.31 60.255 8.54 ;
      RECT 59.565 1.875 59.735 5.165 ;
      RECT 59.565 3.375 59.97 3.705 ;
      RECT 59.565 2.535 59.97 2.865 ;
      RECT 59.565 7.31 59.735 10.6 ;
      RECT 59.565 9.61 59.97 9.94 ;
      RECT 59.565 8.77 59.97 9.1 ;
      RECT 56.84 4.915 57.355 5.085 ;
      RECT 57.185 4.525 57.355 5.085 ;
      RECT 57.29 4.445 57.46 4.775 ;
      RECT 57.08 3.835 57.355 4.245 ;
      RECT 56.96 3.835 57.355 4.045 ;
      RECT 55.43 4.445 55.6 4.805 ;
      RECT 55.43 4.525 56.77 4.695 ;
      RECT 56.6 4.355 56.77 4.695 ;
      RECT 55.16 3.875 55.33 4.245 ;
      RECT 54.68 3.875 55.33 4.145 ;
      RECT 54.6 3.875 55.41 4.045 ;
      RECT 53.96 3.115 54.13 3.405 ;
      RECT 53.96 3.115 55.2 3.285 ;
      RECT 54.68 3.455 54.85 3.665 ;
      RECT 54.32 3.455 54.85 3.625 ;
      RECT 54.47 10.15 54.64 10.6 ;
      RECT 54.525 8.37 54.695 10.32 ;
      RECT 54.47 7.31 54.64 8.54 ;
      RECT 53.95 7.31 54.12 10.6 ;
      RECT 53.95 9.61 54.355 9.94 ;
      RECT 53.95 8.77 54.355 9.1 ;
      RECT 53.72 4.525 54.21 4.695 ;
      RECT 53.72 4.355 53.89 4.695 ;
      RECT 53 4.525 53.17 5.085 ;
      RECT 52.89 4.525 53.22 4.695 ;
      RECT 52.96 3.135 53.13 3.405 ;
      RECT 53 3.055 53.17 3.385 ;
      RECT 52.865 3.135 53.17 3.355 ;
      RECT 51.44 4.525 51.73 5.085 ;
      RECT 51.56 4.445 51.73 5.085 ;
      RECT 51.2 3.875 51.57 4.045 ;
      RECT 51.2 3.235 51.37 4.045 ;
      RECT 51.08 3.235 51.37 3.405 ;
      RECT 47.665 3.04 47.835 4.23 ;
      RECT 47.665 3.04 48.135 3.21 ;
      RECT 47.665 9.265 48.135 9.435 ;
      RECT 47.665 8.245 47.835 9.435 ;
      RECT 46.675 3.04 46.845 4.23 ;
      RECT 46.675 3.04 47.145 3.21 ;
      RECT 46.675 9.265 47.145 9.435 ;
      RECT 46.675 8.245 46.845 9.435 ;
      RECT 44.825 3.935 44.995 5.165 ;
      RECT 44.88 2.155 45.05 4.105 ;
      RECT 44.825 1.875 44.995 2.325 ;
      RECT 44.825 10.15 44.995 10.6 ;
      RECT 44.88 8.37 45.05 10.32 ;
      RECT 44.825 7.31 44.995 8.54 ;
      RECT 44.305 1.875 44.475 5.165 ;
      RECT 44.305 3.375 44.71 3.705 ;
      RECT 44.305 2.535 44.71 2.865 ;
      RECT 44.305 7.31 44.475 10.6 ;
      RECT 44.305 9.61 44.71 9.94 ;
      RECT 44.305 8.77 44.71 9.1 ;
      RECT 41.58 4.915 42.095 5.085 ;
      RECT 41.925 4.525 42.095 5.085 ;
      RECT 42.03 4.445 42.2 4.775 ;
      RECT 41.82 3.835 42.095 4.245 ;
      RECT 41.7 3.835 42.095 4.045 ;
      RECT 40.17 4.445 40.34 4.805 ;
      RECT 40.17 4.525 41.51 4.695 ;
      RECT 41.34 4.355 41.51 4.695 ;
      RECT 39.9 3.875 40.07 4.245 ;
      RECT 39.42 3.875 40.07 4.145 ;
      RECT 39.34 3.875 40.15 4.045 ;
      RECT 38.7 3.115 38.87 3.405 ;
      RECT 38.7 3.115 39.94 3.285 ;
      RECT 39.42 3.455 39.59 3.665 ;
      RECT 39.06 3.455 39.59 3.625 ;
      RECT 39.21 10.15 39.38 10.6 ;
      RECT 39.265 8.37 39.435 10.32 ;
      RECT 39.21 7.31 39.38 8.54 ;
      RECT 38.69 7.31 38.86 10.6 ;
      RECT 38.69 9.61 39.095 9.94 ;
      RECT 38.69 8.77 39.095 9.1 ;
      RECT 38.46 4.525 38.95 4.695 ;
      RECT 38.46 4.355 38.63 4.695 ;
      RECT 37.74 4.525 37.91 5.085 ;
      RECT 37.63 4.525 37.96 4.695 ;
      RECT 37.7 3.135 37.87 3.405 ;
      RECT 37.74 3.055 37.91 3.385 ;
      RECT 37.605 3.135 37.91 3.355 ;
      RECT 36.18 4.525 36.47 5.085 ;
      RECT 36.3 4.445 36.47 5.085 ;
      RECT 35.94 3.875 36.31 4.045 ;
      RECT 35.94 3.235 36.11 4.045 ;
      RECT 35.82 3.235 36.11 3.405 ;
      RECT 32.405 3.04 32.575 4.23 ;
      RECT 32.405 3.04 32.875 3.21 ;
      RECT 32.405 9.265 32.875 9.435 ;
      RECT 32.405 8.245 32.575 9.435 ;
      RECT 31.415 3.04 31.585 4.23 ;
      RECT 31.415 3.04 31.885 3.21 ;
      RECT 31.415 9.265 31.885 9.435 ;
      RECT 31.415 8.245 31.585 9.435 ;
      RECT 29.565 3.935 29.735 5.165 ;
      RECT 29.62 2.155 29.79 4.105 ;
      RECT 29.565 1.875 29.735 2.325 ;
      RECT 29.565 10.15 29.735 10.6 ;
      RECT 29.62 8.37 29.79 10.32 ;
      RECT 29.565 7.31 29.735 8.54 ;
      RECT 29.045 1.875 29.215 5.165 ;
      RECT 29.045 3.375 29.45 3.705 ;
      RECT 29.045 2.535 29.45 2.865 ;
      RECT 29.045 7.31 29.215 10.6 ;
      RECT 29.045 9.61 29.45 9.94 ;
      RECT 29.045 8.77 29.45 9.1 ;
      RECT 26.32 4.915 26.835 5.085 ;
      RECT 26.665 4.525 26.835 5.085 ;
      RECT 26.77 4.445 26.94 4.775 ;
      RECT 26.56 3.835 26.835 4.245 ;
      RECT 26.44 3.835 26.835 4.045 ;
      RECT 24.91 4.445 25.08 4.805 ;
      RECT 24.91 4.525 26.25 4.695 ;
      RECT 26.08 4.355 26.25 4.695 ;
      RECT 24.64 3.875 24.81 4.245 ;
      RECT 24.16 3.875 24.81 4.145 ;
      RECT 24.08 3.875 24.89 4.045 ;
      RECT 23.44 3.115 23.61 3.405 ;
      RECT 23.44 3.115 24.68 3.285 ;
      RECT 24.16 3.455 24.33 3.665 ;
      RECT 23.8 3.455 24.33 3.625 ;
      RECT 23.95 10.15 24.12 10.6 ;
      RECT 24.005 8.37 24.175 10.32 ;
      RECT 23.95 7.31 24.12 8.54 ;
      RECT 23.43 7.31 23.6 10.6 ;
      RECT 23.43 9.61 23.835 9.94 ;
      RECT 23.43 8.77 23.835 9.1 ;
      RECT 23.2 4.525 23.69 4.695 ;
      RECT 23.2 4.355 23.37 4.695 ;
      RECT 22.48 4.525 22.65 5.085 ;
      RECT 22.37 4.525 22.7 4.695 ;
      RECT 22.44 3.135 22.61 3.405 ;
      RECT 22.48 3.055 22.65 3.385 ;
      RECT 22.345 3.135 22.65 3.355 ;
      RECT 20.92 4.525 21.21 5.085 ;
      RECT 21.04 4.445 21.21 5.085 ;
      RECT 20.68 3.875 21.05 4.045 ;
      RECT 20.68 3.235 20.85 4.045 ;
      RECT 20.56 3.235 20.85 3.405 ;
      RECT 17.145 3.04 17.315 4.23 ;
      RECT 17.145 3.04 17.615 3.21 ;
      RECT 17.145 9.265 17.615 9.435 ;
      RECT 17.145 8.245 17.315 9.435 ;
      RECT 16.155 3.04 16.325 4.23 ;
      RECT 16.155 3.04 16.625 3.21 ;
      RECT 16.155 9.265 16.625 9.435 ;
      RECT 16.155 8.245 16.325 9.435 ;
      RECT 14.305 3.935 14.475 5.165 ;
      RECT 14.36 2.155 14.53 4.105 ;
      RECT 14.305 1.875 14.475 2.325 ;
      RECT 14.305 10.15 14.475 10.6 ;
      RECT 14.36 8.37 14.53 10.32 ;
      RECT 14.305 7.31 14.475 8.54 ;
      RECT 13.785 1.875 13.955 5.165 ;
      RECT 13.785 3.375 14.19 3.705 ;
      RECT 13.785 2.535 14.19 2.865 ;
      RECT 13.785 7.31 13.955 10.6 ;
      RECT 13.785 9.61 14.19 9.94 ;
      RECT 13.785 8.77 14.19 9.1 ;
      RECT 11.06 4.915 11.575 5.085 ;
      RECT 11.405 4.525 11.575 5.085 ;
      RECT 11.51 4.445 11.68 4.775 ;
      RECT 11.3 3.835 11.575 4.245 ;
      RECT 11.18 3.835 11.575 4.045 ;
      RECT 9.65 4.445 9.82 4.805 ;
      RECT 9.65 4.525 10.99 4.695 ;
      RECT 10.82 4.355 10.99 4.695 ;
      RECT 9.38 3.875 9.55 4.245 ;
      RECT 8.9 3.875 9.55 4.145 ;
      RECT 8.82 3.875 9.63 4.045 ;
      RECT 8.18 3.115 8.35 3.405 ;
      RECT 8.18 3.115 9.42 3.285 ;
      RECT 8.9 3.455 9.07 3.665 ;
      RECT 8.54 3.455 9.07 3.625 ;
      RECT 8.69 10.15 8.86 10.6 ;
      RECT 8.745 8.37 8.915 10.32 ;
      RECT 8.69 7.31 8.86 8.54 ;
      RECT 8.17 7.31 8.34 10.6 ;
      RECT 8.17 9.61 8.575 9.94 ;
      RECT 8.17 8.77 8.575 9.1 ;
      RECT 7.94 4.525 8.43 4.695 ;
      RECT 7.94 4.355 8.11 4.695 ;
      RECT 7.22 4.525 7.39 5.085 ;
      RECT 7.11 4.525 7.44 4.695 ;
      RECT 7.18 3.135 7.35 3.405 ;
      RECT 7.22 3.055 7.39 3.385 ;
      RECT 7.085 3.135 7.39 3.355 ;
      RECT 5.66 4.525 5.95 5.085 ;
      RECT 5.78 4.445 5.95 5.085 ;
      RECT 5.42 3.875 5.79 4.045 ;
      RECT 5.42 3.235 5.59 4.045 ;
      RECT 5.3 3.235 5.59 3.405 ;
      RECT 1.175 10.15 1.345 10.6 ;
      RECT 1.23 8.37 1.4 10.32 ;
      RECT 1.175 7.31 1.345 8.54 ;
      RECT 0.655 7.31 0.825 10.6 ;
      RECT 0.655 9.61 1.06 9.94 ;
      RECT 0.655 8.77 1.06 9.1 ;
      RECT 78.555 7.315 78.725 8.785 ;
      RECT 78.555 10.095 78.725 10.605 ;
      RECT 77.565 1.87 77.735 2.38 ;
      RECT 77.565 3.69 77.735 5.16 ;
      RECT 77.565 7.315 77.735 8.785 ;
      RECT 77.565 10.095 77.735 10.605 ;
      RECT 76.205 1.875 76.375 5.165 ;
      RECT 76.205 7.31 76.375 10.6 ;
      RECT 75.775 1.875 75.945 2.385 ;
      RECT 75.775 2.955 75.945 5.165 ;
      RECT 75.775 7.31 75.945 9.52 ;
      RECT 75.775 10.09 75.945 10.6 ;
      RECT 72.1 3.055 72.27 3.405 ;
      RECT 71.86 3.795 72.03 4.125 ;
      RECT 71.38 3.795 71.55 4.245 ;
      RECT 71.14 3.055 71.31 3.405 ;
      RECT 70.9 3.795 71.07 4.125 ;
      RECT 70.59 7.31 70.76 10.6 ;
      RECT 70.16 7.31 70.33 9.52 ;
      RECT 70.16 10.09 70.33 10.6 ;
      RECT 70.15 4.785 70.32 5.115 ;
      RECT 69.46 3.795 69.63 4.245 ;
      RECT 68.98 3.795 69.15 4.125 ;
      RECT 68.5 3.795 68.67 4.125 ;
      RECT 68.02 3.795 68.19 4.245 ;
      RECT 67.78 4.785 67.95 5.115 ;
      RECT 67.54 3.795 67.71 4.525 ;
      RECT 67.06 3.795 67.23 4.125 ;
      RECT 66.82 3.055 66.99 3.405 ;
      RECT 66.34 4.355 66.51 4.775 ;
      RECT 66.1 3.795 66.27 4.125 ;
      RECT 65.86 4.445 66.03 4.805 ;
      RECT 65.62 3.795 65.79 4.245 ;
      RECT 65.14 3.795 65.31 4.245 ;
      RECT 64.93 4.445 65.1 4.805 ;
      RECT 63.295 7.315 63.465 8.785 ;
      RECT 63.295 10.095 63.465 10.605 ;
      RECT 62.305 1.87 62.475 2.38 ;
      RECT 62.305 3.69 62.475 5.16 ;
      RECT 62.305 7.315 62.475 8.785 ;
      RECT 62.305 10.095 62.475 10.605 ;
      RECT 60.945 1.875 61.115 5.165 ;
      RECT 60.945 7.31 61.115 10.6 ;
      RECT 60.515 1.875 60.685 2.385 ;
      RECT 60.515 2.955 60.685 5.165 ;
      RECT 60.515 7.31 60.685 9.52 ;
      RECT 60.515 10.09 60.685 10.6 ;
      RECT 56.84 3.055 57.01 3.405 ;
      RECT 56.6 3.795 56.77 4.125 ;
      RECT 56.12 3.795 56.29 4.245 ;
      RECT 55.88 3.055 56.05 3.405 ;
      RECT 55.64 3.795 55.81 4.125 ;
      RECT 55.33 7.31 55.5 10.6 ;
      RECT 54.9 7.31 55.07 9.52 ;
      RECT 54.9 10.09 55.07 10.6 ;
      RECT 54.89 4.785 55.06 5.115 ;
      RECT 54.2 3.795 54.37 4.245 ;
      RECT 53.72 3.795 53.89 4.125 ;
      RECT 53.24 3.795 53.41 4.125 ;
      RECT 52.76 3.795 52.93 4.245 ;
      RECT 52.52 4.785 52.69 5.115 ;
      RECT 52.28 3.795 52.45 4.525 ;
      RECT 51.8 3.795 51.97 4.125 ;
      RECT 51.56 3.055 51.73 3.405 ;
      RECT 51.08 4.355 51.25 4.775 ;
      RECT 50.84 3.795 51.01 4.125 ;
      RECT 50.6 4.445 50.77 4.805 ;
      RECT 50.36 3.795 50.53 4.245 ;
      RECT 49.88 3.795 50.05 4.245 ;
      RECT 49.67 3.055 49.84 3.405 ;
      RECT 49.67 4.445 49.84 4.805 ;
      RECT 48.035 7.315 48.205 8.785 ;
      RECT 48.035 10.095 48.205 10.605 ;
      RECT 47.045 1.87 47.215 2.38 ;
      RECT 47.045 3.69 47.215 5.16 ;
      RECT 47.045 7.315 47.215 8.785 ;
      RECT 47.045 10.095 47.215 10.605 ;
      RECT 45.685 1.875 45.855 5.165 ;
      RECT 45.685 7.31 45.855 10.6 ;
      RECT 45.255 1.875 45.425 2.385 ;
      RECT 45.255 2.955 45.425 5.165 ;
      RECT 45.255 7.31 45.425 9.52 ;
      RECT 45.255 10.09 45.425 10.6 ;
      RECT 41.58 3.055 41.75 3.405 ;
      RECT 41.34 3.795 41.51 4.125 ;
      RECT 40.86 3.795 41.03 4.245 ;
      RECT 40.62 3.055 40.79 3.405 ;
      RECT 40.38 3.795 40.55 4.125 ;
      RECT 40.07 7.31 40.24 10.6 ;
      RECT 39.64 7.31 39.81 9.52 ;
      RECT 39.64 10.09 39.81 10.6 ;
      RECT 39.63 4.785 39.8 5.115 ;
      RECT 38.94 3.795 39.11 4.245 ;
      RECT 38.46 3.795 38.63 4.125 ;
      RECT 37.98 3.795 38.15 4.125 ;
      RECT 37.5 3.795 37.67 4.245 ;
      RECT 37.26 4.785 37.43 5.115 ;
      RECT 37.02 3.795 37.19 4.525 ;
      RECT 36.54 3.795 36.71 4.125 ;
      RECT 36.3 3.055 36.47 3.405 ;
      RECT 35.82 4.355 35.99 4.775 ;
      RECT 35.58 3.795 35.75 4.125 ;
      RECT 35.34 4.445 35.51 4.805 ;
      RECT 35.1 3.795 35.27 4.245 ;
      RECT 34.62 3.795 34.79 4.245 ;
      RECT 34.41 3.055 34.58 3.405 ;
      RECT 34.41 4.445 34.58 4.805 ;
      RECT 32.775 7.315 32.945 8.785 ;
      RECT 32.775 10.095 32.945 10.605 ;
      RECT 31.785 1.87 31.955 2.38 ;
      RECT 31.785 3.69 31.955 5.16 ;
      RECT 31.785 7.315 31.955 8.785 ;
      RECT 31.785 10.095 31.955 10.605 ;
      RECT 30.425 1.875 30.595 5.165 ;
      RECT 30.425 7.31 30.595 10.6 ;
      RECT 29.995 1.875 30.165 2.385 ;
      RECT 29.995 2.955 30.165 5.165 ;
      RECT 29.995 7.31 30.165 9.52 ;
      RECT 29.995 10.09 30.165 10.6 ;
      RECT 26.32 3.055 26.49 3.405 ;
      RECT 26.08 3.795 26.25 4.125 ;
      RECT 25.6 3.795 25.77 4.245 ;
      RECT 25.36 3.055 25.53 3.405 ;
      RECT 25.12 3.795 25.29 4.125 ;
      RECT 24.81 7.31 24.98 10.6 ;
      RECT 24.38 7.31 24.55 9.52 ;
      RECT 24.38 10.09 24.55 10.6 ;
      RECT 24.37 4.785 24.54 5.115 ;
      RECT 23.68 3.795 23.85 4.245 ;
      RECT 23.2 3.795 23.37 4.125 ;
      RECT 22.72 3.795 22.89 4.125 ;
      RECT 22.24 3.795 22.41 4.245 ;
      RECT 22 4.785 22.17 5.115 ;
      RECT 21.76 3.795 21.93 4.525 ;
      RECT 21.28 3.795 21.45 4.125 ;
      RECT 21.04 3.055 21.21 3.405 ;
      RECT 20.56 4.355 20.73 4.775 ;
      RECT 20.32 3.795 20.49 4.125 ;
      RECT 20.08 4.445 20.25 4.805 ;
      RECT 19.84 3.795 20.01 4.245 ;
      RECT 19.36 3.795 19.53 4.245 ;
      RECT 19.15 3.055 19.32 3.405 ;
      RECT 19.15 4.445 19.32 4.805 ;
      RECT 17.515 7.315 17.685 8.785 ;
      RECT 17.515 10.095 17.685 10.605 ;
      RECT 16.525 1.87 16.695 2.38 ;
      RECT 16.525 3.69 16.695 5.16 ;
      RECT 16.525 7.315 16.695 8.785 ;
      RECT 16.525 10.095 16.695 10.605 ;
      RECT 15.165 1.875 15.335 5.165 ;
      RECT 15.165 7.31 15.335 10.6 ;
      RECT 14.735 1.875 14.905 2.385 ;
      RECT 14.735 2.955 14.905 5.165 ;
      RECT 14.735 7.31 14.905 9.52 ;
      RECT 14.735 10.09 14.905 10.6 ;
      RECT 11.06 3.055 11.23 3.405 ;
      RECT 10.82 3.795 10.99 4.125 ;
      RECT 10.34 3.795 10.51 4.245 ;
      RECT 10.1 3.055 10.27 3.405 ;
      RECT 9.86 3.795 10.03 4.125 ;
      RECT 9.55 7.31 9.72 10.6 ;
      RECT 9.12 7.31 9.29 9.52 ;
      RECT 9.12 10.09 9.29 10.6 ;
      RECT 9.11 4.785 9.28 5.115 ;
      RECT 8.42 3.795 8.59 4.245 ;
      RECT 7.94 3.795 8.11 4.125 ;
      RECT 7.46 3.795 7.63 4.125 ;
      RECT 6.98 3.795 7.15 4.245 ;
      RECT 6.74 4.785 6.91 5.115 ;
      RECT 6.5 3.795 6.67 4.525 ;
      RECT 6.02 3.795 6.19 4.125 ;
      RECT 5.78 3.055 5.95 3.405 ;
      RECT 5.3 4.355 5.47 4.775 ;
      RECT 5.06 3.795 5.23 4.125 ;
      RECT 4.82 4.445 4.99 4.805 ;
      RECT 4.58 3.795 4.75 4.245 ;
      RECT 4.1 3.795 4.27 4.245 ;
      RECT 3.89 3.055 4.06 3.405 ;
      RECT 3.89 4.445 4.06 4.805 ;
      RECT 1.605 7.31 1.775 9.52 ;
      RECT 1.605 10.09 1.775 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r1 ;
  SIZE 79.125 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 17.54 1.865 17.71 2.375 ;
        RECT 17.54 3.685 17.71 5.155 ;
      LAYER met1 ;
        RECT 17.48 3.655 17.77 3.885 ;
        RECT 17.48 2.175 17.77 2.405 ;
        RECT 17.54 2.175 17.71 3.885 ;
      LAYER mcon ;
        RECT 17.54 3.685 17.71 3.855 ;
        RECT 17.54 2.205 17.71 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 32.8 1.865 32.97 2.375 ;
        RECT 32.8 3.685 32.97 5.155 ;
      LAYER met1 ;
        RECT 32.74 3.655 33.03 3.885 ;
        RECT 32.74 2.175 33.03 2.405 ;
        RECT 32.8 2.175 32.97 3.885 ;
      LAYER mcon ;
        RECT 32.8 3.685 32.97 3.855 ;
        RECT 32.8 2.205 32.97 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 48.06 1.865 48.23 2.375 ;
        RECT 48.06 3.685 48.23 5.155 ;
      LAYER met1 ;
        RECT 48 3.655 48.29 3.885 ;
        RECT 48 2.175 48.29 2.405 ;
        RECT 48.06 2.175 48.23 3.885 ;
      LAYER mcon ;
        RECT 48.06 3.685 48.23 3.855 ;
        RECT 48.06 2.205 48.23 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 63.32 1.865 63.49 2.375 ;
        RECT 63.32 3.685 63.49 5.155 ;
      LAYER met1 ;
        RECT 63.26 3.655 63.55 3.885 ;
        RECT 63.26 2.175 63.55 2.405 ;
        RECT 63.32 2.175 63.49 3.885 ;
      LAYER mcon ;
        RECT 63.32 3.685 63.49 3.855 ;
        RECT 63.32 2.205 63.49 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 78.58 1.865 78.75 2.375 ;
        RECT 78.58 3.685 78.75 5.155 ;
      LAYER met1 ;
        RECT 78.52 3.655 78.81 3.885 ;
        RECT 78.52 2.175 78.81 2.405 ;
        RECT 78.58 2.175 78.75 3.885 ;
      LAYER mcon ;
        RECT 78.58 3.685 78.75 3.855 ;
        RECT 78.58 2.205 78.75 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 13.31 4 13.65 4.35 ;
        RECT 13.305 8.15 13.645 8.5 ;
        RECT 13.385 4 13.56 8.5 ;
      LAYER li1 ;
        RECT 13.39 2.955 13.56 4.23 ;
        RECT 13.39 8.235 13.56 9.51 ;
        RECT 7.755 8.235 7.925 9.51 ;
      LAYER met1 ;
        RECT 13.31 4.06 13.79 4.23 ;
        RECT 13.31 4 13.65 4.35 ;
        RECT 7.695 8.235 13.79 8.405 ;
        RECT 13.305 8.15 13.645 8.5 ;
        RECT 7.695 8.205 7.985 8.435 ;
      LAYER via1 ;
        RECT 13.405 8.25 13.555 8.4 ;
        RECT 13.41 4.1 13.56 4.25 ;
      LAYER mcon ;
        RECT 7.755 8.235 7.925 8.405 ;
        RECT 13.39 8.235 13.56 8.405 ;
        RECT 13.39 4.06 13.56 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 28.57 4 28.91 4.35 ;
        RECT 28.565 8.15 28.905 8.5 ;
        RECT 28.645 4 28.82 8.5 ;
      LAYER li1 ;
        RECT 28.65 2.955 28.82 4.23 ;
        RECT 28.65 8.235 28.82 9.51 ;
        RECT 23.015 8.235 23.185 9.51 ;
      LAYER met1 ;
        RECT 28.57 4.06 29.05 4.23 ;
        RECT 28.57 4 28.91 4.35 ;
        RECT 22.955 8.235 29.05 8.405 ;
        RECT 28.565 8.15 28.905 8.5 ;
        RECT 22.955 8.205 23.245 8.435 ;
      LAYER via1 ;
        RECT 28.665 8.25 28.815 8.4 ;
        RECT 28.67 4.1 28.82 4.25 ;
      LAYER mcon ;
        RECT 23.015 8.235 23.185 8.405 ;
        RECT 28.65 8.235 28.82 8.405 ;
        RECT 28.65 4.06 28.82 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 43.83 4 44.17 4.35 ;
        RECT 43.825 8.15 44.165 8.5 ;
        RECT 43.905 4 44.08 8.5 ;
      LAYER li1 ;
        RECT 43.91 2.955 44.08 4.23 ;
        RECT 43.91 8.235 44.08 9.51 ;
        RECT 38.275 8.235 38.445 9.51 ;
      LAYER met1 ;
        RECT 43.83 4.06 44.31 4.23 ;
        RECT 43.83 4 44.17 4.35 ;
        RECT 38.215 8.235 44.31 8.405 ;
        RECT 43.825 8.15 44.165 8.5 ;
        RECT 38.215 8.205 38.505 8.435 ;
      LAYER via1 ;
        RECT 43.925 8.25 44.075 8.4 ;
        RECT 43.93 4.1 44.08 4.25 ;
      LAYER mcon ;
        RECT 38.275 8.235 38.445 8.405 ;
        RECT 43.91 8.235 44.08 8.405 ;
        RECT 43.91 4.06 44.08 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 59.09 4 59.43 4.35 ;
        RECT 59.085 8.15 59.425 8.5 ;
        RECT 59.165 4 59.34 8.5 ;
      LAYER li1 ;
        RECT 59.17 2.955 59.34 4.23 ;
        RECT 59.17 8.235 59.34 9.51 ;
        RECT 53.535 8.235 53.705 9.51 ;
      LAYER met1 ;
        RECT 59.09 4.06 59.57 4.23 ;
        RECT 59.09 4 59.43 4.35 ;
        RECT 53.475 8.235 59.57 8.405 ;
        RECT 59.085 8.15 59.425 8.5 ;
        RECT 53.475 8.205 53.765 8.435 ;
      LAYER via1 ;
        RECT 59.185 8.25 59.335 8.4 ;
        RECT 59.19 4.1 59.34 4.25 ;
      LAYER mcon ;
        RECT 53.535 8.235 53.705 8.405 ;
        RECT 59.17 8.235 59.34 8.405 ;
        RECT 59.17 4.06 59.34 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 74.35 4 74.69 4.35 ;
        RECT 74.345 8.15 74.685 8.5 ;
        RECT 74.425 4 74.6 8.5 ;
      LAYER li1 ;
        RECT 74.43 2.955 74.6 4.23 ;
        RECT 74.43 8.235 74.6 9.51 ;
        RECT 68.795 8.235 68.965 9.51 ;
      LAYER met1 ;
        RECT 74.35 4.06 74.83 4.23 ;
        RECT 74.35 4 74.69 4.35 ;
        RECT 68.735 8.235 74.83 8.405 ;
        RECT 74.345 8.15 74.685 8.5 ;
        RECT 68.735 8.205 69.025 8.435 ;
      LAYER via1 ;
        RECT 74.445 8.25 74.595 8.4 ;
        RECT 74.45 4.1 74.6 4.25 ;
      LAYER mcon ;
        RECT 68.795 8.235 68.965 8.405 ;
        RECT 74.43 8.235 74.6 8.405 ;
        RECT 74.43 4.06 74.6 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.26 8.235 0.43 9.51 ;
      LAYER met1 ;
        RECT 0.2 8.235 0.66 8.405 ;
        RECT 0.2 8.205 0.49 8.435 ;
      LAYER mcon ;
        RECT 0.26 8.235 0.43 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.025 5.435 79.125 7.035 ;
        RECT 64.615 5.43 79.125 7.035 ;
        RECT 76.99 5.425 78.97 7.04 ;
        RECT 78.15 4.695 78.32 7.77 ;
        RECT 77.16 4.695 77.33 7.77 ;
        RECT 74.42 4.7 74.59 7.765 ;
        RECT 71.645 4.93 71.815 7.035 ;
        RECT 69.725 4.93 69.895 7.035 ;
        RECT 68.785 4.93 68.955 7.765 ;
        RECT 67.325 4.93 67.495 7.035 ;
        RECT 65.405 4.93 65.575 7.035 ;
        RECT 49.355 5.43 63.865 7.035 ;
        RECT 61.73 5.425 63.71 7.04 ;
        RECT 62.89 4.695 63.06 7.77 ;
        RECT 61.9 4.695 62.07 7.77 ;
        RECT 59.16 4.7 59.33 7.765 ;
        RECT 56.385 4.93 56.555 7.035 ;
        RECT 54.465 4.93 54.635 7.035 ;
        RECT 53.525 4.93 53.695 7.765 ;
        RECT 52.065 4.93 52.235 7.035 ;
        RECT 50.145 4.93 50.315 7.035 ;
        RECT 34.095 5.43 48.605 7.035 ;
        RECT 46.47 5.425 48.45 7.04 ;
        RECT 47.63 4.695 47.8 7.77 ;
        RECT 46.64 4.695 46.81 7.77 ;
        RECT 43.9 4.7 44.07 7.765 ;
        RECT 41.125 4.93 41.295 7.035 ;
        RECT 39.205 4.93 39.375 7.035 ;
        RECT 38.265 4.93 38.435 7.765 ;
        RECT 36.805 4.93 36.975 7.035 ;
        RECT 34.885 4.93 35.055 7.035 ;
        RECT 18.835 5.43 33.345 7.035 ;
        RECT 31.21 5.425 33.19 7.04 ;
        RECT 32.37 4.695 32.54 7.77 ;
        RECT 31.38 4.695 31.55 7.77 ;
        RECT 28.64 4.7 28.81 7.765 ;
        RECT 25.865 4.93 26.035 7.035 ;
        RECT 23.945 4.93 24.115 7.035 ;
        RECT 23.005 4.93 23.175 7.765 ;
        RECT 21.545 4.93 21.715 7.035 ;
        RECT 19.625 4.93 19.795 7.035 ;
        RECT 3.575 5.43 18.085 7.035 ;
        RECT 15.95 5.425 17.93 7.04 ;
        RECT 17.11 4.695 17.28 7.77 ;
        RECT 16.12 4.695 16.29 7.77 ;
        RECT 13.38 4.7 13.55 7.765 ;
        RECT 10.605 4.93 10.775 7.035 ;
        RECT 8.685 4.93 8.855 7.035 ;
        RECT 7.745 4.93 7.915 7.765 ;
        RECT 6.285 4.93 6.455 7.035 ;
        RECT 4.365 4.93 4.535 7.035 ;
        RECT 2.06 5.435 2.23 10.595 ;
        RECT 0.25 5.435 0.42 7.765 ;
      LAYER met1 ;
        RECT 0.025 5.435 79.125 7.035 ;
        RECT 64.615 5.43 79.125 7.035 ;
        RECT 76.99 5.425 78.97 7.04 ;
        RECT 64.615 5.275 73.355 7.035 ;
        RECT 49.355 5.43 63.865 7.035 ;
        RECT 61.73 5.425 63.71 7.04 ;
        RECT 49.355 5.275 58.095 7.035 ;
        RECT 34.095 5.43 48.605 7.035 ;
        RECT 46.47 5.425 48.45 7.04 ;
        RECT 34.095 5.275 42.835 7.035 ;
        RECT 18.835 5.43 33.345 7.035 ;
        RECT 31.21 5.425 33.19 7.04 ;
        RECT 18.835 5.275 27.575 7.035 ;
        RECT 3.575 5.43 18.085 7.035 ;
        RECT 15.95 5.425 17.93 7.04 ;
        RECT 3.575 5.275 12.315 7.035 ;
        RECT 2 8.945 2.29 9.175 ;
        RECT 1.83 8.975 2.29 9.145 ;
      LAYER mcon ;
        RECT 2.06 8.975 2.23 9.145 ;
        RECT 2.37 6.835 2.54 7.005 ;
        RECT 3.72 5.43 3.89 5.6 ;
        RECT 4.18 5.43 4.35 5.6 ;
        RECT 4.64 5.43 4.81 5.6 ;
        RECT 5.1 5.43 5.27 5.6 ;
        RECT 5.56 5.43 5.73 5.6 ;
        RECT 6.02 5.43 6.19 5.6 ;
        RECT 6.48 5.43 6.65 5.6 ;
        RECT 6.94 5.43 7.11 5.6 ;
        RECT 7.4 5.43 7.57 5.6 ;
        RECT 7.86 5.43 8.03 5.6 ;
        RECT 8.32 5.43 8.49 5.6 ;
        RECT 8.78 5.43 8.95 5.6 ;
        RECT 9.24 5.43 9.41 5.6 ;
        RECT 9.7 5.43 9.87 5.6 ;
        RECT 9.865 6.835 10.035 7.005 ;
        RECT 10.16 5.43 10.33 5.6 ;
        RECT 10.62 5.43 10.79 5.6 ;
        RECT 11.08 5.43 11.25 5.6 ;
        RECT 11.54 5.43 11.71 5.6 ;
        RECT 12 5.43 12.17 5.6 ;
        RECT 15.5 6.835 15.67 7.005 ;
        RECT 15.5 5.46 15.67 5.63 ;
        RECT 16.2 6.84 16.37 7.01 ;
        RECT 16.2 5.455 16.37 5.625 ;
        RECT 17.19 6.84 17.36 7.01 ;
        RECT 17.19 5.455 17.36 5.625 ;
        RECT 18.98 5.43 19.15 5.6 ;
        RECT 19.44 5.43 19.61 5.6 ;
        RECT 19.9 5.43 20.07 5.6 ;
        RECT 20.36 5.43 20.53 5.6 ;
        RECT 20.82 5.43 20.99 5.6 ;
        RECT 21.28 5.43 21.45 5.6 ;
        RECT 21.74 5.43 21.91 5.6 ;
        RECT 22.2 5.43 22.37 5.6 ;
        RECT 22.66 5.43 22.83 5.6 ;
        RECT 23.12 5.43 23.29 5.6 ;
        RECT 23.58 5.43 23.75 5.6 ;
        RECT 24.04 5.43 24.21 5.6 ;
        RECT 24.5 5.43 24.67 5.6 ;
        RECT 24.96 5.43 25.13 5.6 ;
        RECT 25.125 6.835 25.295 7.005 ;
        RECT 25.42 5.43 25.59 5.6 ;
        RECT 25.88 5.43 26.05 5.6 ;
        RECT 26.34 5.43 26.51 5.6 ;
        RECT 26.8 5.43 26.97 5.6 ;
        RECT 27.26 5.43 27.43 5.6 ;
        RECT 30.76 6.835 30.93 7.005 ;
        RECT 30.76 5.46 30.93 5.63 ;
        RECT 31.46 6.84 31.63 7.01 ;
        RECT 31.46 5.455 31.63 5.625 ;
        RECT 32.45 6.84 32.62 7.01 ;
        RECT 32.45 5.455 32.62 5.625 ;
        RECT 34.24 5.43 34.41 5.6 ;
        RECT 34.7 5.43 34.87 5.6 ;
        RECT 35.16 5.43 35.33 5.6 ;
        RECT 35.62 5.43 35.79 5.6 ;
        RECT 36.08 5.43 36.25 5.6 ;
        RECT 36.54 5.43 36.71 5.6 ;
        RECT 37 5.43 37.17 5.6 ;
        RECT 37.46 5.43 37.63 5.6 ;
        RECT 37.92 5.43 38.09 5.6 ;
        RECT 38.38 5.43 38.55 5.6 ;
        RECT 38.84 5.43 39.01 5.6 ;
        RECT 39.3 5.43 39.47 5.6 ;
        RECT 39.76 5.43 39.93 5.6 ;
        RECT 40.22 5.43 40.39 5.6 ;
        RECT 40.385 6.835 40.555 7.005 ;
        RECT 40.68 5.43 40.85 5.6 ;
        RECT 41.14 5.43 41.31 5.6 ;
        RECT 41.6 5.43 41.77 5.6 ;
        RECT 42.06 5.43 42.23 5.6 ;
        RECT 42.52 5.43 42.69 5.6 ;
        RECT 46.02 6.835 46.19 7.005 ;
        RECT 46.02 5.46 46.19 5.63 ;
        RECT 46.72 6.84 46.89 7.01 ;
        RECT 46.72 5.455 46.89 5.625 ;
        RECT 47.71 6.84 47.88 7.01 ;
        RECT 47.71 5.455 47.88 5.625 ;
        RECT 49.5 5.43 49.67 5.6 ;
        RECT 49.96 5.43 50.13 5.6 ;
        RECT 50.42 5.43 50.59 5.6 ;
        RECT 50.88 5.43 51.05 5.6 ;
        RECT 51.34 5.43 51.51 5.6 ;
        RECT 51.8 5.43 51.97 5.6 ;
        RECT 52.26 5.43 52.43 5.6 ;
        RECT 52.72 5.43 52.89 5.6 ;
        RECT 53.18 5.43 53.35 5.6 ;
        RECT 53.64 5.43 53.81 5.6 ;
        RECT 54.1 5.43 54.27 5.6 ;
        RECT 54.56 5.43 54.73 5.6 ;
        RECT 55.02 5.43 55.19 5.6 ;
        RECT 55.48 5.43 55.65 5.6 ;
        RECT 55.645 6.835 55.815 7.005 ;
        RECT 55.94 5.43 56.11 5.6 ;
        RECT 56.4 5.43 56.57 5.6 ;
        RECT 56.86 5.43 57.03 5.6 ;
        RECT 57.32 5.43 57.49 5.6 ;
        RECT 57.78 5.43 57.95 5.6 ;
        RECT 61.28 6.835 61.45 7.005 ;
        RECT 61.28 5.46 61.45 5.63 ;
        RECT 61.98 6.84 62.15 7.01 ;
        RECT 61.98 5.455 62.15 5.625 ;
        RECT 62.97 6.84 63.14 7.01 ;
        RECT 62.97 5.455 63.14 5.625 ;
        RECT 64.76 5.43 64.93 5.6 ;
        RECT 65.22 5.43 65.39 5.6 ;
        RECT 65.68 5.43 65.85 5.6 ;
        RECT 66.14 5.43 66.31 5.6 ;
        RECT 66.6 5.43 66.77 5.6 ;
        RECT 67.06 5.43 67.23 5.6 ;
        RECT 67.52 5.43 67.69 5.6 ;
        RECT 67.98 5.43 68.15 5.6 ;
        RECT 68.44 5.43 68.61 5.6 ;
        RECT 68.9 5.43 69.07 5.6 ;
        RECT 69.36 5.43 69.53 5.6 ;
        RECT 69.82 5.43 69.99 5.6 ;
        RECT 70.28 5.43 70.45 5.6 ;
        RECT 70.74 5.43 70.91 5.6 ;
        RECT 70.905 6.835 71.075 7.005 ;
        RECT 71.2 5.43 71.37 5.6 ;
        RECT 71.66 5.43 71.83 5.6 ;
        RECT 72.12 5.43 72.29 5.6 ;
        RECT 72.58 5.43 72.75 5.6 ;
        RECT 73.04 5.43 73.21 5.6 ;
        RECT 76.54 6.835 76.71 7.005 ;
        RECT 76.54 5.46 76.71 5.63 ;
        RECT 77.24 6.84 77.41 7.01 ;
        RECT 77.24 5.455 77.41 5.625 ;
        RECT 78.23 6.84 78.4 7.01 ;
        RECT 78.23 5.455 78.4 5.625 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.035 10.865 79.125 12.465 ;
        RECT 78.15 10.24 78.32 12.465 ;
        RECT 77.16 10.24 77.33 12.465 ;
        RECT 74.42 10.235 74.59 12.465 ;
        RECT 68.785 10.235 68.955 12.465 ;
        RECT 62.89 10.24 63.06 12.465 ;
        RECT 61.9 10.24 62.07 12.465 ;
        RECT 59.16 10.235 59.33 12.465 ;
        RECT 53.525 10.235 53.695 12.465 ;
        RECT 47.63 10.24 47.8 12.465 ;
        RECT 46.64 10.24 46.81 12.465 ;
        RECT 43.9 10.235 44.07 12.465 ;
        RECT 38.265 10.235 38.435 12.465 ;
        RECT 32.37 10.24 32.54 12.465 ;
        RECT 31.38 10.24 31.55 12.465 ;
        RECT 28.64 10.235 28.81 12.465 ;
        RECT 23.005 10.235 23.175 12.465 ;
        RECT 17.11 10.24 17.28 12.465 ;
        RECT 16.12 10.24 16.29 12.465 ;
        RECT 13.38 10.235 13.55 12.465 ;
        RECT 7.745 10.235 7.915 12.465 ;
        RECT 0.25 10.235 0.42 12.465 ;
        RECT 69.79 8.365 69.96 10.315 ;
        RECT 69.735 10.145 69.905 10.595 ;
        RECT 69.735 7.305 69.905 8.535 ;
        RECT 54.53 8.365 54.7 10.315 ;
        RECT 54.475 10.145 54.645 10.595 ;
        RECT 54.475 7.305 54.645 8.535 ;
        RECT 39.27 8.365 39.44 10.315 ;
        RECT 39.215 10.145 39.385 10.595 ;
        RECT 39.215 7.305 39.385 8.535 ;
        RECT 24.01 8.365 24.18 10.315 ;
        RECT 23.955 10.145 24.125 10.595 ;
        RECT 23.955 7.305 24.125 8.535 ;
        RECT 8.75 8.365 8.92 10.315 ;
        RECT 8.695 10.145 8.865 10.595 ;
        RECT 8.695 7.305 8.865 8.535 ;
      LAYER met1 ;
        RECT 0.035 10.865 79.125 12.465 ;
        RECT 69.73 8.575 70.02 8.805 ;
        RECT 69.56 8.605 69.73 12.465 ;
        RECT 54.47 8.575 54.76 8.805 ;
        RECT 54.3 8.605 54.47 12.465 ;
        RECT 39.21 8.575 39.5 8.805 ;
        RECT 39.04 8.605 39.21 12.465 ;
        RECT 23.95 8.575 24.24 8.805 ;
        RECT 23.78 8.605 23.95 12.465 ;
        RECT 8.69 8.575 8.98 8.805 ;
        RECT 8.52 8.605 8.69 12.465 ;
      LAYER mcon ;
        RECT 0.33 10.895 0.5 11.065 ;
        RECT 1.01 10.895 1.18 11.065 ;
        RECT 1.69 10.895 1.86 11.065 ;
        RECT 2.37 10.895 2.54 11.065 ;
        RECT 7.825 10.895 7.995 11.065 ;
        RECT 8.505 10.895 8.675 11.065 ;
        RECT 8.75 8.605 8.92 8.775 ;
        RECT 9.185 10.895 9.355 11.065 ;
        RECT 9.865 10.895 10.035 11.065 ;
        RECT 13.46 10.895 13.63 11.065 ;
        RECT 14.14 10.895 14.31 11.065 ;
        RECT 14.82 10.895 14.99 11.065 ;
        RECT 15.5 10.895 15.67 11.065 ;
        RECT 16.2 10.9 16.37 11.07 ;
        RECT 17.19 10.9 17.36 11.07 ;
        RECT 23.085 10.895 23.255 11.065 ;
        RECT 23.765 10.895 23.935 11.065 ;
        RECT 24.01 8.605 24.18 8.775 ;
        RECT 24.445 10.895 24.615 11.065 ;
        RECT 25.125 10.895 25.295 11.065 ;
        RECT 28.72 10.895 28.89 11.065 ;
        RECT 29.4 10.895 29.57 11.065 ;
        RECT 30.08 10.895 30.25 11.065 ;
        RECT 30.76 10.895 30.93 11.065 ;
        RECT 31.46 10.9 31.63 11.07 ;
        RECT 32.45 10.9 32.62 11.07 ;
        RECT 38.345 10.895 38.515 11.065 ;
        RECT 39.025 10.895 39.195 11.065 ;
        RECT 39.27 8.605 39.44 8.775 ;
        RECT 39.705 10.895 39.875 11.065 ;
        RECT 40.385 10.895 40.555 11.065 ;
        RECT 43.98 10.895 44.15 11.065 ;
        RECT 44.66 10.895 44.83 11.065 ;
        RECT 45.34 10.895 45.51 11.065 ;
        RECT 46.02 10.895 46.19 11.065 ;
        RECT 46.72 10.9 46.89 11.07 ;
        RECT 47.71 10.9 47.88 11.07 ;
        RECT 53.605 10.895 53.775 11.065 ;
        RECT 54.285 10.895 54.455 11.065 ;
        RECT 54.53 8.605 54.7 8.775 ;
        RECT 54.965 10.895 55.135 11.065 ;
        RECT 55.645 10.895 55.815 11.065 ;
        RECT 59.24 10.895 59.41 11.065 ;
        RECT 59.92 10.895 60.09 11.065 ;
        RECT 60.6 10.895 60.77 11.065 ;
        RECT 61.28 10.895 61.45 11.065 ;
        RECT 61.98 10.9 62.15 11.07 ;
        RECT 62.97 10.9 63.14 11.07 ;
        RECT 68.865 10.895 69.035 11.065 ;
        RECT 69.545 10.895 69.715 11.065 ;
        RECT 69.79 8.605 69.96 8.775 ;
        RECT 70.225 10.895 70.395 11.065 ;
        RECT 70.905 10.895 71.075 11.065 ;
        RECT 74.5 10.895 74.67 11.065 ;
        RECT 75.18 10.895 75.35 11.065 ;
        RECT 75.86 10.895 76.03 11.065 ;
        RECT 76.54 10.895 76.71 11.065 ;
        RECT 77.24 10.9 77.41 11.07 ;
        RECT 78.23 10.9 78.4 11.07 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 70.065 9.345 70.435 9.715 ;
      RECT 70.1 5.565 70.4 9.715 ;
      RECT 65.91 5.565 70.4 6.86 ;
      RECT 69.09 3.15 69.39 6.86 ;
      RECT 65.91 3.73 66.21 6.86 ;
      RECT 69.045 4.055 69.39 4.785 ;
      RECT 65.805 3.31 66.135 4.04 ;
      RECT 68.685 3.15 69.415 3.48 ;
      RECT 54.805 9.345 55.175 9.715 ;
      RECT 54.84 5.565 55.14 9.715 ;
      RECT 50.65 5.565 55.14 6.86 ;
      RECT 53.83 3.15 54.13 6.86 ;
      RECT 50.65 3.73 50.95 6.86 ;
      RECT 53.785 4.055 54.13 4.785 ;
      RECT 50.545 3.31 50.875 4.04 ;
      RECT 53.425 3.15 54.155 3.48 ;
      RECT 39.545 9.345 39.915 9.715 ;
      RECT 39.58 5.565 39.88 9.715 ;
      RECT 35.39 5.565 39.88 6.86 ;
      RECT 38.57 3.15 38.87 6.86 ;
      RECT 35.39 3.73 35.69 6.86 ;
      RECT 38.525 4.055 38.87 4.785 ;
      RECT 35.285 3.31 35.615 4.04 ;
      RECT 38.165 3.15 38.895 3.48 ;
      RECT 24.285 9.345 24.655 9.715 ;
      RECT 24.32 5.565 24.62 9.715 ;
      RECT 20.13 5.565 24.62 6.86 ;
      RECT 23.31 3.15 23.61 6.86 ;
      RECT 20.13 3.73 20.43 6.86 ;
      RECT 23.265 4.055 23.61 4.785 ;
      RECT 20.025 3.31 20.355 4.04 ;
      RECT 22.905 3.15 23.635 3.48 ;
      RECT 9.025 9.345 9.395 9.715 ;
      RECT 9.06 5.565 9.36 9.715 ;
      RECT 4.87 5.565 9.36 6.86 ;
      RECT 8.05 3.15 8.35 6.86 ;
      RECT 4.87 3.73 5.17 6.86 ;
      RECT 8.005 4.055 8.35 4.785 ;
      RECT 4.765 3.31 5.095 4.04 ;
      RECT 7.645 3.15 8.375 3.48 ;
      RECT 72.165 3.31 72.495 4.04 ;
      RECT 70.965 4.175 71.295 4.905 ;
      RECT 70.125 3.15 70.855 3.48 ;
      RECT 67.725 3.15 68.055 3.88 ;
      RECT 66.525 3.31 66.855 4.04 ;
      RECT 56.905 3.31 57.235 4.04 ;
      RECT 55.705 4.175 56.035 4.905 ;
      RECT 54.865 3.15 55.595 3.48 ;
      RECT 52.465 3.15 52.795 3.88 ;
      RECT 51.265 3.31 51.595 4.04 ;
      RECT 41.645 3.31 41.975 4.04 ;
      RECT 40.445 4.175 40.775 4.905 ;
      RECT 39.605 3.15 40.335 3.48 ;
      RECT 37.205 3.15 37.535 3.88 ;
      RECT 36.005 3.31 36.335 4.04 ;
      RECT 26.385 3.31 26.715 4.04 ;
      RECT 25.185 4.175 25.515 4.905 ;
      RECT 24.345 3.15 25.075 3.48 ;
      RECT 21.945 3.15 22.275 3.88 ;
      RECT 20.745 3.31 21.075 4.04 ;
      RECT 11.125 3.31 11.455 4.04 ;
      RECT 9.925 4.175 10.255 4.905 ;
      RECT 9.085 3.15 9.815 3.48 ;
      RECT 6.685 3.15 7.015 3.88 ;
      RECT 5.485 3.31 5.815 4.04 ;
    LAYER via2 ;
      RECT 72.23 3.775 72.43 3.975 ;
      RECT 71.03 4.335 71.23 4.535 ;
      RECT 70.19 3.215 70.39 3.415 ;
      RECT 70.15 9.43 70.35 9.63 ;
      RECT 69.11 4.12 69.31 4.32 ;
      RECT 68.75 3.215 68.95 3.415 ;
      RECT 67.79 3.215 67.99 3.415 ;
      RECT 66.59 3.775 66.79 3.975 ;
      RECT 65.87 3.775 66.07 3.975 ;
      RECT 56.97 3.775 57.17 3.975 ;
      RECT 55.77 4.335 55.97 4.535 ;
      RECT 54.93 3.215 55.13 3.415 ;
      RECT 54.89 9.43 55.09 9.63 ;
      RECT 53.85 4.12 54.05 4.32 ;
      RECT 53.49 3.215 53.69 3.415 ;
      RECT 52.53 3.215 52.73 3.415 ;
      RECT 51.33 3.775 51.53 3.975 ;
      RECT 50.61 3.775 50.81 3.975 ;
      RECT 41.71 3.775 41.91 3.975 ;
      RECT 40.51 4.335 40.71 4.535 ;
      RECT 39.67 3.215 39.87 3.415 ;
      RECT 39.63 9.43 39.83 9.63 ;
      RECT 38.59 4.12 38.79 4.32 ;
      RECT 38.23 3.215 38.43 3.415 ;
      RECT 37.27 3.215 37.47 3.415 ;
      RECT 36.07 3.775 36.27 3.975 ;
      RECT 35.35 3.775 35.55 3.975 ;
      RECT 26.45 3.775 26.65 3.975 ;
      RECT 25.25 4.335 25.45 4.535 ;
      RECT 24.41 3.215 24.61 3.415 ;
      RECT 24.37 9.43 24.57 9.63 ;
      RECT 23.33 4.12 23.53 4.32 ;
      RECT 22.97 3.215 23.17 3.415 ;
      RECT 22.01 3.215 22.21 3.415 ;
      RECT 20.81 3.775 21.01 3.975 ;
      RECT 20.09 3.775 20.29 3.975 ;
      RECT 11.19 3.775 11.39 3.975 ;
      RECT 9.99 4.335 10.19 4.535 ;
      RECT 9.15 3.215 9.35 3.415 ;
      RECT 9.11 9.43 9.31 9.63 ;
      RECT 8.07 4.12 8.27 4.32 ;
      RECT 7.71 3.215 7.91 3.415 ;
      RECT 6.75 3.215 6.95 3.415 ;
      RECT 5.55 3.775 5.75 3.975 ;
      RECT 4.83 3.775 5.03 3.975 ;
    LAYER met2 ;
      RECT 1.26 10.69 78.755 10.86 ;
      RECT 78.585 9.565 78.755 10.86 ;
      RECT 1.26 8.545 1.43 10.86 ;
      RECT 78.555 9.565 78.905 9.915 ;
      RECT 1.195 8.545 1.485 8.895 ;
      RECT 75.395 8.51 75.715 8.835 ;
      RECT 75.425 7.985 75.595 8.835 ;
      RECT 75.425 7.985 75.6 8.335 ;
      RECT 75.425 7.985 76.4 8.16 ;
      RECT 76.225 3.26 76.4 8.16 ;
      RECT 76.17 3.26 76.52 3.61 ;
      RECT 76.195 8.945 76.52 9.27 ;
      RECT 75.08 9.035 76.52 9.205 ;
      RECT 75.08 3.69 75.24 9.205 ;
      RECT 75.395 3.66 75.715 3.98 ;
      RECT 75.08 3.69 75.715 3.86 ;
      RECT 73.79 4 74.13 4.35 ;
      RECT 73.185 4.065 74.13 4.265 ;
      RECT 73.185 4.06 73.4 4.265 ;
      RECT 73.2 3.635 73.4 4.265 ;
      RECT 72.19 3.635 72.47 4.015 ;
      RECT 73.88 3.995 74.05 4.35 ;
      RECT 72.185 3.635 72.47 3.968 ;
      RECT 72.165 3.635 72.47 3.945 ;
      RECT 72.155 3.635 72.47 3.925 ;
      RECT 72.145 3.635 72.47 3.91 ;
      RECT 72.12 3.635 72.47 3.883 ;
      RECT 72.11 3.635 72.47 3.858 ;
      RECT 72.065 3.59 72.345 3.85 ;
      RECT 72.065 3.635 73.4 3.835 ;
      RECT 72.065 3.63 72.39 3.85 ;
      RECT 72.065 3.622 72.385 3.85 ;
      RECT 72.065 3.612 72.38 3.85 ;
      RECT 72.065 3.6 72.375 3.85 ;
      RECT 70.99 4.295 71.27 4.575 ;
      RECT 70.99 4.295 71.305 4.555 ;
      RECT 63.27 8.945 63.62 9.295 ;
      RECT 70.735 8.9 71.085 9.25 ;
      RECT 63.27 8.975 71.085 9.175 ;
      RECT 71.025 3.715 71.075 3.975 ;
      RECT 70.815 3.715 70.82 3.975 ;
      RECT 70.01 3.27 70.04 3.53 ;
      RECT 69.78 3.27 69.855 3.53 ;
      RECT 71 3.665 71.025 3.975 ;
      RECT 70.995 3.622 71 3.975 ;
      RECT 70.99 3.605 70.995 3.975 ;
      RECT 70.985 3.592 70.99 3.975 ;
      RECT 70.91 3.475 70.985 3.975 ;
      RECT 70.865 3.292 70.91 3.975 ;
      RECT 70.86 3.22 70.865 3.975 ;
      RECT 70.845 3.195 70.86 3.975 ;
      RECT 70.82 3.157 70.845 3.975 ;
      RECT 70.81 3.137 70.82 3.697 ;
      RECT 70.795 3.129 70.81 3.652 ;
      RECT 70.79 3.121 70.795 3.623 ;
      RECT 70.785 3.118 70.79 3.603 ;
      RECT 70.78 3.115 70.785 3.583 ;
      RECT 70.775 3.112 70.78 3.563 ;
      RECT 70.745 3.101 70.775 3.5 ;
      RECT 70.725 3.086 70.745 3.415 ;
      RECT 70.72 3.078 70.725 3.378 ;
      RECT 70.71 3.072 70.72 3.345 ;
      RECT 70.695 3.064 70.71 3.305 ;
      RECT 70.69 3.057 70.695 3.265 ;
      RECT 70.685 3.054 70.69 3.243 ;
      RECT 70.68 3.051 70.685 3.23 ;
      RECT 70.675 3.05 70.68 3.22 ;
      RECT 70.66 3.044 70.675 3.21 ;
      RECT 70.635 3.031 70.66 3.195 ;
      RECT 70.585 3.006 70.635 3.166 ;
      RECT 70.57 2.985 70.585 3.141 ;
      RECT 70.56 2.978 70.57 3.13 ;
      RECT 70.505 2.959 70.56 3.103 ;
      RECT 70.48 2.937 70.505 3.076 ;
      RECT 70.475 2.93 70.48 3.071 ;
      RECT 70.46 2.93 70.475 3.069 ;
      RECT 70.435 2.922 70.46 3.065 ;
      RECT 70.42 2.92 70.435 3.061 ;
      RECT 70.39 2.92 70.42 3.058 ;
      RECT 70.38 2.92 70.39 3.053 ;
      RECT 70.335 2.92 70.38 3.051 ;
      RECT 70.306 2.92 70.335 3.052 ;
      RECT 70.22 2.92 70.306 3.054 ;
      RECT 70.206 2.921 70.22 3.056 ;
      RECT 70.12 2.922 70.206 3.058 ;
      RECT 70.105 2.923 70.12 3.068 ;
      RECT 70.1 2.924 70.105 3.077 ;
      RECT 70.08 2.927 70.1 3.087 ;
      RECT 70.065 2.935 70.08 3.102 ;
      RECT 70.045 2.953 70.065 3.117 ;
      RECT 70.035 2.965 70.045 3.14 ;
      RECT 70.025 2.974 70.035 3.17 ;
      RECT 70.01 2.986 70.025 3.215 ;
      RECT 69.955 3.019 70.01 3.53 ;
      RECT 69.95 3.047 69.955 3.53 ;
      RECT 69.93 3.062 69.95 3.53 ;
      RECT 69.895 3.122 69.93 3.53 ;
      RECT 69.893 3.172 69.895 3.53 ;
      RECT 69.89 3.18 69.893 3.53 ;
      RECT 69.88 3.195 69.89 3.53 ;
      RECT 69.875 3.207 69.88 3.53 ;
      RECT 69.865 3.232 69.875 3.53 ;
      RECT 69.855 3.26 69.865 3.53 ;
      RECT 67.76 4.765 67.81 5.025 ;
      RECT 70.67 4.315 70.73 4.575 ;
      RECT 70.655 4.315 70.67 4.585 ;
      RECT 70.636 4.315 70.655 4.618 ;
      RECT 70.55 4.315 70.636 4.743 ;
      RECT 70.47 4.315 70.55 4.925 ;
      RECT 70.465 4.552 70.47 5.01 ;
      RECT 70.44 4.622 70.465 5.038 ;
      RECT 70.435 4.692 70.44 5.065 ;
      RECT 70.415 4.764 70.435 5.087 ;
      RECT 70.41 4.831 70.415 5.11 ;
      RECT 70.4 4.86 70.41 5.125 ;
      RECT 70.39 4.882 70.4 5.142 ;
      RECT 70.385 4.892 70.39 5.153 ;
      RECT 70.38 4.9 70.385 5.161 ;
      RECT 70.37 4.908 70.38 5.173 ;
      RECT 70.365 4.92 70.37 5.183 ;
      RECT 70.36 4.928 70.365 5.188 ;
      RECT 70.34 4.946 70.36 5.198 ;
      RECT 70.335 4.963 70.34 5.205 ;
      RECT 70.33 4.971 70.335 5.206 ;
      RECT 70.325 4.982 70.33 5.208 ;
      RECT 70.285 5.02 70.325 5.218 ;
      RECT 70.28 5.055 70.285 5.229 ;
      RECT 70.275 5.06 70.28 5.232 ;
      RECT 70.25 5.07 70.275 5.239 ;
      RECT 70.24 5.084 70.25 5.248 ;
      RECT 70.22 5.096 70.24 5.251 ;
      RECT 70.17 5.115 70.22 5.255 ;
      RECT 70.125 5.13 70.17 5.26 ;
      RECT 70.06 5.133 70.125 5.266 ;
      RECT 70.045 5.131 70.06 5.273 ;
      RECT 70.015 5.13 70.045 5.273 ;
      RECT 69.976 5.129 70.015 5.269 ;
      RECT 69.89 5.126 69.976 5.265 ;
      RECT 69.873 5.124 69.89 5.262 ;
      RECT 69.787 5.122 69.873 5.259 ;
      RECT 69.701 5.119 69.787 5.253 ;
      RECT 69.615 5.115 69.701 5.248 ;
      RECT 69.537 5.112 69.615 5.244 ;
      RECT 69.451 5.109 69.537 5.242 ;
      RECT 69.365 5.106 69.451 5.239 ;
      RECT 69.307 5.104 69.365 5.236 ;
      RECT 69.221 5.101 69.307 5.234 ;
      RECT 69.135 5.097 69.221 5.232 ;
      RECT 69.049 5.094 69.135 5.229 ;
      RECT 68.963 5.09 69.049 5.227 ;
      RECT 68.877 5.086 68.963 5.224 ;
      RECT 68.791 5.083 68.877 5.222 ;
      RECT 68.705 5.079 68.791 5.219 ;
      RECT 68.619 5.076 68.705 5.217 ;
      RECT 68.533 5.072 68.619 5.214 ;
      RECT 68.447 5.069 68.533 5.212 ;
      RECT 68.361 5.065 68.447 5.209 ;
      RECT 68.275 5.062 68.361 5.207 ;
      RECT 68.265 5.06 68.275 5.203 ;
      RECT 68.26 5.06 68.265 5.201 ;
      RECT 68.22 5.055 68.26 5.195 ;
      RECT 68.206 5.046 68.22 5.188 ;
      RECT 68.12 5.016 68.206 5.173 ;
      RECT 68.1 4.982 68.12 5.158 ;
      RECT 68.03 4.951 68.1 5.145 ;
      RECT 68.025 4.926 68.03 5.134 ;
      RECT 68.02 4.92 68.025 5.132 ;
      RECT 67.951 4.765 68.02 5.12 ;
      RECT 67.865 4.765 67.951 5.094 ;
      RECT 67.84 4.765 67.865 5.073 ;
      RECT 67.835 4.765 67.84 5.063 ;
      RECT 67.83 4.765 67.835 5.055 ;
      RECT 67.81 4.765 67.83 5.038 ;
      RECT 70.23 3.335 70.49 3.595 ;
      RECT 70.215 3.335 70.49 3.498 ;
      RECT 70.185 3.335 70.49 3.473 ;
      RECT 70.15 3.175 70.43 3.455 ;
      RECT 70.12 4.665 70.18 4.925 ;
      RECT 69.145 3.355 69.2 3.615 ;
      RECT 70.08 4.622 70.12 4.925 ;
      RECT 70.051 4.543 70.08 4.925 ;
      RECT 69.965 4.415 70.051 4.925 ;
      RECT 69.945 4.295 69.965 4.925 ;
      RECT 69.92 4.246 69.945 4.925 ;
      RECT 69.915 4.211 69.92 4.775 ;
      RECT 69.885 4.171 69.915 4.713 ;
      RECT 69.86 4.108 69.885 4.628 ;
      RECT 69.85 4.07 69.86 4.565 ;
      RECT 69.835 4.045 69.85 4.526 ;
      RECT 69.792 4.003 69.835 4.432 ;
      RECT 69.79 3.976 69.792 4.359 ;
      RECT 69.785 3.971 69.79 4.35 ;
      RECT 69.78 3.964 69.785 4.325 ;
      RECT 69.775 3.958 69.78 4.31 ;
      RECT 69.77 3.952 69.775 4.298 ;
      RECT 69.76 3.943 69.77 4.28 ;
      RECT 69.755 3.934 69.76 4.258 ;
      RECT 69.73 3.915 69.755 4.208 ;
      RECT 69.725 3.896 69.73 4.158 ;
      RECT 69.71 3.882 69.725 4.118 ;
      RECT 69.705 3.868 69.71 4.085 ;
      RECT 69.7 3.861 69.705 4.078 ;
      RECT 69.685 3.848 69.7 4.07 ;
      RECT 69.64 3.81 69.685 4.043 ;
      RECT 69.61 3.763 69.64 4.008 ;
      RECT 69.59 3.732 69.61 3.985 ;
      RECT 69.51 3.665 69.59 3.938 ;
      RECT 69.48 3.595 69.51 3.885 ;
      RECT 69.475 3.572 69.48 3.868 ;
      RECT 69.445 3.55 69.475 3.853 ;
      RECT 69.415 3.509 69.445 3.825 ;
      RECT 69.41 3.484 69.415 3.81 ;
      RECT 69.405 3.478 69.41 3.803 ;
      RECT 69.395 3.355 69.405 3.795 ;
      RECT 69.385 3.355 69.395 3.788 ;
      RECT 69.38 3.355 69.385 3.78 ;
      RECT 69.36 3.355 69.38 3.768 ;
      RECT 69.31 3.355 69.36 3.738 ;
      RECT 69.255 3.355 69.31 3.688 ;
      RECT 69.225 3.355 69.255 3.648 ;
      RECT 69.2 3.355 69.225 3.625 ;
      RECT 69.07 4.08 69.35 4.36 ;
      RECT 69.035 3.995 69.295 4.255 ;
      RECT 69.035 4.077 69.305 4.255 ;
      RECT 67.235 3.45 67.24 3.935 ;
      RECT 67.125 3.635 67.13 3.935 ;
      RECT 67.035 3.675 67.1 3.935 ;
      RECT 68.71 3.175 68.8 3.805 ;
      RECT 68.675 3.225 68.68 3.805 ;
      RECT 68.62 3.25 68.63 3.805 ;
      RECT 68.575 3.25 68.585 3.805 ;
      RECT 68.945 3.175 68.99 3.455 ;
      RECT 67.795 2.905 67.995 3.045 ;
      RECT 68.911 3.175 68.945 3.467 ;
      RECT 68.825 3.175 68.911 3.507 ;
      RECT 68.81 3.175 68.825 3.548 ;
      RECT 68.805 3.175 68.81 3.568 ;
      RECT 68.8 3.175 68.805 3.588 ;
      RECT 68.68 3.217 68.71 3.805 ;
      RECT 68.63 3.237 68.675 3.805 ;
      RECT 68.615 3.252 68.62 3.805 ;
      RECT 68.585 3.252 68.615 3.805 ;
      RECT 68.54 3.237 68.575 3.805 ;
      RECT 68.535 3.225 68.54 3.585 ;
      RECT 68.53 3.222 68.535 3.565 ;
      RECT 68.515 3.212 68.53 3.518 ;
      RECT 68.51 3.205 68.515 3.481 ;
      RECT 68.505 3.202 68.51 3.464 ;
      RECT 68.49 3.192 68.505 3.42 ;
      RECT 68.485 3.183 68.49 3.38 ;
      RECT 68.48 3.179 68.485 3.365 ;
      RECT 68.47 3.173 68.48 3.348 ;
      RECT 68.43 3.154 68.47 3.323 ;
      RECT 68.425 3.136 68.43 3.303 ;
      RECT 68.415 3.13 68.425 3.298 ;
      RECT 68.385 3.114 68.415 3.285 ;
      RECT 68.37 3.096 68.385 3.268 ;
      RECT 68.355 3.084 68.37 3.255 ;
      RECT 68.35 3.076 68.355 3.248 ;
      RECT 68.32 3.062 68.35 3.235 ;
      RECT 68.315 3.047 68.32 3.223 ;
      RECT 68.305 3.041 68.315 3.215 ;
      RECT 68.285 3.029 68.305 3.203 ;
      RECT 68.275 3.017 68.285 3.19 ;
      RECT 68.245 3.001 68.275 3.175 ;
      RECT 68.225 2.981 68.245 3.158 ;
      RECT 68.22 2.971 68.225 3.148 ;
      RECT 68.195 2.959 68.22 3.135 ;
      RECT 68.19 2.947 68.195 3.123 ;
      RECT 68.185 2.942 68.19 3.119 ;
      RECT 68.17 2.935 68.185 3.111 ;
      RECT 68.16 2.922 68.17 3.101 ;
      RECT 68.155 2.92 68.16 3.095 ;
      RECT 68.13 2.913 68.155 3.084 ;
      RECT 68.125 2.906 68.13 3.073 ;
      RECT 68.1 2.905 68.125 3.06 ;
      RECT 68.081 2.905 68.1 3.05 ;
      RECT 67.995 2.905 68.081 3.047 ;
      RECT 67.765 2.905 67.795 3.05 ;
      RECT 67.725 2.912 67.765 3.063 ;
      RECT 67.7 2.922 67.725 3.076 ;
      RECT 67.685 2.931 67.7 3.086 ;
      RECT 67.655 2.936 67.685 3.105 ;
      RECT 67.65 2.942 67.655 3.123 ;
      RECT 67.63 2.952 67.65 3.138 ;
      RECT 67.62 2.965 67.63 3.158 ;
      RECT 67.605 2.977 67.62 3.175 ;
      RECT 67.6 2.987 67.605 3.185 ;
      RECT 67.595 2.992 67.6 3.19 ;
      RECT 67.585 3 67.595 3.203 ;
      RECT 67.535 3.032 67.585 3.24 ;
      RECT 67.52 3.067 67.535 3.281 ;
      RECT 67.515 3.077 67.52 3.296 ;
      RECT 67.51 3.082 67.515 3.303 ;
      RECT 67.485 3.098 67.51 3.323 ;
      RECT 67.47 3.119 67.485 3.348 ;
      RECT 67.445 3.14 67.47 3.373 ;
      RECT 67.435 3.159 67.445 3.396 ;
      RECT 67.41 3.177 67.435 3.419 ;
      RECT 67.395 3.197 67.41 3.443 ;
      RECT 67.39 3.207 67.395 3.455 ;
      RECT 67.375 3.219 67.39 3.475 ;
      RECT 67.365 3.234 67.375 3.515 ;
      RECT 67.36 3.242 67.365 3.543 ;
      RECT 67.35 3.252 67.36 3.563 ;
      RECT 67.345 3.265 67.35 3.588 ;
      RECT 67.34 3.278 67.345 3.608 ;
      RECT 67.335 3.284 67.34 3.63 ;
      RECT 67.325 3.293 67.335 3.65 ;
      RECT 67.32 3.313 67.325 3.673 ;
      RECT 67.315 3.319 67.32 3.693 ;
      RECT 67.31 3.326 67.315 3.715 ;
      RECT 67.305 3.337 67.31 3.728 ;
      RECT 67.295 3.347 67.305 3.753 ;
      RECT 67.275 3.372 67.295 3.935 ;
      RECT 67.245 3.412 67.275 3.935 ;
      RECT 67.24 3.442 67.245 3.935 ;
      RECT 67.215 3.47 67.235 3.935 ;
      RECT 67.185 3.515 67.215 3.935 ;
      RECT 67.18 3.542 67.185 3.935 ;
      RECT 67.16 3.56 67.18 3.935 ;
      RECT 67.15 3.585 67.16 3.935 ;
      RECT 67.145 3.597 67.15 3.935 ;
      RECT 67.13 3.62 67.145 3.935 ;
      RECT 67.11 3.647 67.125 3.935 ;
      RECT 67.1 3.67 67.11 3.935 ;
      RECT 68.89 4.555 68.97 4.815 ;
      RECT 68.125 3.775 68.195 4.035 ;
      RECT 68.856 4.522 68.89 4.815 ;
      RECT 68.77 4.425 68.856 4.815 ;
      RECT 68.75 4.337 68.77 4.815 ;
      RECT 68.74 4.307 68.75 4.815 ;
      RECT 68.73 4.287 68.74 4.815 ;
      RECT 68.71 4.274 68.73 4.815 ;
      RECT 68.695 4.264 68.71 4.643 ;
      RECT 68.69 4.257 68.695 4.598 ;
      RECT 68.68 4.251 68.69 4.588 ;
      RECT 68.67 4.243 68.68 4.57 ;
      RECT 68.665 4.237 68.67 4.558 ;
      RECT 68.655 4.232 68.665 4.545 ;
      RECT 68.635 4.222 68.655 4.518 ;
      RECT 68.595 4.201 68.635 4.47 ;
      RECT 68.58 4.182 68.595 4.428 ;
      RECT 68.555 4.168 68.58 4.398 ;
      RECT 68.545 4.156 68.555 4.365 ;
      RECT 68.54 4.151 68.545 4.355 ;
      RECT 68.51 4.137 68.54 4.335 ;
      RECT 68.5 4.121 68.51 4.308 ;
      RECT 68.495 4.116 68.5 4.298 ;
      RECT 68.47 4.107 68.495 4.278 ;
      RECT 68.46 4.095 68.47 4.258 ;
      RECT 68.39 4.063 68.46 4.233 ;
      RECT 68.385 4.032 68.39 4.21 ;
      RECT 68.336 3.775 68.385 4.193 ;
      RECT 68.25 3.775 68.336 4.152 ;
      RECT 68.195 3.775 68.25 4.08 ;
      RECT 68.285 4.56 68.445 4.82 ;
      RECT 67.81 3.175 67.86 3.86 ;
      RECT 67.6 3.6 67.635 3.86 ;
      RECT 67.915 3.175 67.92 3.635 ;
      RECT 68.005 3.175 68.03 3.455 ;
      RECT 68.28 4.557 68.285 4.82 ;
      RECT 68.245 4.545 68.28 4.82 ;
      RECT 68.185 4.518 68.245 4.82 ;
      RECT 68.18 4.501 68.185 4.674 ;
      RECT 68.175 4.498 68.18 4.661 ;
      RECT 68.155 4.491 68.175 4.648 ;
      RECT 68.12 4.474 68.155 4.63 ;
      RECT 68.08 4.453 68.12 4.61 ;
      RECT 68.075 4.441 68.08 4.598 ;
      RECT 68.035 4.427 68.075 4.584 ;
      RECT 68.015 4.41 68.035 4.566 ;
      RECT 68.005 4.402 68.015 4.558 ;
      RECT 67.99 3.175 68.005 3.473 ;
      RECT 67.975 4.392 68.005 4.545 ;
      RECT 67.96 3.175 67.99 3.518 ;
      RECT 67.965 4.382 67.975 4.532 ;
      RECT 67.935 4.367 67.965 4.519 ;
      RECT 67.92 3.175 67.96 3.585 ;
      RECT 67.92 4.335 67.935 4.505 ;
      RECT 67.915 4.307 67.92 4.499 ;
      RECT 67.91 3.175 67.915 3.64 ;
      RECT 67.9 4.277 67.915 4.493 ;
      RECT 67.905 3.175 67.91 3.653 ;
      RECT 67.895 3.175 67.905 3.673 ;
      RECT 67.86 4.19 67.9 4.478 ;
      RECT 67.86 3.175 67.895 3.713 ;
      RECT 67.855 4.122 67.86 4.466 ;
      RECT 67.84 4.077 67.855 4.461 ;
      RECT 67.835 4.015 67.84 4.456 ;
      RECT 67.81 3.922 67.835 4.449 ;
      RECT 67.805 3.175 67.81 4.441 ;
      RECT 67.79 3.175 67.805 4.428 ;
      RECT 67.77 3.175 67.79 4.385 ;
      RECT 67.76 3.175 67.77 4.335 ;
      RECT 67.755 3.175 67.76 4.308 ;
      RECT 67.75 3.175 67.755 4.286 ;
      RECT 67.745 3.401 67.75 4.269 ;
      RECT 67.74 3.423 67.745 4.247 ;
      RECT 67.735 3.465 67.74 4.23 ;
      RECT 67.705 3.515 67.735 4.174 ;
      RECT 67.7 3.542 67.705 4.116 ;
      RECT 67.685 3.56 67.7 4.08 ;
      RECT 67.68 3.578 67.685 4.044 ;
      RECT 67.674 3.585 67.68 4.025 ;
      RECT 67.67 3.592 67.674 4.008 ;
      RECT 67.665 3.597 67.67 3.977 ;
      RECT 67.655 3.6 67.665 3.952 ;
      RECT 67.645 3.6 67.655 3.918 ;
      RECT 67.64 3.6 67.645 3.895 ;
      RECT 67.635 3.6 67.64 3.875 ;
      RECT 66.55 3.735 66.83 4.015 ;
      RECT 66.55 3.735 66.85 3.91 ;
      RECT 66.64 3.625 66.9 3.885 ;
      RECT 66.605 3.72 66.9 3.885 ;
      RECT 66.73 2.24 66.895 3.885 ;
      RECT 66.63 2.24 67 2.61 ;
      RECT 66.255 4.765 66.515 5.025 ;
      RECT 66.275 4.692 66.455 5.025 ;
      RECT 66.275 4.435 66.45 5.025 ;
      RECT 66.275 4.227 66.44 5.025 ;
      RECT 66.28 4.145 66.44 5.025 ;
      RECT 66.28 3.91 66.43 5.025 ;
      RECT 66.28 3.757 66.425 5.025 ;
      RECT 66.285 3.742 66.425 5.025 ;
      RECT 66.335 3.457 66.425 5.025 ;
      RECT 66.29 3.692 66.425 5.025 ;
      RECT 66.32 3.51 66.425 5.025 ;
      RECT 66.305 3.622 66.425 5.025 ;
      RECT 66.31 3.58 66.425 5.025 ;
      RECT 66.305 3.622 66.44 3.685 ;
      RECT 66.34 3.21 66.445 3.63 ;
      RECT 66.34 3.21 66.46 3.613 ;
      RECT 66.34 3.21 66.495 3.575 ;
      RECT 66.335 3.457 66.545 3.508 ;
      RECT 66.34 3.21 66.6 3.47 ;
      RECT 65.6 3.915 65.86 4.175 ;
      RECT 65.6 3.915 65.87 4.133 ;
      RECT 65.6 3.915 65.956 4.104 ;
      RECT 65.6 3.915 66.025 4.056 ;
      RECT 65.6 3.915 66.06 4.025 ;
      RECT 65.83 3.735 66.11 4.015 ;
      RECT 65.665 3.9 66.11 4.015 ;
      RECT 65.755 3.777 65.86 4.175 ;
      RECT 65.685 3.84 66.11 4.015 ;
      RECT 60.135 8.51 60.455 8.835 ;
      RECT 60.165 7.985 60.335 8.835 ;
      RECT 60.165 7.985 60.34 8.335 ;
      RECT 60.165 7.985 61.14 8.16 ;
      RECT 60.965 3.26 61.14 8.16 ;
      RECT 60.91 3.26 61.26 3.61 ;
      RECT 60.935 8.945 61.26 9.27 ;
      RECT 59.82 9.035 61.26 9.205 ;
      RECT 59.82 3.69 59.98 9.205 ;
      RECT 60.135 3.66 60.455 3.98 ;
      RECT 59.82 3.69 60.455 3.86 ;
      RECT 58.53 4 58.87 4.35 ;
      RECT 57.925 4.065 58.87 4.265 ;
      RECT 57.925 4.06 58.14 4.265 ;
      RECT 57.94 3.635 58.14 4.265 ;
      RECT 56.93 3.635 57.21 4.015 ;
      RECT 58.62 3.995 58.79 4.35 ;
      RECT 56.925 3.635 57.21 3.968 ;
      RECT 56.905 3.635 57.21 3.945 ;
      RECT 56.895 3.635 57.21 3.925 ;
      RECT 56.885 3.635 57.21 3.91 ;
      RECT 56.86 3.635 57.21 3.883 ;
      RECT 56.85 3.635 57.21 3.858 ;
      RECT 56.805 3.59 57.085 3.85 ;
      RECT 56.805 3.635 58.14 3.835 ;
      RECT 56.805 3.63 57.13 3.85 ;
      RECT 56.805 3.622 57.125 3.85 ;
      RECT 56.805 3.612 57.12 3.85 ;
      RECT 56.805 3.6 57.115 3.85 ;
      RECT 55.73 4.295 56.01 4.575 ;
      RECT 55.73 4.295 56.045 4.555 ;
      RECT 48.01 8.945 48.36 9.295 ;
      RECT 55.475 8.9 55.825 9.25 ;
      RECT 48.01 8.975 55.825 9.175 ;
      RECT 55.765 3.715 55.815 3.975 ;
      RECT 55.555 3.715 55.56 3.975 ;
      RECT 54.75 3.27 54.78 3.53 ;
      RECT 54.52 3.27 54.595 3.53 ;
      RECT 55.74 3.665 55.765 3.975 ;
      RECT 55.735 3.622 55.74 3.975 ;
      RECT 55.73 3.605 55.735 3.975 ;
      RECT 55.725 3.592 55.73 3.975 ;
      RECT 55.65 3.475 55.725 3.975 ;
      RECT 55.605 3.292 55.65 3.975 ;
      RECT 55.6 3.22 55.605 3.975 ;
      RECT 55.585 3.195 55.6 3.975 ;
      RECT 55.56 3.157 55.585 3.975 ;
      RECT 55.55 3.137 55.56 3.697 ;
      RECT 55.535 3.129 55.55 3.652 ;
      RECT 55.53 3.121 55.535 3.623 ;
      RECT 55.525 3.118 55.53 3.603 ;
      RECT 55.52 3.115 55.525 3.583 ;
      RECT 55.515 3.112 55.52 3.563 ;
      RECT 55.485 3.101 55.515 3.5 ;
      RECT 55.465 3.086 55.485 3.415 ;
      RECT 55.46 3.078 55.465 3.378 ;
      RECT 55.45 3.072 55.46 3.345 ;
      RECT 55.435 3.064 55.45 3.305 ;
      RECT 55.43 3.057 55.435 3.265 ;
      RECT 55.425 3.054 55.43 3.243 ;
      RECT 55.42 3.051 55.425 3.23 ;
      RECT 55.415 3.05 55.42 3.22 ;
      RECT 55.4 3.044 55.415 3.21 ;
      RECT 55.375 3.031 55.4 3.195 ;
      RECT 55.325 3.006 55.375 3.166 ;
      RECT 55.31 2.985 55.325 3.141 ;
      RECT 55.3 2.978 55.31 3.13 ;
      RECT 55.245 2.959 55.3 3.103 ;
      RECT 55.22 2.937 55.245 3.076 ;
      RECT 55.215 2.93 55.22 3.071 ;
      RECT 55.2 2.93 55.215 3.069 ;
      RECT 55.175 2.922 55.2 3.065 ;
      RECT 55.16 2.92 55.175 3.061 ;
      RECT 55.13 2.92 55.16 3.058 ;
      RECT 55.12 2.92 55.13 3.053 ;
      RECT 55.075 2.92 55.12 3.051 ;
      RECT 55.046 2.92 55.075 3.052 ;
      RECT 54.96 2.92 55.046 3.054 ;
      RECT 54.946 2.921 54.96 3.056 ;
      RECT 54.86 2.922 54.946 3.058 ;
      RECT 54.845 2.923 54.86 3.068 ;
      RECT 54.84 2.924 54.845 3.077 ;
      RECT 54.82 2.927 54.84 3.087 ;
      RECT 54.805 2.935 54.82 3.102 ;
      RECT 54.785 2.953 54.805 3.117 ;
      RECT 54.775 2.965 54.785 3.14 ;
      RECT 54.765 2.974 54.775 3.17 ;
      RECT 54.75 2.986 54.765 3.215 ;
      RECT 54.695 3.019 54.75 3.53 ;
      RECT 54.69 3.047 54.695 3.53 ;
      RECT 54.67 3.062 54.69 3.53 ;
      RECT 54.635 3.122 54.67 3.53 ;
      RECT 54.633 3.172 54.635 3.53 ;
      RECT 54.63 3.18 54.633 3.53 ;
      RECT 54.62 3.195 54.63 3.53 ;
      RECT 54.615 3.207 54.62 3.53 ;
      RECT 54.605 3.232 54.615 3.53 ;
      RECT 54.595 3.26 54.605 3.53 ;
      RECT 52.5 4.765 52.55 5.025 ;
      RECT 55.41 4.315 55.47 4.575 ;
      RECT 55.395 4.315 55.41 4.585 ;
      RECT 55.376 4.315 55.395 4.618 ;
      RECT 55.29 4.315 55.376 4.743 ;
      RECT 55.21 4.315 55.29 4.925 ;
      RECT 55.205 4.552 55.21 5.01 ;
      RECT 55.18 4.622 55.205 5.038 ;
      RECT 55.175 4.692 55.18 5.065 ;
      RECT 55.155 4.764 55.175 5.087 ;
      RECT 55.15 4.831 55.155 5.11 ;
      RECT 55.14 4.86 55.15 5.125 ;
      RECT 55.13 4.882 55.14 5.142 ;
      RECT 55.125 4.892 55.13 5.153 ;
      RECT 55.12 4.9 55.125 5.161 ;
      RECT 55.11 4.908 55.12 5.173 ;
      RECT 55.105 4.92 55.11 5.183 ;
      RECT 55.1 4.928 55.105 5.188 ;
      RECT 55.08 4.946 55.1 5.198 ;
      RECT 55.075 4.963 55.08 5.205 ;
      RECT 55.07 4.971 55.075 5.206 ;
      RECT 55.065 4.982 55.07 5.208 ;
      RECT 55.025 5.02 55.065 5.218 ;
      RECT 55.02 5.055 55.025 5.229 ;
      RECT 55.015 5.06 55.02 5.232 ;
      RECT 54.99 5.07 55.015 5.239 ;
      RECT 54.98 5.084 54.99 5.248 ;
      RECT 54.96 5.096 54.98 5.251 ;
      RECT 54.91 5.115 54.96 5.255 ;
      RECT 54.865 5.13 54.91 5.26 ;
      RECT 54.8 5.133 54.865 5.266 ;
      RECT 54.785 5.131 54.8 5.273 ;
      RECT 54.755 5.13 54.785 5.273 ;
      RECT 54.716 5.129 54.755 5.269 ;
      RECT 54.63 5.126 54.716 5.265 ;
      RECT 54.613 5.124 54.63 5.262 ;
      RECT 54.527 5.122 54.613 5.259 ;
      RECT 54.441 5.119 54.527 5.253 ;
      RECT 54.355 5.115 54.441 5.248 ;
      RECT 54.277 5.112 54.355 5.244 ;
      RECT 54.191 5.109 54.277 5.242 ;
      RECT 54.105 5.106 54.191 5.239 ;
      RECT 54.047 5.104 54.105 5.236 ;
      RECT 53.961 5.101 54.047 5.234 ;
      RECT 53.875 5.097 53.961 5.232 ;
      RECT 53.789 5.094 53.875 5.229 ;
      RECT 53.703 5.09 53.789 5.227 ;
      RECT 53.617 5.086 53.703 5.224 ;
      RECT 53.531 5.083 53.617 5.222 ;
      RECT 53.445 5.079 53.531 5.219 ;
      RECT 53.359 5.076 53.445 5.217 ;
      RECT 53.273 5.072 53.359 5.214 ;
      RECT 53.187 5.069 53.273 5.212 ;
      RECT 53.101 5.065 53.187 5.209 ;
      RECT 53.015 5.062 53.101 5.207 ;
      RECT 53.005 5.06 53.015 5.203 ;
      RECT 53 5.06 53.005 5.201 ;
      RECT 52.96 5.055 53 5.195 ;
      RECT 52.946 5.046 52.96 5.188 ;
      RECT 52.86 5.016 52.946 5.173 ;
      RECT 52.84 4.982 52.86 5.158 ;
      RECT 52.77 4.951 52.84 5.145 ;
      RECT 52.765 4.926 52.77 5.134 ;
      RECT 52.76 4.92 52.765 5.132 ;
      RECT 52.691 4.765 52.76 5.12 ;
      RECT 52.605 4.765 52.691 5.094 ;
      RECT 52.58 4.765 52.605 5.073 ;
      RECT 52.575 4.765 52.58 5.063 ;
      RECT 52.57 4.765 52.575 5.055 ;
      RECT 52.55 4.765 52.57 5.038 ;
      RECT 54.97 3.335 55.23 3.595 ;
      RECT 54.955 3.335 55.23 3.498 ;
      RECT 54.925 3.335 55.23 3.473 ;
      RECT 54.89 3.175 55.17 3.455 ;
      RECT 54.86 4.665 54.92 4.925 ;
      RECT 53.885 3.355 53.94 3.615 ;
      RECT 54.82 4.622 54.86 4.925 ;
      RECT 54.791 4.543 54.82 4.925 ;
      RECT 54.705 4.415 54.791 4.925 ;
      RECT 54.685 4.295 54.705 4.925 ;
      RECT 54.66 4.246 54.685 4.925 ;
      RECT 54.655 4.211 54.66 4.775 ;
      RECT 54.625 4.171 54.655 4.713 ;
      RECT 54.6 4.108 54.625 4.628 ;
      RECT 54.59 4.07 54.6 4.565 ;
      RECT 54.575 4.045 54.59 4.526 ;
      RECT 54.532 4.003 54.575 4.432 ;
      RECT 54.53 3.976 54.532 4.359 ;
      RECT 54.525 3.971 54.53 4.35 ;
      RECT 54.52 3.964 54.525 4.325 ;
      RECT 54.515 3.958 54.52 4.31 ;
      RECT 54.51 3.952 54.515 4.298 ;
      RECT 54.5 3.943 54.51 4.28 ;
      RECT 54.495 3.934 54.5 4.258 ;
      RECT 54.47 3.915 54.495 4.208 ;
      RECT 54.465 3.896 54.47 4.158 ;
      RECT 54.45 3.882 54.465 4.118 ;
      RECT 54.445 3.868 54.45 4.085 ;
      RECT 54.44 3.861 54.445 4.078 ;
      RECT 54.425 3.848 54.44 4.07 ;
      RECT 54.38 3.81 54.425 4.043 ;
      RECT 54.35 3.763 54.38 4.008 ;
      RECT 54.33 3.732 54.35 3.985 ;
      RECT 54.25 3.665 54.33 3.938 ;
      RECT 54.22 3.595 54.25 3.885 ;
      RECT 54.215 3.572 54.22 3.868 ;
      RECT 54.185 3.55 54.215 3.853 ;
      RECT 54.155 3.509 54.185 3.825 ;
      RECT 54.15 3.484 54.155 3.81 ;
      RECT 54.145 3.478 54.15 3.803 ;
      RECT 54.135 3.355 54.145 3.795 ;
      RECT 54.125 3.355 54.135 3.788 ;
      RECT 54.12 3.355 54.125 3.78 ;
      RECT 54.1 3.355 54.12 3.768 ;
      RECT 54.05 3.355 54.1 3.738 ;
      RECT 53.995 3.355 54.05 3.688 ;
      RECT 53.965 3.355 53.995 3.648 ;
      RECT 53.94 3.355 53.965 3.625 ;
      RECT 53.81 4.08 54.09 4.36 ;
      RECT 53.775 3.995 54.035 4.255 ;
      RECT 53.775 4.077 54.045 4.255 ;
      RECT 51.975 3.45 51.98 3.935 ;
      RECT 51.865 3.635 51.87 3.935 ;
      RECT 51.775 3.675 51.84 3.935 ;
      RECT 53.45 3.175 53.54 3.805 ;
      RECT 53.415 3.225 53.42 3.805 ;
      RECT 53.36 3.25 53.37 3.805 ;
      RECT 53.315 3.25 53.325 3.805 ;
      RECT 53.685 3.175 53.73 3.455 ;
      RECT 52.535 2.905 52.735 3.045 ;
      RECT 53.651 3.175 53.685 3.467 ;
      RECT 53.565 3.175 53.651 3.507 ;
      RECT 53.55 3.175 53.565 3.548 ;
      RECT 53.545 3.175 53.55 3.568 ;
      RECT 53.54 3.175 53.545 3.588 ;
      RECT 53.42 3.217 53.45 3.805 ;
      RECT 53.37 3.237 53.415 3.805 ;
      RECT 53.355 3.252 53.36 3.805 ;
      RECT 53.325 3.252 53.355 3.805 ;
      RECT 53.28 3.237 53.315 3.805 ;
      RECT 53.275 3.225 53.28 3.585 ;
      RECT 53.27 3.222 53.275 3.565 ;
      RECT 53.255 3.212 53.27 3.518 ;
      RECT 53.25 3.205 53.255 3.481 ;
      RECT 53.245 3.202 53.25 3.464 ;
      RECT 53.23 3.192 53.245 3.42 ;
      RECT 53.225 3.183 53.23 3.38 ;
      RECT 53.22 3.179 53.225 3.365 ;
      RECT 53.21 3.173 53.22 3.348 ;
      RECT 53.17 3.154 53.21 3.323 ;
      RECT 53.165 3.136 53.17 3.303 ;
      RECT 53.155 3.13 53.165 3.298 ;
      RECT 53.125 3.114 53.155 3.285 ;
      RECT 53.11 3.096 53.125 3.268 ;
      RECT 53.095 3.084 53.11 3.255 ;
      RECT 53.09 3.076 53.095 3.248 ;
      RECT 53.06 3.062 53.09 3.235 ;
      RECT 53.055 3.047 53.06 3.223 ;
      RECT 53.045 3.041 53.055 3.215 ;
      RECT 53.025 3.029 53.045 3.203 ;
      RECT 53.015 3.017 53.025 3.19 ;
      RECT 52.985 3.001 53.015 3.175 ;
      RECT 52.965 2.981 52.985 3.158 ;
      RECT 52.96 2.971 52.965 3.148 ;
      RECT 52.935 2.959 52.96 3.135 ;
      RECT 52.93 2.947 52.935 3.123 ;
      RECT 52.925 2.942 52.93 3.119 ;
      RECT 52.91 2.935 52.925 3.111 ;
      RECT 52.9 2.922 52.91 3.101 ;
      RECT 52.895 2.92 52.9 3.095 ;
      RECT 52.87 2.913 52.895 3.084 ;
      RECT 52.865 2.906 52.87 3.073 ;
      RECT 52.84 2.905 52.865 3.06 ;
      RECT 52.821 2.905 52.84 3.05 ;
      RECT 52.735 2.905 52.821 3.047 ;
      RECT 52.505 2.905 52.535 3.05 ;
      RECT 52.465 2.912 52.505 3.063 ;
      RECT 52.44 2.922 52.465 3.076 ;
      RECT 52.425 2.931 52.44 3.086 ;
      RECT 52.395 2.936 52.425 3.105 ;
      RECT 52.39 2.942 52.395 3.123 ;
      RECT 52.37 2.952 52.39 3.138 ;
      RECT 52.36 2.965 52.37 3.158 ;
      RECT 52.345 2.977 52.36 3.175 ;
      RECT 52.34 2.987 52.345 3.185 ;
      RECT 52.335 2.992 52.34 3.19 ;
      RECT 52.325 3 52.335 3.203 ;
      RECT 52.275 3.032 52.325 3.24 ;
      RECT 52.26 3.067 52.275 3.281 ;
      RECT 52.255 3.077 52.26 3.296 ;
      RECT 52.25 3.082 52.255 3.303 ;
      RECT 52.225 3.098 52.25 3.323 ;
      RECT 52.21 3.119 52.225 3.348 ;
      RECT 52.185 3.14 52.21 3.373 ;
      RECT 52.175 3.159 52.185 3.396 ;
      RECT 52.15 3.177 52.175 3.419 ;
      RECT 52.135 3.197 52.15 3.443 ;
      RECT 52.13 3.207 52.135 3.455 ;
      RECT 52.115 3.219 52.13 3.475 ;
      RECT 52.105 3.234 52.115 3.515 ;
      RECT 52.1 3.242 52.105 3.543 ;
      RECT 52.09 3.252 52.1 3.563 ;
      RECT 52.085 3.265 52.09 3.588 ;
      RECT 52.08 3.278 52.085 3.608 ;
      RECT 52.075 3.284 52.08 3.63 ;
      RECT 52.065 3.293 52.075 3.65 ;
      RECT 52.06 3.313 52.065 3.673 ;
      RECT 52.055 3.319 52.06 3.693 ;
      RECT 52.05 3.326 52.055 3.715 ;
      RECT 52.045 3.337 52.05 3.728 ;
      RECT 52.035 3.347 52.045 3.753 ;
      RECT 52.015 3.372 52.035 3.935 ;
      RECT 51.985 3.412 52.015 3.935 ;
      RECT 51.98 3.442 51.985 3.935 ;
      RECT 51.955 3.47 51.975 3.935 ;
      RECT 51.925 3.515 51.955 3.935 ;
      RECT 51.92 3.542 51.925 3.935 ;
      RECT 51.9 3.56 51.92 3.935 ;
      RECT 51.89 3.585 51.9 3.935 ;
      RECT 51.885 3.597 51.89 3.935 ;
      RECT 51.87 3.62 51.885 3.935 ;
      RECT 51.85 3.647 51.865 3.935 ;
      RECT 51.84 3.67 51.85 3.935 ;
      RECT 53.63 4.555 53.71 4.815 ;
      RECT 52.865 3.775 52.935 4.035 ;
      RECT 53.596 4.522 53.63 4.815 ;
      RECT 53.51 4.425 53.596 4.815 ;
      RECT 53.49 4.337 53.51 4.815 ;
      RECT 53.48 4.307 53.49 4.815 ;
      RECT 53.47 4.287 53.48 4.815 ;
      RECT 53.45 4.274 53.47 4.815 ;
      RECT 53.435 4.264 53.45 4.643 ;
      RECT 53.43 4.257 53.435 4.598 ;
      RECT 53.42 4.251 53.43 4.588 ;
      RECT 53.41 4.243 53.42 4.57 ;
      RECT 53.405 4.237 53.41 4.558 ;
      RECT 53.395 4.232 53.405 4.545 ;
      RECT 53.375 4.222 53.395 4.518 ;
      RECT 53.335 4.201 53.375 4.47 ;
      RECT 53.32 4.182 53.335 4.428 ;
      RECT 53.295 4.168 53.32 4.398 ;
      RECT 53.285 4.156 53.295 4.365 ;
      RECT 53.28 4.151 53.285 4.355 ;
      RECT 53.25 4.137 53.28 4.335 ;
      RECT 53.24 4.121 53.25 4.308 ;
      RECT 53.235 4.116 53.24 4.298 ;
      RECT 53.21 4.107 53.235 4.278 ;
      RECT 53.2 4.095 53.21 4.258 ;
      RECT 53.13 4.063 53.2 4.233 ;
      RECT 53.125 4.032 53.13 4.21 ;
      RECT 53.076 3.775 53.125 4.193 ;
      RECT 52.99 3.775 53.076 4.152 ;
      RECT 52.935 3.775 52.99 4.08 ;
      RECT 53.025 4.56 53.185 4.82 ;
      RECT 52.55 3.175 52.6 3.86 ;
      RECT 52.34 3.6 52.375 3.86 ;
      RECT 52.655 3.175 52.66 3.635 ;
      RECT 52.745 3.175 52.77 3.455 ;
      RECT 53.02 4.557 53.025 4.82 ;
      RECT 52.985 4.545 53.02 4.82 ;
      RECT 52.925 4.518 52.985 4.82 ;
      RECT 52.92 4.501 52.925 4.674 ;
      RECT 52.915 4.498 52.92 4.661 ;
      RECT 52.895 4.491 52.915 4.648 ;
      RECT 52.86 4.474 52.895 4.63 ;
      RECT 52.82 4.453 52.86 4.61 ;
      RECT 52.815 4.441 52.82 4.598 ;
      RECT 52.775 4.427 52.815 4.584 ;
      RECT 52.755 4.41 52.775 4.566 ;
      RECT 52.745 4.402 52.755 4.558 ;
      RECT 52.73 3.175 52.745 3.473 ;
      RECT 52.715 4.392 52.745 4.545 ;
      RECT 52.7 3.175 52.73 3.518 ;
      RECT 52.705 4.382 52.715 4.532 ;
      RECT 52.675 4.367 52.705 4.519 ;
      RECT 52.66 3.175 52.7 3.585 ;
      RECT 52.66 4.335 52.675 4.505 ;
      RECT 52.655 4.307 52.66 4.499 ;
      RECT 52.65 3.175 52.655 3.64 ;
      RECT 52.64 4.277 52.655 4.493 ;
      RECT 52.645 3.175 52.65 3.653 ;
      RECT 52.635 3.175 52.645 3.673 ;
      RECT 52.6 4.19 52.64 4.478 ;
      RECT 52.6 3.175 52.635 3.713 ;
      RECT 52.595 4.122 52.6 4.466 ;
      RECT 52.58 4.077 52.595 4.461 ;
      RECT 52.575 4.015 52.58 4.456 ;
      RECT 52.55 3.922 52.575 4.449 ;
      RECT 52.545 3.175 52.55 4.441 ;
      RECT 52.53 3.175 52.545 4.428 ;
      RECT 52.51 3.175 52.53 4.385 ;
      RECT 52.5 3.175 52.51 4.335 ;
      RECT 52.495 3.175 52.5 4.308 ;
      RECT 52.49 3.175 52.495 4.286 ;
      RECT 52.485 3.401 52.49 4.269 ;
      RECT 52.48 3.423 52.485 4.247 ;
      RECT 52.475 3.465 52.48 4.23 ;
      RECT 52.445 3.515 52.475 4.174 ;
      RECT 52.44 3.542 52.445 4.116 ;
      RECT 52.425 3.56 52.44 4.08 ;
      RECT 52.42 3.578 52.425 4.044 ;
      RECT 52.414 3.585 52.42 4.025 ;
      RECT 52.41 3.592 52.414 4.008 ;
      RECT 52.405 3.597 52.41 3.977 ;
      RECT 52.395 3.6 52.405 3.952 ;
      RECT 52.385 3.6 52.395 3.918 ;
      RECT 52.38 3.6 52.385 3.895 ;
      RECT 52.375 3.6 52.38 3.875 ;
      RECT 51.29 3.735 51.57 4.015 ;
      RECT 51.29 3.735 51.59 3.91 ;
      RECT 51.38 3.625 51.64 3.885 ;
      RECT 51.345 3.72 51.64 3.885 ;
      RECT 51.47 2.24 51.635 3.885 ;
      RECT 51.37 2.24 51.74 2.61 ;
      RECT 50.995 4.765 51.255 5.025 ;
      RECT 51.015 4.692 51.195 5.025 ;
      RECT 51.015 4.435 51.19 5.025 ;
      RECT 51.015 4.227 51.18 5.025 ;
      RECT 51.02 4.145 51.18 5.025 ;
      RECT 51.02 3.91 51.17 5.025 ;
      RECT 51.02 3.757 51.165 5.025 ;
      RECT 51.025 3.742 51.165 5.025 ;
      RECT 51.075 3.457 51.165 5.025 ;
      RECT 51.03 3.692 51.165 5.025 ;
      RECT 51.06 3.51 51.165 5.025 ;
      RECT 51.045 3.622 51.165 5.025 ;
      RECT 51.05 3.58 51.165 5.025 ;
      RECT 51.045 3.622 51.18 3.685 ;
      RECT 51.08 3.21 51.185 3.63 ;
      RECT 51.08 3.21 51.2 3.613 ;
      RECT 51.08 3.21 51.235 3.575 ;
      RECT 51.075 3.457 51.285 3.508 ;
      RECT 51.08 3.21 51.34 3.47 ;
      RECT 50.34 3.915 50.6 4.175 ;
      RECT 50.34 3.915 50.61 4.133 ;
      RECT 50.34 3.915 50.696 4.104 ;
      RECT 50.34 3.915 50.765 4.056 ;
      RECT 50.34 3.915 50.8 4.025 ;
      RECT 50.57 3.735 50.85 4.015 ;
      RECT 50.405 3.9 50.85 4.015 ;
      RECT 50.495 3.777 50.6 4.175 ;
      RECT 50.425 3.84 50.85 4.015 ;
      RECT 44.875 8.51 45.195 8.835 ;
      RECT 44.905 7.985 45.075 8.835 ;
      RECT 44.905 7.985 45.08 8.335 ;
      RECT 44.905 7.985 45.88 8.16 ;
      RECT 45.705 3.26 45.88 8.16 ;
      RECT 45.65 3.26 46 3.61 ;
      RECT 45.675 8.945 46 9.27 ;
      RECT 44.56 9.035 46 9.205 ;
      RECT 44.56 3.69 44.72 9.205 ;
      RECT 44.875 3.66 45.195 3.98 ;
      RECT 44.56 3.69 45.195 3.86 ;
      RECT 43.27 4 43.61 4.35 ;
      RECT 42.665 4.065 43.61 4.265 ;
      RECT 42.665 4.06 42.88 4.265 ;
      RECT 42.68 3.635 42.88 4.265 ;
      RECT 41.67 3.635 41.95 4.015 ;
      RECT 43.36 3.995 43.53 4.35 ;
      RECT 41.665 3.635 41.95 3.968 ;
      RECT 41.645 3.635 41.95 3.945 ;
      RECT 41.635 3.635 41.95 3.925 ;
      RECT 41.625 3.635 41.95 3.91 ;
      RECT 41.6 3.635 41.95 3.883 ;
      RECT 41.59 3.635 41.95 3.858 ;
      RECT 41.545 3.59 41.825 3.85 ;
      RECT 41.545 3.635 42.88 3.835 ;
      RECT 41.545 3.63 41.87 3.85 ;
      RECT 41.545 3.622 41.865 3.85 ;
      RECT 41.545 3.612 41.86 3.85 ;
      RECT 41.545 3.6 41.855 3.85 ;
      RECT 40.47 4.295 40.75 4.575 ;
      RECT 40.47 4.295 40.785 4.555 ;
      RECT 32.795 8.95 33.145 9.3 ;
      RECT 40.215 8.905 40.565 9.255 ;
      RECT 32.795 8.98 40.565 9.18 ;
      RECT 40.505 3.715 40.555 3.975 ;
      RECT 40.295 3.715 40.3 3.975 ;
      RECT 39.49 3.27 39.52 3.53 ;
      RECT 39.26 3.27 39.335 3.53 ;
      RECT 40.48 3.665 40.505 3.975 ;
      RECT 40.475 3.622 40.48 3.975 ;
      RECT 40.47 3.605 40.475 3.975 ;
      RECT 40.465 3.592 40.47 3.975 ;
      RECT 40.39 3.475 40.465 3.975 ;
      RECT 40.345 3.292 40.39 3.975 ;
      RECT 40.34 3.22 40.345 3.975 ;
      RECT 40.325 3.195 40.34 3.975 ;
      RECT 40.3 3.157 40.325 3.975 ;
      RECT 40.29 3.137 40.3 3.697 ;
      RECT 40.275 3.129 40.29 3.652 ;
      RECT 40.27 3.121 40.275 3.623 ;
      RECT 40.265 3.118 40.27 3.603 ;
      RECT 40.26 3.115 40.265 3.583 ;
      RECT 40.255 3.112 40.26 3.563 ;
      RECT 40.225 3.101 40.255 3.5 ;
      RECT 40.205 3.086 40.225 3.415 ;
      RECT 40.2 3.078 40.205 3.378 ;
      RECT 40.19 3.072 40.2 3.345 ;
      RECT 40.175 3.064 40.19 3.305 ;
      RECT 40.17 3.057 40.175 3.265 ;
      RECT 40.165 3.054 40.17 3.243 ;
      RECT 40.16 3.051 40.165 3.23 ;
      RECT 40.155 3.05 40.16 3.22 ;
      RECT 40.14 3.044 40.155 3.21 ;
      RECT 40.115 3.031 40.14 3.195 ;
      RECT 40.065 3.006 40.115 3.166 ;
      RECT 40.05 2.985 40.065 3.141 ;
      RECT 40.04 2.978 40.05 3.13 ;
      RECT 39.985 2.959 40.04 3.103 ;
      RECT 39.96 2.937 39.985 3.076 ;
      RECT 39.955 2.93 39.96 3.071 ;
      RECT 39.94 2.93 39.955 3.069 ;
      RECT 39.915 2.922 39.94 3.065 ;
      RECT 39.9 2.92 39.915 3.061 ;
      RECT 39.87 2.92 39.9 3.058 ;
      RECT 39.86 2.92 39.87 3.053 ;
      RECT 39.815 2.92 39.86 3.051 ;
      RECT 39.786 2.92 39.815 3.052 ;
      RECT 39.7 2.92 39.786 3.054 ;
      RECT 39.686 2.921 39.7 3.056 ;
      RECT 39.6 2.922 39.686 3.058 ;
      RECT 39.585 2.923 39.6 3.068 ;
      RECT 39.58 2.924 39.585 3.077 ;
      RECT 39.56 2.927 39.58 3.087 ;
      RECT 39.545 2.935 39.56 3.102 ;
      RECT 39.525 2.953 39.545 3.117 ;
      RECT 39.515 2.965 39.525 3.14 ;
      RECT 39.505 2.974 39.515 3.17 ;
      RECT 39.49 2.986 39.505 3.215 ;
      RECT 39.435 3.019 39.49 3.53 ;
      RECT 39.43 3.047 39.435 3.53 ;
      RECT 39.41 3.062 39.43 3.53 ;
      RECT 39.375 3.122 39.41 3.53 ;
      RECT 39.373 3.172 39.375 3.53 ;
      RECT 39.37 3.18 39.373 3.53 ;
      RECT 39.36 3.195 39.37 3.53 ;
      RECT 39.355 3.207 39.36 3.53 ;
      RECT 39.345 3.232 39.355 3.53 ;
      RECT 39.335 3.26 39.345 3.53 ;
      RECT 37.24 4.765 37.29 5.025 ;
      RECT 40.15 4.315 40.21 4.575 ;
      RECT 40.135 4.315 40.15 4.585 ;
      RECT 40.116 4.315 40.135 4.618 ;
      RECT 40.03 4.315 40.116 4.743 ;
      RECT 39.95 4.315 40.03 4.925 ;
      RECT 39.945 4.552 39.95 5.01 ;
      RECT 39.92 4.622 39.945 5.038 ;
      RECT 39.915 4.692 39.92 5.065 ;
      RECT 39.895 4.764 39.915 5.087 ;
      RECT 39.89 4.831 39.895 5.11 ;
      RECT 39.88 4.86 39.89 5.125 ;
      RECT 39.87 4.882 39.88 5.142 ;
      RECT 39.865 4.892 39.87 5.153 ;
      RECT 39.86 4.9 39.865 5.161 ;
      RECT 39.85 4.908 39.86 5.173 ;
      RECT 39.845 4.92 39.85 5.183 ;
      RECT 39.84 4.928 39.845 5.188 ;
      RECT 39.82 4.946 39.84 5.198 ;
      RECT 39.815 4.963 39.82 5.205 ;
      RECT 39.81 4.971 39.815 5.206 ;
      RECT 39.805 4.982 39.81 5.208 ;
      RECT 39.765 5.02 39.805 5.218 ;
      RECT 39.76 5.055 39.765 5.229 ;
      RECT 39.755 5.06 39.76 5.232 ;
      RECT 39.73 5.07 39.755 5.239 ;
      RECT 39.72 5.084 39.73 5.248 ;
      RECT 39.7 5.096 39.72 5.251 ;
      RECT 39.65 5.115 39.7 5.255 ;
      RECT 39.605 5.13 39.65 5.26 ;
      RECT 39.54 5.133 39.605 5.266 ;
      RECT 39.525 5.131 39.54 5.273 ;
      RECT 39.495 5.13 39.525 5.273 ;
      RECT 39.456 5.129 39.495 5.269 ;
      RECT 39.37 5.126 39.456 5.265 ;
      RECT 39.353 5.124 39.37 5.262 ;
      RECT 39.267 5.122 39.353 5.259 ;
      RECT 39.181 5.119 39.267 5.253 ;
      RECT 39.095 5.115 39.181 5.248 ;
      RECT 39.017 5.112 39.095 5.244 ;
      RECT 38.931 5.109 39.017 5.242 ;
      RECT 38.845 5.106 38.931 5.239 ;
      RECT 38.787 5.104 38.845 5.236 ;
      RECT 38.701 5.101 38.787 5.234 ;
      RECT 38.615 5.097 38.701 5.232 ;
      RECT 38.529 5.094 38.615 5.229 ;
      RECT 38.443 5.09 38.529 5.227 ;
      RECT 38.357 5.086 38.443 5.224 ;
      RECT 38.271 5.083 38.357 5.222 ;
      RECT 38.185 5.079 38.271 5.219 ;
      RECT 38.099 5.076 38.185 5.217 ;
      RECT 38.013 5.072 38.099 5.214 ;
      RECT 37.927 5.069 38.013 5.212 ;
      RECT 37.841 5.065 37.927 5.209 ;
      RECT 37.755 5.062 37.841 5.207 ;
      RECT 37.745 5.06 37.755 5.203 ;
      RECT 37.74 5.06 37.745 5.201 ;
      RECT 37.7 5.055 37.74 5.195 ;
      RECT 37.686 5.046 37.7 5.188 ;
      RECT 37.6 5.016 37.686 5.173 ;
      RECT 37.58 4.982 37.6 5.158 ;
      RECT 37.51 4.951 37.58 5.145 ;
      RECT 37.505 4.926 37.51 5.134 ;
      RECT 37.5 4.92 37.505 5.132 ;
      RECT 37.431 4.765 37.5 5.12 ;
      RECT 37.345 4.765 37.431 5.094 ;
      RECT 37.32 4.765 37.345 5.073 ;
      RECT 37.315 4.765 37.32 5.063 ;
      RECT 37.31 4.765 37.315 5.055 ;
      RECT 37.29 4.765 37.31 5.038 ;
      RECT 39.71 3.335 39.97 3.595 ;
      RECT 39.695 3.335 39.97 3.498 ;
      RECT 39.665 3.335 39.97 3.473 ;
      RECT 39.63 3.175 39.91 3.455 ;
      RECT 39.6 4.665 39.66 4.925 ;
      RECT 38.625 3.355 38.68 3.615 ;
      RECT 39.56 4.622 39.6 4.925 ;
      RECT 39.531 4.543 39.56 4.925 ;
      RECT 39.445 4.415 39.531 4.925 ;
      RECT 39.425 4.295 39.445 4.925 ;
      RECT 39.4 4.246 39.425 4.925 ;
      RECT 39.395 4.211 39.4 4.775 ;
      RECT 39.365 4.171 39.395 4.713 ;
      RECT 39.34 4.108 39.365 4.628 ;
      RECT 39.33 4.07 39.34 4.565 ;
      RECT 39.315 4.045 39.33 4.526 ;
      RECT 39.272 4.003 39.315 4.432 ;
      RECT 39.27 3.976 39.272 4.359 ;
      RECT 39.265 3.971 39.27 4.35 ;
      RECT 39.26 3.964 39.265 4.325 ;
      RECT 39.255 3.958 39.26 4.31 ;
      RECT 39.25 3.952 39.255 4.298 ;
      RECT 39.24 3.943 39.25 4.28 ;
      RECT 39.235 3.934 39.24 4.258 ;
      RECT 39.21 3.915 39.235 4.208 ;
      RECT 39.205 3.896 39.21 4.158 ;
      RECT 39.19 3.882 39.205 4.118 ;
      RECT 39.185 3.868 39.19 4.085 ;
      RECT 39.18 3.861 39.185 4.078 ;
      RECT 39.165 3.848 39.18 4.07 ;
      RECT 39.12 3.81 39.165 4.043 ;
      RECT 39.09 3.763 39.12 4.008 ;
      RECT 39.07 3.732 39.09 3.985 ;
      RECT 38.99 3.665 39.07 3.938 ;
      RECT 38.96 3.595 38.99 3.885 ;
      RECT 38.955 3.572 38.96 3.868 ;
      RECT 38.925 3.55 38.955 3.853 ;
      RECT 38.895 3.509 38.925 3.825 ;
      RECT 38.89 3.484 38.895 3.81 ;
      RECT 38.885 3.478 38.89 3.803 ;
      RECT 38.875 3.355 38.885 3.795 ;
      RECT 38.865 3.355 38.875 3.788 ;
      RECT 38.86 3.355 38.865 3.78 ;
      RECT 38.84 3.355 38.86 3.768 ;
      RECT 38.79 3.355 38.84 3.738 ;
      RECT 38.735 3.355 38.79 3.688 ;
      RECT 38.705 3.355 38.735 3.648 ;
      RECT 38.68 3.355 38.705 3.625 ;
      RECT 38.55 4.08 38.83 4.36 ;
      RECT 38.515 3.995 38.775 4.255 ;
      RECT 38.515 4.077 38.785 4.255 ;
      RECT 36.715 3.45 36.72 3.935 ;
      RECT 36.605 3.635 36.61 3.935 ;
      RECT 36.515 3.675 36.58 3.935 ;
      RECT 38.19 3.175 38.28 3.805 ;
      RECT 38.155 3.225 38.16 3.805 ;
      RECT 38.1 3.25 38.11 3.805 ;
      RECT 38.055 3.25 38.065 3.805 ;
      RECT 38.425 3.175 38.47 3.455 ;
      RECT 37.275 2.905 37.475 3.045 ;
      RECT 38.391 3.175 38.425 3.467 ;
      RECT 38.305 3.175 38.391 3.507 ;
      RECT 38.29 3.175 38.305 3.548 ;
      RECT 38.285 3.175 38.29 3.568 ;
      RECT 38.28 3.175 38.285 3.588 ;
      RECT 38.16 3.217 38.19 3.805 ;
      RECT 38.11 3.237 38.155 3.805 ;
      RECT 38.095 3.252 38.1 3.805 ;
      RECT 38.065 3.252 38.095 3.805 ;
      RECT 38.02 3.237 38.055 3.805 ;
      RECT 38.015 3.225 38.02 3.585 ;
      RECT 38.01 3.222 38.015 3.565 ;
      RECT 37.995 3.212 38.01 3.518 ;
      RECT 37.99 3.205 37.995 3.481 ;
      RECT 37.985 3.202 37.99 3.464 ;
      RECT 37.97 3.192 37.985 3.42 ;
      RECT 37.965 3.183 37.97 3.38 ;
      RECT 37.96 3.179 37.965 3.365 ;
      RECT 37.95 3.173 37.96 3.348 ;
      RECT 37.91 3.154 37.95 3.323 ;
      RECT 37.905 3.136 37.91 3.303 ;
      RECT 37.895 3.13 37.905 3.298 ;
      RECT 37.865 3.114 37.895 3.285 ;
      RECT 37.85 3.096 37.865 3.268 ;
      RECT 37.835 3.084 37.85 3.255 ;
      RECT 37.83 3.076 37.835 3.248 ;
      RECT 37.8 3.062 37.83 3.235 ;
      RECT 37.795 3.047 37.8 3.223 ;
      RECT 37.785 3.041 37.795 3.215 ;
      RECT 37.765 3.029 37.785 3.203 ;
      RECT 37.755 3.017 37.765 3.19 ;
      RECT 37.725 3.001 37.755 3.175 ;
      RECT 37.705 2.981 37.725 3.158 ;
      RECT 37.7 2.971 37.705 3.148 ;
      RECT 37.675 2.959 37.7 3.135 ;
      RECT 37.67 2.947 37.675 3.123 ;
      RECT 37.665 2.942 37.67 3.119 ;
      RECT 37.65 2.935 37.665 3.111 ;
      RECT 37.64 2.922 37.65 3.101 ;
      RECT 37.635 2.92 37.64 3.095 ;
      RECT 37.61 2.913 37.635 3.084 ;
      RECT 37.605 2.906 37.61 3.073 ;
      RECT 37.58 2.905 37.605 3.06 ;
      RECT 37.561 2.905 37.58 3.05 ;
      RECT 37.475 2.905 37.561 3.047 ;
      RECT 37.245 2.905 37.275 3.05 ;
      RECT 37.205 2.912 37.245 3.063 ;
      RECT 37.18 2.922 37.205 3.076 ;
      RECT 37.165 2.931 37.18 3.086 ;
      RECT 37.135 2.936 37.165 3.105 ;
      RECT 37.13 2.942 37.135 3.123 ;
      RECT 37.11 2.952 37.13 3.138 ;
      RECT 37.1 2.965 37.11 3.158 ;
      RECT 37.085 2.977 37.1 3.175 ;
      RECT 37.08 2.987 37.085 3.185 ;
      RECT 37.075 2.992 37.08 3.19 ;
      RECT 37.065 3 37.075 3.203 ;
      RECT 37.015 3.032 37.065 3.24 ;
      RECT 37 3.067 37.015 3.281 ;
      RECT 36.995 3.077 37 3.296 ;
      RECT 36.99 3.082 36.995 3.303 ;
      RECT 36.965 3.098 36.99 3.323 ;
      RECT 36.95 3.119 36.965 3.348 ;
      RECT 36.925 3.14 36.95 3.373 ;
      RECT 36.915 3.159 36.925 3.396 ;
      RECT 36.89 3.177 36.915 3.419 ;
      RECT 36.875 3.197 36.89 3.443 ;
      RECT 36.87 3.207 36.875 3.455 ;
      RECT 36.855 3.219 36.87 3.475 ;
      RECT 36.845 3.234 36.855 3.515 ;
      RECT 36.84 3.242 36.845 3.543 ;
      RECT 36.83 3.252 36.84 3.563 ;
      RECT 36.825 3.265 36.83 3.588 ;
      RECT 36.82 3.278 36.825 3.608 ;
      RECT 36.815 3.284 36.82 3.63 ;
      RECT 36.805 3.293 36.815 3.65 ;
      RECT 36.8 3.313 36.805 3.673 ;
      RECT 36.795 3.319 36.8 3.693 ;
      RECT 36.79 3.326 36.795 3.715 ;
      RECT 36.785 3.337 36.79 3.728 ;
      RECT 36.775 3.347 36.785 3.753 ;
      RECT 36.755 3.372 36.775 3.935 ;
      RECT 36.725 3.412 36.755 3.935 ;
      RECT 36.72 3.442 36.725 3.935 ;
      RECT 36.695 3.47 36.715 3.935 ;
      RECT 36.665 3.515 36.695 3.935 ;
      RECT 36.66 3.542 36.665 3.935 ;
      RECT 36.64 3.56 36.66 3.935 ;
      RECT 36.63 3.585 36.64 3.935 ;
      RECT 36.625 3.597 36.63 3.935 ;
      RECT 36.61 3.62 36.625 3.935 ;
      RECT 36.59 3.647 36.605 3.935 ;
      RECT 36.58 3.67 36.59 3.935 ;
      RECT 38.37 4.555 38.45 4.815 ;
      RECT 37.605 3.775 37.675 4.035 ;
      RECT 38.336 4.522 38.37 4.815 ;
      RECT 38.25 4.425 38.336 4.815 ;
      RECT 38.23 4.337 38.25 4.815 ;
      RECT 38.22 4.307 38.23 4.815 ;
      RECT 38.21 4.287 38.22 4.815 ;
      RECT 38.19 4.274 38.21 4.815 ;
      RECT 38.175 4.264 38.19 4.643 ;
      RECT 38.17 4.257 38.175 4.598 ;
      RECT 38.16 4.251 38.17 4.588 ;
      RECT 38.15 4.243 38.16 4.57 ;
      RECT 38.145 4.237 38.15 4.558 ;
      RECT 38.135 4.232 38.145 4.545 ;
      RECT 38.115 4.222 38.135 4.518 ;
      RECT 38.075 4.201 38.115 4.47 ;
      RECT 38.06 4.182 38.075 4.428 ;
      RECT 38.035 4.168 38.06 4.398 ;
      RECT 38.025 4.156 38.035 4.365 ;
      RECT 38.02 4.151 38.025 4.355 ;
      RECT 37.99 4.137 38.02 4.335 ;
      RECT 37.98 4.121 37.99 4.308 ;
      RECT 37.975 4.116 37.98 4.298 ;
      RECT 37.95 4.107 37.975 4.278 ;
      RECT 37.94 4.095 37.95 4.258 ;
      RECT 37.87 4.063 37.94 4.233 ;
      RECT 37.865 4.032 37.87 4.21 ;
      RECT 37.816 3.775 37.865 4.193 ;
      RECT 37.73 3.775 37.816 4.152 ;
      RECT 37.675 3.775 37.73 4.08 ;
      RECT 37.765 4.56 37.925 4.82 ;
      RECT 37.29 3.175 37.34 3.86 ;
      RECT 37.08 3.6 37.115 3.86 ;
      RECT 37.395 3.175 37.4 3.635 ;
      RECT 37.485 3.175 37.51 3.455 ;
      RECT 37.76 4.557 37.765 4.82 ;
      RECT 37.725 4.545 37.76 4.82 ;
      RECT 37.665 4.518 37.725 4.82 ;
      RECT 37.66 4.501 37.665 4.674 ;
      RECT 37.655 4.498 37.66 4.661 ;
      RECT 37.635 4.491 37.655 4.648 ;
      RECT 37.6 4.474 37.635 4.63 ;
      RECT 37.56 4.453 37.6 4.61 ;
      RECT 37.555 4.441 37.56 4.598 ;
      RECT 37.515 4.427 37.555 4.584 ;
      RECT 37.495 4.41 37.515 4.566 ;
      RECT 37.485 4.402 37.495 4.558 ;
      RECT 37.47 3.175 37.485 3.473 ;
      RECT 37.455 4.392 37.485 4.545 ;
      RECT 37.44 3.175 37.47 3.518 ;
      RECT 37.445 4.382 37.455 4.532 ;
      RECT 37.415 4.367 37.445 4.519 ;
      RECT 37.4 3.175 37.44 3.585 ;
      RECT 37.4 4.335 37.415 4.505 ;
      RECT 37.395 4.307 37.4 4.499 ;
      RECT 37.39 3.175 37.395 3.64 ;
      RECT 37.38 4.277 37.395 4.493 ;
      RECT 37.385 3.175 37.39 3.653 ;
      RECT 37.375 3.175 37.385 3.673 ;
      RECT 37.34 4.19 37.38 4.478 ;
      RECT 37.34 3.175 37.375 3.713 ;
      RECT 37.335 4.122 37.34 4.466 ;
      RECT 37.32 4.077 37.335 4.461 ;
      RECT 37.315 4.015 37.32 4.456 ;
      RECT 37.29 3.922 37.315 4.449 ;
      RECT 37.285 3.175 37.29 4.441 ;
      RECT 37.27 3.175 37.285 4.428 ;
      RECT 37.25 3.175 37.27 4.385 ;
      RECT 37.24 3.175 37.25 4.335 ;
      RECT 37.235 3.175 37.24 4.308 ;
      RECT 37.23 3.175 37.235 4.286 ;
      RECT 37.225 3.401 37.23 4.269 ;
      RECT 37.22 3.423 37.225 4.247 ;
      RECT 37.215 3.465 37.22 4.23 ;
      RECT 37.185 3.515 37.215 4.174 ;
      RECT 37.18 3.542 37.185 4.116 ;
      RECT 37.165 3.56 37.18 4.08 ;
      RECT 37.16 3.578 37.165 4.044 ;
      RECT 37.154 3.585 37.16 4.025 ;
      RECT 37.15 3.592 37.154 4.008 ;
      RECT 37.145 3.597 37.15 3.977 ;
      RECT 37.135 3.6 37.145 3.952 ;
      RECT 37.125 3.6 37.135 3.918 ;
      RECT 37.12 3.6 37.125 3.895 ;
      RECT 37.115 3.6 37.12 3.875 ;
      RECT 36.03 3.735 36.31 4.015 ;
      RECT 36.03 3.735 36.33 3.91 ;
      RECT 36.12 3.625 36.38 3.885 ;
      RECT 36.085 3.72 36.38 3.885 ;
      RECT 36.21 2.24 36.375 3.885 ;
      RECT 36.11 2.24 36.48 2.61 ;
      RECT 35.735 4.765 35.995 5.025 ;
      RECT 35.755 4.692 35.935 5.025 ;
      RECT 35.755 4.435 35.93 5.025 ;
      RECT 35.755 4.227 35.92 5.025 ;
      RECT 35.76 4.145 35.92 5.025 ;
      RECT 35.76 3.91 35.91 5.025 ;
      RECT 35.76 3.757 35.905 5.025 ;
      RECT 35.765 3.742 35.905 5.025 ;
      RECT 35.815 3.457 35.905 5.025 ;
      RECT 35.77 3.692 35.905 5.025 ;
      RECT 35.8 3.51 35.905 5.025 ;
      RECT 35.785 3.622 35.905 5.025 ;
      RECT 35.79 3.58 35.905 5.025 ;
      RECT 35.785 3.622 35.92 3.685 ;
      RECT 35.82 3.21 35.925 3.63 ;
      RECT 35.82 3.21 35.94 3.613 ;
      RECT 35.82 3.21 35.975 3.575 ;
      RECT 35.815 3.457 36.025 3.508 ;
      RECT 35.82 3.21 36.08 3.47 ;
      RECT 35.08 3.915 35.34 4.175 ;
      RECT 35.08 3.915 35.35 4.133 ;
      RECT 35.08 3.915 35.436 4.104 ;
      RECT 35.08 3.915 35.505 4.056 ;
      RECT 35.08 3.915 35.54 4.025 ;
      RECT 35.31 3.735 35.59 4.015 ;
      RECT 35.145 3.9 35.59 4.015 ;
      RECT 35.235 3.777 35.34 4.175 ;
      RECT 35.165 3.84 35.59 4.015 ;
      RECT 29.615 8.51 29.935 8.835 ;
      RECT 29.645 7.985 29.815 8.835 ;
      RECT 29.645 7.985 29.82 8.335 ;
      RECT 29.645 7.985 30.62 8.16 ;
      RECT 30.445 3.26 30.62 8.16 ;
      RECT 30.39 3.26 30.74 3.61 ;
      RECT 30.415 8.945 30.74 9.27 ;
      RECT 29.3 9.035 30.74 9.205 ;
      RECT 29.3 3.69 29.46 9.205 ;
      RECT 29.615 3.66 29.935 3.98 ;
      RECT 29.3 3.69 29.935 3.86 ;
      RECT 28.01 4 28.35 4.35 ;
      RECT 27.405 4.065 28.35 4.265 ;
      RECT 27.405 4.06 27.62 4.265 ;
      RECT 27.42 3.635 27.62 4.265 ;
      RECT 26.41 3.635 26.69 4.015 ;
      RECT 28.1 3.995 28.27 4.35 ;
      RECT 26.405 3.635 26.69 3.968 ;
      RECT 26.385 3.635 26.69 3.945 ;
      RECT 26.375 3.635 26.69 3.925 ;
      RECT 26.365 3.635 26.69 3.91 ;
      RECT 26.34 3.635 26.69 3.883 ;
      RECT 26.33 3.635 26.69 3.858 ;
      RECT 26.285 3.59 26.565 3.85 ;
      RECT 26.285 3.635 27.62 3.835 ;
      RECT 26.285 3.63 26.61 3.85 ;
      RECT 26.285 3.622 26.605 3.85 ;
      RECT 26.285 3.612 26.6 3.85 ;
      RECT 26.285 3.6 26.595 3.85 ;
      RECT 25.21 4.295 25.49 4.575 ;
      RECT 25.21 4.295 25.525 4.555 ;
      RECT 17.535 8.945 17.885 9.295 ;
      RECT 24.955 8.9 25.305 9.25 ;
      RECT 17.535 8.975 25.305 9.175 ;
      RECT 25.245 3.715 25.295 3.975 ;
      RECT 25.035 3.715 25.04 3.975 ;
      RECT 24.23 3.27 24.26 3.53 ;
      RECT 24 3.27 24.075 3.53 ;
      RECT 25.22 3.665 25.245 3.975 ;
      RECT 25.215 3.622 25.22 3.975 ;
      RECT 25.21 3.605 25.215 3.975 ;
      RECT 25.205 3.592 25.21 3.975 ;
      RECT 25.13 3.475 25.205 3.975 ;
      RECT 25.085 3.292 25.13 3.975 ;
      RECT 25.08 3.22 25.085 3.975 ;
      RECT 25.065 3.195 25.08 3.975 ;
      RECT 25.04 3.157 25.065 3.975 ;
      RECT 25.03 3.137 25.04 3.697 ;
      RECT 25.015 3.129 25.03 3.652 ;
      RECT 25.01 3.121 25.015 3.623 ;
      RECT 25.005 3.118 25.01 3.603 ;
      RECT 25 3.115 25.005 3.583 ;
      RECT 24.995 3.112 25 3.563 ;
      RECT 24.965 3.101 24.995 3.5 ;
      RECT 24.945 3.086 24.965 3.415 ;
      RECT 24.94 3.078 24.945 3.378 ;
      RECT 24.93 3.072 24.94 3.345 ;
      RECT 24.915 3.064 24.93 3.305 ;
      RECT 24.91 3.057 24.915 3.265 ;
      RECT 24.905 3.054 24.91 3.243 ;
      RECT 24.9 3.051 24.905 3.23 ;
      RECT 24.895 3.05 24.9 3.22 ;
      RECT 24.88 3.044 24.895 3.21 ;
      RECT 24.855 3.031 24.88 3.195 ;
      RECT 24.805 3.006 24.855 3.166 ;
      RECT 24.79 2.985 24.805 3.141 ;
      RECT 24.78 2.978 24.79 3.13 ;
      RECT 24.725 2.959 24.78 3.103 ;
      RECT 24.7 2.937 24.725 3.076 ;
      RECT 24.695 2.93 24.7 3.071 ;
      RECT 24.68 2.93 24.695 3.069 ;
      RECT 24.655 2.922 24.68 3.065 ;
      RECT 24.64 2.92 24.655 3.061 ;
      RECT 24.61 2.92 24.64 3.058 ;
      RECT 24.6 2.92 24.61 3.053 ;
      RECT 24.555 2.92 24.6 3.051 ;
      RECT 24.526 2.92 24.555 3.052 ;
      RECT 24.44 2.92 24.526 3.054 ;
      RECT 24.426 2.921 24.44 3.056 ;
      RECT 24.34 2.922 24.426 3.058 ;
      RECT 24.325 2.923 24.34 3.068 ;
      RECT 24.32 2.924 24.325 3.077 ;
      RECT 24.3 2.927 24.32 3.087 ;
      RECT 24.285 2.935 24.3 3.102 ;
      RECT 24.265 2.953 24.285 3.117 ;
      RECT 24.255 2.965 24.265 3.14 ;
      RECT 24.245 2.974 24.255 3.17 ;
      RECT 24.23 2.986 24.245 3.215 ;
      RECT 24.175 3.019 24.23 3.53 ;
      RECT 24.17 3.047 24.175 3.53 ;
      RECT 24.15 3.062 24.17 3.53 ;
      RECT 24.115 3.122 24.15 3.53 ;
      RECT 24.113 3.172 24.115 3.53 ;
      RECT 24.11 3.18 24.113 3.53 ;
      RECT 24.1 3.195 24.11 3.53 ;
      RECT 24.095 3.207 24.1 3.53 ;
      RECT 24.085 3.232 24.095 3.53 ;
      RECT 24.075 3.26 24.085 3.53 ;
      RECT 21.98 4.765 22.03 5.025 ;
      RECT 24.89 4.315 24.95 4.575 ;
      RECT 24.875 4.315 24.89 4.585 ;
      RECT 24.856 4.315 24.875 4.618 ;
      RECT 24.77 4.315 24.856 4.743 ;
      RECT 24.69 4.315 24.77 4.925 ;
      RECT 24.685 4.552 24.69 5.01 ;
      RECT 24.66 4.622 24.685 5.038 ;
      RECT 24.655 4.692 24.66 5.065 ;
      RECT 24.635 4.764 24.655 5.087 ;
      RECT 24.63 4.831 24.635 5.11 ;
      RECT 24.62 4.86 24.63 5.125 ;
      RECT 24.61 4.882 24.62 5.142 ;
      RECT 24.605 4.892 24.61 5.153 ;
      RECT 24.6 4.9 24.605 5.161 ;
      RECT 24.59 4.908 24.6 5.173 ;
      RECT 24.585 4.92 24.59 5.183 ;
      RECT 24.58 4.928 24.585 5.188 ;
      RECT 24.56 4.946 24.58 5.198 ;
      RECT 24.555 4.963 24.56 5.205 ;
      RECT 24.55 4.971 24.555 5.206 ;
      RECT 24.545 4.982 24.55 5.208 ;
      RECT 24.505 5.02 24.545 5.218 ;
      RECT 24.5 5.055 24.505 5.229 ;
      RECT 24.495 5.06 24.5 5.232 ;
      RECT 24.47 5.07 24.495 5.239 ;
      RECT 24.46 5.084 24.47 5.248 ;
      RECT 24.44 5.096 24.46 5.251 ;
      RECT 24.39 5.115 24.44 5.255 ;
      RECT 24.345 5.13 24.39 5.26 ;
      RECT 24.28 5.133 24.345 5.266 ;
      RECT 24.265 5.131 24.28 5.273 ;
      RECT 24.235 5.13 24.265 5.273 ;
      RECT 24.196 5.129 24.235 5.269 ;
      RECT 24.11 5.126 24.196 5.265 ;
      RECT 24.093 5.124 24.11 5.262 ;
      RECT 24.007 5.122 24.093 5.259 ;
      RECT 23.921 5.119 24.007 5.253 ;
      RECT 23.835 5.115 23.921 5.248 ;
      RECT 23.757 5.112 23.835 5.244 ;
      RECT 23.671 5.109 23.757 5.242 ;
      RECT 23.585 5.106 23.671 5.239 ;
      RECT 23.527 5.104 23.585 5.236 ;
      RECT 23.441 5.101 23.527 5.234 ;
      RECT 23.355 5.097 23.441 5.232 ;
      RECT 23.269 5.094 23.355 5.229 ;
      RECT 23.183 5.09 23.269 5.227 ;
      RECT 23.097 5.086 23.183 5.224 ;
      RECT 23.011 5.083 23.097 5.222 ;
      RECT 22.925 5.079 23.011 5.219 ;
      RECT 22.839 5.076 22.925 5.217 ;
      RECT 22.753 5.072 22.839 5.214 ;
      RECT 22.667 5.069 22.753 5.212 ;
      RECT 22.581 5.065 22.667 5.209 ;
      RECT 22.495 5.062 22.581 5.207 ;
      RECT 22.485 5.06 22.495 5.203 ;
      RECT 22.48 5.06 22.485 5.201 ;
      RECT 22.44 5.055 22.48 5.195 ;
      RECT 22.426 5.046 22.44 5.188 ;
      RECT 22.34 5.016 22.426 5.173 ;
      RECT 22.32 4.982 22.34 5.158 ;
      RECT 22.25 4.951 22.32 5.145 ;
      RECT 22.245 4.926 22.25 5.134 ;
      RECT 22.24 4.92 22.245 5.132 ;
      RECT 22.171 4.765 22.24 5.12 ;
      RECT 22.085 4.765 22.171 5.094 ;
      RECT 22.06 4.765 22.085 5.073 ;
      RECT 22.055 4.765 22.06 5.063 ;
      RECT 22.05 4.765 22.055 5.055 ;
      RECT 22.03 4.765 22.05 5.038 ;
      RECT 24.45 3.335 24.71 3.595 ;
      RECT 24.435 3.335 24.71 3.498 ;
      RECT 24.405 3.335 24.71 3.473 ;
      RECT 24.37 3.175 24.65 3.455 ;
      RECT 24.34 4.665 24.4 4.925 ;
      RECT 23.365 3.355 23.42 3.615 ;
      RECT 24.3 4.622 24.34 4.925 ;
      RECT 24.271 4.543 24.3 4.925 ;
      RECT 24.185 4.415 24.271 4.925 ;
      RECT 24.165 4.295 24.185 4.925 ;
      RECT 24.14 4.246 24.165 4.925 ;
      RECT 24.135 4.211 24.14 4.775 ;
      RECT 24.105 4.171 24.135 4.713 ;
      RECT 24.08 4.108 24.105 4.628 ;
      RECT 24.07 4.07 24.08 4.565 ;
      RECT 24.055 4.045 24.07 4.526 ;
      RECT 24.012 4.003 24.055 4.432 ;
      RECT 24.01 3.976 24.012 4.359 ;
      RECT 24.005 3.971 24.01 4.35 ;
      RECT 24 3.964 24.005 4.325 ;
      RECT 23.995 3.958 24 4.31 ;
      RECT 23.99 3.952 23.995 4.298 ;
      RECT 23.98 3.943 23.99 4.28 ;
      RECT 23.975 3.934 23.98 4.258 ;
      RECT 23.95 3.915 23.975 4.208 ;
      RECT 23.945 3.896 23.95 4.158 ;
      RECT 23.93 3.882 23.945 4.118 ;
      RECT 23.925 3.868 23.93 4.085 ;
      RECT 23.92 3.861 23.925 4.078 ;
      RECT 23.905 3.848 23.92 4.07 ;
      RECT 23.86 3.81 23.905 4.043 ;
      RECT 23.83 3.763 23.86 4.008 ;
      RECT 23.81 3.732 23.83 3.985 ;
      RECT 23.73 3.665 23.81 3.938 ;
      RECT 23.7 3.595 23.73 3.885 ;
      RECT 23.695 3.572 23.7 3.868 ;
      RECT 23.665 3.55 23.695 3.853 ;
      RECT 23.635 3.509 23.665 3.825 ;
      RECT 23.63 3.484 23.635 3.81 ;
      RECT 23.625 3.478 23.63 3.803 ;
      RECT 23.615 3.355 23.625 3.795 ;
      RECT 23.605 3.355 23.615 3.788 ;
      RECT 23.6 3.355 23.605 3.78 ;
      RECT 23.58 3.355 23.6 3.768 ;
      RECT 23.53 3.355 23.58 3.738 ;
      RECT 23.475 3.355 23.53 3.688 ;
      RECT 23.445 3.355 23.475 3.648 ;
      RECT 23.42 3.355 23.445 3.625 ;
      RECT 23.29 4.08 23.57 4.36 ;
      RECT 23.255 3.995 23.515 4.255 ;
      RECT 23.255 4.077 23.525 4.255 ;
      RECT 21.455 3.45 21.46 3.935 ;
      RECT 21.345 3.635 21.35 3.935 ;
      RECT 21.255 3.675 21.32 3.935 ;
      RECT 22.93 3.175 23.02 3.805 ;
      RECT 22.895 3.225 22.9 3.805 ;
      RECT 22.84 3.25 22.85 3.805 ;
      RECT 22.795 3.25 22.805 3.805 ;
      RECT 23.165 3.175 23.21 3.455 ;
      RECT 22.015 2.905 22.215 3.045 ;
      RECT 23.131 3.175 23.165 3.467 ;
      RECT 23.045 3.175 23.131 3.507 ;
      RECT 23.03 3.175 23.045 3.548 ;
      RECT 23.025 3.175 23.03 3.568 ;
      RECT 23.02 3.175 23.025 3.588 ;
      RECT 22.9 3.217 22.93 3.805 ;
      RECT 22.85 3.237 22.895 3.805 ;
      RECT 22.835 3.252 22.84 3.805 ;
      RECT 22.805 3.252 22.835 3.805 ;
      RECT 22.76 3.237 22.795 3.805 ;
      RECT 22.755 3.225 22.76 3.585 ;
      RECT 22.75 3.222 22.755 3.565 ;
      RECT 22.735 3.212 22.75 3.518 ;
      RECT 22.73 3.205 22.735 3.481 ;
      RECT 22.725 3.202 22.73 3.464 ;
      RECT 22.71 3.192 22.725 3.42 ;
      RECT 22.705 3.183 22.71 3.38 ;
      RECT 22.7 3.179 22.705 3.365 ;
      RECT 22.69 3.173 22.7 3.348 ;
      RECT 22.65 3.154 22.69 3.323 ;
      RECT 22.645 3.136 22.65 3.303 ;
      RECT 22.635 3.13 22.645 3.298 ;
      RECT 22.605 3.114 22.635 3.285 ;
      RECT 22.59 3.096 22.605 3.268 ;
      RECT 22.575 3.084 22.59 3.255 ;
      RECT 22.57 3.076 22.575 3.248 ;
      RECT 22.54 3.062 22.57 3.235 ;
      RECT 22.535 3.047 22.54 3.223 ;
      RECT 22.525 3.041 22.535 3.215 ;
      RECT 22.505 3.029 22.525 3.203 ;
      RECT 22.495 3.017 22.505 3.19 ;
      RECT 22.465 3.001 22.495 3.175 ;
      RECT 22.445 2.981 22.465 3.158 ;
      RECT 22.44 2.971 22.445 3.148 ;
      RECT 22.415 2.959 22.44 3.135 ;
      RECT 22.41 2.947 22.415 3.123 ;
      RECT 22.405 2.942 22.41 3.119 ;
      RECT 22.39 2.935 22.405 3.111 ;
      RECT 22.38 2.922 22.39 3.101 ;
      RECT 22.375 2.92 22.38 3.095 ;
      RECT 22.35 2.913 22.375 3.084 ;
      RECT 22.345 2.906 22.35 3.073 ;
      RECT 22.32 2.905 22.345 3.06 ;
      RECT 22.301 2.905 22.32 3.05 ;
      RECT 22.215 2.905 22.301 3.047 ;
      RECT 21.985 2.905 22.015 3.05 ;
      RECT 21.945 2.912 21.985 3.063 ;
      RECT 21.92 2.922 21.945 3.076 ;
      RECT 21.905 2.931 21.92 3.086 ;
      RECT 21.875 2.936 21.905 3.105 ;
      RECT 21.87 2.942 21.875 3.123 ;
      RECT 21.85 2.952 21.87 3.138 ;
      RECT 21.84 2.965 21.85 3.158 ;
      RECT 21.825 2.977 21.84 3.175 ;
      RECT 21.82 2.987 21.825 3.185 ;
      RECT 21.815 2.992 21.82 3.19 ;
      RECT 21.805 3 21.815 3.203 ;
      RECT 21.755 3.032 21.805 3.24 ;
      RECT 21.74 3.067 21.755 3.281 ;
      RECT 21.735 3.077 21.74 3.296 ;
      RECT 21.73 3.082 21.735 3.303 ;
      RECT 21.705 3.098 21.73 3.323 ;
      RECT 21.69 3.119 21.705 3.348 ;
      RECT 21.665 3.14 21.69 3.373 ;
      RECT 21.655 3.159 21.665 3.396 ;
      RECT 21.63 3.177 21.655 3.419 ;
      RECT 21.615 3.197 21.63 3.443 ;
      RECT 21.61 3.207 21.615 3.455 ;
      RECT 21.595 3.219 21.61 3.475 ;
      RECT 21.585 3.234 21.595 3.515 ;
      RECT 21.58 3.242 21.585 3.543 ;
      RECT 21.57 3.252 21.58 3.563 ;
      RECT 21.565 3.265 21.57 3.588 ;
      RECT 21.56 3.278 21.565 3.608 ;
      RECT 21.555 3.284 21.56 3.63 ;
      RECT 21.545 3.293 21.555 3.65 ;
      RECT 21.54 3.313 21.545 3.673 ;
      RECT 21.535 3.319 21.54 3.693 ;
      RECT 21.53 3.326 21.535 3.715 ;
      RECT 21.525 3.337 21.53 3.728 ;
      RECT 21.515 3.347 21.525 3.753 ;
      RECT 21.495 3.372 21.515 3.935 ;
      RECT 21.465 3.412 21.495 3.935 ;
      RECT 21.46 3.442 21.465 3.935 ;
      RECT 21.435 3.47 21.455 3.935 ;
      RECT 21.405 3.515 21.435 3.935 ;
      RECT 21.4 3.542 21.405 3.935 ;
      RECT 21.38 3.56 21.4 3.935 ;
      RECT 21.37 3.585 21.38 3.935 ;
      RECT 21.365 3.597 21.37 3.935 ;
      RECT 21.35 3.62 21.365 3.935 ;
      RECT 21.33 3.647 21.345 3.935 ;
      RECT 21.32 3.67 21.33 3.935 ;
      RECT 23.11 4.555 23.19 4.815 ;
      RECT 22.345 3.775 22.415 4.035 ;
      RECT 23.076 4.522 23.11 4.815 ;
      RECT 22.99 4.425 23.076 4.815 ;
      RECT 22.97 4.337 22.99 4.815 ;
      RECT 22.96 4.307 22.97 4.815 ;
      RECT 22.95 4.287 22.96 4.815 ;
      RECT 22.93 4.274 22.95 4.815 ;
      RECT 22.915 4.264 22.93 4.643 ;
      RECT 22.91 4.257 22.915 4.598 ;
      RECT 22.9 4.251 22.91 4.588 ;
      RECT 22.89 4.243 22.9 4.57 ;
      RECT 22.885 4.237 22.89 4.558 ;
      RECT 22.875 4.232 22.885 4.545 ;
      RECT 22.855 4.222 22.875 4.518 ;
      RECT 22.815 4.201 22.855 4.47 ;
      RECT 22.8 4.182 22.815 4.428 ;
      RECT 22.775 4.168 22.8 4.398 ;
      RECT 22.765 4.156 22.775 4.365 ;
      RECT 22.76 4.151 22.765 4.355 ;
      RECT 22.73 4.137 22.76 4.335 ;
      RECT 22.72 4.121 22.73 4.308 ;
      RECT 22.715 4.116 22.72 4.298 ;
      RECT 22.69 4.107 22.715 4.278 ;
      RECT 22.68 4.095 22.69 4.258 ;
      RECT 22.61 4.063 22.68 4.233 ;
      RECT 22.605 4.032 22.61 4.21 ;
      RECT 22.556 3.775 22.605 4.193 ;
      RECT 22.47 3.775 22.556 4.152 ;
      RECT 22.415 3.775 22.47 4.08 ;
      RECT 22.505 4.56 22.665 4.82 ;
      RECT 22.03 3.175 22.08 3.86 ;
      RECT 21.82 3.6 21.855 3.86 ;
      RECT 22.135 3.175 22.14 3.635 ;
      RECT 22.225 3.175 22.25 3.455 ;
      RECT 22.5 4.557 22.505 4.82 ;
      RECT 22.465 4.545 22.5 4.82 ;
      RECT 22.405 4.518 22.465 4.82 ;
      RECT 22.4 4.501 22.405 4.674 ;
      RECT 22.395 4.498 22.4 4.661 ;
      RECT 22.375 4.491 22.395 4.648 ;
      RECT 22.34 4.474 22.375 4.63 ;
      RECT 22.3 4.453 22.34 4.61 ;
      RECT 22.295 4.441 22.3 4.598 ;
      RECT 22.255 4.427 22.295 4.584 ;
      RECT 22.235 4.41 22.255 4.566 ;
      RECT 22.225 4.402 22.235 4.558 ;
      RECT 22.21 3.175 22.225 3.473 ;
      RECT 22.195 4.392 22.225 4.545 ;
      RECT 22.18 3.175 22.21 3.518 ;
      RECT 22.185 4.382 22.195 4.532 ;
      RECT 22.155 4.367 22.185 4.519 ;
      RECT 22.14 3.175 22.18 3.585 ;
      RECT 22.14 4.335 22.155 4.505 ;
      RECT 22.135 4.307 22.14 4.499 ;
      RECT 22.13 3.175 22.135 3.64 ;
      RECT 22.12 4.277 22.135 4.493 ;
      RECT 22.125 3.175 22.13 3.653 ;
      RECT 22.115 3.175 22.125 3.673 ;
      RECT 22.08 4.19 22.12 4.478 ;
      RECT 22.08 3.175 22.115 3.713 ;
      RECT 22.075 4.122 22.08 4.466 ;
      RECT 22.06 4.077 22.075 4.461 ;
      RECT 22.055 4.015 22.06 4.456 ;
      RECT 22.03 3.922 22.055 4.449 ;
      RECT 22.025 3.175 22.03 4.441 ;
      RECT 22.01 3.175 22.025 4.428 ;
      RECT 21.99 3.175 22.01 4.385 ;
      RECT 21.98 3.175 21.99 4.335 ;
      RECT 21.975 3.175 21.98 4.308 ;
      RECT 21.97 3.175 21.975 4.286 ;
      RECT 21.965 3.401 21.97 4.269 ;
      RECT 21.96 3.423 21.965 4.247 ;
      RECT 21.955 3.465 21.96 4.23 ;
      RECT 21.925 3.515 21.955 4.174 ;
      RECT 21.92 3.542 21.925 4.116 ;
      RECT 21.905 3.56 21.92 4.08 ;
      RECT 21.9 3.578 21.905 4.044 ;
      RECT 21.894 3.585 21.9 4.025 ;
      RECT 21.89 3.592 21.894 4.008 ;
      RECT 21.885 3.597 21.89 3.977 ;
      RECT 21.875 3.6 21.885 3.952 ;
      RECT 21.865 3.6 21.875 3.918 ;
      RECT 21.86 3.6 21.865 3.895 ;
      RECT 21.855 3.6 21.86 3.875 ;
      RECT 20.77 3.735 21.05 4.015 ;
      RECT 20.77 3.735 21.07 3.91 ;
      RECT 20.86 3.625 21.12 3.885 ;
      RECT 20.825 3.72 21.12 3.885 ;
      RECT 20.95 2.24 21.115 3.885 ;
      RECT 20.85 2.24 21.22 2.61 ;
      RECT 20.475 4.765 20.735 5.025 ;
      RECT 20.495 4.692 20.675 5.025 ;
      RECT 20.495 4.435 20.67 5.025 ;
      RECT 20.495 4.227 20.66 5.025 ;
      RECT 20.5 4.145 20.66 5.025 ;
      RECT 20.5 3.91 20.65 5.025 ;
      RECT 20.5 3.757 20.645 5.025 ;
      RECT 20.505 3.742 20.645 5.025 ;
      RECT 20.555 3.457 20.645 5.025 ;
      RECT 20.51 3.692 20.645 5.025 ;
      RECT 20.54 3.51 20.645 5.025 ;
      RECT 20.525 3.622 20.645 5.025 ;
      RECT 20.53 3.58 20.645 5.025 ;
      RECT 20.525 3.622 20.66 3.685 ;
      RECT 20.56 3.21 20.665 3.63 ;
      RECT 20.56 3.21 20.68 3.613 ;
      RECT 20.56 3.21 20.715 3.575 ;
      RECT 20.555 3.457 20.765 3.508 ;
      RECT 20.56 3.21 20.82 3.47 ;
      RECT 19.82 3.915 20.08 4.175 ;
      RECT 19.82 3.915 20.09 4.133 ;
      RECT 19.82 3.915 20.176 4.104 ;
      RECT 19.82 3.915 20.245 4.056 ;
      RECT 19.82 3.915 20.28 4.025 ;
      RECT 20.05 3.735 20.33 4.015 ;
      RECT 19.885 3.9 20.33 4.015 ;
      RECT 19.975 3.777 20.08 4.175 ;
      RECT 19.905 3.84 20.33 4.015 ;
      RECT 14.355 8.51 14.675 8.835 ;
      RECT 14.385 7.985 14.555 8.835 ;
      RECT 14.385 7.985 14.56 8.335 ;
      RECT 14.385 7.985 15.36 8.16 ;
      RECT 15.185 3.26 15.36 8.16 ;
      RECT 15.13 3.26 15.48 3.61 ;
      RECT 15.155 8.945 15.48 9.27 ;
      RECT 14.04 9.035 15.48 9.205 ;
      RECT 14.04 3.69 14.2 9.205 ;
      RECT 14.355 3.66 14.675 3.98 ;
      RECT 14.04 3.69 14.675 3.86 ;
      RECT 12.75 4 13.09 4.35 ;
      RECT 12.145 4.065 13.09 4.265 ;
      RECT 12.145 4.06 12.36 4.265 ;
      RECT 12.16 3.635 12.36 4.265 ;
      RECT 11.15 3.635 11.43 4.015 ;
      RECT 12.84 3.995 13.01 4.35 ;
      RECT 11.145 3.635 11.43 3.968 ;
      RECT 11.125 3.635 11.43 3.945 ;
      RECT 11.115 3.635 11.43 3.925 ;
      RECT 11.105 3.635 11.43 3.91 ;
      RECT 11.08 3.635 11.43 3.883 ;
      RECT 11.07 3.635 11.43 3.858 ;
      RECT 11.025 3.59 11.305 3.85 ;
      RECT 11.025 3.635 12.36 3.835 ;
      RECT 11.025 3.63 11.35 3.85 ;
      RECT 11.025 3.622 11.345 3.85 ;
      RECT 11.025 3.612 11.34 3.85 ;
      RECT 11.025 3.6 11.335 3.85 ;
      RECT 9.95 4.295 10.23 4.575 ;
      RECT 9.95 4.295 10.265 4.555 ;
      RECT 1.57 9.285 1.86 9.635 ;
      RECT 1.57 9.345 2.9 9.515 ;
      RECT 2.73 8.975 2.9 9.515 ;
      RECT 9.695 8.895 10.045 9.245 ;
      RECT 2.73 8.975 10.045 9.145 ;
      RECT 9.985 3.715 10.035 3.975 ;
      RECT 9.775 3.715 9.78 3.975 ;
      RECT 8.97 3.27 9 3.53 ;
      RECT 8.74 3.27 8.815 3.53 ;
      RECT 9.96 3.665 9.985 3.975 ;
      RECT 9.955 3.622 9.96 3.975 ;
      RECT 9.95 3.605 9.955 3.975 ;
      RECT 9.945 3.592 9.95 3.975 ;
      RECT 9.87 3.475 9.945 3.975 ;
      RECT 9.825 3.292 9.87 3.975 ;
      RECT 9.82 3.22 9.825 3.975 ;
      RECT 9.805 3.195 9.82 3.975 ;
      RECT 9.78 3.157 9.805 3.975 ;
      RECT 9.77 3.137 9.78 3.697 ;
      RECT 9.755 3.129 9.77 3.652 ;
      RECT 9.75 3.121 9.755 3.623 ;
      RECT 9.745 3.118 9.75 3.603 ;
      RECT 9.74 3.115 9.745 3.583 ;
      RECT 9.735 3.112 9.74 3.563 ;
      RECT 9.705 3.101 9.735 3.5 ;
      RECT 9.685 3.086 9.705 3.415 ;
      RECT 9.68 3.078 9.685 3.378 ;
      RECT 9.67 3.072 9.68 3.345 ;
      RECT 9.655 3.064 9.67 3.305 ;
      RECT 9.65 3.057 9.655 3.265 ;
      RECT 9.645 3.054 9.65 3.243 ;
      RECT 9.64 3.051 9.645 3.23 ;
      RECT 9.635 3.05 9.64 3.22 ;
      RECT 9.62 3.044 9.635 3.21 ;
      RECT 9.595 3.031 9.62 3.195 ;
      RECT 9.545 3.006 9.595 3.166 ;
      RECT 9.53 2.985 9.545 3.141 ;
      RECT 9.52 2.978 9.53 3.13 ;
      RECT 9.465 2.959 9.52 3.103 ;
      RECT 9.44 2.937 9.465 3.076 ;
      RECT 9.435 2.93 9.44 3.071 ;
      RECT 9.42 2.93 9.435 3.069 ;
      RECT 9.395 2.922 9.42 3.065 ;
      RECT 9.38 2.92 9.395 3.061 ;
      RECT 9.35 2.92 9.38 3.058 ;
      RECT 9.34 2.92 9.35 3.053 ;
      RECT 9.295 2.92 9.34 3.051 ;
      RECT 9.266 2.92 9.295 3.052 ;
      RECT 9.18 2.92 9.266 3.054 ;
      RECT 9.166 2.921 9.18 3.056 ;
      RECT 9.08 2.922 9.166 3.058 ;
      RECT 9.065 2.923 9.08 3.068 ;
      RECT 9.06 2.924 9.065 3.077 ;
      RECT 9.04 2.927 9.06 3.087 ;
      RECT 9.025 2.935 9.04 3.102 ;
      RECT 9.005 2.953 9.025 3.117 ;
      RECT 8.995 2.965 9.005 3.14 ;
      RECT 8.985 2.974 8.995 3.17 ;
      RECT 8.97 2.986 8.985 3.215 ;
      RECT 8.915 3.019 8.97 3.53 ;
      RECT 8.91 3.047 8.915 3.53 ;
      RECT 8.89 3.062 8.91 3.53 ;
      RECT 8.855 3.122 8.89 3.53 ;
      RECT 8.853 3.172 8.855 3.53 ;
      RECT 8.85 3.18 8.853 3.53 ;
      RECT 8.84 3.195 8.85 3.53 ;
      RECT 8.835 3.207 8.84 3.53 ;
      RECT 8.825 3.232 8.835 3.53 ;
      RECT 8.815 3.26 8.825 3.53 ;
      RECT 6.72 4.765 6.77 5.025 ;
      RECT 9.63 4.315 9.69 4.575 ;
      RECT 9.615 4.315 9.63 4.585 ;
      RECT 9.596 4.315 9.615 4.618 ;
      RECT 9.51 4.315 9.596 4.743 ;
      RECT 9.43 4.315 9.51 4.925 ;
      RECT 9.425 4.552 9.43 5.01 ;
      RECT 9.4 4.622 9.425 5.038 ;
      RECT 9.395 4.692 9.4 5.065 ;
      RECT 9.375 4.764 9.395 5.087 ;
      RECT 9.37 4.831 9.375 5.11 ;
      RECT 9.36 4.86 9.37 5.125 ;
      RECT 9.35 4.882 9.36 5.142 ;
      RECT 9.345 4.892 9.35 5.153 ;
      RECT 9.34 4.9 9.345 5.161 ;
      RECT 9.33 4.908 9.34 5.173 ;
      RECT 9.325 4.92 9.33 5.183 ;
      RECT 9.32 4.928 9.325 5.188 ;
      RECT 9.3 4.946 9.32 5.198 ;
      RECT 9.295 4.963 9.3 5.205 ;
      RECT 9.29 4.971 9.295 5.206 ;
      RECT 9.285 4.982 9.29 5.208 ;
      RECT 9.245 5.02 9.285 5.218 ;
      RECT 9.24 5.055 9.245 5.229 ;
      RECT 9.235 5.06 9.24 5.232 ;
      RECT 9.21 5.07 9.235 5.239 ;
      RECT 9.2 5.084 9.21 5.248 ;
      RECT 9.18 5.096 9.2 5.251 ;
      RECT 9.13 5.115 9.18 5.255 ;
      RECT 9.085 5.13 9.13 5.26 ;
      RECT 9.02 5.133 9.085 5.266 ;
      RECT 9.005 5.131 9.02 5.273 ;
      RECT 8.975 5.13 9.005 5.273 ;
      RECT 8.936 5.129 8.975 5.269 ;
      RECT 8.85 5.126 8.936 5.265 ;
      RECT 8.833 5.124 8.85 5.262 ;
      RECT 8.747 5.122 8.833 5.259 ;
      RECT 8.661 5.119 8.747 5.253 ;
      RECT 8.575 5.115 8.661 5.248 ;
      RECT 8.497 5.112 8.575 5.244 ;
      RECT 8.411 5.109 8.497 5.242 ;
      RECT 8.325 5.106 8.411 5.239 ;
      RECT 8.267 5.104 8.325 5.236 ;
      RECT 8.181 5.101 8.267 5.234 ;
      RECT 8.095 5.097 8.181 5.232 ;
      RECT 8.009 5.094 8.095 5.229 ;
      RECT 7.923 5.09 8.009 5.227 ;
      RECT 7.837 5.086 7.923 5.224 ;
      RECT 7.751 5.083 7.837 5.222 ;
      RECT 7.665 5.079 7.751 5.219 ;
      RECT 7.579 5.076 7.665 5.217 ;
      RECT 7.493 5.072 7.579 5.214 ;
      RECT 7.407 5.069 7.493 5.212 ;
      RECT 7.321 5.065 7.407 5.209 ;
      RECT 7.235 5.062 7.321 5.207 ;
      RECT 7.225 5.06 7.235 5.203 ;
      RECT 7.22 5.06 7.225 5.201 ;
      RECT 7.18 5.055 7.22 5.195 ;
      RECT 7.166 5.046 7.18 5.188 ;
      RECT 7.08 5.016 7.166 5.173 ;
      RECT 7.06 4.982 7.08 5.158 ;
      RECT 6.99 4.951 7.06 5.145 ;
      RECT 6.985 4.926 6.99 5.134 ;
      RECT 6.98 4.92 6.985 5.132 ;
      RECT 6.911 4.765 6.98 5.12 ;
      RECT 6.825 4.765 6.911 5.094 ;
      RECT 6.8 4.765 6.825 5.073 ;
      RECT 6.795 4.765 6.8 5.063 ;
      RECT 6.79 4.765 6.795 5.055 ;
      RECT 6.77 4.765 6.79 5.038 ;
      RECT 9.19 3.335 9.45 3.595 ;
      RECT 9.175 3.335 9.45 3.498 ;
      RECT 9.145 3.335 9.45 3.473 ;
      RECT 9.11 3.175 9.39 3.455 ;
      RECT 9.08 4.665 9.14 4.925 ;
      RECT 8.105 3.355 8.16 3.615 ;
      RECT 9.04 4.622 9.08 4.925 ;
      RECT 9.011 4.543 9.04 4.925 ;
      RECT 8.925 4.415 9.011 4.925 ;
      RECT 8.905 4.295 8.925 4.925 ;
      RECT 8.88 4.246 8.905 4.925 ;
      RECT 8.875 4.211 8.88 4.775 ;
      RECT 8.845 4.171 8.875 4.713 ;
      RECT 8.82 4.108 8.845 4.628 ;
      RECT 8.81 4.07 8.82 4.565 ;
      RECT 8.795 4.045 8.81 4.526 ;
      RECT 8.752 4.003 8.795 4.432 ;
      RECT 8.75 3.976 8.752 4.359 ;
      RECT 8.745 3.971 8.75 4.35 ;
      RECT 8.74 3.964 8.745 4.325 ;
      RECT 8.735 3.958 8.74 4.31 ;
      RECT 8.73 3.952 8.735 4.298 ;
      RECT 8.72 3.943 8.73 4.28 ;
      RECT 8.715 3.934 8.72 4.258 ;
      RECT 8.69 3.915 8.715 4.208 ;
      RECT 8.685 3.896 8.69 4.158 ;
      RECT 8.67 3.882 8.685 4.118 ;
      RECT 8.665 3.868 8.67 4.085 ;
      RECT 8.66 3.861 8.665 4.078 ;
      RECT 8.645 3.848 8.66 4.07 ;
      RECT 8.6 3.81 8.645 4.043 ;
      RECT 8.57 3.763 8.6 4.008 ;
      RECT 8.55 3.732 8.57 3.985 ;
      RECT 8.47 3.665 8.55 3.938 ;
      RECT 8.44 3.595 8.47 3.885 ;
      RECT 8.435 3.572 8.44 3.868 ;
      RECT 8.405 3.55 8.435 3.853 ;
      RECT 8.375 3.509 8.405 3.825 ;
      RECT 8.37 3.484 8.375 3.81 ;
      RECT 8.365 3.478 8.37 3.803 ;
      RECT 8.355 3.355 8.365 3.795 ;
      RECT 8.345 3.355 8.355 3.788 ;
      RECT 8.34 3.355 8.345 3.78 ;
      RECT 8.32 3.355 8.34 3.768 ;
      RECT 8.27 3.355 8.32 3.738 ;
      RECT 8.215 3.355 8.27 3.688 ;
      RECT 8.185 3.355 8.215 3.648 ;
      RECT 8.16 3.355 8.185 3.625 ;
      RECT 8.03 4.08 8.31 4.36 ;
      RECT 7.995 3.995 8.255 4.255 ;
      RECT 7.995 4.077 8.265 4.255 ;
      RECT 6.195 3.45 6.2 3.935 ;
      RECT 6.085 3.635 6.09 3.935 ;
      RECT 5.995 3.675 6.06 3.935 ;
      RECT 7.67 3.175 7.76 3.805 ;
      RECT 7.635 3.225 7.64 3.805 ;
      RECT 7.58 3.25 7.59 3.805 ;
      RECT 7.535 3.25 7.545 3.805 ;
      RECT 7.905 3.175 7.95 3.455 ;
      RECT 6.755 2.905 6.955 3.045 ;
      RECT 7.871 3.175 7.905 3.467 ;
      RECT 7.785 3.175 7.871 3.507 ;
      RECT 7.77 3.175 7.785 3.548 ;
      RECT 7.765 3.175 7.77 3.568 ;
      RECT 7.76 3.175 7.765 3.588 ;
      RECT 7.64 3.217 7.67 3.805 ;
      RECT 7.59 3.237 7.635 3.805 ;
      RECT 7.575 3.252 7.58 3.805 ;
      RECT 7.545 3.252 7.575 3.805 ;
      RECT 7.5 3.237 7.535 3.805 ;
      RECT 7.495 3.225 7.5 3.585 ;
      RECT 7.49 3.222 7.495 3.565 ;
      RECT 7.475 3.212 7.49 3.518 ;
      RECT 7.47 3.205 7.475 3.481 ;
      RECT 7.465 3.202 7.47 3.464 ;
      RECT 7.45 3.192 7.465 3.42 ;
      RECT 7.445 3.183 7.45 3.38 ;
      RECT 7.44 3.179 7.445 3.365 ;
      RECT 7.43 3.173 7.44 3.348 ;
      RECT 7.39 3.154 7.43 3.323 ;
      RECT 7.385 3.136 7.39 3.303 ;
      RECT 7.375 3.13 7.385 3.298 ;
      RECT 7.345 3.114 7.375 3.285 ;
      RECT 7.33 3.096 7.345 3.268 ;
      RECT 7.315 3.084 7.33 3.255 ;
      RECT 7.31 3.076 7.315 3.248 ;
      RECT 7.28 3.062 7.31 3.235 ;
      RECT 7.275 3.047 7.28 3.223 ;
      RECT 7.265 3.041 7.275 3.215 ;
      RECT 7.245 3.029 7.265 3.203 ;
      RECT 7.235 3.017 7.245 3.19 ;
      RECT 7.205 3.001 7.235 3.175 ;
      RECT 7.185 2.981 7.205 3.158 ;
      RECT 7.18 2.971 7.185 3.148 ;
      RECT 7.155 2.959 7.18 3.135 ;
      RECT 7.15 2.947 7.155 3.123 ;
      RECT 7.145 2.942 7.15 3.119 ;
      RECT 7.13 2.935 7.145 3.111 ;
      RECT 7.12 2.922 7.13 3.101 ;
      RECT 7.115 2.92 7.12 3.095 ;
      RECT 7.09 2.913 7.115 3.084 ;
      RECT 7.085 2.906 7.09 3.073 ;
      RECT 7.06 2.905 7.085 3.06 ;
      RECT 7.041 2.905 7.06 3.05 ;
      RECT 6.955 2.905 7.041 3.047 ;
      RECT 6.725 2.905 6.755 3.05 ;
      RECT 6.685 2.912 6.725 3.063 ;
      RECT 6.66 2.922 6.685 3.076 ;
      RECT 6.645 2.931 6.66 3.086 ;
      RECT 6.615 2.936 6.645 3.105 ;
      RECT 6.61 2.942 6.615 3.123 ;
      RECT 6.59 2.952 6.61 3.138 ;
      RECT 6.58 2.965 6.59 3.158 ;
      RECT 6.565 2.977 6.58 3.175 ;
      RECT 6.56 2.987 6.565 3.185 ;
      RECT 6.555 2.992 6.56 3.19 ;
      RECT 6.545 3 6.555 3.203 ;
      RECT 6.495 3.032 6.545 3.24 ;
      RECT 6.48 3.067 6.495 3.281 ;
      RECT 6.475 3.077 6.48 3.296 ;
      RECT 6.47 3.082 6.475 3.303 ;
      RECT 6.445 3.098 6.47 3.323 ;
      RECT 6.43 3.119 6.445 3.348 ;
      RECT 6.405 3.14 6.43 3.373 ;
      RECT 6.395 3.159 6.405 3.396 ;
      RECT 6.37 3.177 6.395 3.419 ;
      RECT 6.355 3.197 6.37 3.443 ;
      RECT 6.35 3.207 6.355 3.455 ;
      RECT 6.335 3.219 6.35 3.475 ;
      RECT 6.325 3.234 6.335 3.515 ;
      RECT 6.32 3.242 6.325 3.543 ;
      RECT 6.31 3.252 6.32 3.563 ;
      RECT 6.305 3.265 6.31 3.588 ;
      RECT 6.3 3.278 6.305 3.608 ;
      RECT 6.295 3.284 6.3 3.63 ;
      RECT 6.285 3.293 6.295 3.65 ;
      RECT 6.28 3.313 6.285 3.673 ;
      RECT 6.275 3.319 6.28 3.693 ;
      RECT 6.27 3.326 6.275 3.715 ;
      RECT 6.265 3.337 6.27 3.728 ;
      RECT 6.255 3.347 6.265 3.753 ;
      RECT 6.235 3.372 6.255 3.935 ;
      RECT 6.205 3.412 6.235 3.935 ;
      RECT 6.2 3.442 6.205 3.935 ;
      RECT 6.175 3.47 6.195 3.935 ;
      RECT 6.145 3.515 6.175 3.935 ;
      RECT 6.14 3.542 6.145 3.935 ;
      RECT 6.12 3.56 6.14 3.935 ;
      RECT 6.11 3.585 6.12 3.935 ;
      RECT 6.105 3.597 6.11 3.935 ;
      RECT 6.09 3.62 6.105 3.935 ;
      RECT 6.07 3.647 6.085 3.935 ;
      RECT 6.06 3.67 6.07 3.935 ;
      RECT 7.85 4.555 7.93 4.815 ;
      RECT 7.085 3.775 7.155 4.035 ;
      RECT 7.816 4.522 7.85 4.815 ;
      RECT 7.73 4.425 7.816 4.815 ;
      RECT 7.71 4.337 7.73 4.815 ;
      RECT 7.7 4.307 7.71 4.815 ;
      RECT 7.69 4.287 7.7 4.815 ;
      RECT 7.67 4.274 7.69 4.815 ;
      RECT 7.655 4.264 7.67 4.643 ;
      RECT 7.65 4.257 7.655 4.598 ;
      RECT 7.64 4.251 7.65 4.588 ;
      RECT 7.63 4.243 7.64 4.57 ;
      RECT 7.625 4.237 7.63 4.558 ;
      RECT 7.615 4.232 7.625 4.545 ;
      RECT 7.595 4.222 7.615 4.518 ;
      RECT 7.555 4.201 7.595 4.47 ;
      RECT 7.54 4.182 7.555 4.428 ;
      RECT 7.515 4.168 7.54 4.398 ;
      RECT 7.505 4.156 7.515 4.365 ;
      RECT 7.5 4.151 7.505 4.355 ;
      RECT 7.47 4.137 7.5 4.335 ;
      RECT 7.46 4.121 7.47 4.308 ;
      RECT 7.455 4.116 7.46 4.298 ;
      RECT 7.43 4.107 7.455 4.278 ;
      RECT 7.42 4.095 7.43 4.258 ;
      RECT 7.35 4.063 7.42 4.233 ;
      RECT 7.345 4.032 7.35 4.21 ;
      RECT 7.296 3.775 7.345 4.193 ;
      RECT 7.21 3.775 7.296 4.152 ;
      RECT 7.155 3.775 7.21 4.08 ;
      RECT 7.245 4.56 7.405 4.82 ;
      RECT 6.77 3.175 6.82 3.86 ;
      RECT 6.56 3.6 6.595 3.86 ;
      RECT 6.875 3.175 6.88 3.635 ;
      RECT 6.965 3.175 6.99 3.455 ;
      RECT 7.24 4.557 7.245 4.82 ;
      RECT 7.205 4.545 7.24 4.82 ;
      RECT 7.145 4.518 7.205 4.82 ;
      RECT 7.14 4.501 7.145 4.674 ;
      RECT 7.135 4.498 7.14 4.661 ;
      RECT 7.115 4.491 7.135 4.648 ;
      RECT 7.08 4.474 7.115 4.63 ;
      RECT 7.04 4.453 7.08 4.61 ;
      RECT 7.035 4.441 7.04 4.598 ;
      RECT 6.995 4.427 7.035 4.584 ;
      RECT 6.975 4.41 6.995 4.566 ;
      RECT 6.965 4.402 6.975 4.558 ;
      RECT 6.95 3.175 6.965 3.473 ;
      RECT 6.935 4.392 6.965 4.545 ;
      RECT 6.92 3.175 6.95 3.518 ;
      RECT 6.925 4.382 6.935 4.532 ;
      RECT 6.895 4.367 6.925 4.519 ;
      RECT 6.88 3.175 6.92 3.585 ;
      RECT 6.88 4.335 6.895 4.505 ;
      RECT 6.875 4.307 6.88 4.499 ;
      RECT 6.87 3.175 6.875 3.64 ;
      RECT 6.86 4.277 6.875 4.493 ;
      RECT 6.865 3.175 6.87 3.653 ;
      RECT 6.855 3.175 6.865 3.673 ;
      RECT 6.82 4.19 6.86 4.478 ;
      RECT 6.82 3.175 6.855 3.713 ;
      RECT 6.815 4.122 6.82 4.466 ;
      RECT 6.8 4.077 6.815 4.461 ;
      RECT 6.795 4.015 6.8 4.456 ;
      RECT 6.77 3.922 6.795 4.449 ;
      RECT 6.765 3.175 6.77 4.441 ;
      RECT 6.75 3.175 6.765 4.428 ;
      RECT 6.73 3.175 6.75 4.385 ;
      RECT 6.72 3.175 6.73 4.335 ;
      RECT 6.715 3.175 6.72 4.308 ;
      RECT 6.71 3.175 6.715 4.286 ;
      RECT 6.705 3.401 6.71 4.269 ;
      RECT 6.7 3.423 6.705 4.247 ;
      RECT 6.695 3.465 6.7 4.23 ;
      RECT 6.665 3.515 6.695 4.174 ;
      RECT 6.66 3.542 6.665 4.116 ;
      RECT 6.645 3.56 6.66 4.08 ;
      RECT 6.64 3.578 6.645 4.044 ;
      RECT 6.634 3.585 6.64 4.025 ;
      RECT 6.63 3.592 6.634 4.008 ;
      RECT 6.625 3.597 6.63 3.977 ;
      RECT 6.615 3.6 6.625 3.952 ;
      RECT 6.605 3.6 6.615 3.918 ;
      RECT 6.6 3.6 6.605 3.895 ;
      RECT 6.595 3.6 6.6 3.875 ;
      RECT 5.51 3.735 5.79 4.015 ;
      RECT 5.51 3.735 5.81 3.91 ;
      RECT 5.6 3.625 5.86 3.885 ;
      RECT 5.565 3.72 5.86 3.885 ;
      RECT 5.69 2.24 5.855 3.885 ;
      RECT 5.59 2.24 5.96 2.61 ;
      RECT 5.215 4.765 5.475 5.025 ;
      RECT 5.235 4.692 5.415 5.025 ;
      RECT 5.235 4.435 5.41 5.025 ;
      RECT 5.235 4.227 5.4 5.025 ;
      RECT 5.24 4.145 5.4 5.025 ;
      RECT 5.24 3.91 5.39 5.025 ;
      RECT 5.24 3.757 5.385 5.025 ;
      RECT 5.245 3.742 5.385 5.025 ;
      RECT 5.295 3.457 5.385 5.025 ;
      RECT 5.25 3.692 5.385 5.025 ;
      RECT 5.28 3.51 5.385 5.025 ;
      RECT 5.265 3.622 5.385 5.025 ;
      RECT 5.27 3.58 5.385 5.025 ;
      RECT 5.265 3.622 5.4 3.685 ;
      RECT 5.3 3.21 5.405 3.63 ;
      RECT 5.3 3.21 5.42 3.613 ;
      RECT 5.3 3.21 5.455 3.575 ;
      RECT 5.295 3.457 5.505 3.508 ;
      RECT 5.3 3.21 5.56 3.47 ;
      RECT 4.56 3.915 4.82 4.175 ;
      RECT 4.56 3.915 4.83 4.133 ;
      RECT 4.56 3.915 4.916 4.104 ;
      RECT 4.56 3.915 4.985 4.056 ;
      RECT 4.56 3.915 5.02 4.025 ;
      RECT 4.79 3.735 5.07 4.015 ;
      RECT 4.625 3.9 5.07 4.015 ;
      RECT 4.715 3.777 4.82 4.175 ;
      RECT 4.645 3.84 5.07 4.015 ;
      RECT 70.065 9.345 70.435 9.715 ;
      RECT 54.805 9.345 55.175 9.715 ;
      RECT 39.545 9.345 39.915 9.715 ;
      RECT 24.285 9.345 24.655 9.715 ;
      RECT 9.025 9.345 9.395 9.715 ;
    LAYER via1 ;
      RECT 78.655 9.665 78.805 9.815 ;
      RECT 76.285 9.03 76.435 9.18 ;
      RECT 76.27 3.36 76.42 3.51 ;
      RECT 75.48 3.745 75.63 3.895 ;
      RECT 75.48 8.615 75.63 8.765 ;
      RECT 73.89 4.1 74.04 4.25 ;
      RECT 72.12 3.645 72.27 3.795 ;
      RECT 71.1 4.35 71.25 4.5 ;
      RECT 70.87 3.77 71.02 3.92 ;
      RECT 70.835 9 70.985 9.15 ;
      RECT 70.525 4.37 70.675 4.52 ;
      RECT 70.285 3.39 70.435 3.54 ;
      RECT 70.175 9.455 70.325 9.605 ;
      RECT 69.975 4.72 70.125 4.87 ;
      RECT 69.835 3.325 69.985 3.475 ;
      RECT 69.2 3.41 69.35 3.56 ;
      RECT 69.09 4.05 69.24 4.2 ;
      RECT 68.765 4.61 68.915 4.76 ;
      RECT 68.595 3.6 68.745 3.75 ;
      RECT 68.24 4.615 68.39 4.765 ;
      RECT 68.18 3.83 68.33 3.98 ;
      RECT 67.815 4.82 67.965 4.97 ;
      RECT 67.655 3.655 67.805 3.805 ;
      RECT 67.09 3.73 67.24 3.88 ;
      RECT 66.74 2.35 66.89 2.5 ;
      RECT 66.695 3.68 66.845 3.83 ;
      RECT 66.395 3.265 66.545 3.415 ;
      RECT 66.31 4.82 66.46 4.97 ;
      RECT 65.655 3.97 65.805 4.12 ;
      RECT 63.37 9.045 63.52 9.195 ;
      RECT 61.025 9.03 61.175 9.18 ;
      RECT 61.01 3.36 61.16 3.51 ;
      RECT 60.22 3.745 60.37 3.895 ;
      RECT 60.22 8.615 60.37 8.765 ;
      RECT 58.63 4.1 58.78 4.25 ;
      RECT 56.86 3.645 57.01 3.795 ;
      RECT 55.84 4.35 55.99 4.5 ;
      RECT 55.61 3.77 55.76 3.92 ;
      RECT 55.575 9 55.725 9.15 ;
      RECT 55.265 4.37 55.415 4.52 ;
      RECT 55.025 3.39 55.175 3.54 ;
      RECT 54.915 9.455 55.065 9.605 ;
      RECT 54.715 4.72 54.865 4.87 ;
      RECT 54.575 3.325 54.725 3.475 ;
      RECT 53.94 3.41 54.09 3.56 ;
      RECT 53.83 4.05 53.98 4.2 ;
      RECT 53.505 4.61 53.655 4.76 ;
      RECT 53.335 3.6 53.485 3.75 ;
      RECT 52.98 4.615 53.13 4.765 ;
      RECT 52.92 3.83 53.07 3.98 ;
      RECT 52.555 4.82 52.705 4.97 ;
      RECT 52.395 3.655 52.545 3.805 ;
      RECT 51.83 3.73 51.98 3.88 ;
      RECT 51.48 2.35 51.63 2.5 ;
      RECT 51.435 3.68 51.585 3.83 ;
      RECT 51.135 3.265 51.285 3.415 ;
      RECT 51.05 4.82 51.2 4.97 ;
      RECT 50.395 3.97 50.545 4.12 ;
      RECT 48.11 9.045 48.26 9.195 ;
      RECT 45.765 9.03 45.915 9.18 ;
      RECT 45.75 3.36 45.9 3.51 ;
      RECT 44.96 3.745 45.11 3.895 ;
      RECT 44.96 8.615 45.11 8.765 ;
      RECT 43.37 4.1 43.52 4.25 ;
      RECT 41.6 3.645 41.75 3.795 ;
      RECT 40.58 4.35 40.73 4.5 ;
      RECT 40.35 3.77 40.5 3.92 ;
      RECT 40.315 9.005 40.465 9.155 ;
      RECT 40.005 4.37 40.155 4.52 ;
      RECT 39.765 3.39 39.915 3.54 ;
      RECT 39.655 9.455 39.805 9.605 ;
      RECT 39.455 4.72 39.605 4.87 ;
      RECT 39.315 3.325 39.465 3.475 ;
      RECT 38.68 3.41 38.83 3.56 ;
      RECT 38.57 4.05 38.72 4.2 ;
      RECT 38.245 4.61 38.395 4.76 ;
      RECT 38.075 3.6 38.225 3.75 ;
      RECT 37.72 4.615 37.87 4.765 ;
      RECT 37.66 3.83 37.81 3.98 ;
      RECT 37.295 4.82 37.445 4.97 ;
      RECT 37.135 3.655 37.285 3.805 ;
      RECT 36.57 3.73 36.72 3.88 ;
      RECT 36.22 2.35 36.37 2.5 ;
      RECT 36.175 3.68 36.325 3.83 ;
      RECT 35.875 3.265 36.025 3.415 ;
      RECT 35.79 4.82 35.94 4.97 ;
      RECT 35.135 3.97 35.285 4.12 ;
      RECT 32.895 9.05 33.045 9.2 ;
      RECT 30.505 9.03 30.655 9.18 ;
      RECT 30.49 3.36 30.64 3.51 ;
      RECT 29.7 3.745 29.85 3.895 ;
      RECT 29.7 8.615 29.85 8.765 ;
      RECT 28.11 4.1 28.26 4.25 ;
      RECT 26.34 3.645 26.49 3.795 ;
      RECT 25.32 4.35 25.47 4.5 ;
      RECT 25.09 3.77 25.24 3.92 ;
      RECT 25.055 9 25.205 9.15 ;
      RECT 24.745 4.37 24.895 4.52 ;
      RECT 24.505 3.39 24.655 3.54 ;
      RECT 24.395 9.455 24.545 9.605 ;
      RECT 24.195 4.72 24.345 4.87 ;
      RECT 24.055 3.325 24.205 3.475 ;
      RECT 23.42 3.41 23.57 3.56 ;
      RECT 23.31 4.05 23.46 4.2 ;
      RECT 22.985 4.61 23.135 4.76 ;
      RECT 22.815 3.6 22.965 3.75 ;
      RECT 22.46 4.615 22.61 4.765 ;
      RECT 22.4 3.83 22.55 3.98 ;
      RECT 22.035 4.82 22.185 4.97 ;
      RECT 21.875 3.655 22.025 3.805 ;
      RECT 21.31 3.73 21.46 3.88 ;
      RECT 20.96 2.35 21.11 2.5 ;
      RECT 20.915 3.68 21.065 3.83 ;
      RECT 20.615 3.265 20.765 3.415 ;
      RECT 20.53 4.82 20.68 4.97 ;
      RECT 19.875 3.97 20.025 4.12 ;
      RECT 17.635 9.045 17.785 9.195 ;
      RECT 15.245 9.03 15.395 9.18 ;
      RECT 15.23 3.36 15.38 3.51 ;
      RECT 14.44 3.745 14.59 3.895 ;
      RECT 14.44 8.615 14.59 8.765 ;
      RECT 12.85 4.1 13 4.25 ;
      RECT 11.08 3.645 11.23 3.795 ;
      RECT 10.06 4.35 10.21 4.5 ;
      RECT 9.83 3.77 9.98 3.92 ;
      RECT 9.795 8.995 9.945 9.145 ;
      RECT 9.485 4.37 9.635 4.52 ;
      RECT 9.245 3.39 9.395 3.54 ;
      RECT 9.135 9.455 9.285 9.605 ;
      RECT 8.935 4.72 9.085 4.87 ;
      RECT 8.795 3.325 8.945 3.475 ;
      RECT 8.16 3.41 8.31 3.56 ;
      RECT 8.05 4.05 8.2 4.2 ;
      RECT 7.725 4.61 7.875 4.76 ;
      RECT 7.555 3.6 7.705 3.75 ;
      RECT 7.2 4.615 7.35 4.765 ;
      RECT 7.14 3.83 7.29 3.98 ;
      RECT 6.775 4.82 6.925 4.97 ;
      RECT 6.615 3.655 6.765 3.805 ;
      RECT 6.05 3.73 6.2 3.88 ;
      RECT 5.7 2.35 5.85 2.5 ;
      RECT 5.655 3.68 5.805 3.83 ;
      RECT 5.355 3.265 5.505 3.415 ;
      RECT 5.27 4.82 5.42 4.97 ;
      RECT 4.615 3.97 4.765 4.12 ;
      RECT 1.64 9.385 1.79 9.535 ;
      RECT 1.265 8.645 1.415 8.795 ;
    LAYER met1 ;
      RECT 64.615 0 73.355 3.035 ;
      RECT 49.355 0 58.095 3.035 ;
      RECT 34.095 0 42.835 3.035 ;
      RECT 18.835 0 27.575 3.035 ;
      RECT 3.575 0 12.315 3.035 ;
      RECT 0.03 0 79.125 1.6 ;
      RECT 78.52 10.06 78.81 10.29 ;
      RECT 78.58 8.58 78.75 10.29 ;
      RECT 78.555 9.565 78.905 9.915 ;
      RECT 78.52 8.58 78.81 8.81 ;
      RECT 78.115 3.69 78.22 4.26 ;
      RECT 78.115 4.025 78.44 4.255 ;
      RECT 78.115 4.055 78.61 4.225 ;
      RECT 78.115 3.69 78.305 4.255 ;
      RECT 77.53 3.655 77.82 3.885 ;
      RECT 77.53 3.69 78.305 3.86 ;
      RECT 77.59 2.175 77.76 3.885 ;
      RECT 77.53 2.175 77.82 2.405 ;
      RECT 77.53 10.06 77.82 10.29 ;
      RECT 77.59 8.58 77.76 10.29 ;
      RECT 77.53 8.58 77.82 8.81 ;
      RECT 77.53 8.615 78.38 8.775 ;
      RECT 78.215 8.21 78.38 8.775 ;
      RECT 77.53 8.61 77.925 8.775 ;
      RECT 78.15 8.21 78.44 8.44 ;
      RECT 78.15 8.24 78.61 8.41 ;
      RECT 77.16 4.025 77.45 4.255 ;
      RECT 77.16 4.055 77.62 4.225 ;
      RECT 77.225 2.95 77.39 4.255 ;
      RECT 75.74 2.92 76.03 3.15 ;
      RECT 75.74 2.95 77.39 3.12 ;
      RECT 75.8 2.18 75.97 3.15 ;
      RECT 75.74 2.18 76.03 2.41 ;
      RECT 75.74 10.055 76.03 10.285 ;
      RECT 75.8 9.315 75.97 10.285 ;
      RECT 75.8 9.41 77.39 9.58 ;
      RECT 77.22 8.21 77.39 9.58 ;
      RECT 75.74 9.315 76.03 9.545 ;
      RECT 77.16 8.21 77.45 8.44 ;
      RECT 77.16 8.24 77.62 8.41 ;
      RECT 73.79 4 74.13 4.35 ;
      RECT 73.88 3.32 74.05 4.35 ;
      RECT 76.17 3.26 76.52 3.61 ;
      RECT 73.88 3.32 76.52 3.49 ;
      RECT 76.195 8.945 76.52 9.27 ;
      RECT 70.735 8.9 71.085 9.25 ;
      RECT 76.17 8.945 76.52 9.175 ;
      RECT 70.535 8.945 71.085 9.175 ;
      RECT 70.365 8.975 76.52 9.145 ;
      RECT 75.395 3.66 75.715 3.98 ;
      RECT 75.365 3.66 75.715 3.89 ;
      RECT 75.195 3.69 75.715 3.86 ;
      RECT 75.395 8.545 75.715 8.835 ;
      RECT 75.365 8.575 75.715 8.805 ;
      RECT 75.195 8.605 75.715 8.775 ;
      RECT 71.085 4.28 71.235 4.555 ;
      RECT 71.625 3.36 71.63 3.58 ;
      RECT 72.775 3.56 72.79 3.758 ;
      RECT 72.74 3.552 72.775 3.765 ;
      RECT 72.71 3.545 72.74 3.765 ;
      RECT 72.655 3.51 72.71 3.765 ;
      RECT 72.59 3.447 72.655 3.765 ;
      RECT 72.585 3.412 72.59 3.763 ;
      RECT 72.58 3.407 72.585 3.755 ;
      RECT 72.575 3.402 72.58 3.741 ;
      RECT 72.57 3.399 72.575 3.734 ;
      RECT 72.525 3.389 72.57 3.685 ;
      RECT 72.505 3.376 72.525 3.62 ;
      RECT 72.5 3.371 72.505 3.593 ;
      RECT 72.495 3.37 72.5 3.586 ;
      RECT 72.49 3.369 72.495 3.579 ;
      RECT 72.405 3.354 72.49 3.525 ;
      RECT 72.375 3.335 72.405 3.475 ;
      RECT 72.295 3.318 72.375 3.46 ;
      RECT 72.26 3.305 72.295 3.445 ;
      RECT 72.252 3.305 72.26 3.44 ;
      RECT 72.166 3.306 72.252 3.44 ;
      RECT 72.08 3.308 72.166 3.44 ;
      RECT 72.055 3.309 72.08 3.444 ;
      RECT 71.98 3.315 72.055 3.459 ;
      RECT 71.897 3.327 71.98 3.483 ;
      RECT 71.811 3.34 71.897 3.509 ;
      RECT 71.725 3.353 71.811 3.535 ;
      RECT 71.69 3.362 71.725 3.554 ;
      RECT 71.64 3.362 71.69 3.567 ;
      RECT 71.63 3.36 71.64 3.578 ;
      RECT 71.615 3.357 71.625 3.58 ;
      RECT 71.6 3.349 71.615 3.588 ;
      RECT 71.585 3.341 71.6 3.608 ;
      RECT 71.58 3.336 71.585 3.665 ;
      RECT 71.565 3.331 71.58 3.738 ;
      RECT 71.56 3.326 71.565 3.78 ;
      RECT 71.555 3.324 71.56 3.808 ;
      RECT 71.55 3.322 71.555 3.83 ;
      RECT 71.54 3.318 71.55 3.873 ;
      RECT 71.535 3.315 71.54 3.898 ;
      RECT 71.53 3.313 71.535 3.918 ;
      RECT 71.525 3.311 71.53 3.942 ;
      RECT 71.52 3.307 71.525 3.965 ;
      RECT 71.515 3.303 71.52 3.988 ;
      RECT 71.48 3.293 71.515 4.095 ;
      RECT 71.475 3.283 71.48 4.193 ;
      RECT 71.47 3.281 71.475 4.22 ;
      RECT 71.465 3.28 71.47 4.24 ;
      RECT 71.46 3.272 71.465 4.26 ;
      RECT 71.455 3.267 71.46 4.295 ;
      RECT 71.45 3.265 71.455 4.313 ;
      RECT 71.445 3.265 71.45 4.338 ;
      RECT 71.44 3.265 71.445 4.36 ;
      RECT 71.405 3.265 71.44 4.403 ;
      RECT 71.38 3.265 71.405 4.432 ;
      RECT 71.37 3.265 71.38 3.618 ;
      RECT 71.373 3.675 71.38 4.442 ;
      RECT 71.37 3.732 71.373 4.445 ;
      RECT 71.365 3.265 71.37 3.59 ;
      RECT 71.365 3.782 71.37 4.448 ;
      RECT 71.355 3.265 71.365 3.58 ;
      RECT 71.36 3.835 71.365 4.451 ;
      RECT 71.355 3.92 71.36 4.455 ;
      RECT 71.345 3.265 71.355 3.568 ;
      RECT 71.35 3.967 71.355 4.459 ;
      RECT 71.345 4.042 71.35 4.463 ;
      RECT 71.31 3.265 71.345 3.543 ;
      RECT 71.335 4.125 71.345 4.468 ;
      RECT 71.325 4.192 71.335 4.475 ;
      RECT 71.32 4.22 71.325 4.48 ;
      RECT 71.31 4.233 71.32 4.486 ;
      RECT 71.265 3.265 71.31 3.5 ;
      RECT 71.305 4.238 71.31 4.493 ;
      RECT 71.265 4.255 71.305 4.555 ;
      RECT 71.26 3.267 71.265 3.473 ;
      RECT 71.235 4.275 71.265 4.555 ;
      RECT 71.255 3.272 71.26 3.445 ;
      RECT 71.045 4.284 71.085 4.555 ;
      RECT 71.02 4.292 71.045 4.525 ;
      RECT 70.975 4.3 71.02 4.525 ;
      RECT 70.96 4.305 70.975 4.52 ;
      RECT 70.95 4.305 70.96 4.514 ;
      RECT 70.94 4.312 70.95 4.511 ;
      RECT 70.935 4.35 70.94 4.5 ;
      RECT 70.93 4.412 70.935 4.478 ;
      RECT 72.2 4.287 72.385 4.51 ;
      RECT 72.2 4.302 72.39 4.506 ;
      RECT 72.19 3.575 72.275 4.505 ;
      RECT 72.19 4.302 72.395 4.499 ;
      RECT 72.185 4.31 72.395 4.498 ;
      RECT 72.39 4.03 72.71 4.35 ;
      RECT 72.185 4.202 72.355 4.293 ;
      RECT 72.18 4.202 72.355 4.275 ;
      RECT 72.17 4.01 72.305 4.25 ;
      RECT 72.165 4.01 72.305 4.195 ;
      RECT 72.125 3.59 72.295 4.095 ;
      RECT 72.11 3.59 72.295 3.965 ;
      RECT 72.105 3.59 72.295 3.918 ;
      RECT 72.1 3.59 72.295 3.898 ;
      RECT 72.095 3.59 72.295 3.873 ;
      RECT 72.065 3.59 72.325 3.85 ;
      RECT 72.075 3.587 72.285 3.85 ;
      RECT 72.2 3.582 72.285 4.51 ;
      RECT 72.085 3.575 72.275 3.85 ;
      RECT 72.08 3.58 72.275 3.85 ;
      RECT 70.91 3.792 71.095 4.005 ;
      RECT 70.91 3.8 71.105 3.998 ;
      RECT 70.89 3.8 71.105 3.995 ;
      RECT 70.885 3.8 71.105 3.98 ;
      RECT 70.815 3.715 71.075 3.975 ;
      RECT 70.815 3.86 71.11 3.888 ;
      RECT 70.47 4.315 70.73 4.575 ;
      RECT 70.495 4.26 70.69 4.575 ;
      RECT 70.49 4.009 70.67 4.303 ;
      RECT 70.49 4.015 70.68 4.303 ;
      RECT 70.47 4.017 70.68 4.248 ;
      RECT 70.465 4.027 70.68 4.115 ;
      RECT 70.495 4.007 70.67 4.575 ;
      RECT 70.581 4.005 70.67 4.575 ;
      RECT 70.44 3.225 70.475 3.595 ;
      RECT 70.23 3.335 70.235 3.595 ;
      RECT 70.475 3.232 70.49 3.595 ;
      RECT 70.365 3.225 70.44 3.673 ;
      RECT 70.355 3.225 70.365 3.758 ;
      RECT 70.33 3.225 70.355 3.793 ;
      RECT 70.29 3.225 70.33 3.861 ;
      RECT 70.28 3.232 70.29 3.913 ;
      RECT 70.25 3.335 70.28 3.954 ;
      RECT 70.245 3.335 70.25 3.993 ;
      RECT 70.235 3.335 70.245 4.013 ;
      RECT 70.23 3.63 70.235 4.05 ;
      RECT 70.225 3.647 70.23 4.07 ;
      RECT 70.21 3.71 70.225 4.11 ;
      RECT 70.205 3.753 70.21 4.145 ;
      RECT 70.2 3.761 70.205 4.158 ;
      RECT 70.19 3.775 70.2 4.18 ;
      RECT 70.165 3.81 70.19 4.245 ;
      RECT 70.155 3.845 70.165 4.308 ;
      RECT 70.135 3.875 70.155 4.369 ;
      RECT 70.12 3.911 70.135 4.436 ;
      RECT 70.11 3.939 70.12 4.475 ;
      RECT 70.1 3.961 70.11 4.495 ;
      RECT 70.095 3.971 70.1 4.506 ;
      RECT 70.09 3.98 70.095 4.509 ;
      RECT 70.08 3.998 70.09 4.513 ;
      RECT 70.07 4.016 70.08 4.514 ;
      RECT 70.045 4.055 70.07 4.511 ;
      RECT 70.025 4.097 70.045 4.508 ;
      RECT 70.01 4.135 70.025 4.507 ;
      RECT 69.975 4.17 70.01 4.504 ;
      RECT 69.97 4.192 69.975 4.502 ;
      RECT 69.905 4.232 69.97 4.499 ;
      RECT 69.9 4.272 69.905 4.495 ;
      RECT 69.885 4.282 69.9 4.486 ;
      RECT 69.875 4.402 69.885 4.471 ;
      RECT 70.355 4.815 70.365 5.075 ;
      RECT 70.355 4.818 70.375 5.074 ;
      RECT 70.345 4.808 70.355 5.073 ;
      RECT 70.335 4.823 70.415 5.069 ;
      RECT 70.32 4.802 70.335 5.067 ;
      RECT 70.295 4.827 70.42 5.063 ;
      RECT 70.28 4.787 70.295 5.058 ;
      RECT 70.28 4.829 70.43 5.057 ;
      RECT 70.28 4.837 70.445 5.05 ;
      RECT 70.22 4.774 70.28 5.04 ;
      RECT 70.21 4.761 70.22 5.022 ;
      RECT 70.185 4.751 70.21 5.012 ;
      RECT 70.18 4.741 70.185 5.004 ;
      RECT 70.115 4.837 70.445 4.986 ;
      RECT 70.03 4.837 70.445 4.948 ;
      RECT 69.92 4.665 70.18 4.925 ;
      RECT 70.295 4.795 70.32 5.063 ;
      RECT 70.335 4.805 70.345 5.069 ;
      RECT 69.92 4.813 70.36 4.925 ;
      RECT 70.105 10.055 70.395 10.285 ;
      RECT 70.165 9.315 70.335 10.285 ;
      RECT 70.065 9.345 70.435 9.715 ;
      RECT 70.105 9.315 70.395 9.715 ;
      RECT 69.135 4.57 69.165 4.87 ;
      RECT 68.91 4.555 68.915 4.83 ;
      RECT 68.71 4.555 68.865 4.815 ;
      RECT 70.01 3.27 70.04 3.53 ;
      RECT 70 3.27 70.01 3.638 ;
      RECT 69.98 3.27 70 3.648 ;
      RECT 69.965 3.27 69.98 3.66 ;
      RECT 69.91 3.27 69.965 3.71 ;
      RECT 69.895 3.27 69.91 3.758 ;
      RECT 69.865 3.27 69.895 3.793 ;
      RECT 69.81 3.27 69.865 3.855 ;
      RECT 69.79 3.27 69.81 3.923 ;
      RECT 69.785 3.27 69.79 3.953 ;
      RECT 69.78 3.27 69.785 3.965 ;
      RECT 69.775 3.387 69.78 3.983 ;
      RECT 69.755 3.405 69.775 4.008 ;
      RECT 69.735 3.432 69.755 4.058 ;
      RECT 69.73 3.452 69.735 4.089 ;
      RECT 69.725 3.46 69.73 4.106 ;
      RECT 69.71 3.486 69.725 4.135 ;
      RECT 69.695 3.528 69.71 4.17 ;
      RECT 69.69 3.557 69.695 4.193 ;
      RECT 69.685 3.572 69.69 4.206 ;
      RECT 69.68 3.595 69.685 4.217 ;
      RECT 69.67 3.615 69.68 4.235 ;
      RECT 69.66 3.645 69.67 4.258 ;
      RECT 69.655 3.667 69.66 4.278 ;
      RECT 69.65 3.682 69.655 4.293 ;
      RECT 69.635 3.712 69.65 4.32 ;
      RECT 69.63 3.742 69.635 4.346 ;
      RECT 69.625 3.76 69.63 4.358 ;
      RECT 69.615 3.79 69.625 4.377 ;
      RECT 69.605 3.815 69.615 4.402 ;
      RECT 69.6 3.835 69.605 4.421 ;
      RECT 69.595 3.852 69.6 4.434 ;
      RECT 69.585 3.878 69.595 4.453 ;
      RECT 69.575 3.916 69.585 4.48 ;
      RECT 69.57 3.942 69.575 4.5 ;
      RECT 69.565 3.952 69.57 4.51 ;
      RECT 69.56 3.965 69.565 4.525 ;
      RECT 69.555 3.98 69.56 4.535 ;
      RECT 69.55 4.002 69.555 4.55 ;
      RECT 69.545 4.02 69.55 4.561 ;
      RECT 69.54 4.03 69.545 4.572 ;
      RECT 69.535 4.038 69.54 4.584 ;
      RECT 69.53 4.046 69.535 4.595 ;
      RECT 69.525 4.072 69.53 4.608 ;
      RECT 69.515 4.1 69.525 4.621 ;
      RECT 69.51 4.13 69.515 4.63 ;
      RECT 69.505 4.145 69.51 4.637 ;
      RECT 69.49 4.17 69.505 4.644 ;
      RECT 69.485 4.192 69.49 4.65 ;
      RECT 69.48 4.217 69.485 4.653 ;
      RECT 69.471 4.245 69.48 4.657 ;
      RECT 69.465 4.262 69.471 4.662 ;
      RECT 69.46 4.28 69.465 4.666 ;
      RECT 69.455 4.292 69.46 4.669 ;
      RECT 69.45 4.313 69.455 4.673 ;
      RECT 69.445 4.331 69.45 4.676 ;
      RECT 69.44 4.345 69.445 4.679 ;
      RECT 69.435 4.362 69.44 4.682 ;
      RECT 69.43 4.375 69.435 4.685 ;
      RECT 69.405 4.412 69.43 4.693 ;
      RECT 69.4 4.457 69.405 4.702 ;
      RECT 69.395 4.485 69.4 4.705 ;
      RECT 69.385 4.505 69.395 4.709 ;
      RECT 69.38 4.525 69.385 4.714 ;
      RECT 69.375 4.54 69.38 4.717 ;
      RECT 69.355 4.55 69.375 4.724 ;
      RECT 69.29 4.557 69.355 4.75 ;
      RECT 69.255 4.56 69.29 4.778 ;
      RECT 69.24 4.563 69.255 4.793 ;
      RECT 69.23 4.564 69.24 4.808 ;
      RECT 69.22 4.565 69.23 4.825 ;
      RECT 69.215 4.565 69.22 4.84 ;
      RECT 69.21 4.565 69.215 4.848 ;
      RECT 69.195 4.566 69.21 4.863 ;
      RECT 69.165 4.568 69.195 4.87 ;
      RECT 69.055 4.575 69.135 4.87 ;
      RECT 69.01 4.58 69.055 4.87 ;
      RECT 69 4.581 69.01 4.86 ;
      RECT 68.99 4.582 69 4.853 ;
      RECT 68.97 4.584 68.99 4.848 ;
      RECT 68.96 4.555 68.97 4.843 ;
      RECT 68.915 4.555 68.96 4.835 ;
      RECT 68.885 4.555 68.91 4.825 ;
      RECT 68.865 4.555 68.885 4.818 ;
      RECT 69.145 3.355 69.405 3.615 ;
      RECT 69.025 3.37 69.035 3.535 ;
      RECT 69.01 3.37 69.015 3.53 ;
      RECT 66.375 3.21 66.56 3.5 ;
      RECT 68.19 3.335 68.205 3.49 ;
      RECT 66.34 3.21 66.365 3.47 ;
      RECT 68.755 3.26 68.76 3.402 ;
      RECT 68.67 3.255 68.695 3.395 ;
      RECT 69.07 3.372 69.145 3.565 ;
      RECT 69.055 3.37 69.07 3.548 ;
      RECT 69.035 3.37 69.055 3.54 ;
      RECT 69.015 3.37 69.025 3.533 ;
      RECT 68.97 3.365 69.01 3.523 ;
      RECT 68.93 3.34 68.97 3.508 ;
      RECT 68.915 3.315 68.93 3.498 ;
      RECT 68.91 3.309 68.915 3.496 ;
      RECT 68.875 3.301 68.91 3.479 ;
      RECT 68.87 3.294 68.875 3.467 ;
      RECT 68.85 3.289 68.87 3.455 ;
      RECT 68.84 3.283 68.85 3.44 ;
      RECT 68.82 3.278 68.84 3.425 ;
      RECT 68.81 3.273 68.82 3.418 ;
      RECT 68.805 3.271 68.81 3.413 ;
      RECT 68.8 3.27 68.805 3.41 ;
      RECT 68.76 3.265 68.8 3.406 ;
      RECT 68.74 3.259 68.755 3.401 ;
      RECT 68.705 3.256 68.74 3.398 ;
      RECT 68.695 3.255 68.705 3.396 ;
      RECT 68.635 3.255 68.67 3.393 ;
      RECT 68.59 3.255 68.635 3.393 ;
      RECT 68.54 3.255 68.59 3.396 ;
      RECT 68.525 3.257 68.54 3.398 ;
      RECT 68.51 3.26 68.525 3.399 ;
      RECT 68.5 3.265 68.51 3.4 ;
      RECT 68.47 3.27 68.5 3.405 ;
      RECT 68.46 3.276 68.47 3.413 ;
      RECT 68.45 3.278 68.46 3.417 ;
      RECT 68.44 3.282 68.45 3.421 ;
      RECT 68.415 3.288 68.44 3.429 ;
      RECT 68.405 3.293 68.415 3.437 ;
      RECT 68.39 3.297 68.405 3.441 ;
      RECT 68.355 3.303 68.39 3.449 ;
      RECT 68.335 3.308 68.355 3.459 ;
      RECT 68.305 3.315 68.335 3.468 ;
      RECT 68.26 3.324 68.305 3.482 ;
      RECT 68.255 3.329 68.26 3.493 ;
      RECT 68.235 3.332 68.255 3.494 ;
      RECT 68.205 3.335 68.235 3.492 ;
      RECT 68.17 3.335 68.19 3.488 ;
      RECT 68.1 3.335 68.17 3.479 ;
      RECT 68.085 3.332 68.1 3.471 ;
      RECT 68.045 3.325 68.085 3.466 ;
      RECT 68.02 3.315 68.045 3.459 ;
      RECT 68.015 3.309 68.02 3.456 ;
      RECT 67.975 3.303 68.015 3.453 ;
      RECT 67.96 3.296 67.975 3.448 ;
      RECT 67.94 3.292 67.96 3.443 ;
      RECT 67.925 3.287 67.94 3.439 ;
      RECT 67.91 3.282 67.925 3.437 ;
      RECT 67.895 3.278 67.91 3.436 ;
      RECT 67.88 3.276 67.895 3.432 ;
      RECT 67.87 3.274 67.88 3.427 ;
      RECT 67.855 3.271 67.87 3.423 ;
      RECT 67.845 3.269 67.855 3.418 ;
      RECT 67.825 3.266 67.845 3.414 ;
      RECT 67.78 3.265 67.825 3.412 ;
      RECT 67.72 3.267 67.78 3.413 ;
      RECT 67.7 3.269 67.72 3.415 ;
      RECT 67.67 3.272 67.7 3.416 ;
      RECT 67.62 3.277 67.67 3.418 ;
      RECT 67.615 3.28 67.62 3.42 ;
      RECT 67.605 3.282 67.615 3.423 ;
      RECT 67.6 3.284 67.605 3.426 ;
      RECT 67.55 3.287 67.6 3.433 ;
      RECT 67.53 3.291 67.55 3.445 ;
      RECT 67.52 3.294 67.53 3.451 ;
      RECT 67.51 3.295 67.52 3.454 ;
      RECT 67.471 3.298 67.51 3.456 ;
      RECT 67.385 3.305 67.471 3.459 ;
      RECT 67.311 3.315 67.385 3.463 ;
      RECT 67.225 3.326 67.311 3.468 ;
      RECT 67.21 3.333 67.225 3.47 ;
      RECT 67.155 3.337 67.21 3.471 ;
      RECT 67.141 3.34 67.155 3.473 ;
      RECT 67.055 3.34 67.141 3.475 ;
      RECT 67.015 3.337 67.055 3.478 ;
      RECT 66.991 3.333 67.015 3.48 ;
      RECT 66.905 3.323 66.991 3.483 ;
      RECT 66.875 3.312 66.905 3.484 ;
      RECT 66.856 3.308 66.875 3.483 ;
      RECT 66.77 3.301 66.856 3.48 ;
      RECT 66.71 3.29 66.77 3.477 ;
      RECT 66.69 3.282 66.71 3.475 ;
      RECT 66.655 3.277 66.69 3.474 ;
      RECT 66.63 3.272 66.655 3.473 ;
      RECT 66.6 3.267 66.63 3.472 ;
      RECT 66.575 3.21 66.6 3.471 ;
      RECT 66.56 3.21 66.575 3.495 ;
      RECT 66.365 3.21 66.375 3.495 ;
      RECT 68.14 4.23 68.145 4.37 ;
      RECT 67.8 4.23 67.835 4.368 ;
      RECT 67.375 4.215 67.39 4.36 ;
      RECT 69.205 3.995 69.295 4.255 ;
      RECT 69.035 3.86 69.135 4.255 ;
      RECT 66.07 3.835 66.15 4.045 ;
      RECT 69.16 3.972 69.205 4.255 ;
      RECT 69.15 3.942 69.16 4.255 ;
      RECT 69.135 3.865 69.15 4.255 ;
      RECT 68.95 3.86 69.035 4.22 ;
      RECT 68.945 3.862 68.95 4.215 ;
      RECT 68.94 3.867 68.945 4.215 ;
      RECT 68.905 3.967 68.94 4.215 ;
      RECT 68.895 3.995 68.905 4.215 ;
      RECT 68.885 4.01 68.895 4.215 ;
      RECT 68.875 4.022 68.885 4.215 ;
      RECT 68.87 4.032 68.875 4.215 ;
      RECT 68.855 4.042 68.87 4.217 ;
      RECT 68.85 4.057 68.855 4.219 ;
      RECT 68.835 4.07 68.85 4.221 ;
      RECT 68.83 4.085 68.835 4.224 ;
      RECT 68.81 4.095 68.83 4.228 ;
      RECT 68.795 4.105 68.81 4.231 ;
      RECT 68.76 4.112 68.795 4.236 ;
      RECT 68.716 4.119 68.76 4.244 ;
      RECT 68.63 4.131 68.716 4.257 ;
      RECT 68.605 4.142 68.63 4.268 ;
      RECT 68.575 4.147 68.605 4.273 ;
      RECT 68.54 4.152 68.575 4.281 ;
      RECT 68.51 4.157 68.54 4.288 ;
      RECT 68.485 4.162 68.51 4.293 ;
      RECT 68.42 4.169 68.485 4.302 ;
      RECT 68.35 4.182 68.42 4.318 ;
      RECT 68.32 4.192 68.35 4.33 ;
      RECT 68.295 4.197 68.32 4.337 ;
      RECT 68.24 4.204 68.295 4.345 ;
      RECT 68.235 4.211 68.24 4.35 ;
      RECT 68.23 4.213 68.235 4.351 ;
      RECT 68.215 4.215 68.23 4.353 ;
      RECT 68.21 4.215 68.215 4.356 ;
      RECT 68.145 4.222 68.21 4.363 ;
      RECT 68.11 4.232 68.14 4.373 ;
      RECT 68.093 4.235 68.11 4.375 ;
      RECT 68.007 4.234 68.093 4.374 ;
      RECT 67.921 4.232 68.007 4.371 ;
      RECT 67.835 4.231 67.921 4.369 ;
      RECT 67.734 4.229 67.8 4.368 ;
      RECT 67.648 4.226 67.734 4.366 ;
      RECT 67.562 4.222 67.648 4.364 ;
      RECT 67.476 4.219 67.562 4.363 ;
      RECT 67.39 4.216 67.476 4.361 ;
      RECT 67.29 4.215 67.375 4.358 ;
      RECT 67.24 4.213 67.29 4.356 ;
      RECT 67.22 4.21 67.24 4.354 ;
      RECT 67.2 4.208 67.22 4.351 ;
      RECT 67.175 4.204 67.2 4.348 ;
      RECT 67.13 4.198 67.175 4.343 ;
      RECT 67.09 4.192 67.13 4.335 ;
      RECT 67.065 4.187 67.09 4.328 ;
      RECT 67.01 4.18 67.065 4.32 ;
      RECT 66.986 4.173 67.01 4.313 ;
      RECT 66.9 4.164 66.986 4.303 ;
      RECT 66.87 4.156 66.9 4.293 ;
      RECT 66.84 4.152 66.87 4.288 ;
      RECT 66.835 4.149 66.84 4.285 ;
      RECT 66.83 4.148 66.835 4.285 ;
      RECT 66.755 4.141 66.83 4.278 ;
      RECT 66.716 4.132 66.755 4.267 ;
      RECT 66.63 4.122 66.716 4.255 ;
      RECT 66.59 4.112 66.63 4.243 ;
      RECT 66.551 4.107 66.59 4.236 ;
      RECT 66.465 4.097 66.551 4.225 ;
      RECT 66.425 4.085 66.465 4.214 ;
      RECT 66.39 4.07 66.425 4.207 ;
      RECT 66.38 4.06 66.39 4.204 ;
      RECT 66.36 4.045 66.38 4.202 ;
      RECT 66.33 4.015 66.36 4.198 ;
      RECT 66.32 3.995 66.33 4.193 ;
      RECT 66.315 3.987 66.32 4.19 ;
      RECT 66.31 3.98 66.315 4.188 ;
      RECT 66.295 3.967 66.31 4.181 ;
      RECT 66.29 3.957 66.295 4.173 ;
      RECT 66.285 3.95 66.29 4.168 ;
      RECT 66.28 3.945 66.285 4.164 ;
      RECT 66.265 3.932 66.28 4.156 ;
      RECT 66.26 3.842 66.265 4.145 ;
      RECT 66.255 3.837 66.26 4.138 ;
      RECT 66.18 3.835 66.255 4.098 ;
      RECT 66.15 3.835 66.18 4.053 ;
      RECT 66.055 3.84 66.07 4.04 ;
      RECT 68.54 3.545 68.8 3.805 ;
      RECT 68.525 3.533 68.705 3.77 ;
      RECT 68.52 3.534 68.705 3.768 ;
      RECT 68.505 3.538 68.715 3.758 ;
      RECT 68.5 3.543 68.72 3.728 ;
      RECT 68.505 3.54 68.72 3.758 ;
      RECT 68.52 3.535 68.715 3.768 ;
      RECT 68.54 3.532 68.705 3.805 ;
      RECT 68.54 3.531 68.695 3.805 ;
      RECT 68.565 3.53 68.695 3.805 ;
      RECT 68.125 3.775 68.385 4.035 ;
      RECT 68 3.82 68.385 4.03 ;
      RECT 67.99 3.825 68.385 4.025 ;
      RECT 68.005 4.765 68.02 5.075 ;
      RECT 66.6 4.535 66.61 4.665 ;
      RECT 66.38 4.53 66.485 4.665 ;
      RECT 66.295 4.535 66.345 4.665 ;
      RECT 64.845 3.27 64.85 4.375 ;
      RECT 68.1 4.857 68.105 4.993 ;
      RECT 68.095 4.852 68.1 5.053 ;
      RECT 68.09 4.85 68.095 5.066 ;
      RECT 68.075 4.847 68.09 5.068 ;
      RECT 68.07 4.842 68.075 5.07 ;
      RECT 68.065 4.838 68.07 5.073 ;
      RECT 68.05 4.833 68.065 5.075 ;
      RECT 68.02 4.825 68.05 5.075 ;
      RECT 67.981 4.765 68.005 5.075 ;
      RECT 67.895 4.765 67.981 5.072 ;
      RECT 67.865 4.765 67.895 5.065 ;
      RECT 67.84 4.765 67.865 5.058 ;
      RECT 67.815 4.765 67.84 5.05 ;
      RECT 67.8 4.765 67.815 5.043 ;
      RECT 67.775 4.765 67.8 5.035 ;
      RECT 67.76 4.765 67.775 5.028 ;
      RECT 67.72 4.775 67.76 5.017 ;
      RECT 67.71 4.77 67.72 5.007 ;
      RECT 67.706 4.769 67.71 5.004 ;
      RECT 67.62 4.761 67.706 4.987 ;
      RECT 67.587 4.75 67.62 4.964 ;
      RECT 67.501 4.739 67.587 4.942 ;
      RECT 67.415 4.723 67.501 4.911 ;
      RECT 67.345 4.708 67.415 4.883 ;
      RECT 67.335 4.701 67.345 4.87 ;
      RECT 67.305 4.698 67.335 4.86 ;
      RECT 67.28 4.694 67.305 4.853 ;
      RECT 67.265 4.691 67.28 4.848 ;
      RECT 67.26 4.69 67.265 4.843 ;
      RECT 67.23 4.685 67.26 4.836 ;
      RECT 67.225 4.68 67.23 4.831 ;
      RECT 67.21 4.677 67.225 4.826 ;
      RECT 67.205 4.672 67.21 4.821 ;
      RECT 67.185 4.667 67.205 4.818 ;
      RECT 67.17 4.662 67.185 4.81 ;
      RECT 67.155 4.656 67.17 4.805 ;
      RECT 67.125 4.647 67.155 4.798 ;
      RECT 67.12 4.64 67.125 4.79 ;
      RECT 67.115 4.638 67.12 4.788 ;
      RECT 67.11 4.637 67.115 4.785 ;
      RECT 67.07 4.63 67.11 4.778 ;
      RECT 67.056 4.62 67.07 4.768 ;
      RECT 67.005 4.609 67.056 4.756 ;
      RECT 66.98 4.595 67.005 4.742 ;
      RECT 66.955 4.584 66.98 4.734 ;
      RECT 66.935 4.573 66.955 4.728 ;
      RECT 66.925 4.567 66.935 4.723 ;
      RECT 66.92 4.565 66.925 4.719 ;
      RECT 66.9 4.56 66.92 4.714 ;
      RECT 66.87 4.55 66.9 4.704 ;
      RECT 66.865 4.542 66.87 4.697 ;
      RECT 66.85 4.54 66.865 4.693 ;
      RECT 66.83 4.54 66.85 4.688 ;
      RECT 66.825 4.539 66.83 4.686 ;
      RECT 66.82 4.539 66.825 4.683 ;
      RECT 66.78 4.538 66.82 4.678 ;
      RECT 66.755 4.537 66.78 4.673 ;
      RECT 66.695 4.536 66.755 4.67 ;
      RECT 66.61 4.535 66.695 4.668 ;
      RECT 66.571 4.534 66.6 4.665 ;
      RECT 66.485 4.532 66.571 4.665 ;
      RECT 66.345 4.532 66.38 4.665 ;
      RECT 66.255 4.536 66.295 4.668 ;
      RECT 66.24 4.539 66.255 4.675 ;
      RECT 66.23 4.54 66.24 4.682 ;
      RECT 66.205 4.543 66.23 4.687 ;
      RECT 66.2 4.545 66.205 4.69 ;
      RECT 66.15 4.547 66.2 4.691 ;
      RECT 66.111 4.551 66.15 4.693 ;
      RECT 66.025 4.553 66.111 4.696 ;
      RECT 66.007 4.555 66.025 4.698 ;
      RECT 65.921 4.558 66.007 4.7 ;
      RECT 65.835 4.562 65.921 4.703 ;
      RECT 65.798 4.566 65.835 4.706 ;
      RECT 65.712 4.569 65.798 4.709 ;
      RECT 65.626 4.573 65.712 4.712 ;
      RECT 65.54 4.578 65.626 4.716 ;
      RECT 65.52 4.58 65.54 4.719 ;
      RECT 65.5 4.579 65.52 4.72 ;
      RECT 65.451 4.576 65.5 4.721 ;
      RECT 65.365 4.571 65.451 4.724 ;
      RECT 65.315 4.566 65.365 4.726 ;
      RECT 65.291 4.564 65.315 4.727 ;
      RECT 65.205 4.559 65.291 4.729 ;
      RECT 65.18 4.555 65.205 4.728 ;
      RECT 65.17 4.552 65.18 4.726 ;
      RECT 65.16 4.545 65.17 4.723 ;
      RECT 65.155 4.525 65.16 4.718 ;
      RECT 65.145 4.495 65.155 4.713 ;
      RECT 65.13 4.365 65.145 4.704 ;
      RECT 65.125 4.357 65.13 4.697 ;
      RECT 65.105 4.35 65.125 4.689 ;
      RECT 65.1 4.332 65.105 4.681 ;
      RECT 65.09 4.312 65.1 4.676 ;
      RECT 65.085 4.285 65.09 4.672 ;
      RECT 65.08 4.262 65.085 4.669 ;
      RECT 65.06 4.22 65.08 4.661 ;
      RECT 65.025 4.135 65.06 4.645 ;
      RECT 65.02 4.067 65.025 4.633 ;
      RECT 65.005 4.037 65.02 4.627 ;
      RECT 65 3.282 65.005 3.528 ;
      RECT 64.99 4.007 65.005 4.618 ;
      RECT 64.995 3.277 65 3.56 ;
      RECT 64.99 3.272 64.995 3.603 ;
      RECT 64.985 3.27 64.99 3.638 ;
      RECT 64.97 3.97 64.99 4.608 ;
      RECT 64.98 3.27 64.985 3.675 ;
      RECT 64.965 3.27 64.98 3.773 ;
      RECT 64.965 3.943 64.97 4.601 ;
      RECT 64.96 3.27 64.965 3.848 ;
      RECT 64.96 3.931 64.965 4.598 ;
      RECT 64.955 3.27 64.96 3.88 ;
      RECT 64.955 3.91 64.96 4.595 ;
      RECT 64.95 3.27 64.955 4.592 ;
      RECT 64.915 3.27 64.95 4.578 ;
      RECT 64.9 3.27 64.915 4.56 ;
      RECT 64.88 3.27 64.9 4.55 ;
      RECT 64.855 3.27 64.88 4.533 ;
      RECT 64.85 3.27 64.855 4.483 ;
      RECT 64.84 3.27 64.845 4.313 ;
      RECT 64.835 3.27 64.84 4.22 ;
      RECT 64.83 3.27 64.835 4.133 ;
      RECT 64.825 3.27 64.83 4.065 ;
      RECT 64.82 3.27 64.825 4.008 ;
      RECT 64.81 3.27 64.82 3.903 ;
      RECT 64.805 3.27 64.81 3.775 ;
      RECT 64.8 3.27 64.805 3.693 ;
      RECT 64.795 3.272 64.8 3.61 ;
      RECT 64.79 3.277 64.795 3.543 ;
      RECT 64.785 3.282 64.79 3.47 ;
      RECT 67.6 3.6 67.86 3.86 ;
      RECT 67.62 3.567 67.83 3.86 ;
      RECT 67.62 3.565 67.82 3.86 ;
      RECT 67.63 3.552 67.82 3.86 ;
      RECT 67.63 3.55 67.745 3.86 ;
      RECT 67.105 3.675 67.28 3.955 ;
      RECT 67.1 3.675 67.28 3.953 ;
      RECT 67.1 3.675 67.295 3.95 ;
      RECT 67.09 3.675 67.295 3.948 ;
      RECT 67.035 3.675 67.295 3.935 ;
      RECT 67.035 3.75 67.3 3.913 ;
      RECT 66.58 3.687 66.6 3.93 ;
      RECT 66.58 3.687 66.64 3.929 ;
      RECT 66.575 3.689 66.64 3.928 ;
      RECT 66.575 3.689 66.726 3.927 ;
      RECT 66.575 3.689 66.795 3.926 ;
      RECT 66.575 3.689 66.815 3.918 ;
      RECT 66.555 3.692 66.815 3.916 ;
      RECT 66.54 3.702 66.815 3.901 ;
      RECT 66.54 3.702 66.83 3.9 ;
      RECT 66.535 3.711 66.83 3.892 ;
      RECT 66.535 3.711 66.835 3.888 ;
      RECT 66.64 3.625 66.9 3.885 ;
      RECT 66.53 3.713 66.9 3.77 ;
      RECT 66.6 3.68 66.9 3.885 ;
      RECT 66.565 4.873 66.57 5.08 ;
      RECT 66.515 4.867 66.565 5.079 ;
      RECT 66.482 4.881 66.575 5.078 ;
      RECT 66.396 4.881 66.575 5.077 ;
      RECT 66.31 4.881 66.575 5.076 ;
      RECT 66.31 4.98 66.58 5.073 ;
      RECT 66.305 4.98 66.58 5.068 ;
      RECT 66.3 4.98 66.58 5.05 ;
      RECT 66.295 4.98 66.58 5.033 ;
      RECT 66.255 4.765 66.515 5.025 ;
      RECT 65.715 3.915 65.801 4.329 ;
      RECT 65.715 3.915 65.84 4.326 ;
      RECT 65.715 3.915 65.86 4.316 ;
      RECT 65.67 3.915 65.86 4.313 ;
      RECT 65.67 4.067 65.87 4.303 ;
      RECT 65.67 4.088 65.875 4.297 ;
      RECT 65.67 4.106 65.88 4.293 ;
      RECT 65.67 4.126 65.89 4.288 ;
      RECT 65.645 4.126 65.89 4.285 ;
      RECT 65.635 4.126 65.89 4.263 ;
      RECT 65.635 4.142 65.895 4.233 ;
      RECT 65.6 3.915 65.86 4.22 ;
      RECT 65.6 4.154 65.9 4.175 ;
      RECT 63.26 10.06 63.55 10.29 ;
      RECT 63.32 8.58 63.49 10.29 ;
      RECT 63.27 8.945 63.62 9.295 ;
      RECT 63.26 8.58 63.55 8.81 ;
      RECT 62.855 3.69 62.96 4.26 ;
      RECT 62.855 4.025 63.18 4.255 ;
      RECT 62.855 4.055 63.35 4.225 ;
      RECT 62.855 3.69 63.045 4.255 ;
      RECT 62.27 3.655 62.56 3.885 ;
      RECT 62.27 3.69 63.045 3.86 ;
      RECT 62.33 2.175 62.5 3.885 ;
      RECT 62.27 2.175 62.56 2.405 ;
      RECT 62.27 10.06 62.56 10.29 ;
      RECT 62.33 8.58 62.5 10.29 ;
      RECT 62.27 8.58 62.56 8.81 ;
      RECT 62.27 8.615 63.12 8.775 ;
      RECT 62.955 8.21 63.12 8.775 ;
      RECT 62.27 8.61 62.665 8.775 ;
      RECT 62.89 8.21 63.18 8.44 ;
      RECT 62.89 8.24 63.35 8.41 ;
      RECT 61.9 4.025 62.19 4.255 ;
      RECT 61.9 4.055 62.36 4.225 ;
      RECT 61.965 2.95 62.13 4.255 ;
      RECT 60.48 2.92 60.77 3.15 ;
      RECT 60.48 2.95 62.13 3.12 ;
      RECT 60.54 2.18 60.71 3.15 ;
      RECT 60.48 2.18 60.77 2.41 ;
      RECT 60.48 10.055 60.77 10.285 ;
      RECT 60.54 9.315 60.71 10.285 ;
      RECT 60.54 9.41 62.13 9.58 ;
      RECT 61.96 8.21 62.13 9.58 ;
      RECT 60.48 9.315 60.77 9.545 ;
      RECT 61.9 8.21 62.19 8.44 ;
      RECT 61.9 8.24 62.36 8.41 ;
      RECT 58.53 4 58.87 4.35 ;
      RECT 58.62 3.32 58.79 4.35 ;
      RECT 60.91 3.26 61.26 3.61 ;
      RECT 58.62 3.32 61.26 3.49 ;
      RECT 60.935 8.945 61.26 9.27 ;
      RECT 55.475 8.9 55.825 9.25 ;
      RECT 60.91 8.945 61.26 9.175 ;
      RECT 55.275 8.945 55.825 9.175 ;
      RECT 55.105 8.975 61.26 9.145 ;
      RECT 60.135 3.66 60.455 3.98 ;
      RECT 60.105 3.66 60.455 3.89 ;
      RECT 59.935 3.69 60.455 3.86 ;
      RECT 60.135 8.545 60.455 8.835 ;
      RECT 60.105 8.575 60.455 8.805 ;
      RECT 59.935 8.605 60.455 8.775 ;
      RECT 55.825 4.28 55.975 4.555 ;
      RECT 56.365 3.36 56.37 3.58 ;
      RECT 57.515 3.56 57.53 3.758 ;
      RECT 57.48 3.552 57.515 3.765 ;
      RECT 57.45 3.545 57.48 3.765 ;
      RECT 57.395 3.51 57.45 3.765 ;
      RECT 57.33 3.447 57.395 3.765 ;
      RECT 57.325 3.412 57.33 3.763 ;
      RECT 57.32 3.407 57.325 3.755 ;
      RECT 57.315 3.402 57.32 3.741 ;
      RECT 57.31 3.399 57.315 3.734 ;
      RECT 57.265 3.389 57.31 3.685 ;
      RECT 57.245 3.376 57.265 3.62 ;
      RECT 57.24 3.371 57.245 3.593 ;
      RECT 57.235 3.37 57.24 3.586 ;
      RECT 57.23 3.369 57.235 3.579 ;
      RECT 57.145 3.354 57.23 3.525 ;
      RECT 57.115 3.335 57.145 3.475 ;
      RECT 57.035 3.318 57.115 3.46 ;
      RECT 57 3.305 57.035 3.445 ;
      RECT 56.992 3.305 57 3.44 ;
      RECT 56.906 3.306 56.992 3.44 ;
      RECT 56.82 3.308 56.906 3.44 ;
      RECT 56.795 3.309 56.82 3.444 ;
      RECT 56.72 3.315 56.795 3.459 ;
      RECT 56.637 3.327 56.72 3.483 ;
      RECT 56.551 3.34 56.637 3.509 ;
      RECT 56.465 3.353 56.551 3.535 ;
      RECT 56.43 3.362 56.465 3.554 ;
      RECT 56.38 3.362 56.43 3.567 ;
      RECT 56.37 3.36 56.38 3.578 ;
      RECT 56.355 3.357 56.365 3.58 ;
      RECT 56.34 3.349 56.355 3.588 ;
      RECT 56.325 3.341 56.34 3.608 ;
      RECT 56.32 3.336 56.325 3.665 ;
      RECT 56.305 3.331 56.32 3.738 ;
      RECT 56.3 3.326 56.305 3.78 ;
      RECT 56.295 3.324 56.3 3.808 ;
      RECT 56.29 3.322 56.295 3.83 ;
      RECT 56.28 3.318 56.29 3.873 ;
      RECT 56.275 3.315 56.28 3.898 ;
      RECT 56.27 3.313 56.275 3.918 ;
      RECT 56.265 3.311 56.27 3.942 ;
      RECT 56.26 3.307 56.265 3.965 ;
      RECT 56.255 3.303 56.26 3.988 ;
      RECT 56.22 3.293 56.255 4.095 ;
      RECT 56.215 3.283 56.22 4.193 ;
      RECT 56.21 3.281 56.215 4.22 ;
      RECT 56.205 3.28 56.21 4.24 ;
      RECT 56.2 3.272 56.205 4.26 ;
      RECT 56.195 3.267 56.2 4.295 ;
      RECT 56.19 3.265 56.195 4.313 ;
      RECT 56.185 3.265 56.19 4.338 ;
      RECT 56.18 3.265 56.185 4.36 ;
      RECT 56.145 3.265 56.18 4.403 ;
      RECT 56.12 3.265 56.145 4.432 ;
      RECT 56.11 3.265 56.12 3.618 ;
      RECT 56.113 3.675 56.12 4.442 ;
      RECT 56.11 3.732 56.113 4.445 ;
      RECT 56.105 3.265 56.11 3.59 ;
      RECT 56.105 3.782 56.11 4.448 ;
      RECT 56.095 3.265 56.105 3.58 ;
      RECT 56.1 3.835 56.105 4.451 ;
      RECT 56.095 3.92 56.1 4.455 ;
      RECT 56.085 3.265 56.095 3.568 ;
      RECT 56.09 3.967 56.095 4.459 ;
      RECT 56.085 4.042 56.09 4.463 ;
      RECT 56.05 3.265 56.085 3.543 ;
      RECT 56.075 4.125 56.085 4.468 ;
      RECT 56.065 4.192 56.075 4.475 ;
      RECT 56.06 4.22 56.065 4.48 ;
      RECT 56.05 4.233 56.06 4.486 ;
      RECT 56.005 3.265 56.05 3.5 ;
      RECT 56.045 4.238 56.05 4.493 ;
      RECT 56.005 4.255 56.045 4.555 ;
      RECT 56 3.267 56.005 3.473 ;
      RECT 55.975 4.275 56.005 4.555 ;
      RECT 55.995 3.272 56 3.445 ;
      RECT 55.785 4.284 55.825 4.555 ;
      RECT 55.76 4.292 55.785 4.525 ;
      RECT 55.715 4.3 55.76 4.525 ;
      RECT 55.7 4.305 55.715 4.52 ;
      RECT 55.69 4.305 55.7 4.514 ;
      RECT 55.68 4.312 55.69 4.511 ;
      RECT 55.675 4.35 55.68 4.5 ;
      RECT 55.67 4.412 55.675 4.478 ;
      RECT 56.94 4.287 57.125 4.51 ;
      RECT 56.94 4.302 57.13 4.506 ;
      RECT 56.93 3.575 57.015 4.505 ;
      RECT 56.93 4.302 57.135 4.499 ;
      RECT 56.925 4.31 57.135 4.498 ;
      RECT 57.13 4.03 57.45 4.35 ;
      RECT 56.925 4.202 57.095 4.293 ;
      RECT 56.92 4.202 57.095 4.275 ;
      RECT 56.91 4.01 57.045 4.25 ;
      RECT 56.905 4.01 57.045 4.195 ;
      RECT 56.865 3.59 57.035 4.095 ;
      RECT 56.85 3.59 57.035 3.965 ;
      RECT 56.845 3.59 57.035 3.918 ;
      RECT 56.84 3.59 57.035 3.898 ;
      RECT 56.835 3.59 57.035 3.873 ;
      RECT 56.805 3.59 57.065 3.85 ;
      RECT 56.815 3.587 57.025 3.85 ;
      RECT 56.94 3.582 57.025 4.51 ;
      RECT 56.825 3.575 57.015 3.85 ;
      RECT 56.82 3.58 57.015 3.85 ;
      RECT 55.65 3.792 55.835 4.005 ;
      RECT 55.65 3.8 55.845 3.998 ;
      RECT 55.63 3.8 55.845 3.995 ;
      RECT 55.625 3.8 55.845 3.98 ;
      RECT 55.555 3.715 55.815 3.975 ;
      RECT 55.555 3.86 55.85 3.888 ;
      RECT 55.21 4.315 55.47 4.575 ;
      RECT 55.235 4.26 55.43 4.575 ;
      RECT 55.23 4.009 55.41 4.303 ;
      RECT 55.23 4.015 55.42 4.303 ;
      RECT 55.21 4.017 55.42 4.248 ;
      RECT 55.205 4.027 55.42 4.115 ;
      RECT 55.235 4.007 55.41 4.575 ;
      RECT 55.321 4.005 55.41 4.575 ;
      RECT 55.18 3.225 55.215 3.595 ;
      RECT 54.97 3.335 54.975 3.595 ;
      RECT 55.215 3.232 55.23 3.595 ;
      RECT 55.105 3.225 55.18 3.673 ;
      RECT 55.095 3.225 55.105 3.758 ;
      RECT 55.07 3.225 55.095 3.793 ;
      RECT 55.03 3.225 55.07 3.861 ;
      RECT 55.02 3.232 55.03 3.913 ;
      RECT 54.99 3.335 55.02 3.954 ;
      RECT 54.985 3.335 54.99 3.993 ;
      RECT 54.975 3.335 54.985 4.013 ;
      RECT 54.97 3.63 54.975 4.05 ;
      RECT 54.965 3.647 54.97 4.07 ;
      RECT 54.95 3.71 54.965 4.11 ;
      RECT 54.945 3.753 54.95 4.145 ;
      RECT 54.94 3.761 54.945 4.158 ;
      RECT 54.93 3.775 54.94 4.18 ;
      RECT 54.905 3.81 54.93 4.245 ;
      RECT 54.895 3.845 54.905 4.308 ;
      RECT 54.875 3.875 54.895 4.369 ;
      RECT 54.86 3.911 54.875 4.436 ;
      RECT 54.85 3.939 54.86 4.475 ;
      RECT 54.84 3.961 54.85 4.495 ;
      RECT 54.835 3.971 54.84 4.506 ;
      RECT 54.83 3.98 54.835 4.509 ;
      RECT 54.82 3.998 54.83 4.513 ;
      RECT 54.81 4.016 54.82 4.514 ;
      RECT 54.785 4.055 54.81 4.511 ;
      RECT 54.765 4.097 54.785 4.508 ;
      RECT 54.75 4.135 54.765 4.507 ;
      RECT 54.715 4.17 54.75 4.504 ;
      RECT 54.71 4.192 54.715 4.502 ;
      RECT 54.645 4.232 54.71 4.499 ;
      RECT 54.64 4.272 54.645 4.495 ;
      RECT 54.625 4.282 54.64 4.486 ;
      RECT 54.615 4.402 54.625 4.471 ;
      RECT 55.095 4.815 55.105 5.075 ;
      RECT 55.095 4.818 55.115 5.074 ;
      RECT 55.085 4.808 55.095 5.073 ;
      RECT 55.075 4.823 55.155 5.069 ;
      RECT 55.06 4.802 55.075 5.067 ;
      RECT 55.035 4.827 55.16 5.063 ;
      RECT 55.02 4.787 55.035 5.058 ;
      RECT 55.02 4.829 55.17 5.057 ;
      RECT 55.02 4.837 55.185 5.05 ;
      RECT 54.96 4.774 55.02 5.04 ;
      RECT 54.95 4.761 54.96 5.022 ;
      RECT 54.925 4.751 54.95 5.012 ;
      RECT 54.92 4.741 54.925 5.004 ;
      RECT 54.855 4.837 55.185 4.986 ;
      RECT 54.77 4.837 55.185 4.948 ;
      RECT 54.66 4.665 54.92 4.925 ;
      RECT 55.035 4.795 55.06 5.063 ;
      RECT 55.075 4.805 55.085 5.069 ;
      RECT 54.66 4.813 55.1 4.925 ;
      RECT 54.845 10.055 55.135 10.285 ;
      RECT 54.905 9.315 55.075 10.285 ;
      RECT 54.805 9.345 55.175 9.715 ;
      RECT 54.845 9.315 55.135 9.715 ;
      RECT 53.875 4.57 53.905 4.87 ;
      RECT 53.65 4.555 53.655 4.83 ;
      RECT 53.45 4.555 53.605 4.815 ;
      RECT 54.75 3.27 54.78 3.53 ;
      RECT 54.74 3.27 54.75 3.638 ;
      RECT 54.72 3.27 54.74 3.648 ;
      RECT 54.705 3.27 54.72 3.66 ;
      RECT 54.65 3.27 54.705 3.71 ;
      RECT 54.635 3.27 54.65 3.758 ;
      RECT 54.605 3.27 54.635 3.793 ;
      RECT 54.55 3.27 54.605 3.855 ;
      RECT 54.53 3.27 54.55 3.923 ;
      RECT 54.525 3.27 54.53 3.953 ;
      RECT 54.52 3.27 54.525 3.965 ;
      RECT 54.515 3.387 54.52 3.983 ;
      RECT 54.495 3.405 54.515 4.008 ;
      RECT 54.475 3.432 54.495 4.058 ;
      RECT 54.47 3.452 54.475 4.089 ;
      RECT 54.465 3.46 54.47 4.106 ;
      RECT 54.45 3.486 54.465 4.135 ;
      RECT 54.435 3.528 54.45 4.17 ;
      RECT 54.43 3.557 54.435 4.193 ;
      RECT 54.425 3.572 54.43 4.206 ;
      RECT 54.42 3.595 54.425 4.217 ;
      RECT 54.41 3.615 54.42 4.235 ;
      RECT 54.4 3.645 54.41 4.258 ;
      RECT 54.395 3.667 54.4 4.278 ;
      RECT 54.39 3.682 54.395 4.293 ;
      RECT 54.375 3.712 54.39 4.32 ;
      RECT 54.37 3.742 54.375 4.346 ;
      RECT 54.365 3.76 54.37 4.358 ;
      RECT 54.355 3.79 54.365 4.377 ;
      RECT 54.345 3.815 54.355 4.402 ;
      RECT 54.34 3.835 54.345 4.421 ;
      RECT 54.335 3.852 54.34 4.434 ;
      RECT 54.325 3.878 54.335 4.453 ;
      RECT 54.315 3.916 54.325 4.48 ;
      RECT 54.31 3.942 54.315 4.5 ;
      RECT 54.305 3.952 54.31 4.51 ;
      RECT 54.3 3.965 54.305 4.525 ;
      RECT 54.295 3.98 54.3 4.535 ;
      RECT 54.29 4.002 54.295 4.55 ;
      RECT 54.285 4.02 54.29 4.561 ;
      RECT 54.28 4.03 54.285 4.572 ;
      RECT 54.275 4.038 54.28 4.584 ;
      RECT 54.27 4.046 54.275 4.595 ;
      RECT 54.265 4.072 54.27 4.608 ;
      RECT 54.255 4.1 54.265 4.621 ;
      RECT 54.25 4.13 54.255 4.63 ;
      RECT 54.245 4.145 54.25 4.637 ;
      RECT 54.23 4.17 54.245 4.644 ;
      RECT 54.225 4.192 54.23 4.65 ;
      RECT 54.22 4.217 54.225 4.653 ;
      RECT 54.211 4.245 54.22 4.657 ;
      RECT 54.205 4.262 54.211 4.662 ;
      RECT 54.2 4.28 54.205 4.666 ;
      RECT 54.195 4.292 54.2 4.669 ;
      RECT 54.19 4.313 54.195 4.673 ;
      RECT 54.185 4.331 54.19 4.676 ;
      RECT 54.18 4.345 54.185 4.679 ;
      RECT 54.175 4.362 54.18 4.682 ;
      RECT 54.17 4.375 54.175 4.685 ;
      RECT 54.145 4.412 54.17 4.693 ;
      RECT 54.14 4.457 54.145 4.702 ;
      RECT 54.135 4.485 54.14 4.705 ;
      RECT 54.125 4.505 54.135 4.709 ;
      RECT 54.12 4.525 54.125 4.714 ;
      RECT 54.115 4.54 54.12 4.717 ;
      RECT 54.095 4.55 54.115 4.724 ;
      RECT 54.03 4.557 54.095 4.75 ;
      RECT 53.995 4.56 54.03 4.778 ;
      RECT 53.98 4.563 53.995 4.793 ;
      RECT 53.97 4.564 53.98 4.808 ;
      RECT 53.96 4.565 53.97 4.825 ;
      RECT 53.955 4.565 53.96 4.84 ;
      RECT 53.95 4.565 53.955 4.848 ;
      RECT 53.935 4.566 53.95 4.863 ;
      RECT 53.905 4.568 53.935 4.87 ;
      RECT 53.795 4.575 53.875 4.87 ;
      RECT 53.75 4.58 53.795 4.87 ;
      RECT 53.74 4.581 53.75 4.86 ;
      RECT 53.73 4.582 53.74 4.853 ;
      RECT 53.71 4.584 53.73 4.848 ;
      RECT 53.7 4.555 53.71 4.843 ;
      RECT 53.655 4.555 53.7 4.835 ;
      RECT 53.625 4.555 53.65 4.825 ;
      RECT 53.605 4.555 53.625 4.818 ;
      RECT 53.885 3.355 54.145 3.615 ;
      RECT 53.765 3.37 53.775 3.535 ;
      RECT 53.75 3.37 53.755 3.53 ;
      RECT 51.115 3.21 51.3 3.5 ;
      RECT 52.93 3.335 52.945 3.49 ;
      RECT 51.08 3.21 51.105 3.47 ;
      RECT 53.495 3.26 53.5 3.402 ;
      RECT 53.41 3.255 53.435 3.395 ;
      RECT 53.81 3.372 53.885 3.565 ;
      RECT 53.795 3.37 53.81 3.548 ;
      RECT 53.775 3.37 53.795 3.54 ;
      RECT 53.755 3.37 53.765 3.533 ;
      RECT 53.71 3.365 53.75 3.523 ;
      RECT 53.67 3.34 53.71 3.508 ;
      RECT 53.655 3.315 53.67 3.498 ;
      RECT 53.65 3.309 53.655 3.496 ;
      RECT 53.615 3.301 53.65 3.479 ;
      RECT 53.61 3.294 53.615 3.467 ;
      RECT 53.59 3.289 53.61 3.455 ;
      RECT 53.58 3.283 53.59 3.44 ;
      RECT 53.56 3.278 53.58 3.425 ;
      RECT 53.55 3.273 53.56 3.418 ;
      RECT 53.545 3.271 53.55 3.413 ;
      RECT 53.54 3.27 53.545 3.41 ;
      RECT 53.5 3.265 53.54 3.406 ;
      RECT 53.48 3.259 53.495 3.401 ;
      RECT 53.445 3.256 53.48 3.398 ;
      RECT 53.435 3.255 53.445 3.396 ;
      RECT 53.375 3.255 53.41 3.393 ;
      RECT 53.33 3.255 53.375 3.393 ;
      RECT 53.28 3.255 53.33 3.396 ;
      RECT 53.265 3.257 53.28 3.398 ;
      RECT 53.25 3.26 53.265 3.399 ;
      RECT 53.24 3.265 53.25 3.4 ;
      RECT 53.21 3.27 53.24 3.405 ;
      RECT 53.2 3.276 53.21 3.413 ;
      RECT 53.19 3.278 53.2 3.417 ;
      RECT 53.18 3.282 53.19 3.421 ;
      RECT 53.155 3.288 53.18 3.429 ;
      RECT 53.145 3.293 53.155 3.437 ;
      RECT 53.13 3.297 53.145 3.441 ;
      RECT 53.095 3.303 53.13 3.449 ;
      RECT 53.075 3.308 53.095 3.459 ;
      RECT 53.045 3.315 53.075 3.468 ;
      RECT 53 3.324 53.045 3.482 ;
      RECT 52.995 3.329 53 3.493 ;
      RECT 52.975 3.332 52.995 3.494 ;
      RECT 52.945 3.335 52.975 3.492 ;
      RECT 52.91 3.335 52.93 3.488 ;
      RECT 52.84 3.335 52.91 3.479 ;
      RECT 52.825 3.332 52.84 3.471 ;
      RECT 52.785 3.325 52.825 3.466 ;
      RECT 52.76 3.315 52.785 3.459 ;
      RECT 52.755 3.309 52.76 3.456 ;
      RECT 52.715 3.303 52.755 3.453 ;
      RECT 52.7 3.296 52.715 3.448 ;
      RECT 52.68 3.292 52.7 3.443 ;
      RECT 52.665 3.287 52.68 3.439 ;
      RECT 52.65 3.282 52.665 3.437 ;
      RECT 52.635 3.278 52.65 3.436 ;
      RECT 52.62 3.276 52.635 3.432 ;
      RECT 52.61 3.274 52.62 3.427 ;
      RECT 52.595 3.271 52.61 3.423 ;
      RECT 52.585 3.269 52.595 3.418 ;
      RECT 52.565 3.266 52.585 3.414 ;
      RECT 52.52 3.265 52.565 3.412 ;
      RECT 52.46 3.267 52.52 3.413 ;
      RECT 52.44 3.269 52.46 3.415 ;
      RECT 52.41 3.272 52.44 3.416 ;
      RECT 52.36 3.277 52.41 3.418 ;
      RECT 52.355 3.28 52.36 3.42 ;
      RECT 52.345 3.282 52.355 3.423 ;
      RECT 52.34 3.284 52.345 3.426 ;
      RECT 52.29 3.287 52.34 3.433 ;
      RECT 52.27 3.291 52.29 3.445 ;
      RECT 52.26 3.294 52.27 3.451 ;
      RECT 52.25 3.295 52.26 3.454 ;
      RECT 52.211 3.298 52.25 3.456 ;
      RECT 52.125 3.305 52.211 3.459 ;
      RECT 52.051 3.315 52.125 3.463 ;
      RECT 51.965 3.326 52.051 3.468 ;
      RECT 51.95 3.333 51.965 3.47 ;
      RECT 51.895 3.337 51.95 3.471 ;
      RECT 51.881 3.34 51.895 3.473 ;
      RECT 51.795 3.34 51.881 3.475 ;
      RECT 51.755 3.337 51.795 3.478 ;
      RECT 51.731 3.333 51.755 3.48 ;
      RECT 51.645 3.323 51.731 3.483 ;
      RECT 51.615 3.312 51.645 3.484 ;
      RECT 51.596 3.308 51.615 3.483 ;
      RECT 51.51 3.301 51.596 3.48 ;
      RECT 51.45 3.29 51.51 3.477 ;
      RECT 51.43 3.282 51.45 3.475 ;
      RECT 51.395 3.277 51.43 3.474 ;
      RECT 51.37 3.272 51.395 3.473 ;
      RECT 51.34 3.267 51.37 3.472 ;
      RECT 51.315 3.21 51.34 3.471 ;
      RECT 51.3 3.21 51.315 3.495 ;
      RECT 51.105 3.21 51.115 3.495 ;
      RECT 52.88 4.23 52.885 4.37 ;
      RECT 52.54 4.23 52.575 4.368 ;
      RECT 52.115 4.215 52.13 4.36 ;
      RECT 53.945 3.995 54.035 4.255 ;
      RECT 53.775 3.86 53.875 4.255 ;
      RECT 50.81 3.835 50.89 4.045 ;
      RECT 53.9 3.972 53.945 4.255 ;
      RECT 53.89 3.942 53.9 4.255 ;
      RECT 53.875 3.865 53.89 4.255 ;
      RECT 53.69 3.86 53.775 4.22 ;
      RECT 53.685 3.862 53.69 4.215 ;
      RECT 53.68 3.867 53.685 4.215 ;
      RECT 53.645 3.967 53.68 4.215 ;
      RECT 53.635 3.995 53.645 4.215 ;
      RECT 53.625 4.01 53.635 4.215 ;
      RECT 53.615 4.022 53.625 4.215 ;
      RECT 53.61 4.032 53.615 4.215 ;
      RECT 53.595 4.042 53.61 4.217 ;
      RECT 53.59 4.057 53.595 4.219 ;
      RECT 53.575 4.07 53.59 4.221 ;
      RECT 53.57 4.085 53.575 4.224 ;
      RECT 53.55 4.095 53.57 4.228 ;
      RECT 53.535 4.105 53.55 4.231 ;
      RECT 53.5 4.112 53.535 4.236 ;
      RECT 53.456 4.119 53.5 4.244 ;
      RECT 53.37 4.131 53.456 4.257 ;
      RECT 53.345 4.142 53.37 4.268 ;
      RECT 53.315 4.147 53.345 4.273 ;
      RECT 53.28 4.152 53.315 4.281 ;
      RECT 53.25 4.157 53.28 4.288 ;
      RECT 53.225 4.162 53.25 4.293 ;
      RECT 53.16 4.169 53.225 4.302 ;
      RECT 53.09 4.182 53.16 4.318 ;
      RECT 53.06 4.192 53.09 4.33 ;
      RECT 53.035 4.197 53.06 4.337 ;
      RECT 52.98 4.204 53.035 4.345 ;
      RECT 52.975 4.211 52.98 4.35 ;
      RECT 52.97 4.213 52.975 4.351 ;
      RECT 52.955 4.215 52.97 4.353 ;
      RECT 52.95 4.215 52.955 4.356 ;
      RECT 52.885 4.222 52.95 4.363 ;
      RECT 52.85 4.232 52.88 4.373 ;
      RECT 52.833 4.235 52.85 4.375 ;
      RECT 52.747 4.234 52.833 4.374 ;
      RECT 52.661 4.232 52.747 4.371 ;
      RECT 52.575 4.231 52.661 4.369 ;
      RECT 52.474 4.229 52.54 4.368 ;
      RECT 52.388 4.226 52.474 4.366 ;
      RECT 52.302 4.222 52.388 4.364 ;
      RECT 52.216 4.219 52.302 4.363 ;
      RECT 52.13 4.216 52.216 4.361 ;
      RECT 52.03 4.215 52.115 4.358 ;
      RECT 51.98 4.213 52.03 4.356 ;
      RECT 51.96 4.21 51.98 4.354 ;
      RECT 51.94 4.208 51.96 4.351 ;
      RECT 51.915 4.204 51.94 4.348 ;
      RECT 51.87 4.198 51.915 4.343 ;
      RECT 51.83 4.192 51.87 4.335 ;
      RECT 51.805 4.187 51.83 4.328 ;
      RECT 51.75 4.18 51.805 4.32 ;
      RECT 51.726 4.173 51.75 4.313 ;
      RECT 51.64 4.164 51.726 4.303 ;
      RECT 51.61 4.156 51.64 4.293 ;
      RECT 51.58 4.152 51.61 4.288 ;
      RECT 51.575 4.149 51.58 4.285 ;
      RECT 51.57 4.148 51.575 4.285 ;
      RECT 51.495 4.141 51.57 4.278 ;
      RECT 51.456 4.132 51.495 4.267 ;
      RECT 51.37 4.122 51.456 4.255 ;
      RECT 51.33 4.112 51.37 4.243 ;
      RECT 51.291 4.107 51.33 4.236 ;
      RECT 51.205 4.097 51.291 4.225 ;
      RECT 51.165 4.085 51.205 4.214 ;
      RECT 51.13 4.07 51.165 4.207 ;
      RECT 51.12 4.06 51.13 4.204 ;
      RECT 51.1 4.045 51.12 4.202 ;
      RECT 51.07 4.015 51.1 4.198 ;
      RECT 51.06 3.995 51.07 4.193 ;
      RECT 51.055 3.987 51.06 4.19 ;
      RECT 51.05 3.98 51.055 4.188 ;
      RECT 51.035 3.967 51.05 4.181 ;
      RECT 51.03 3.957 51.035 4.173 ;
      RECT 51.025 3.95 51.03 4.168 ;
      RECT 51.02 3.945 51.025 4.164 ;
      RECT 51.005 3.932 51.02 4.156 ;
      RECT 51 3.842 51.005 4.145 ;
      RECT 50.995 3.837 51 4.138 ;
      RECT 50.92 3.835 50.995 4.098 ;
      RECT 50.89 3.835 50.92 4.053 ;
      RECT 50.795 3.84 50.81 4.04 ;
      RECT 53.28 3.545 53.54 3.805 ;
      RECT 53.265 3.533 53.445 3.77 ;
      RECT 53.26 3.534 53.445 3.768 ;
      RECT 53.245 3.538 53.455 3.758 ;
      RECT 53.24 3.543 53.46 3.728 ;
      RECT 53.245 3.54 53.46 3.758 ;
      RECT 53.26 3.535 53.455 3.768 ;
      RECT 53.28 3.532 53.445 3.805 ;
      RECT 53.28 3.531 53.435 3.805 ;
      RECT 53.305 3.53 53.435 3.805 ;
      RECT 52.865 3.775 53.125 4.035 ;
      RECT 52.74 3.82 53.125 4.03 ;
      RECT 52.73 3.825 53.125 4.025 ;
      RECT 52.745 4.765 52.76 5.075 ;
      RECT 51.34 4.535 51.35 4.665 ;
      RECT 51.12 4.53 51.225 4.665 ;
      RECT 51.035 4.535 51.085 4.665 ;
      RECT 49.585 3.27 49.59 4.375 ;
      RECT 52.84 4.857 52.845 4.993 ;
      RECT 52.835 4.852 52.84 5.053 ;
      RECT 52.83 4.85 52.835 5.066 ;
      RECT 52.815 4.847 52.83 5.068 ;
      RECT 52.81 4.842 52.815 5.07 ;
      RECT 52.805 4.838 52.81 5.073 ;
      RECT 52.79 4.833 52.805 5.075 ;
      RECT 52.76 4.825 52.79 5.075 ;
      RECT 52.721 4.765 52.745 5.075 ;
      RECT 52.635 4.765 52.721 5.072 ;
      RECT 52.605 4.765 52.635 5.065 ;
      RECT 52.58 4.765 52.605 5.058 ;
      RECT 52.555 4.765 52.58 5.05 ;
      RECT 52.54 4.765 52.555 5.043 ;
      RECT 52.515 4.765 52.54 5.035 ;
      RECT 52.5 4.765 52.515 5.028 ;
      RECT 52.46 4.775 52.5 5.017 ;
      RECT 52.45 4.77 52.46 5.007 ;
      RECT 52.446 4.769 52.45 5.004 ;
      RECT 52.36 4.761 52.446 4.987 ;
      RECT 52.327 4.75 52.36 4.964 ;
      RECT 52.241 4.739 52.327 4.942 ;
      RECT 52.155 4.723 52.241 4.911 ;
      RECT 52.085 4.708 52.155 4.883 ;
      RECT 52.075 4.701 52.085 4.87 ;
      RECT 52.045 4.698 52.075 4.86 ;
      RECT 52.02 4.694 52.045 4.853 ;
      RECT 52.005 4.691 52.02 4.848 ;
      RECT 52 4.69 52.005 4.843 ;
      RECT 51.97 4.685 52 4.836 ;
      RECT 51.965 4.68 51.97 4.831 ;
      RECT 51.95 4.677 51.965 4.826 ;
      RECT 51.945 4.672 51.95 4.821 ;
      RECT 51.925 4.667 51.945 4.818 ;
      RECT 51.91 4.662 51.925 4.81 ;
      RECT 51.895 4.656 51.91 4.805 ;
      RECT 51.865 4.647 51.895 4.798 ;
      RECT 51.86 4.64 51.865 4.79 ;
      RECT 51.855 4.638 51.86 4.788 ;
      RECT 51.85 4.637 51.855 4.785 ;
      RECT 51.81 4.63 51.85 4.778 ;
      RECT 51.796 4.62 51.81 4.768 ;
      RECT 51.745 4.609 51.796 4.756 ;
      RECT 51.72 4.595 51.745 4.742 ;
      RECT 51.695 4.584 51.72 4.734 ;
      RECT 51.675 4.573 51.695 4.728 ;
      RECT 51.665 4.567 51.675 4.723 ;
      RECT 51.66 4.565 51.665 4.719 ;
      RECT 51.64 4.56 51.66 4.714 ;
      RECT 51.61 4.55 51.64 4.704 ;
      RECT 51.605 4.542 51.61 4.697 ;
      RECT 51.59 4.54 51.605 4.693 ;
      RECT 51.57 4.54 51.59 4.688 ;
      RECT 51.565 4.539 51.57 4.686 ;
      RECT 51.56 4.539 51.565 4.683 ;
      RECT 51.52 4.538 51.56 4.678 ;
      RECT 51.495 4.537 51.52 4.673 ;
      RECT 51.435 4.536 51.495 4.67 ;
      RECT 51.35 4.535 51.435 4.668 ;
      RECT 51.311 4.534 51.34 4.665 ;
      RECT 51.225 4.532 51.311 4.665 ;
      RECT 51.085 4.532 51.12 4.665 ;
      RECT 50.995 4.536 51.035 4.668 ;
      RECT 50.98 4.539 50.995 4.675 ;
      RECT 50.97 4.54 50.98 4.682 ;
      RECT 50.945 4.543 50.97 4.687 ;
      RECT 50.94 4.545 50.945 4.69 ;
      RECT 50.89 4.547 50.94 4.691 ;
      RECT 50.851 4.551 50.89 4.693 ;
      RECT 50.765 4.553 50.851 4.696 ;
      RECT 50.747 4.555 50.765 4.698 ;
      RECT 50.661 4.558 50.747 4.7 ;
      RECT 50.575 4.562 50.661 4.703 ;
      RECT 50.538 4.566 50.575 4.706 ;
      RECT 50.452 4.569 50.538 4.709 ;
      RECT 50.366 4.573 50.452 4.712 ;
      RECT 50.28 4.578 50.366 4.716 ;
      RECT 50.26 4.58 50.28 4.719 ;
      RECT 50.24 4.579 50.26 4.72 ;
      RECT 50.191 4.576 50.24 4.721 ;
      RECT 50.105 4.571 50.191 4.724 ;
      RECT 50.055 4.566 50.105 4.726 ;
      RECT 50.031 4.564 50.055 4.727 ;
      RECT 49.945 4.559 50.031 4.729 ;
      RECT 49.92 4.555 49.945 4.728 ;
      RECT 49.91 4.552 49.92 4.726 ;
      RECT 49.9 4.545 49.91 4.723 ;
      RECT 49.895 4.525 49.9 4.718 ;
      RECT 49.885 4.495 49.895 4.713 ;
      RECT 49.87 4.365 49.885 4.704 ;
      RECT 49.865 4.357 49.87 4.697 ;
      RECT 49.845 4.35 49.865 4.689 ;
      RECT 49.84 4.332 49.845 4.681 ;
      RECT 49.83 4.312 49.84 4.676 ;
      RECT 49.825 4.285 49.83 4.672 ;
      RECT 49.82 4.262 49.825 4.669 ;
      RECT 49.8 4.22 49.82 4.661 ;
      RECT 49.765 4.135 49.8 4.645 ;
      RECT 49.76 4.067 49.765 4.633 ;
      RECT 49.745 4.037 49.76 4.627 ;
      RECT 49.74 3.282 49.745 3.528 ;
      RECT 49.73 4.007 49.745 4.618 ;
      RECT 49.735 3.277 49.74 3.56 ;
      RECT 49.73 3.272 49.735 3.603 ;
      RECT 49.725 3.27 49.73 3.638 ;
      RECT 49.71 3.97 49.73 4.608 ;
      RECT 49.72 3.27 49.725 3.675 ;
      RECT 49.705 3.27 49.72 3.773 ;
      RECT 49.705 3.943 49.71 4.601 ;
      RECT 49.7 3.27 49.705 3.848 ;
      RECT 49.7 3.931 49.705 4.598 ;
      RECT 49.695 3.27 49.7 3.88 ;
      RECT 49.695 3.91 49.7 4.595 ;
      RECT 49.69 3.27 49.695 4.592 ;
      RECT 49.655 3.27 49.69 4.578 ;
      RECT 49.64 3.27 49.655 4.56 ;
      RECT 49.62 3.27 49.64 4.55 ;
      RECT 49.595 3.27 49.62 4.533 ;
      RECT 49.59 3.27 49.595 4.483 ;
      RECT 49.58 3.27 49.585 4.313 ;
      RECT 49.575 3.27 49.58 4.22 ;
      RECT 49.57 3.27 49.575 4.133 ;
      RECT 49.565 3.27 49.57 4.065 ;
      RECT 49.56 3.27 49.565 4.008 ;
      RECT 49.55 3.27 49.56 3.903 ;
      RECT 49.545 3.27 49.55 3.775 ;
      RECT 49.54 3.27 49.545 3.693 ;
      RECT 49.535 3.272 49.54 3.61 ;
      RECT 49.53 3.277 49.535 3.543 ;
      RECT 49.525 3.282 49.53 3.47 ;
      RECT 52.34 3.6 52.6 3.86 ;
      RECT 52.36 3.567 52.57 3.86 ;
      RECT 52.36 3.565 52.56 3.86 ;
      RECT 52.37 3.552 52.56 3.86 ;
      RECT 52.37 3.55 52.485 3.86 ;
      RECT 51.845 3.675 52.02 3.955 ;
      RECT 51.84 3.675 52.02 3.953 ;
      RECT 51.84 3.675 52.035 3.95 ;
      RECT 51.83 3.675 52.035 3.948 ;
      RECT 51.775 3.675 52.035 3.935 ;
      RECT 51.775 3.75 52.04 3.913 ;
      RECT 51.32 3.687 51.34 3.93 ;
      RECT 51.32 3.687 51.38 3.929 ;
      RECT 51.315 3.689 51.38 3.928 ;
      RECT 51.315 3.689 51.466 3.927 ;
      RECT 51.315 3.689 51.535 3.926 ;
      RECT 51.315 3.689 51.555 3.918 ;
      RECT 51.295 3.692 51.555 3.916 ;
      RECT 51.28 3.702 51.555 3.901 ;
      RECT 51.28 3.702 51.57 3.9 ;
      RECT 51.275 3.711 51.57 3.892 ;
      RECT 51.275 3.711 51.575 3.888 ;
      RECT 51.38 3.625 51.64 3.885 ;
      RECT 51.27 3.713 51.64 3.77 ;
      RECT 51.34 3.68 51.64 3.885 ;
      RECT 51.305 4.873 51.31 5.08 ;
      RECT 51.255 4.867 51.305 5.079 ;
      RECT 51.222 4.881 51.315 5.078 ;
      RECT 51.136 4.881 51.315 5.077 ;
      RECT 51.05 4.881 51.315 5.076 ;
      RECT 51.05 4.98 51.32 5.073 ;
      RECT 51.045 4.98 51.32 5.068 ;
      RECT 51.04 4.98 51.32 5.05 ;
      RECT 51.035 4.98 51.32 5.033 ;
      RECT 50.995 4.765 51.255 5.025 ;
      RECT 50.455 3.915 50.541 4.329 ;
      RECT 50.455 3.915 50.58 4.326 ;
      RECT 50.455 3.915 50.6 4.316 ;
      RECT 50.41 3.915 50.6 4.313 ;
      RECT 50.41 4.067 50.61 4.303 ;
      RECT 50.41 4.088 50.615 4.297 ;
      RECT 50.41 4.106 50.62 4.293 ;
      RECT 50.41 4.126 50.63 4.288 ;
      RECT 50.385 4.126 50.63 4.285 ;
      RECT 50.375 4.126 50.63 4.263 ;
      RECT 50.375 4.142 50.635 4.233 ;
      RECT 50.34 3.915 50.6 4.22 ;
      RECT 50.34 4.154 50.64 4.175 ;
      RECT 48 10.06 48.29 10.29 ;
      RECT 48.06 8.58 48.23 10.29 ;
      RECT 48.01 8.945 48.36 9.295 ;
      RECT 48 8.58 48.29 8.81 ;
      RECT 47.595 3.69 47.7 4.26 ;
      RECT 47.595 4.025 47.92 4.255 ;
      RECT 47.595 4.055 48.09 4.225 ;
      RECT 47.595 3.69 47.785 4.255 ;
      RECT 47.01 3.655 47.3 3.885 ;
      RECT 47.01 3.69 47.785 3.86 ;
      RECT 47.07 2.175 47.24 3.885 ;
      RECT 47.01 2.175 47.3 2.405 ;
      RECT 47.01 10.06 47.3 10.29 ;
      RECT 47.07 8.58 47.24 10.29 ;
      RECT 47.01 8.58 47.3 8.81 ;
      RECT 47.01 8.615 47.86 8.775 ;
      RECT 47.695 8.21 47.86 8.775 ;
      RECT 47.01 8.61 47.405 8.775 ;
      RECT 47.63 8.21 47.92 8.44 ;
      RECT 47.63 8.24 48.09 8.41 ;
      RECT 46.64 4.025 46.93 4.255 ;
      RECT 46.64 4.055 47.1 4.225 ;
      RECT 46.705 2.95 46.87 4.255 ;
      RECT 45.22 2.92 45.51 3.15 ;
      RECT 45.22 2.95 46.87 3.12 ;
      RECT 45.28 2.18 45.45 3.15 ;
      RECT 45.22 2.18 45.51 2.41 ;
      RECT 45.22 10.055 45.51 10.285 ;
      RECT 45.28 9.315 45.45 10.285 ;
      RECT 45.28 9.41 46.87 9.58 ;
      RECT 46.7 8.21 46.87 9.58 ;
      RECT 45.22 9.315 45.51 9.545 ;
      RECT 46.64 8.21 46.93 8.44 ;
      RECT 46.64 8.24 47.1 8.41 ;
      RECT 43.27 4 43.61 4.35 ;
      RECT 43.36 3.32 43.53 4.35 ;
      RECT 45.65 3.26 46 3.61 ;
      RECT 43.36 3.32 46 3.49 ;
      RECT 45.675 8.945 46 9.27 ;
      RECT 40.215 8.905 40.565 9.255 ;
      RECT 45.65 8.945 46 9.175 ;
      RECT 40.015 8.945 40.565 9.175 ;
      RECT 39.845 8.975 46 9.145 ;
      RECT 44.875 3.66 45.195 3.98 ;
      RECT 44.845 3.66 45.195 3.89 ;
      RECT 44.675 3.69 45.195 3.86 ;
      RECT 44.875 8.545 45.195 8.835 ;
      RECT 44.845 8.575 45.195 8.805 ;
      RECT 44.675 8.605 45.195 8.775 ;
      RECT 40.565 4.28 40.715 4.555 ;
      RECT 41.105 3.36 41.11 3.58 ;
      RECT 42.255 3.56 42.27 3.758 ;
      RECT 42.22 3.552 42.255 3.765 ;
      RECT 42.19 3.545 42.22 3.765 ;
      RECT 42.135 3.51 42.19 3.765 ;
      RECT 42.07 3.447 42.135 3.765 ;
      RECT 42.065 3.412 42.07 3.763 ;
      RECT 42.06 3.407 42.065 3.755 ;
      RECT 42.055 3.402 42.06 3.741 ;
      RECT 42.05 3.399 42.055 3.734 ;
      RECT 42.005 3.389 42.05 3.685 ;
      RECT 41.985 3.376 42.005 3.62 ;
      RECT 41.98 3.371 41.985 3.593 ;
      RECT 41.975 3.37 41.98 3.586 ;
      RECT 41.97 3.369 41.975 3.579 ;
      RECT 41.885 3.354 41.97 3.525 ;
      RECT 41.855 3.335 41.885 3.475 ;
      RECT 41.775 3.318 41.855 3.46 ;
      RECT 41.74 3.305 41.775 3.445 ;
      RECT 41.732 3.305 41.74 3.44 ;
      RECT 41.646 3.306 41.732 3.44 ;
      RECT 41.56 3.308 41.646 3.44 ;
      RECT 41.535 3.309 41.56 3.444 ;
      RECT 41.46 3.315 41.535 3.459 ;
      RECT 41.377 3.327 41.46 3.483 ;
      RECT 41.291 3.34 41.377 3.509 ;
      RECT 41.205 3.353 41.291 3.535 ;
      RECT 41.17 3.362 41.205 3.554 ;
      RECT 41.12 3.362 41.17 3.567 ;
      RECT 41.11 3.36 41.12 3.578 ;
      RECT 41.095 3.357 41.105 3.58 ;
      RECT 41.08 3.349 41.095 3.588 ;
      RECT 41.065 3.341 41.08 3.608 ;
      RECT 41.06 3.336 41.065 3.665 ;
      RECT 41.045 3.331 41.06 3.738 ;
      RECT 41.04 3.326 41.045 3.78 ;
      RECT 41.035 3.324 41.04 3.808 ;
      RECT 41.03 3.322 41.035 3.83 ;
      RECT 41.02 3.318 41.03 3.873 ;
      RECT 41.015 3.315 41.02 3.898 ;
      RECT 41.01 3.313 41.015 3.918 ;
      RECT 41.005 3.311 41.01 3.942 ;
      RECT 41 3.307 41.005 3.965 ;
      RECT 40.995 3.303 41 3.988 ;
      RECT 40.96 3.293 40.995 4.095 ;
      RECT 40.955 3.283 40.96 4.193 ;
      RECT 40.95 3.281 40.955 4.22 ;
      RECT 40.945 3.28 40.95 4.24 ;
      RECT 40.94 3.272 40.945 4.26 ;
      RECT 40.935 3.267 40.94 4.295 ;
      RECT 40.93 3.265 40.935 4.313 ;
      RECT 40.925 3.265 40.93 4.338 ;
      RECT 40.92 3.265 40.925 4.36 ;
      RECT 40.885 3.265 40.92 4.403 ;
      RECT 40.86 3.265 40.885 4.432 ;
      RECT 40.85 3.265 40.86 3.618 ;
      RECT 40.853 3.675 40.86 4.442 ;
      RECT 40.85 3.732 40.853 4.445 ;
      RECT 40.845 3.265 40.85 3.59 ;
      RECT 40.845 3.782 40.85 4.448 ;
      RECT 40.835 3.265 40.845 3.58 ;
      RECT 40.84 3.835 40.845 4.451 ;
      RECT 40.835 3.92 40.84 4.455 ;
      RECT 40.825 3.265 40.835 3.568 ;
      RECT 40.83 3.967 40.835 4.459 ;
      RECT 40.825 4.042 40.83 4.463 ;
      RECT 40.79 3.265 40.825 3.543 ;
      RECT 40.815 4.125 40.825 4.468 ;
      RECT 40.805 4.192 40.815 4.475 ;
      RECT 40.8 4.22 40.805 4.48 ;
      RECT 40.79 4.233 40.8 4.486 ;
      RECT 40.745 3.265 40.79 3.5 ;
      RECT 40.785 4.238 40.79 4.493 ;
      RECT 40.745 4.255 40.785 4.555 ;
      RECT 40.74 3.267 40.745 3.473 ;
      RECT 40.715 4.275 40.745 4.555 ;
      RECT 40.735 3.272 40.74 3.445 ;
      RECT 40.525 4.284 40.565 4.555 ;
      RECT 40.5 4.292 40.525 4.525 ;
      RECT 40.455 4.3 40.5 4.525 ;
      RECT 40.44 4.305 40.455 4.52 ;
      RECT 40.43 4.305 40.44 4.514 ;
      RECT 40.42 4.312 40.43 4.511 ;
      RECT 40.415 4.35 40.42 4.5 ;
      RECT 40.41 4.412 40.415 4.478 ;
      RECT 41.68 4.287 41.865 4.51 ;
      RECT 41.68 4.302 41.87 4.506 ;
      RECT 41.67 3.575 41.755 4.505 ;
      RECT 41.67 4.302 41.875 4.499 ;
      RECT 41.665 4.31 41.875 4.498 ;
      RECT 41.87 4.03 42.19 4.35 ;
      RECT 41.665 4.202 41.835 4.293 ;
      RECT 41.66 4.202 41.835 4.275 ;
      RECT 41.65 4.01 41.785 4.25 ;
      RECT 41.645 4.01 41.785 4.195 ;
      RECT 41.605 3.59 41.775 4.095 ;
      RECT 41.59 3.59 41.775 3.965 ;
      RECT 41.585 3.59 41.775 3.918 ;
      RECT 41.58 3.59 41.775 3.898 ;
      RECT 41.575 3.59 41.775 3.873 ;
      RECT 41.545 3.59 41.805 3.85 ;
      RECT 41.555 3.587 41.765 3.85 ;
      RECT 41.68 3.582 41.765 4.51 ;
      RECT 41.565 3.575 41.755 3.85 ;
      RECT 41.56 3.58 41.755 3.85 ;
      RECT 40.39 3.792 40.575 4.005 ;
      RECT 40.39 3.8 40.585 3.998 ;
      RECT 40.37 3.8 40.585 3.995 ;
      RECT 40.365 3.8 40.585 3.98 ;
      RECT 40.295 3.715 40.555 3.975 ;
      RECT 40.295 3.86 40.59 3.888 ;
      RECT 39.95 4.315 40.21 4.575 ;
      RECT 39.975 4.26 40.17 4.575 ;
      RECT 39.97 4.009 40.15 4.303 ;
      RECT 39.97 4.015 40.16 4.303 ;
      RECT 39.95 4.017 40.16 4.248 ;
      RECT 39.945 4.027 40.16 4.115 ;
      RECT 39.975 4.007 40.15 4.575 ;
      RECT 40.061 4.005 40.15 4.575 ;
      RECT 39.92 3.225 39.955 3.595 ;
      RECT 39.71 3.335 39.715 3.595 ;
      RECT 39.955 3.232 39.97 3.595 ;
      RECT 39.845 3.225 39.92 3.673 ;
      RECT 39.835 3.225 39.845 3.758 ;
      RECT 39.81 3.225 39.835 3.793 ;
      RECT 39.77 3.225 39.81 3.861 ;
      RECT 39.76 3.232 39.77 3.913 ;
      RECT 39.73 3.335 39.76 3.954 ;
      RECT 39.725 3.335 39.73 3.993 ;
      RECT 39.715 3.335 39.725 4.013 ;
      RECT 39.71 3.63 39.715 4.05 ;
      RECT 39.705 3.647 39.71 4.07 ;
      RECT 39.69 3.71 39.705 4.11 ;
      RECT 39.685 3.753 39.69 4.145 ;
      RECT 39.68 3.761 39.685 4.158 ;
      RECT 39.67 3.775 39.68 4.18 ;
      RECT 39.645 3.81 39.67 4.245 ;
      RECT 39.635 3.845 39.645 4.308 ;
      RECT 39.615 3.875 39.635 4.369 ;
      RECT 39.6 3.911 39.615 4.436 ;
      RECT 39.59 3.939 39.6 4.475 ;
      RECT 39.58 3.961 39.59 4.495 ;
      RECT 39.575 3.971 39.58 4.506 ;
      RECT 39.57 3.98 39.575 4.509 ;
      RECT 39.56 3.998 39.57 4.513 ;
      RECT 39.55 4.016 39.56 4.514 ;
      RECT 39.525 4.055 39.55 4.511 ;
      RECT 39.505 4.097 39.525 4.508 ;
      RECT 39.49 4.135 39.505 4.507 ;
      RECT 39.455 4.17 39.49 4.504 ;
      RECT 39.45 4.192 39.455 4.502 ;
      RECT 39.385 4.232 39.45 4.499 ;
      RECT 39.38 4.272 39.385 4.495 ;
      RECT 39.365 4.282 39.38 4.486 ;
      RECT 39.355 4.402 39.365 4.471 ;
      RECT 39.835 4.815 39.845 5.075 ;
      RECT 39.835 4.818 39.855 5.074 ;
      RECT 39.825 4.808 39.835 5.073 ;
      RECT 39.815 4.823 39.895 5.069 ;
      RECT 39.8 4.802 39.815 5.067 ;
      RECT 39.775 4.827 39.9 5.063 ;
      RECT 39.76 4.787 39.775 5.058 ;
      RECT 39.76 4.829 39.91 5.057 ;
      RECT 39.76 4.837 39.925 5.05 ;
      RECT 39.7 4.774 39.76 5.04 ;
      RECT 39.69 4.761 39.7 5.022 ;
      RECT 39.665 4.751 39.69 5.012 ;
      RECT 39.66 4.741 39.665 5.004 ;
      RECT 39.595 4.837 39.925 4.986 ;
      RECT 39.51 4.837 39.925 4.948 ;
      RECT 39.4 4.665 39.66 4.925 ;
      RECT 39.775 4.795 39.8 5.063 ;
      RECT 39.815 4.805 39.825 5.069 ;
      RECT 39.4 4.813 39.84 4.925 ;
      RECT 39.585 10.055 39.875 10.285 ;
      RECT 39.645 9.315 39.815 10.285 ;
      RECT 39.545 9.345 39.915 9.715 ;
      RECT 39.585 9.315 39.875 9.715 ;
      RECT 38.615 4.57 38.645 4.87 ;
      RECT 38.39 4.555 38.395 4.83 ;
      RECT 38.19 4.555 38.345 4.815 ;
      RECT 39.49 3.27 39.52 3.53 ;
      RECT 39.48 3.27 39.49 3.638 ;
      RECT 39.46 3.27 39.48 3.648 ;
      RECT 39.445 3.27 39.46 3.66 ;
      RECT 39.39 3.27 39.445 3.71 ;
      RECT 39.375 3.27 39.39 3.758 ;
      RECT 39.345 3.27 39.375 3.793 ;
      RECT 39.29 3.27 39.345 3.855 ;
      RECT 39.27 3.27 39.29 3.923 ;
      RECT 39.265 3.27 39.27 3.953 ;
      RECT 39.26 3.27 39.265 3.965 ;
      RECT 39.255 3.387 39.26 3.983 ;
      RECT 39.235 3.405 39.255 4.008 ;
      RECT 39.215 3.432 39.235 4.058 ;
      RECT 39.21 3.452 39.215 4.089 ;
      RECT 39.205 3.46 39.21 4.106 ;
      RECT 39.19 3.486 39.205 4.135 ;
      RECT 39.175 3.528 39.19 4.17 ;
      RECT 39.17 3.557 39.175 4.193 ;
      RECT 39.165 3.572 39.17 4.206 ;
      RECT 39.16 3.595 39.165 4.217 ;
      RECT 39.15 3.615 39.16 4.235 ;
      RECT 39.14 3.645 39.15 4.258 ;
      RECT 39.135 3.667 39.14 4.278 ;
      RECT 39.13 3.682 39.135 4.293 ;
      RECT 39.115 3.712 39.13 4.32 ;
      RECT 39.11 3.742 39.115 4.346 ;
      RECT 39.105 3.76 39.11 4.358 ;
      RECT 39.095 3.79 39.105 4.377 ;
      RECT 39.085 3.815 39.095 4.402 ;
      RECT 39.08 3.835 39.085 4.421 ;
      RECT 39.075 3.852 39.08 4.434 ;
      RECT 39.065 3.878 39.075 4.453 ;
      RECT 39.055 3.916 39.065 4.48 ;
      RECT 39.05 3.942 39.055 4.5 ;
      RECT 39.045 3.952 39.05 4.51 ;
      RECT 39.04 3.965 39.045 4.525 ;
      RECT 39.035 3.98 39.04 4.535 ;
      RECT 39.03 4.002 39.035 4.55 ;
      RECT 39.025 4.02 39.03 4.561 ;
      RECT 39.02 4.03 39.025 4.572 ;
      RECT 39.015 4.038 39.02 4.584 ;
      RECT 39.01 4.046 39.015 4.595 ;
      RECT 39.005 4.072 39.01 4.608 ;
      RECT 38.995 4.1 39.005 4.621 ;
      RECT 38.99 4.13 38.995 4.63 ;
      RECT 38.985 4.145 38.99 4.637 ;
      RECT 38.97 4.17 38.985 4.644 ;
      RECT 38.965 4.192 38.97 4.65 ;
      RECT 38.96 4.217 38.965 4.653 ;
      RECT 38.951 4.245 38.96 4.657 ;
      RECT 38.945 4.262 38.951 4.662 ;
      RECT 38.94 4.28 38.945 4.666 ;
      RECT 38.935 4.292 38.94 4.669 ;
      RECT 38.93 4.313 38.935 4.673 ;
      RECT 38.925 4.331 38.93 4.676 ;
      RECT 38.92 4.345 38.925 4.679 ;
      RECT 38.915 4.362 38.92 4.682 ;
      RECT 38.91 4.375 38.915 4.685 ;
      RECT 38.885 4.412 38.91 4.693 ;
      RECT 38.88 4.457 38.885 4.702 ;
      RECT 38.875 4.485 38.88 4.705 ;
      RECT 38.865 4.505 38.875 4.709 ;
      RECT 38.86 4.525 38.865 4.714 ;
      RECT 38.855 4.54 38.86 4.717 ;
      RECT 38.835 4.55 38.855 4.724 ;
      RECT 38.77 4.557 38.835 4.75 ;
      RECT 38.735 4.56 38.77 4.778 ;
      RECT 38.72 4.563 38.735 4.793 ;
      RECT 38.71 4.564 38.72 4.808 ;
      RECT 38.7 4.565 38.71 4.825 ;
      RECT 38.695 4.565 38.7 4.84 ;
      RECT 38.69 4.565 38.695 4.848 ;
      RECT 38.675 4.566 38.69 4.863 ;
      RECT 38.645 4.568 38.675 4.87 ;
      RECT 38.535 4.575 38.615 4.87 ;
      RECT 38.49 4.58 38.535 4.87 ;
      RECT 38.48 4.581 38.49 4.86 ;
      RECT 38.47 4.582 38.48 4.853 ;
      RECT 38.45 4.584 38.47 4.848 ;
      RECT 38.44 4.555 38.45 4.843 ;
      RECT 38.395 4.555 38.44 4.835 ;
      RECT 38.365 4.555 38.39 4.825 ;
      RECT 38.345 4.555 38.365 4.818 ;
      RECT 38.625 3.355 38.885 3.615 ;
      RECT 38.505 3.37 38.515 3.535 ;
      RECT 38.49 3.37 38.495 3.53 ;
      RECT 35.855 3.21 36.04 3.5 ;
      RECT 37.67 3.335 37.685 3.49 ;
      RECT 35.82 3.21 35.845 3.47 ;
      RECT 38.235 3.26 38.24 3.402 ;
      RECT 38.15 3.255 38.175 3.395 ;
      RECT 38.55 3.372 38.625 3.565 ;
      RECT 38.535 3.37 38.55 3.548 ;
      RECT 38.515 3.37 38.535 3.54 ;
      RECT 38.495 3.37 38.505 3.533 ;
      RECT 38.45 3.365 38.49 3.523 ;
      RECT 38.41 3.34 38.45 3.508 ;
      RECT 38.395 3.315 38.41 3.498 ;
      RECT 38.39 3.309 38.395 3.496 ;
      RECT 38.355 3.301 38.39 3.479 ;
      RECT 38.35 3.294 38.355 3.467 ;
      RECT 38.33 3.289 38.35 3.455 ;
      RECT 38.32 3.283 38.33 3.44 ;
      RECT 38.3 3.278 38.32 3.425 ;
      RECT 38.29 3.273 38.3 3.418 ;
      RECT 38.285 3.271 38.29 3.413 ;
      RECT 38.28 3.27 38.285 3.41 ;
      RECT 38.24 3.265 38.28 3.406 ;
      RECT 38.22 3.259 38.235 3.401 ;
      RECT 38.185 3.256 38.22 3.398 ;
      RECT 38.175 3.255 38.185 3.396 ;
      RECT 38.115 3.255 38.15 3.393 ;
      RECT 38.07 3.255 38.115 3.393 ;
      RECT 38.02 3.255 38.07 3.396 ;
      RECT 38.005 3.257 38.02 3.398 ;
      RECT 37.99 3.26 38.005 3.399 ;
      RECT 37.98 3.265 37.99 3.4 ;
      RECT 37.95 3.27 37.98 3.405 ;
      RECT 37.94 3.276 37.95 3.413 ;
      RECT 37.93 3.278 37.94 3.417 ;
      RECT 37.92 3.282 37.93 3.421 ;
      RECT 37.895 3.288 37.92 3.429 ;
      RECT 37.885 3.293 37.895 3.437 ;
      RECT 37.87 3.297 37.885 3.441 ;
      RECT 37.835 3.303 37.87 3.449 ;
      RECT 37.815 3.308 37.835 3.459 ;
      RECT 37.785 3.315 37.815 3.468 ;
      RECT 37.74 3.324 37.785 3.482 ;
      RECT 37.735 3.329 37.74 3.493 ;
      RECT 37.715 3.332 37.735 3.494 ;
      RECT 37.685 3.335 37.715 3.492 ;
      RECT 37.65 3.335 37.67 3.488 ;
      RECT 37.58 3.335 37.65 3.479 ;
      RECT 37.565 3.332 37.58 3.471 ;
      RECT 37.525 3.325 37.565 3.466 ;
      RECT 37.5 3.315 37.525 3.459 ;
      RECT 37.495 3.309 37.5 3.456 ;
      RECT 37.455 3.303 37.495 3.453 ;
      RECT 37.44 3.296 37.455 3.448 ;
      RECT 37.42 3.292 37.44 3.443 ;
      RECT 37.405 3.287 37.42 3.439 ;
      RECT 37.39 3.282 37.405 3.437 ;
      RECT 37.375 3.278 37.39 3.436 ;
      RECT 37.36 3.276 37.375 3.432 ;
      RECT 37.35 3.274 37.36 3.427 ;
      RECT 37.335 3.271 37.35 3.423 ;
      RECT 37.325 3.269 37.335 3.418 ;
      RECT 37.305 3.266 37.325 3.414 ;
      RECT 37.26 3.265 37.305 3.412 ;
      RECT 37.2 3.267 37.26 3.413 ;
      RECT 37.18 3.269 37.2 3.415 ;
      RECT 37.15 3.272 37.18 3.416 ;
      RECT 37.1 3.277 37.15 3.418 ;
      RECT 37.095 3.28 37.1 3.42 ;
      RECT 37.085 3.282 37.095 3.423 ;
      RECT 37.08 3.284 37.085 3.426 ;
      RECT 37.03 3.287 37.08 3.433 ;
      RECT 37.01 3.291 37.03 3.445 ;
      RECT 37 3.294 37.01 3.451 ;
      RECT 36.99 3.295 37 3.454 ;
      RECT 36.951 3.298 36.99 3.456 ;
      RECT 36.865 3.305 36.951 3.459 ;
      RECT 36.791 3.315 36.865 3.463 ;
      RECT 36.705 3.326 36.791 3.468 ;
      RECT 36.69 3.333 36.705 3.47 ;
      RECT 36.635 3.337 36.69 3.471 ;
      RECT 36.621 3.34 36.635 3.473 ;
      RECT 36.535 3.34 36.621 3.475 ;
      RECT 36.495 3.337 36.535 3.478 ;
      RECT 36.471 3.333 36.495 3.48 ;
      RECT 36.385 3.323 36.471 3.483 ;
      RECT 36.355 3.312 36.385 3.484 ;
      RECT 36.336 3.308 36.355 3.483 ;
      RECT 36.25 3.301 36.336 3.48 ;
      RECT 36.19 3.29 36.25 3.477 ;
      RECT 36.17 3.282 36.19 3.475 ;
      RECT 36.135 3.277 36.17 3.474 ;
      RECT 36.11 3.272 36.135 3.473 ;
      RECT 36.08 3.267 36.11 3.472 ;
      RECT 36.055 3.21 36.08 3.471 ;
      RECT 36.04 3.21 36.055 3.495 ;
      RECT 35.845 3.21 35.855 3.495 ;
      RECT 37.62 4.23 37.625 4.37 ;
      RECT 37.28 4.23 37.315 4.368 ;
      RECT 36.855 4.215 36.87 4.36 ;
      RECT 38.685 3.995 38.775 4.255 ;
      RECT 38.515 3.86 38.615 4.255 ;
      RECT 35.55 3.835 35.63 4.045 ;
      RECT 38.64 3.972 38.685 4.255 ;
      RECT 38.63 3.942 38.64 4.255 ;
      RECT 38.615 3.865 38.63 4.255 ;
      RECT 38.43 3.86 38.515 4.22 ;
      RECT 38.425 3.862 38.43 4.215 ;
      RECT 38.42 3.867 38.425 4.215 ;
      RECT 38.385 3.967 38.42 4.215 ;
      RECT 38.375 3.995 38.385 4.215 ;
      RECT 38.365 4.01 38.375 4.215 ;
      RECT 38.355 4.022 38.365 4.215 ;
      RECT 38.35 4.032 38.355 4.215 ;
      RECT 38.335 4.042 38.35 4.217 ;
      RECT 38.33 4.057 38.335 4.219 ;
      RECT 38.315 4.07 38.33 4.221 ;
      RECT 38.31 4.085 38.315 4.224 ;
      RECT 38.29 4.095 38.31 4.228 ;
      RECT 38.275 4.105 38.29 4.231 ;
      RECT 38.24 4.112 38.275 4.236 ;
      RECT 38.196 4.119 38.24 4.244 ;
      RECT 38.11 4.131 38.196 4.257 ;
      RECT 38.085 4.142 38.11 4.268 ;
      RECT 38.055 4.147 38.085 4.273 ;
      RECT 38.02 4.152 38.055 4.281 ;
      RECT 37.99 4.157 38.02 4.288 ;
      RECT 37.965 4.162 37.99 4.293 ;
      RECT 37.9 4.169 37.965 4.302 ;
      RECT 37.83 4.182 37.9 4.318 ;
      RECT 37.8 4.192 37.83 4.33 ;
      RECT 37.775 4.197 37.8 4.337 ;
      RECT 37.72 4.204 37.775 4.345 ;
      RECT 37.715 4.211 37.72 4.35 ;
      RECT 37.71 4.213 37.715 4.351 ;
      RECT 37.695 4.215 37.71 4.353 ;
      RECT 37.69 4.215 37.695 4.356 ;
      RECT 37.625 4.222 37.69 4.363 ;
      RECT 37.59 4.232 37.62 4.373 ;
      RECT 37.573 4.235 37.59 4.375 ;
      RECT 37.487 4.234 37.573 4.374 ;
      RECT 37.401 4.232 37.487 4.371 ;
      RECT 37.315 4.231 37.401 4.369 ;
      RECT 37.214 4.229 37.28 4.368 ;
      RECT 37.128 4.226 37.214 4.366 ;
      RECT 37.042 4.222 37.128 4.364 ;
      RECT 36.956 4.219 37.042 4.363 ;
      RECT 36.87 4.216 36.956 4.361 ;
      RECT 36.77 4.215 36.855 4.358 ;
      RECT 36.72 4.213 36.77 4.356 ;
      RECT 36.7 4.21 36.72 4.354 ;
      RECT 36.68 4.208 36.7 4.351 ;
      RECT 36.655 4.204 36.68 4.348 ;
      RECT 36.61 4.198 36.655 4.343 ;
      RECT 36.57 4.192 36.61 4.335 ;
      RECT 36.545 4.187 36.57 4.328 ;
      RECT 36.49 4.18 36.545 4.32 ;
      RECT 36.466 4.173 36.49 4.313 ;
      RECT 36.38 4.164 36.466 4.303 ;
      RECT 36.35 4.156 36.38 4.293 ;
      RECT 36.32 4.152 36.35 4.288 ;
      RECT 36.315 4.149 36.32 4.285 ;
      RECT 36.31 4.148 36.315 4.285 ;
      RECT 36.235 4.141 36.31 4.278 ;
      RECT 36.196 4.132 36.235 4.267 ;
      RECT 36.11 4.122 36.196 4.255 ;
      RECT 36.07 4.112 36.11 4.243 ;
      RECT 36.031 4.107 36.07 4.236 ;
      RECT 35.945 4.097 36.031 4.225 ;
      RECT 35.905 4.085 35.945 4.214 ;
      RECT 35.87 4.07 35.905 4.207 ;
      RECT 35.86 4.06 35.87 4.204 ;
      RECT 35.84 4.045 35.86 4.202 ;
      RECT 35.81 4.015 35.84 4.198 ;
      RECT 35.8 3.995 35.81 4.193 ;
      RECT 35.795 3.987 35.8 4.19 ;
      RECT 35.79 3.98 35.795 4.188 ;
      RECT 35.775 3.967 35.79 4.181 ;
      RECT 35.77 3.957 35.775 4.173 ;
      RECT 35.765 3.95 35.77 4.168 ;
      RECT 35.76 3.945 35.765 4.164 ;
      RECT 35.745 3.932 35.76 4.156 ;
      RECT 35.74 3.842 35.745 4.145 ;
      RECT 35.735 3.837 35.74 4.138 ;
      RECT 35.66 3.835 35.735 4.098 ;
      RECT 35.63 3.835 35.66 4.053 ;
      RECT 35.535 3.84 35.55 4.04 ;
      RECT 38.02 3.545 38.28 3.805 ;
      RECT 38.005 3.533 38.185 3.77 ;
      RECT 38 3.534 38.185 3.768 ;
      RECT 37.985 3.538 38.195 3.758 ;
      RECT 37.98 3.543 38.2 3.728 ;
      RECT 37.985 3.54 38.2 3.758 ;
      RECT 38 3.535 38.195 3.768 ;
      RECT 38.02 3.532 38.185 3.805 ;
      RECT 38.02 3.531 38.175 3.805 ;
      RECT 38.045 3.53 38.175 3.805 ;
      RECT 37.605 3.775 37.865 4.035 ;
      RECT 37.48 3.82 37.865 4.03 ;
      RECT 37.47 3.825 37.865 4.025 ;
      RECT 37.485 4.765 37.5 5.075 ;
      RECT 36.08 4.535 36.09 4.665 ;
      RECT 35.86 4.53 35.965 4.665 ;
      RECT 35.775 4.535 35.825 4.665 ;
      RECT 34.325 3.27 34.33 4.375 ;
      RECT 37.58 4.857 37.585 4.993 ;
      RECT 37.575 4.852 37.58 5.053 ;
      RECT 37.57 4.85 37.575 5.066 ;
      RECT 37.555 4.847 37.57 5.068 ;
      RECT 37.55 4.842 37.555 5.07 ;
      RECT 37.545 4.838 37.55 5.073 ;
      RECT 37.53 4.833 37.545 5.075 ;
      RECT 37.5 4.825 37.53 5.075 ;
      RECT 37.461 4.765 37.485 5.075 ;
      RECT 37.375 4.765 37.461 5.072 ;
      RECT 37.345 4.765 37.375 5.065 ;
      RECT 37.32 4.765 37.345 5.058 ;
      RECT 37.295 4.765 37.32 5.05 ;
      RECT 37.28 4.765 37.295 5.043 ;
      RECT 37.255 4.765 37.28 5.035 ;
      RECT 37.24 4.765 37.255 5.028 ;
      RECT 37.2 4.775 37.24 5.017 ;
      RECT 37.19 4.77 37.2 5.007 ;
      RECT 37.186 4.769 37.19 5.004 ;
      RECT 37.1 4.761 37.186 4.987 ;
      RECT 37.067 4.75 37.1 4.964 ;
      RECT 36.981 4.739 37.067 4.942 ;
      RECT 36.895 4.723 36.981 4.911 ;
      RECT 36.825 4.708 36.895 4.883 ;
      RECT 36.815 4.701 36.825 4.87 ;
      RECT 36.785 4.698 36.815 4.86 ;
      RECT 36.76 4.694 36.785 4.853 ;
      RECT 36.745 4.691 36.76 4.848 ;
      RECT 36.74 4.69 36.745 4.843 ;
      RECT 36.71 4.685 36.74 4.836 ;
      RECT 36.705 4.68 36.71 4.831 ;
      RECT 36.69 4.677 36.705 4.826 ;
      RECT 36.685 4.672 36.69 4.821 ;
      RECT 36.665 4.667 36.685 4.818 ;
      RECT 36.65 4.662 36.665 4.81 ;
      RECT 36.635 4.656 36.65 4.805 ;
      RECT 36.605 4.647 36.635 4.798 ;
      RECT 36.6 4.64 36.605 4.79 ;
      RECT 36.595 4.638 36.6 4.788 ;
      RECT 36.59 4.637 36.595 4.785 ;
      RECT 36.55 4.63 36.59 4.778 ;
      RECT 36.536 4.62 36.55 4.768 ;
      RECT 36.485 4.609 36.536 4.756 ;
      RECT 36.46 4.595 36.485 4.742 ;
      RECT 36.435 4.584 36.46 4.734 ;
      RECT 36.415 4.573 36.435 4.728 ;
      RECT 36.405 4.567 36.415 4.723 ;
      RECT 36.4 4.565 36.405 4.719 ;
      RECT 36.38 4.56 36.4 4.714 ;
      RECT 36.35 4.55 36.38 4.704 ;
      RECT 36.345 4.542 36.35 4.697 ;
      RECT 36.33 4.54 36.345 4.693 ;
      RECT 36.31 4.54 36.33 4.688 ;
      RECT 36.305 4.539 36.31 4.686 ;
      RECT 36.3 4.539 36.305 4.683 ;
      RECT 36.26 4.538 36.3 4.678 ;
      RECT 36.235 4.537 36.26 4.673 ;
      RECT 36.175 4.536 36.235 4.67 ;
      RECT 36.09 4.535 36.175 4.668 ;
      RECT 36.051 4.534 36.08 4.665 ;
      RECT 35.965 4.532 36.051 4.665 ;
      RECT 35.825 4.532 35.86 4.665 ;
      RECT 35.735 4.536 35.775 4.668 ;
      RECT 35.72 4.539 35.735 4.675 ;
      RECT 35.71 4.54 35.72 4.682 ;
      RECT 35.685 4.543 35.71 4.687 ;
      RECT 35.68 4.545 35.685 4.69 ;
      RECT 35.63 4.547 35.68 4.691 ;
      RECT 35.591 4.551 35.63 4.693 ;
      RECT 35.505 4.553 35.591 4.696 ;
      RECT 35.487 4.555 35.505 4.698 ;
      RECT 35.401 4.558 35.487 4.7 ;
      RECT 35.315 4.562 35.401 4.703 ;
      RECT 35.278 4.566 35.315 4.706 ;
      RECT 35.192 4.569 35.278 4.709 ;
      RECT 35.106 4.573 35.192 4.712 ;
      RECT 35.02 4.578 35.106 4.716 ;
      RECT 35 4.58 35.02 4.719 ;
      RECT 34.98 4.579 35 4.72 ;
      RECT 34.931 4.576 34.98 4.721 ;
      RECT 34.845 4.571 34.931 4.724 ;
      RECT 34.795 4.566 34.845 4.726 ;
      RECT 34.771 4.564 34.795 4.727 ;
      RECT 34.685 4.559 34.771 4.729 ;
      RECT 34.66 4.555 34.685 4.728 ;
      RECT 34.65 4.552 34.66 4.726 ;
      RECT 34.64 4.545 34.65 4.723 ;
      RECT 34.635 4.525 34.64 4.718 ;
      RECT 34.625 4.495 34.635 4.713 ;
      RECT 34.61 4.365 34.625 4.704 ;
      RECT 34.605 4.357 34.61 4.697 ;
      RECT 34.585 4.35 34.605 4.689 ;
      RECT 34.58 4.332 34.585 4.681 ;
      RECT 34.57 4.312 34.58 4.676 ;
      RECT 34.565 4.285 34.57 4.672 ;
      RECT 34.56 4.262 34.565 4.669 ;
      RECT 34.54 4.22 34.56 4.661 ;
      RECT 34.505 4.135 34.54 4.645 ;
      RECT 34.5 4.067 34.505 4.633 ;
      RECT 34.485 4.037 34.5 4.627 ;
      RECT 34.48 3.282 34.485 3.528 ;
      RECT 34.47 4.007 34.485 4.618 ;
      RECT 34.475 3.277 34.48 3.56 ;
      RECT 34.47 3.272 34.475 3.603 ;
      RECT 34.465 3.27 34.47 3.638 ;
      RECT 34.45 3.97 34.47 4.608 ;
      RECT 34.46 3.27 34.465 3.675 ;
      RECT 34.445 3.27 34.46 3.773 ;
      RECT 34.445 3.943 34.45 4.601 ;
      RECT 34.44 3.27 34.445 3.848 ;
      RECT 34.44 3.931 34.445 4.598 ;
      RECT 34.435 3.27 34.44 3.88 ;
      RECT 34.435 3.91 34.44 4.595 ;
      RECT 34.43 3.27 34.435 4.592 ;
      RECT 34.395 3.27 34.43 4.578 ;
      RECT 34.38 3.27 34.395 4.56 ;
      RECT 34.36 3.27 34.38 4.55 ;
      RECT 34.335 3.27 34.36 4.533 ;
      RECT 34.33 3.27 34.335 4.483 ;
      RECT 34.32 3.27 34.325 4.313 ;
      RECT 34.315 3.27 34.32 4.22 ;
      RECT 34.31 3.27 34.315 4.133 ;
      RECT 34.305 3.27 34.31 4.065 ;
      RECT 34.3 3.27 34.305 4.008 ;
      RECT 34.29 3.27 34.3 3.903 ;
      RECT 34.285 3.27 34.29 3.775 ;
      RECT 34.28 3.27 34.285 3.693 ;
      RECT 34.275 3.272 34.28 3.61 ;
      RECT 34.27 3.277 34.275 3.543 ;
      RECT 34.265 3.282 34.27 3.47 ;
      RECT 37.08 3.6 37.34 3.86 ;
      RECT 37.1 3.567 37.31 3.86 ;
      RECT 37.1 3.565 37.3 3.86 ;
      RECT 37.11 3.552 37.3 3.86 ;
      RECT 37.11 3.55 37.225 3.86 ;
      RECT 36.585 3.675 36.76 3.955 ;
      RECT 36.58 3.675 36.76 3.953 ;
      RECT 36.58 3.675 36.775 3.95 ;
      RECT 36.57 3.675 36.775 3.948 ;
      RECT 36.515 3.675 36.775 3.935 ;
      RECT 36.515 3.75 36.78 3.913 ;
      RECT 36.06 3.687 36.08 3.93 ;
      RECT 36.06 3.687 36.12 3.929 ;
      RECT 36.055 3.689 36.12 3.928 ;
      RECT 36.055 3.689 36.206 3.927 ;
      RECT 36.055 3.689 36.275 3.926 ;
      RECT 36.055 3.689 36.295 3.918 ;
      RECT 36.035 3.692 36.295 3.916 ;
      RECT 36.02 3.702 36.295 3.901 ;
      RECT 36.02 3.702 36.31 3.9 ;
      RECT 36.015 3.711 36.31 3.892 ;
      RECT 36.015 3.711 36.315 3.888 ;
      RECT 36.12 3.625 36.38 3.885 ;
      RECT 36.01 3.713 36.38 3.77 ;
      RECT 36.08 3.68 36.38 3.885 ;
      RECT 36.045 4.873 36.05 5.08 ;
      RECT 35.995 4.867 36.045 5.079 ;
      RECT 35.962 4.881 36.055 5.078 ;
      RECT 35.876 4.881 36.055 5.077 ;
      RECT 35.79 4.881 36.055 5.076 ;
      RECT 35.79 4.98 36.06 5.073 ;
      RECT 35.785 4.98 36.06 5.068 ;
      RECT 35.78 4.98 36.06 5.05 ;
      RECT 35.775 4.98 36.06 5.033 ;
      RECT 35.735 4.765 35.995 5.025 ;
      RECT 35.195 3.915 35.281 4.329 ;
      RECT 35.195 3.915 35.32 4.326 ;
      RECT 35.195 3.915 35.34 4.316 ;
      RECT 35.15 3.915 35.34 4.313 ;
      RECT 35.15 4.067 35.35 4.303 ;
      RECT 35.15 4.088 35.355 4.297 ;
      RECT 35.15 4.106 35.36 4.293 ;
      RECT 35.15 4.126 35.37 4.288 ;
      RECT 35.125 4.126 35.37 4.285 ;
      RECT 35.115 4.126 35.37 4.263 ;
      RECT 35.115 4.142 35.375 4.233 ;
      RECT 35.08 3.915 35.34 4.22 ;
      RECT 35.08 4.154 35.38 4.175 ;
      RECT 32.74 10.06 33.03 10.29 ;
      RECT 32.8 8.58 32.97 10.29 ;
      RECT 32.79 8.95 33.145 9.305 ;
      RECT 32.74 8.58 33.03 8.81 ;
      RECT 32.335 3.69 32.44 4.26 ;
      RECT 32.335 4.025 32.66 4.255 ;
      RECT 32.335 4.055 32.83 4.225 ;
      RECT 32.335 3.69 32.525 4.255 ;
      RECT 31.75 3.655 32.04 3.885 ;
      RECT 31.75 3.69 32.525 3.86 ;
      RECT 31.81 2.175 31.98 3.885 ;
      RECT 31.75 2.175 32.04 2.405 ;
      RECT 31.75 10.06 32.04 10.29 ;
      RECT 31.81 8.58 31.98 10.29 ;
      RECT 31.75 8.58 32.04 8.81 ;
      RECT 31.75 8.615 32.6 8.775 ;
      RECT 32.435 8.21 32.6 8.775 ;
      RECT 31.75 8.61 32.145 8.775 ;
      RECT 32.37 8.21 32.66 8.44 ;
      RECT 32.37 8.24 32.83 8.41 ;
      RECT 31.38 4.025 31.67 4.255 ;
      RECT 31.38 4.055 31.84 4.225 ;
      RECT 31.445 2.95 31.61 4.255 ;
      RECT 29.96 2.92 30.25 3.15 ;
      RECT 29.96 2.95 31.61 3.12 ;
      RECT 30.02 2.18 30.19 3.15 ;
      RECT 29.96 2.18 30.25 2.41 ;
      RECT 29.96 10.055 30.25 10.285 ;
      RECT 30.02 9.315 30.19 10.285 ;
      RECT 30.02 9.41 31.61 9.58 ;
      RECT 31.44 8.21 31.61 9.58 ;
      RECT 29.96 9.315 30.25 9.545 ;
      RECT 31.38 8.21 31.67 8.44 ;
      RECT 31.38 8.24 31.84 8.41 ;
      RECT 28.01 4 28.35 4.35 ;
      RECT 28.1 3.32 28.27 4.35 ;
      RECT 30.39 3.26 30.74 3.61 ;
      RECT 28.1 3.32 30.74 3.49 ;
      RECT 30.415 8.945 30.74 9.27 ;
      RECT 24.955 8.9 25.305 9.25 ;
      RECT 30.39 8.945 30.74 9.175 ;
      RECT 24.755 8.945 25.305 9.175 ;
      RECT 24.585 8.975 30.74 9.145 ;
      RECT 29.615 3.66 29.935 3.98 ;
      RECT 29.585 3.66 29.935 3.89 ;
      RECT 29.415 3.69 29.935 3.86 ;
      RECT 29.615 8.545 29.935 8.835 ;
      RECT 29.585 8.575 29.935 8.805 ;
      RECT 29.415 8.605 29.935 8.775 ;
      RECT 25.305 4.28 25.455 4.555 ;
      RECT 25.845 3.36 25.85 3.58 ;
      RECT 26.995 3.56 27.01 3.758 ;
      RECT 26.96 3.552 26.995 3.765 ;
      RECT 26.93 3.545 26.96 3.765 ;
      RECT 26.875 3.51 26.93 3.765 ;
      RECT 26.81 3.447 26.875 3.765 ;
      RECT 26.805 3.412 26.81 3.763 ;
      RECT 26.8 3.407 26.805 3.755 ;
      RECT 26.795 3.402 26.8 3.741 ;
      RECT 26.79 3.399 26.795 3.734 ;
      RECT 26.745 3.389 26.79 3.685 ;
      RECT 26.725 3.376 26.745 3.62 ;
      RECT 26.72 3.371 26.725 3.593 ;
      RECT 26.715 3.37 26.72 3.586 ;
      RECT 26.71 3.369 26.715 3.579 ;
      RECT 26.625 3.354 26.71 3.525 ;
      RECT 26.595 3.335 26.625 3.475 ;
      RECT 26.515 3.318 26.595 3.46 ;
      RECT 26.48 3.305 26.515 3.445 ;
      RECT 26.472 3.305 26.48 3.44 ;
      RECT 26.386 3.306 26.472 3.44 ;
      RECT 26.3 3.308 26.386 3.44 ;
      RECT 26.275 3.309 26.3 3.444 ;
      RECT 26.2 3.315 26.275 3.459 ;
      RECT 26.117 3.327 26.2 3.483 ;
      RECT 26.031 3.34 26.117 3.509 ;
      RECT 25.945 3.353 26.031 3.535 ;
      RECT 25.91 3.362 25.945 3.554 ;
      RECT 25.86 3.362 25.91 3.567 ;
      RECT 25.85 3.36 25.86 3.578 ;
      RECT 25.835 3.357 25.845 3.58 ;
      RECT 25.82 3.349 25.835 3.588 ;
      RECT 25.805 3.341 25.82 3.608 ;
      RECT 25.8 3.336 25.805 3.665 ;
      RECT 25.785 3.331 25.8 3.738 ;
      RECT 25.78 3.326 25.785 3.78 ;
      RECT 25.775 3.324 25.78 3.808 ;
      RECT 25.77 3.322 25.775 3.83 ;
      RECT 25.76 3.318 25.77 3.873 ;
      RECT 25.755 3.315 25.76 3.898 ;
      RECT 25.75 3.313 25.755 3.918 ;
      RECT 25.745 3.311 25.75 3.942 ;
      RECT 25.74 3.307 25.745 3.965 ;
      RECT 25.735 3.303 25.74 3.988 ;
      RECT 25.7 3.293 25.735 4.095 ;
      RECT 25.695 3.283 25.7 4.193 ;
      RECT 25.69 3.281 25.695 4.22 ;
      RECT 25.685 3.28 25.69 4.24 ;
      RECT 25.68 3.272 25.685 4.26 ;
      RECT 25.675 3.267 25.68 4.295 ;
      RECT 25.67 3.265 25.675 4.313 ;
      RECT 25.665 3.265 25.67 4.338 ;
      RECT 25.66 3.265 25.665 4.36 ;
      RECT 25.625 3.265 25.66 4.403 ;
      RECT 25.6 3.265 25.625 4.432 ;
      RECT 25.59 3.265 25.6 3.618 ;
      RECT 25.593 3.675 25.6 4.442 ;
      RECT 25.59 3.732 25.593 4.445 ;
      RECT 25.585 3.265 25.59 3.59 ;
      RECT 25.585 3.782 25.59 4.448 ;
      RECT 25.575 3.265 25.585 3.58 ;
      RECT 25.58 3.835 25.585 4.451 ;
      RECT 25.575 3.92 25.58 4.455 ;
      RECT 25.565 3.265 25.575 3.568 ;
      RECT 25.57 3.967 25.575 4.459 ;
      RECT 25.565 4.042 25.57 4.463 ;
      RECT 25.53 3.265 25.565 3.543 ;
      RECT 25.555 4.125 25.565 4.468 ;
      RECT 25.545 4.192 25.555 4.475 ;
      RECT 25.54 4.22 25.545 4.48 ;
      RECT 25.53 4.233 25.54 4.486 ;
      RECT 25.485 3.265 25.53 3.5 ;
      RECT 25.525 4.238 25.53 4.493 ;
      RECT 25.485 4.255 25.525 4.555 ;
      RECT 25.48 3.267 25.485 3.473 ;
      RECT 25.455 4.275 25.485 4.555 ;
      RECT 25.475 3.272 25.48 3.445 ;
      RECT 25.265 4.284 25.305 4.555 ;
      RECT 25.24 4.292 25.265 4.525 ;
      RECT 25.195 4.3 25.24 4.525 ;
      RECT 25.18 4.305 25.195 4.52 ;
      RECT 25.17 4.305 25.18 4.514 ;
      RECT 25.16 4.312 25.17 4.511 ;
      RECT 25.155 4.35 25.16 4.5 ;
      RECT 25.15 4.412 25.155 4.478 ;
      RECT 26.42 4.287 26.605 4.51 ;
      RECT 26.42 4.302 26.61 4.506 ;
      RECT 26.41 3.575 26.495 4.505 ;
      RECT 26.41 4.302 26.615 4.499 ;
      RECT 26.405 4.31 26.615 4.498 ;
      RECT 26.61 4.03 26.93 4.35 ;
      RECT 26.405 4.202 26.575 4.293 ;
      RECT 26.4 4.202 26.575 4.275 ;
      RECT 26.39 4.01 26.525 4.25 ;
      RECT 26.385 4.01 26.525 4.195 ;
      RECT 26.345 3.59 26.515 4.095 ;
      RECT 26.33 3.59 26.515 3.965 ;
      RECT 26.325 3.59 26.515 3.918 ;
      RECT 26.32 3.59 26.515 3.898 ;
      RECT 26.315 3.59 26.515 3.873 ;
      RECT 26.285 3.59 26.545 3.85 ;
      RECT 26.295 3.587 26.505 3.85 ;
      RECT 26.42 3.582 26.505 4.51 ;
      RECT 26.305 3.575 26.495 3.85 ;
      RECT 26.3 3.58 26.495 3.85 ;
      RECT 25.13 3.792 25.315 4.005 ;
      RECT 25.13 3.8 25.325 3.998 ;
      RECT 25.11 3.8 25.325 3.995 ;
      RECT 25.105 3.8 25.325 3.98 ;
      RECT 25.035 3.715 25.295 3.975 ;
      RECT 25.035 3.86 25.33 3.888 ;
      RECT 24.69 4.315 24.95 4.575 ;
      RECT 24.715 4.26 24.91 4.575 ;
      RECT 24.71 4.009 24.89 4.303 ;
      RECT 24.71 4.015 24.9 4.303 ;
      RECT 24.69 4.017 24.9 4.248 ;
      RECT 24.685 4.027 24.9 4.115 ;
      RECT 24.715 4.007 24.89 4.575 ;
      RECT 24.801 4.005 24.89 4.575 ;
      RECT 24.66 3.225 24.695 3.595 ;
      RECT 24.45 3.335 24.455 3.595 ;
      RECT 24.695 3.232 24.71 3.595 ;
      RECT 24.585 3.225 24.66 3.673 ;
      RECT 24.575 3.225 24.585 3.758 ;
      RECT 24.55 3.225 24.575 3.793 ;
      RECT 24.51 3.225 24.55 3.861 ;
      RECT 24.5 3.232 24.51 3.913 ;
      RECT 24.47 3.335 24.5 3.954 ;
      RECT 24.465 3.335 24.47 3.993 ;
      RECT 24.455 3.335 24.465 4.013 ;
      RECT 24.45 3.63 24.455 4.05 ;
      RECT 24.445 3.647 24.45 4.07 ;
      RECT 24.43 3.71 24.445 4.11 ;
      RECT 24.425 3.753 24.43 4.145 ;
      RECT 24.42 3.761 24.425 4.158 ;
      RECT 24.41 3.775 24.42 4.18 ;
      RECT 24.385 3.81 24.41 4.245 ;
      RECT 24.375 3.845 24.385 4.308 ;
      RECT 24.355 3.875 24.375 4.369 ;
      RECT 24.34 3.911 24.355 4.436 ;
      RECT 24.33 3.939 24.34 4.475 ;
      RECT 24.32 3.961 24.33 4.495 ;
      RECT 24.315 3.971 24.32 4.506 ;
      RECT 24.31 3.98 24.315 4.509 ;
      RECT 24.3 3.998 24.31 4.513 ;
      RECT 24.29 4.016 24.3 4.514 ;
      RECT 24.265 4.055 24.29 4.511 ;
      RECT 24.245 4.097 24.265 4.508 ;
      RECT 24.23 4.135 24.245 4.507 ;
      RECT 24.195 4.17 24.23 4.504 ;
      RECT 24.19 4.192 24.195 4.502 ;
      RECT 24.125 4.232 24.19 4.499 ;
      RECT 24.12 4.272 24.125 4.495 ;
      RECT 24.105 4.282 24.12 4.486 ;
      RECT 24.095 4.402 24.105 4.471 ;
      RECT 24.575 4.815 24.585 5.075 ;
      RECT 24.575 4.818 24.595 5.074 ;
      RECT 24.565 4.808 24.575 5.073 ;
      RECT 24.555 4.823 24.635 5.069 ;
      RECT 24.54 4.802 24.555 5.067 ;
      RECT 24.515 4.827 24.64 5.063 ;
      RECT 24.5 4.787 24.515 5.058 ;
      RECT 24.5 4.829 24.65 5.057 ;
      RECT 24.5 4.837 24.665 5.05 ;
      RECT 24.44 4.774 24.5 5.04 ;
      RECT 24.43 4.761 24.44 5.022 ;
      RECT 24.405 4.751 24.43 5.012 ;
      RECT 24.4 4.741 24.405 5.004 ;
      RECT 24.335 4.837 24.665 4.986 ;
      RECT 24.25 4.837 24.665 4.948 ;
      RECT 24.14 4.665 24.4 4.925 ;
      RECT 24.515 4.795 24.54 5.063 ;
      RECT 24.555 4.805 24.565 5.069 ;
      RECT 24.14 4.813 24.58 4.925 ;
      RECT 24.325 10.055 24.615 10.285 ;
      RECT 24.385 9.315 24.555 10.285 ;
      RECT 24.285 9.345 24.655 9.715 ;
      RECT 24.325 9.315 24.615 9.715 ;
      RECT 23.355 4.57 23.385 4.87 ;
      RECT 23.13 4.555 23.135 4.83 ;
      RECT 22.93 4.555 23.085 4.815 ;
      RECT 24.23 3.27 24.26 3.53 ;
      RECT 24.22 3.27 24.23 3.638 ;
      RECT 24.2 3.27 24.22 3.648 ;
      RECT 24.185 3.27 24.2 3.66 ;
      RECT 24.13 3.27 24.185 3.71 ;
      RECT 24.115 3.27 24.13 3.758 ;
      RECT 24.085 3.27 24.115 3.793 ;
      RECT 24.03 3.27 24.085 3.855 ;
      RECT 24.01 3.27 24.03 3.923 ;
      RECT 24.005 3.27 24.01 3.953 ;
      RECT 24 3.27 24.005 3.965 ;
      RECT 23.995 3.387 24 3.983 ;
      RECT 23.975 3.405 23.995 4.008 ;
      RECT 23.955 3.432 23.975 4.058 ;
      RECT 23.95 3.452 23.955 4.089 ;
      RECT 23.945 3.46 23.95 4.106 ;
      RECT 23.93 3.486 23.945 4.135 ;
      RECT 23.915 3.528 23.93 4.17 ;
      RECT 23.91 3.557 23.915 4.193 ;
      RECT 23.905 3.572 23.91 4.206 ;
      RECT 23.9 3.595 23.905 4.217 ;
      RECT 23.89 3.615 23.9 4.235 ;
      RECT 23.88 3.645 23.89 4.258 ;
      RECT 23.875 3.667 23.88 4.278 ;
      RECT 23.87 3.682 23.875 4.293 ;
      RECT 23.855 3.712 23.87 4.32 ;
      RECT 23.85 3.742 23.855 4.346 ;
      RECT 23.845 3.76 23.85 4.358 ;
      RECT 23.835 3.79 23.845 4.377 ;
      RECT 23.825 3.815 23.835 4.402 ;
      RECT 23.82 3.835 23.825 4.421 ;
      RECT 23.815 3.852 23.82 4.434 ;
      RECT 23.805 3.878 23.815 4.453 ;
      RECT 23.795 3.916 23.805 4.48 ;
      RECT 23.79 3.942 23.795 4.5 ;
      RECT 23.785 3.952 23.79 4.51 ;
      RECT 23.78 3.965 23.785 4.525 ;
      RECT 23.775 3.98 23.78 4.535 ;
      RECT 23.77 4.002 23.775 4.55 ;
      RECT 23.765 4.02 23.77 4.561 ;
      RECT 23.76 4.03 23.765 4.572 ;
      RECT 23.755 4.038 23.76 4.584 ;
      RECT 23.75 4.046 23.755 4.595 ;
      RECT 23.745 4.072 23.75 4.608 ;
      RECT 23.735 4.1 23.745 4.621 ;
      RECT 23.73 4.13 23.735 4.63 ;
      RECT 23.725 4.145 23.73 4.637 ;
      RECT 23.71 4.17 23.725 4.644 ;
      RECT 23.705 4.192 23.71 4.65 ;
      RECT 23.7 4.217 23.705 4.653 ;
      RECT 23.691 4.245 23.7 4.657 ;
      RECT 23.685 4.262 23.691 4.662 ;
      RECT 23.68 4.28 23.685 4.666 ;
      RECT 23.675 4.292 23.68 4.669 ;
      RECT 23.67 4.313 23.675 4.673 ;
      RECT 23.665 4.331 23.67 4.676 ;
      RECT 23.66 4.345 23.665 4.679 ;
      RECT 23.655 4.362 23.66 4.682 ;
      RECT 23.65 4.375 23.655 4.685 ;
      RECT 23.625 4.412 23.65 4.693 ;
      RECT 23.62 4.457 23.625 4.702 ;
      RECT 23.615 4.485 23.62 4.705 ;
      RECT 23.605 4.505 23.615 4.709 ;
      RECT 23.6 4.525 23.605 4.714 ;
      RECT 23.595 4.54 23.6 4.717 ;
      RECT 23.575 4.55 23.595 4.724 ;
      RECT 23.51 4.557 23.575 4.75 ;
      RECT 23.475 4.56 23.51 4.778 ;
      RECT 23.46 4.563 23.475 4.793 ;
      RECT 23.45 4.564 23.46 4.808 ;
      RECT 23.44 4.565 23.45 4.825 ;
      RECT 23.435 4.565 23.44 4.84 ;
      RECT 23.43 4.565 23.435 4.848 ;
      RECT 23.415 4.566 23.43 4.863 ;
      RECT 23.385 4.568 23.415 4.87 ;
      RECT 23.275 4.575 23.355 4.87 ;
      RECT 23.23 4.58 23.275 4.87 ;
      RECT 23.22 4.581 23.23 4.86 ;
      RECT 23.21 4.582 23.22 4.853 ;
      RECT 23.19 4.584 23.21 4.848 ;
      RECT 23.18 4.555 23.19 4.843 ;
      RECT 23.135 4.555 23.18 4.835 ;
      RECT 23.105 4.555 23.13 4.825 ;
      RECT 23.085 4.555 23.105 4.818 ;
      RECT 23.365 3.355 23.625 3.615 ;
      RECT 23.245 3.37 23.255 3.535 ;
      RECT 23.23 3.37 23.235 3.53 ;
      RECT 20.595 3.21 20.78 3.5 ;
      RECT 22.41 3.335 22.425 3.49 ;
      RECT 20.56 3.21 20.585 3.47 ;
      RECT 22.975 3.26 22.98 3.402 ;
      RECT 22.89 3.255 22.915 3.395 ;
      RECT 23.29 3.372 23.365 3.565 ;
      RECT 23.275 3.37 23.29 3.548 ;
      RECT 23.255 3.37 23.275 3.54 ;
      RECT 23.235 3.37 23.245 3.533 ;
      RECT 23.19 3.365 23.23 3.523 ;
      RECT 23.15 3.34 23.19 3.508 ;
      RECT 23.135 3.315 23.15 3.498 ;
      RECT 23.13 3.309 23.135 3.496 ;
      RECT 23.095 3.301 23.13 3.479 ;
      RECT 23.09 3.294 23.095 3.467 ;
      RECT 23.07 3.289 23.09 3.455 ;
      RECT 23.06 3.283 23.07 3.44 ;
      RECT 23.04 3.278 23.06 3.425 ;
      RECT 23.03 3.273 23.04 3.418 ;
      RECT 23.025 3.271 23.03 3.413 ;
      RECT 23.02 3.27 23.025 3.41 ;
      RECT 22.98 3.265 23.02 3.406 ;
      RECT 22.96 3.259 22.975 3.401 ;
      RECT 22.925 3.256 22.96 3.398 ;
      RECT 22.915 3.255 22.925 3.396 ;
      RECT 22.855 3.255 22.89 3.393 ;
      RECT 22.81 3.255 22.855 3.393 ;
      RECT 22.76 3.255 22.81 3.396 ;
      RECT 22.745 3.257 22.76 3.398 ;
      RECT 22.73 3.26 22.745 3.399 ;
      RECT 22.72 3.265 22.73 3.4 ;
      RECT 22.69 3.27 22.72 3.405 ;
      RECT 22.68 3.276 22.69 3.413 ;
      RECT 22.67 3.278 22.68 3.417 ;
      RECT 22.66 3.282 22.67 3.421 ;
      RECT 22.635 3.288 22.66 3.429 ;
      RECT 22.625 3.293 22.635 3.437 ;
      RECT 22.61 3.297 22.625 3.441 ;
      RECT 22.575 3.303 22.61 3.449 ;
      RECT 22.555 3.308 22.575 3.459 ;
      RECT 22.525 3.315 22.555 3.468 ;
      RECT 22.48 3.324 22.525 3.482 ;
      RECT 22.475 3.329 22.48 3.493 ;
      RECT 22.455 3.332 22.475 3.494 ;
      RECT 22.425 3.335 22.455 3.492 ;
      RECT 22.39 3.335 22.41 3.488 ;
      RECT 22.32 3.335 22.39 3.479 ;
      RECT 22.305 3.332 22.32 3.471 ;
      RECT 22.265 3.325 22.305 3.466 ;
      RECT 22.24 3.315 22.265 3.459 ;
      RECT 22.235 3.309 22.24 3.456 ;
      RECT 22.195 3.303 22.235 3.453 ;
      RECT 22.18 3.296 22.195 3.448 ;
      RECT 22.16 3.292 22.18 3.443 ;
      RECT 22.145 3.287 22.16 3.439 ;
      RECT 22.13 3.282 22.145 3.437 ;
      RECT 22.115 3.278 22.13 3.436 ;
      RECT 22.1 3.276 22.115 3.432 ;
      RECT 22.09 3.274 22.1 3.427 ;
      RECT 22.075 3.271 22.09 3.423 ;
      RECT 22.065 3.269 22.075 3.418 ;
      RECT 22.045 3.266 22.065 3.414 ;
      RECT 22 3.265 22.045 3.412 ;
      RECT 21.94 3.267 22 3.413 ;
      RECT 21.92 3.269 21.94 3.415 ;
      RECT 21.89 3.272 21.92 3.416 ;
      RECT 21.84 3.277 21.89 3.418 ;
      RECT 21.835 3.28 21.84 3.42 ;
      RECT 21.825 3.282 21.835 3.423 ;
      RECT 21.82 3.284 21.825 3.426 ;
      RECT 21.77 3.287 21.82 3.433 ;
      RECT 21.75 3.291 21.77 3.445 ;
      RECT 21.74 3.294 21.75 3.451 ;
      RECT 21.73 3.295 21.74 3.454 ;
      RECT 21.691 3.298 21.73 3.456 ;
      RECT 21.605 3.305 21.691 3.459 ;
      RECT 21.531 3.315 21.605 3.463 ;
      RECT 21.445 3.326 21.531 3.468 ;
      RECT 21.43 3.333 21.445 3.47 ;
      RECT 21.375 3.337 21.43 3.471 ;
      RECT 21.361 3.34 21.375 3.473 ;
      RECT 21.275 3.34 21.361 3.475 ;
      RECT 21.235 3.337 21.275 3.478 ;
      RECT 21.211 3.333 21.235 3.48 ;
      RECT 21.125 3.323 21.211 3.483 ;
      RECT 21.095 3.312 21.125 3.484 ;
      RECT 21.076 3.308 21.095 3.483 ;
      RECT 20.99 3.301 21.076 3.48 ;
      RECT 20.93 3.29 20.99 3.477 ;
      RECT 20.91 3.282 20.93 3.475 ;
      RECT 20.875 3.277 20.91 3.474 ;
      RECT 20.85 3.272 20.875 3.473 ;
      RECT 20.82 3.267 20.85 3.472 ;
      RECT 20.795 3.21 20.82 3.471 ;
      RECT 20.78 3.21 20.795 3.495 ;
      RECT 20.585 3.21 20.595 3.495 ;
      RECT 22.36 4.23 22.365 4.37 ;
      RECT 22.02 4.23 22.055 4.368 ;
      RECT 21.595 4.215 21.61 4.36 ;
      RECT 23.425 3.995 23.515 4.255 ;
      RECT 23.255 3.86 23.355 4.255 ;
      RECT 20.29 3.835 20.37 4.045 ;
      RECT 23.38 3.972 23.425 4.255 ;
      RECT 23.37 3.942 23.38 4.255 ;
      RECT 23.355 3.865 23.37 4.255 ;
      RECT 23.17 3.86 23.255 4.22 ;
      RECT 23.165 3.862 23.17 4.215 ;
      RECT 23.16 3.867 23.165 4.215 ;
      RECT 23.125 3.967 23.16 4.215 ;
      RECT 23.115 3.995 23.125 4.215 ;
      RECT 23.105 4.01 23.115 4.215 ;
      RECT 23.095 4.022 23.105 4.215 ;
      RECT 23.09 4.032 23.095 4.215 ;
      RECT 23.075 4.042 23.09 4.217 ;
      RECT 23.07 4.057 23.075 4.219 ;
      RECT 23.055 4.07 23.07 4.221 ;
      RECT 23.05 4.085 23.055 4.224 ;
      RECT 23.03 4.095 23.05 4.228 ;
      RECT 23.015 4.105 23.03 4.231 ;
      RECT 22.98 4.112 23.015 4.236 ;
      RECT 22.936 4.119 22.98 4.244 ;
      RECT 22.85 4.131 22.936 4.257 ;
      RECT 22.825 4.142 22.85 4.268 ;
      RECT 22.795 4.147 22.825 4.273 ;
      RECT 22.76 4.152 22.795 4.281 ;
      RECT 22.73 4.157 22.76 4.288 ;
      RECT 22.705 4.162 22.73 4.293 ;
      RECT 22.64 4.169 22.705 4.302 ;
      RECT 22.57 4.182 22.64 4.318 ;
      RECT 22.54 4.192 22.57 4.33 ;
      RECT 22.515 4.197 22.54 4.337 ;
      RECT 22.46 4.204 22.515 4.345 ;
      RECT 22.455 4.211 22.46 4.35 ;
      RECT 22.45 4.213 22.455 4.351 ;
      RECT 22.435 4.215 22.45 4.353 ;
      RECT 22.43 4.215 22.435 4.356 ;
      RECT 22.365 4.222 22.43 4.363 ;
      RECT 22.33 4.232 22.36 4.373 ;
      RECT 22.313 4.235 22.33 4.375 ;
      RECT 22.227 4.234 22.313 4.374 ;
      RECT 22.141 4.232 22.227 4.371 ;
      RECT 22.055 4.231 22.141 4.369 ;
      RECT 21.954 4.229 22.02 4.368 ;
      RECT 21.868 4.226 21.954 4.366 ;
      RECT 21.782 4.222 21.868 4.364 ;
      RECT 21.696 4.219 21.782 4.363 ;
      RECT 21.61 4.216 21.696 4.361 ;
      RECT 21.51 4.215 21.595 4.358 ;
      RECT 21.46 4.213 21.51 4.356 ;
      RECT 21.44 4.21 21.46 4.354 ;
      RECT 21.42 4.208 21.44 4.351 ;
      RECT 21.395 4.204 21.42 4.348 ;
      RECT 21.35 4.198 21.395 4.343 ;
      RECT 21.31 4.192 21.35 4.335 ;
      RECT 21.285 4.187 21.31 4.328 ;
      RECT 21.23 4.18 21.285 4.32 ;
      RECT 21.206 4.173 21.23 4.313 ;
      RECT 21.12 4.164 21.206 4.303 ;
      RECT 21.09 4.156 21.12 4.293 ;
      RECT 21.06 4.152 21.09 4.288 ;
      RECT 21.055 4.149 21.06 4.285 ;
      RECT 21.05 4.148 21.055 4.285 ;
      RECT 20.975 4.141 21.05 4.278 ;
      RECT 20.936 4.132 20.975 4.267 ;
      RECT 20.85 4.122 20.936 4.255 ;
      RECT 20.81 4.112 20.85 4.243 ;
      RECT 20.771 4.107 20.81 4.236 ;
      RECT 20.685 4.097 20.771 4.225 ;
      RECT 20.645 4.085 20.685 4.214 ;
      RECT 20.61 4.07 20.645 4.207 ;
      RECT 20.6 4.06 20.61 4.204 ;
      RECT 20.58 4.045 20.6 4.202 ;
      RECT 20.55 4.015 20.58 4.198 ;
      RECT 20.54 3.995 20.55 4.193 ;
      RECT 20.535 3.987 20.54 4.19 ;
      RECT 20.53 3.98 20.535 4.188 ;
      RECT 20.515 3.967 20.53 4.181 ;
      RECT 20.51 3.957 20.515 4.173 ;
      RECT 20.505 3.95 20.51 4.168 ;
      RECT 20.5 3.945 20.505 4.164 ;
      RECT 20.485 3.932 20.5 4.156 ;
      RECT 20.48 3.842 20.485 4.145 ;
      RECT 20.475 3.837 20.48 4.138 ;
      RECT 20.4 3.835 20.475 4.098 ;
      RECT 20.37 3.835 20.4 4.053 ;
      RECT 20.275 3.84 20.29 4.04 ;
      RECT 22.76 3.545 23.02 3.805 ;
      RECT 22.745 3.533 22.925 3.77 ;
      RECT 22.74 3.534 22.925 3.768 ;
      RECT 22.725 3.538 22.935 3.758 ;
      RECT 22.72 3.543 22.94 3.728 ;
      RECT 22.725 3.54 22.94 3.758 ;
      RECT 22.74 3.535 22.935 3.768 ;
      RECT 22.76 3.532 22.925 3.805 ;
      RECT 22.76 3.531 22.915 3.805 ;
      RECT 22.785 3.53 22.915 3.805 ;
      RECT 22.345 3.775 22.605 4.035 ;
      RECT 22.22 3.82 22.605 4.03 ;
      RECT 22.21 3.825 22.605 4.025 ;
      RECT 22.225 4.765 22.24 5.075 ;
      RECT 20.82 4.535 20.83 4.665 ;
      RECT 20.6 4.53 20.705 4.665 ;
      RECT 20.515 4.535 20.565 4.665 ;
      RECT 19.065 3.27 19.07 4.375 ;
      RECT 22.32 4.857 22.325 4.993 ;
      RECT 22.315 4.852 22.32 5.053 ;
      RECT 22.31 4.85 22.315 5.066 ;
      RECT 22.295 4.847 22.31 5.068 ;
      RECT 22.29 4.842 22.295 5.07 ;
      RECT 22.285 4.838 22.29 5.073 ;
      RECT 22.27 4.833 22.285 5.075 ;
      RECT 22.24 4.825 22.27 5.075 ;
      RECT 22.201 4.765 22.225 5.075 ;
      RECT 22.115 4.765 22.201 5.072 ;
      RECT 22.085 4.765 22.115 5.065 ;
      RECT 22.06 4.765 22.085 5.058 ;
      RECT 22.035 4.765 22.06 5.05 ;
      RECT 22.02 4.765 22.035 5.043 ;
      RECT 21.995 4.765 22.02 5.035 ;
      RECT 21.98 4.765 21.995 5.028 ;
      RECT 21.94 4.775 21.98 5.017 ;
      RECT 21.93 4.77 21.94 5.007 ;
      RECT 21.926 4.769 21.93 5.004 ;
      RECT 21.84 4.761 21.926 4.987 ;
      RECT 21.807 4.75 21.84 4.964 ;
      RECT 21.721 4.739 21.807 4.942 ;
      RECT 21.635 4.723 21.721 4.911 ;
      RECT 21.565 4.708 21.635 4.883 ;
      RECT 21.555 4.701 21.565 4.87 ;
      RECT 21.525 4.698 21.555 4.86 ;
      RECT 21.5 4.694 21.525 4.853 ;
      RECT 21.485 4.691 21.5 4.848 ;
      RECT 21.48 4.69 21.485 4.843 ;
      RECT 21.45 4.685 21.48 4.836 ;
      RECT 21.445 4.68 21.45 4.831 ;
      RECT 21.43 4.677 21.445 4.826 ;
      RECT 21.425 4.672 21.43 4.821 ;
      RECT 21.405 4.667 21.425 4.818 ;
      RECT 21.39 4.662 21.405 4.81 ;
      RECT 21.375 4.656 21.39 4.805 ;
      RECT 21.345 4.647 21.375 4.798 ;
      RECT 21.34 4.64 21.345 4.79 ;
      RECT 21.335 4.638 21.34 4.788 ;
      RECT 21.33 4.637 21.335 4.785 ;
      RECT 21.29 4.63 21.33 4.778 ;
      RECT 21.276 4.62 21.29 4.768 ;
      RECT 21.225 4.609 21.276 4.756 ;
      RECT 21.2 4.595 21.225 4.742 ;
      RECT 21.175 4.584 21.2 4.734 ;
      RECT 21.155 4.573 21.175 4.728 ;
      RECT 21.145 4.567 21.155 4.723 ;
      RECT 21.14 4.565 21.145 4.719 ;
      RECT 21.12 4.56 21.14 4.714 ;
      RECT 21.09 4.55 21.12 4.704 ;
      RECT 21.085 4.542 21.09 4.697 ;
      RECT 21.07 4.54 21.085 4.693 ;
      RECT 21.05 4.54 21.07 4.688 ;
      RECT 21.045 4.539 21.05 4.686 ;
      RECT 21.04 4.539 21.045 4.683 ;
      RECT 21 4.538 21.04 4.678 ;
      RECT 20.975 4.537 21 4.673 ;
      RECT 20.915 4.536 20.975 4.67 ;
      RECT 20.83 4.535 20.915 4.668 ;
      RECT 20.791 4.534 20.82 4.665 ;
      RECT 20.705 4.532 20.791 4.665 ;
      RECT 20.565 4.532 20.6 4.665 ;
      RECT 20.475 4.536 20.515 4.668 ;
      RECT 20.46 4.539 20.475 4.675 ;
      RECT 20.45 4.54 20.46 4.682 ;
      RECT 20.425 4.543 20.45 4.687 ;
      RECT 20.42 4.545 20.425 4.69 ;
      RECT 20.37 4.547 20.42 4.691 ;
      RECT 20.331 4.551 20.37 4.693 ;
      RECT 20.245 4.553 20.331 4.696 ;
      RECT 20.227 4.555 20.245 4.698 ;
      RECT 20.141 4.558 20.227 4.7 ;
      RECT 20.055 4.562 20.141 4.703 ;
      RECT 20.018 4.566 20.055 4.706 ;
      RECT 19.932 4.569 20.018 4.709 ;
      RECT 19.846 4.573 19.932 4.712 ;
      RECT 19.76 4.578 19.846 4.716 ;
      RECT 19.74 4.58 19.76 4.719 ;
      RECT 19.72 4.579 19.74 4.72 ;
      RECT 19.671 4.576 19.72 4.721 ;
      RECT 19.585 4.571 19.671 4.724 ;
      RECT 19.535 4.566 19.585 4.726 ;
      RECT 19.511 4.564 19.535 4.727 ;
      RECT 19.425 4.559 19.511 4.729 ;
      RECT 19.4 4.555 19.425 4.728 ;
      RECT 19.39 4.552 19.4 4.726 ;
      RECT 19.38 4.545 19.39 4.723 ;
      RECT 19.375 4.525 19.38 4.718 ;
      RECT 19.365 4.495 19.375 4.713 ;
      RECT 19.35 4.365 19.365 4.704 ;
      RECT 19.345 4.357 19.35 4.697 ;
      RECT 19.325 4.35 19.345 4.689 ;
      RECT 19.32 4.332 19.325 4.681 ;
      RECT 19.31 4.312 19.32 4.676 ;
      RECT 19.305 4.285 19.31 4.672 ;
      RECT 19.3 4.262 19.305 4.669 ;
      RECT 19.28 4.22 19.3 4.661 ;
      RECT 19.245 4.135 19.28 4.645 ;
      RECT 19.24 4.067 19.245 4.633 ;
      RECT 19.225 4.037 19.24 4.627 ;
      RECT 19.22 3.282 19.225 3.528 ;
      RECT 19.21 4.007 19.225 4.618 ;
      RECT 19.215 3.277 19.22 3.56 ;
      RECT 19.21 3.272 19.215 3.603 ;
      RECT 19.205 3.27 19.21 3.638 ;
      RECT 19.19 3.97 19.21 4.608 ;
      RECT 19.2 3.27 19.205 3.675 ;
      RECT 19.185 3.27 19.2 3.773 ;
      RECT 19.185 3.943 19.19 4.601 ;
      RECT 19.18 3.27 19.185 3.848 ;
      RECT 19.18 3.931 19.185 4.598 ;
      RECT 19.175 3.27 19.18 3.88 ;
      RECT 19.175 3.91 19.18 4.595 ;
      RECT 19.17 3.27 19.175 4.592 ;
      RECT 19.135 3.27 19.17 4.578 ;
      RECT 19.12 3.27 19.135 4.56 ;
      RECT 19.1 3.27 19.12 4.55 ;
      RECT 19.075 3.27 19.1 4.533 ;
      RECT 19.07 3.27 19.075 4.483 ;
      RECT 19.06 3.27 19.065 4.313 ;
      RECT 19.055 3.27 19.06 4.22 ;
      RECT 19.05 3.27 19.055 4.133 ;
      RECT 19.045 3.27 19.05 4.065 ;
      RECT 19.04 3.27 19.045 4.008 ;
      RECT 19.03 3.27 19.04 3.903 ;
      RECT 19.025 3.27 19.03 3.775 ;
      RECT 19.02 3.27 19.025 3.693 ;
      RECT 19.015 3.272 19.02 3.61 ;
      RECT 19.01 3.277 19.015 3.543 ;
      RECT 19.005 3.282 19.01 3.47 ;
      RECT 21.82 3.6 22.08 3.86 ;
      RECT 21.84 3.567 22.05 3.86 ;
      RECT 21.84 3.565 22.04 3.86 ;
      RECT 21.85 3.552 22.04 3.86 ;
      RECT 21.85 3.55 21.965 3.86 ;
      RECT 21.325 3.675 21.5 3.955 ;
      RECT 21.32 3.675 21.5 3.953 ;
      RECT 21.32 3.675 21.515 3.95 ;
      RECT 21.31 3.675 21.515 3.948 ;
      RECT 21.255 3.675 21.515 3.935 ;
      RECT 21.255 3.75 21.52 3.913 ;
      RECT 20.8 3.687 20.82 3.93 ;
      RECT 20.8 3.687 20.86 3.929 ;
      RECT 20.795 3.689 20.86 3.928 ;
      RECT 20.795 3.689 20.946 3.927 ;
      RECT 20.795 3.689 21.015 3.926 ;
      RECT 20.795 3.689 21.035 3.918 ;
      RECT 20.775 3.692 21.035 3.916 ;
      RECT 20.76 3.702 21.035 3.901 ;
      RECT 20.76 3.702 21.05 3.9 ;
      RECT 20.755 3.711 21.05 3.892 ;
      RECT 20.755 3.711 21.055 3.888 ;
      RECT 20.86 3.625 21.12 3.885 ;
      RECT 20.75 3.713 21.12 3.77 ;
      RECT 20.82 3.68 21.12 3.885 ;
      RECT 20.785 4.873 20.79 5.08 ;
      RECT 20.735 4.867 20.785 5.079 ;
      RECT 20.702 4.881 20.795 5.078 ;
      RECT 20.616 4.881 20.795 5.077 ;
      RECT 20.53 4.881 20.795 5.076 ;
      RECT 20.53 4.98 20.8 5.073 ;
      RECT 20.525 4.98 20.8 5.068 ;
      RECT 20.52 4.98 20.8 5.05 ;
      RECT 20.515 4.98 20.8 5.033 ;
      RECT 20.475 4.765 20.735 5.025 ;
      RECT 19.935 3.915 20.021 4.329 ;
      RECT 19.935 3.915 20.06 4.326 ;
      RECT 19.935 3.915 20.08 4.316 ;
      RECT 19.89 3.915 20.08 4.313 ;
      RECT 19.89 4.067 20.09 4.303 ;
      RECT 19.89 4.088 20.095 4.297 ;
      RECT 19.89 4.106 20.1 4.293 ;
      RECT 19.89 4.126 20.11 4.288 ;
      RECT 19.865 4.126 20.11 4.285 ;
      RECT 19.855 4.126 20.11 4.263 ;
      RECT 19.855 4.142 20.115 4.233 ;
      RECT 19.82 3.915 20.08 4.22 ;
      RECT 19.82 4.154 20.12 4.175 ;
      RECT 17.48 10.06 17.77 10.29 ;
      RECT 17.54 8.58 17.71 10.29 ;
      RECT 17.535 8.945 17.885 9.295 ;
      RECT 17.48 8.58 17.77 8.81 ;
      RECT 17.075 3.69 17.18 4.26 ;
      RECT 17.075 4.025 17.4 4.255 ;
      RECT 17.075 4.055 17.57 4.225 ;
      RECT 17.075 3.69 17.265 4.255 ;
      RECT 16.49 3.655 16.78 3.885 ;
      RECT 16.49 3.69 17.265 3.86 ;
      RECT 16.55 2.175 16.72 3.885 ;
      RECT 16.49 2.175 16.78 2.405 ;
      RECT 16.49 10.06 16.78 10.29 ;
      RECT 16.55 8.58 16.72 10.29 ;
      RECT 16.49 8.58 16.78 8.81 ;
      RECT 16.49 8.615 17.34 8.775 ;
      RECT 17.175 8.21 17.34 8.775 ;
      RECT 16.49 8.61 16.885 8.775 ;
      RECT 17.11 8.21 17.4 8.44 ;
      RECT 17.11 8.24 17.57 8.41 ;
      RECT 16.12 4.025 16.41 4.255 ;
      RECT 16.12 4.055 16.58 4.225 ;
      RECT 16.185 2.95 16.35 4.255 ;
      RECT 14.7 2.92 14.99 3.15 ;
      RECT 14.7 2.95 16.35 3.12 ;
      RECT 14.76 2.18 14.93 3.15 ;
      RECT 14.7 2.18 14.99 2.41 ;
      RECT 14.7 10.055 14.99 10.285 ;
      RECT 14.76 9.315 14.93 10.285 ;
      RECT 14.76 9.41 16.35 9.58 ;
      RECT 16.18 8.21 16.35 9.58 ;
      RECT 14.7 9.315 14.99 9.545 ;
      RECT 16.12 8.21 16.41 8.44 ;
      RECT 16.12 8.24 16.58 8.41 ;
      RECT 12.75 4 13.09 4.35 ;
      RECT 12.84 3.32 13.01 4.35 ;
      RECT 15.13 3.26 15.48 3.61 ;
      RECT 12.84 3.32 15.48 3.49 ;
      RECT 15.155 8.945 15.48 9.27 ;
      RECT 9.695 8.895 10.045 9.245 ;
      RECT 15.13 8.945 15.48 9.175 ;
      RECT 9.495 8.945 10.045 9.175 ;
      RECT 9.325 8.975 15.48 9.145 ;
      RECT 14.355 3.66 14.675 3.98 ;
      RECT 14.325 3.66 14.675 3.89 ;
      RECT 14.155 3.69 14.675 3.86 ;
      RECT 14.355 8.545 14.675 8.835 ;
      RECT 14.325 8.575 14.675 8.805 ;
      RECT 14.155 8.605 14.675 8.775 ;
      RECT 10.045 4.28 10.195 4.555 ;
      RECT 10.585 3.36 10.59 3.58 ;
      RECT 11.735 3.56 11.75 3.758 ;
      RECT 11.7 3.552 11.735 3.765 ;
      RECT 11.67 3.545 11.7 3.765 ;
      RECT 11.615 3.51 11.67 3.765 ;
      RECT 11.55 3.447 11.615 3.765 ;
      RECT 11.545 3.412 11.55 3.763 ;
      RECT 11.54 3.407 11.545 3.755 ;
      RECT 11.535 3.402 11.54 3.741 ;
      RECT 11.53 3.399 11.535 3.734 ;
      RECT 11.485 3.389 11.53 3.685 ;
      RECT 11.465 3.376 11.485 3.62 ;
      RECT 11.46 3.371 11.465 3.593 ;
      RECT 11.455 3.37 11.46 3.586 ;
      RECT 11.45 3.369 11.455 3.579 ;
      RECT 11.365 3.354 11.45 3.525 ;
      RECT 11.335 3.335 11.365 3.475 ;
      RECT 11.255 3.318 11.335 3.46 ;
      RECT 11.22 3.305 11.255 3.445 ;
      RECT 11.212 3.305 11.22 3.44 ;
      RECT 11.126 3.306 11.212 3.44 ;
      RECT 11.04 3.308 11.126 3.44 ;
      RECT 11.015 3.309 11.04 3.444 ;
      RECT 10.94 3.315 11.015 3.459 ;
      RECT 10.857 3.327 10.94 3.483 ;
      RECT 10.771 3.34 10.857 3.509 ;
      RECT 10.685 3.353 10.771 3.535 ;
      RECT 10.65 3.362 10.685 3.554 ;
      RECT 10.6 3.362 10.65 3.567 ;
      RECT 10.59 3.36 10.6 3.578 ;
      RECT 10.575 3.357 10.585 3.58 ;
      RECT 10.56 3.349 10.575 3.588 ;
      RECT 10.545 3.341 10.56 3.608 ;
      RECT 10.54 3.336 10.545 3.665 ;
      RECT 10.525 3.331 10.54 3.738 ;
      RECT 10.52 3.326 10.525 3.78 ;
      RECT 10.515 3.324 10.52 3.808 ;
      RECT 10.51 3.322 10.515 3.83 ;
      RECT 10.5 3.318 10.51 3.873 ;
      RECT 10.495 3.315 10.5 3.898 ;
      RECT 10.49 3.313 10.495 3.918 ;
      RECT 10.485 3.311 10.49 3.942 ;
      RECT 10.48 3.307 10.485 3.965 ;
      RECT 10.475 3.303 10.48 3.988 ;
      RECT 10.44 3.293 10.475 4.095 ;
      RECT 10.435 3.283 10.44 4.193 ;
      RECT 10.43 3.281 10.435 4.22 ;
      RECT 10.425 3.28 10.43 4.24 ;
      RECT 10.42 3.272 10.425 4.26 ;
      RECT 10.415 3.267 10.42 4.295 ;
      RECT 10.41 3.265 10.415 4.313 ;
      RECT 10.405 3.265 10.41 4.338 ;
      RECT 10.4 3.265 10.405 4.36 ;
      RECT 10.365 3.265 10.4 4.403 ;
      RECT 10.34 3.265 10.365 4.432 ;
      RECT 10.33 3.265 10.34 3.618 ;
      RECT 10.333 3.675 10.34 4.442 ;
      RECT 10.33 3.732 10.333 4.445 ;
      RECT 10.325 3.265 10.33 3.59 ;
      RECT 10.325 3.782 10.33 4.448 ;
      RECT 10.315 3.265 10.325 3.58 ;
      RECT 10.32 3.835 10.325 4.451 ;
      RECT 10.315 3.92 10.32 4.455 ;
      RECT 10.305 3.265 10.315 3.568 ;
      RECT 10.31 3.967 10.315 4.459 ;
      RECT 10.305 4.042 10.31 4.463 ;
      RECT 10.27 3.265 10.305 3.543 ;
      RECT 10.295 4.125 10.305 4.468 ;
      RECT 10.285 4.192 10.295 4.475 ;
      RECT 10.28 4.22 10.285 4.48 ;
      RECT 10.27 4.233 10.28 4.486 ;
      RECT 10.225 3.265 10.27 3.5 ;
      RECT 10.265 4.238 10.27 4.493 ;
      RECT 10.225 4.255 10.265 4.555 ;
      RECT 10.22 3.267 10.225 3.473 ;
      RECT 10.195 4.275 10.225 4.555 ;
      RECT 10.215 3.272 10.22 3.445 ;
      RECT 10.005 4.284 10.045 4.555 ;
      RECT 9.98 4.292 10.005 4.525 ;
      RECT 9.935 4.3 9.98 4.525 ;
      RECT 9.92 4.305 9.935 4.52 ;
      RECT 9.91 4.305 9.92 4.514 ;
      RECT 9.9 4.312 9.91 4.511 ;
      RECT 9.895 4.35 9.9 4.5 ;
      RECT 9.89 4.412 9.895 4.478 ;
      RECT 11.16 4.287 11.345 4.51 ;
      RECT 11.16 4.302 11.35 4.506 ;
      RECT 11.15 3.575 11.235 4.505 ;
      RECT 11.15 4.302 11.355 4.499 ;
      RECT 11.145 4.31 11.355 4.498 ;
      RECT 11.35 4.03 11.67 4.35 ;
      RECT 11.145 4.202 11.315 4.293 ;
      RECT 11.14 4.202 11.315 4.275 ;
      RECT 11.13 4.01 11.265 4.25 ;
      RECT 11.125 4.01 11.265 4.195 ;
      RECT 11.085 3.59 11.255 4.095 ;
      RECT 11.07 3.59 11.255 3.965 ;
      RECT 11.065 3.59 11.255 3.918 ;
      RECT 11.06 3.59 11.255 3.898 ;
      RECT 11.055 3.59 11.255 3.873 ;
      RECT 11.025 3.59 11.285 3.85 ;
      RECT 11.035 3.587 11.245 3.85 ;
      RECT 11.16 3.582 11.245 4.51 ;
      RECT 11.045 3.575 11.235 3.85 ;
      RECT 11.04 3.58 11.235 3.85 ;
      RECT 9.87 3.792 10.055 4.005 ;
      RECT 9.87 3.8 10.065 3.998 ;
      RECT 9.85 3.8 10.065 3.995 ;
      RECT 9.845 3.8 10.065 3.98 ;
      RECT 9.775 3.715 10.035 3.975 ;
      RECT 9.775 3.86 10.07 3.888 ;
      RECT 9.43 4.315 9.69 4.575 ;
      RECT 9.455 4.26 9.65 4.575 ;
      RECT 9.45 4.009 9.63 4.303 ;
      RECT 9.45 4.015 9.64 4.303 ;
      RECT 9.43 4.017 9.64 4.248 ;
      RECT 9.425 4.027 9.64 4.115 ;
      RECT 9.455 4.007 9.63 4.575 ;
      RECT 9.541 4.005 9.63 4.575 ;
      RECT 9.4 3.225 9.435 3.595 ;
      RECT 9.19 3.335 9.195 3.595 ;
      RECT 9.435 3.232 9.45 3.595 ;
      RECT 9.325 3.225 9.4 3.673 ;
      RECT 9.315 3.225 9.325 3.758 ;
      RECT 9.29 3.225 9.315 3.793 ;
      RECT 9.25 3.225 9.29 3.861 ;
      RECT 9.24 3.232 9.25 3.913 ;
      RECT 9.21 3.335 9.24 3.954 ;
      RECT 9.205 3.335 9.21 3.993 ;
      RECT 9.195 3.335 9.205 4.013 ;
      RECT 9.19 3.63 9.195 4.05 ;
      RECT 9.185 3.647 9.19 4.07 ;
      RECT 9.17 3.71 9.185 4.11 ;
      RECT 9.165 3.753 9.17 4.145 ;
      RECT 9.16 3.761 9.165 4.158 ;
      RECT 9.15 3.775 9.16 4.18 ;
      RECT 9.125 3.81 9.15 4.245 ;
      RECT 9.115 3.845 9.125 4.308 ;
      RECT 9.095 3.875 9.115 4.369 ;
      RECT 9.08 3.911 9.095 4.436 ;
      RECT 9.07 3.939 9.08 4.475 ;
      RECT 9.06 3.961 9.07 4.495 ;
      RECT 9.055 3.971 9.06 4.506 ;
      RECT 9.05 3.98 9.055 4.509 ;
      RECT 9.04 3.998 9.05 4.513 ;
      RECT 9.03 4.016 9.04 4.514 ;
      RECT 9.005 4.055 9.03 4.511 ;
      RECT 8.985 4.097 9.005 4.508 ;
      RECT 8.97 4.135 8.985 4.507 ;
      RECT 8.935 4.17 8.97 4.504 ;
      RECT 8.93 4.192 8.935 4.502 ;
      RECT 8.865 4.232 8.93 4.499 ;
      RECT 8.86 4.272 8.865 4.495 ;
      RECT 8.845 4.282 8.86 4.486 ;
      RECT 8.835 4.402 8.845 4.471 ;
      RECT 9.315 4.815 9.325 5.075 ;
      RECT 9.315 4.818 9.335 5.074 ;
      RECT 9.305 4.808 9.315 5.073 ;
      RECT 9.295 4.823 9.375 5.069 ;
      RECT 9.28 4.802 9.295 5.067 ;
      RECT 9.255 4.827 9.38 5.063 ;
      RECT 9.24 4.787 9.255 5.058 ;
      RECT 9.24 4.829 9.39 5.057 ;
      RECT 9.24 4.837 9.405 5.05 ;
      RECT 9.18 4.774 9.24 5.04 ;
      RECT 9.17 4.761 9.18 5.022 ;
      RECT 9.145 4.751 9.17 5.012 ;
      RECT 9.14 4.741 9.145 5.004 ;
      RECT 9.075 4.837 9.405 4.986 ;
      RECT 8.99 4.837 9.405 4.948 ;
      RECT 8.88 4.665 9.14 4.925 ;
      RECT 9.255 4.795 9.28 5.063 ;
      RECT 9.295 4.805 9.305 5.069 ;
      RECT 8.88 4.813 9.32 4.925 ;
      RECT 9.065 10.055 9.355 10.285 ;
      RECT 9.125 9.315 9.295 10.285 ;
      RECT 9.025 9.345 9.395 9.715 ;
      RECT 9.065 9.315 9.355 9.715 ;
      RECT 8.095 4.57 8.125 4.87 ;
      RECT 7.87 4.555 7.875 4.83 ;
      RECT 7.67 4.555 7.825 4.815 ;
      RECT 8.97 3.27 9 3.53 ;
      RECT 8.96 3.27 8.97 3.638 ;
      RECT 8.94 3.27 8.96 3.648 ;
      RECT 8.925 3.27 8.94 3.66 ;
      RECT 8.87 3.27 8.925 3.71 ;
      RECT 8.855 3.27 8.87 3.758 ;
      RECT 8.825 3.27 8.855 3.793 ;
      RECT 8.77 3.27 8.825 3.855 ;
      RECT 8.75 3.27 8.77 3.923 ;
      RECT 8.745 3.27 8.75 3.953 ;
      RECT 8.74 3.27 8.745 3.965 ;
      RECT 8.735 3.387 8.74 3.983 ;
      RECT 8.715 3.405 8.735 4.008 ;
      RECT 8.695 3.432 8.715 4.058 ;
      RECT 8.69 3.452 8.695 4.089 ;
      RECT 8.685 3.46 8.69 4.106 ;
      RECT 8.67 3.486 8.685 4.135 ;
      RECT 8.655 3.528 8.67 4.17 ;
      RECT 8.65 3.557 8.655 4.193 ;
      RECT 8.645 3.572 8.65 4.206 ;
      RECT 8.64 3.595 8.645 4.217 ;
      RECT 8.63 3.615 8.64 4.235 ;
      RECT 8.62 3.645 8.63 4.258 ;
      RECT 8.615 3.667 8.62 4.278 ;
      RECT 8.61 3.682 8.615 4.293 ;
      RECT 8.595 3.712 8.61 4.32 ;
      RECT 8.59 3.742 8.595 4.346 ;
      RECT 8.585 3.76 8.59 4.358 ;
      RECT 8.575 3.79 8.585 4.377 ;
      RECT 8.565 3.815 8.575 4.402 ;
      RECT 8.56 3.835 8.565 4.421 ;
      RECT 8.555 3.852 8.56 4.434 ;
      RECT 8.545 3.878 8.555 4.453 ;
      RECT 8.535 3.916 8.545 4.48 ;
      RECT 8.53 3.942 8.535 4.5 ;
      RECT 8.525 3.952 8.53 4.51 ;
      RECT 8.52 3.965 8.525 4.525 ;
      RECT 8.515 3.98 8.52 4.535 ;
      RECT 8.51 4.002 8.515 4.55 ;
      RECT 8.505 4.02 8.51 4.561 ;
      RECT 8.5 4.03 8.505 4.572 ;
      RECT 8.495 4.038 8.5 4.584 ;
      RECT 8.49 4.046 8.495 4.595 ;
      RECT 8.485 4.072 8.49 4.608 ;
      RECT 8.475 4.1 8.485 4.621 ;
      RECT 8.47 4.13 8.475 4.63 ;
      RECT 8.465 4.145 8.47 4.637 ;
      RECT 8.45 4.17 8.465 4.644 ;
      RECT 8.445 4.192 8.45 4.65 ;
      RECT 8.44 4.217 8.445 4.653 ;
      RECT 8.431 4.245 8.44 4.657 ;
      RECT 8.425 4.262 8.431 4.662 ;
      RECT 8.42 4.28 8.425 4.666 ;
      RECT 8.415 4.292 8.42 4.669 ;
      RECT 8.41 4.313 8.415 4.673 ;
      RECT 8.405 4.331 8.41 4.676 ;
      RECT 8.4 4.345 8.405 4.679 ;
      RECT 8.395 4.362 8.4 4.682 ;
      RECT 8.39 4.375 8.395 4.685 ;
      RECT 8.365 4.412 8.39 4.693 ;
      RECT 8.36 4.457 8.365 4.702 ;
      RECT 8.355 4.485 8.36 4.705 ;
      RECT 8.345 4.505 8.355 4.709 ;
      RECT 8.34 4.525 8.345 4.714 ;
      RECT 8.335 4.54 8.34 4.717 ;
      RECT 8.315 4.55 8.335 4.724 ;
      RECT 8.25 4.557 8.315 4.75 ;
      RECT 8.215 4.56 8.25 4.778 ;
      RECT 8.2 4.563 8.215 4.793 ;
      RECT 8.19 4.564 8.2 4.808 ;
      RECT 8.18 4.565 8.19 4.825 ;
      RECT 8.175 4.565 8.18 4.84 ;
      RECT 8.17 4.565 8.175 4.848 ;
      RECT 8.155 4.566 8.17 4.863 ;
      RECT 8.125 4.568 8.155 4.87 ;
      RECT 8.015 4.575 8.095 4.87 ;
      RECT 7.97 4.58 8.015 4.87 ;
      RECT 7.96 4.581 7.97 4.86 ;
      RECT 7.95 4.582 7.96 4.853 ;
      RECT 7.93 4.584 7.95 4.848 ;
      RECT 7.92 4.555 7.93 4.843 ;
      RECT 7.875 4.555 7.92 4.835 ;
      RECT 7.845 4.555 7.87 4.825 ;
      RECT 7.825 4.555 7.845 4.818 ;
      RECT 8.105 3.355 8.365 3.615 ;
      RECT 7.985 3.37 7.995 3.535 ;
      RECT 7.97 3.37 7.975 3.53 ;
      RECT 5.335 3.21 5.52 3.5 ;
      RECT 7.15 3.335 7.165 3.49 ;
      RECT 5.3 3.21 5.325 3.47 ;
      RECT 7.715 3.26 7.72 3.402 ;
      RECT 7.63 3.255 7.655 3.395 ;
      RECT 8.03 3.372 8.105 3.565 ;
      RECT 8.015 3.37 8.03 3.548 ;
      RECT 7.995 3.37 8.015 3.54 ;
      RECT 7.975 3.37 7.985 3.533 ;
      RECT 7.93 3.365 7.97 3.523 ;
      RECT 7.89 3.34 7.93 3.508 ;
      RECT 7.875 3.315 7.89 3.498 ;
      RECT 7.87 3.309 7.875 3.496 ;
      RECT 7.835 3.301 7.87 3.479 ;
      RECT 7.83 3.294 7.835 3.467 ;
      RECT 7.81 3.289 7.83 3.455 ;
      RECT 7.8 3.283 7.81 3.44 ;
      RECT 7.78 3.278 7.8 3.425 ;
      RECT 7.77 3.273 7.78 3.418 ;
      RECT 7.765 3.271 7.77 3.413 ;
      RECT 7.76 3.27 7.765 3.41 ;
      RECT 7.72 3.265 7.76 3.406 ;
      RECT 7.7 3.259 7.715 3.401 ;
      RECT 7.665 3.256 7.7 3.398 ;
      RECT 7.655 3.255 7.665 3.396 ;
      RECT 7.595 3.255 7.63 3.393 ;
      RECT 7.55 3.255 7.595 3.393 ;
      RECT 7.5 3.255 7.55 3.396 ;
      RECT 7.485 3.257 7.5 3.398 ;
      RECT 7.47 3.26 7.485 3.399 ;
      RECT 7.46 3.265 7.47 3.4 ;
      RECT 7.43 3.27 7.46 3.405 ;
      RECT 7.42 3.276 7.43 3.413 ;
      RECT 7.41 3.278 7.42 3.417 ;
      RECT 7.4 3.282 7.41 3.421 ;
      RECT 7.375 3.288 7.4 3.429 ;
      RECT 7.365 3.293 7.375 3.437 ;
      RECT 7.35 3.297 7.365 3.441 ;
      RECT 7.315 3.303 7.35 3.449 ;
      RECT 7.295 3.308 7.315 3.459 ;
      RECT 7.265 3.315 7.295 3.468 ;
      RECT 7.22 3.324 7.265 3.482 ;
      RECT 7.215 3.329 7.22 3.493 ;
      RECT 7.195 3.332 7.215 3.494 ;
      RECT 7.165 3.335 7.195 3.492 ;
      RECT 7.13 3.335 7.15 3.488 ;
      RECT 7.06 3.335 7.13 3.479 ;
      RECT 7.045 3.332 7.06 3.471 ;
      RECT 7.005 3.325 7.045 3.466 ;
      RECT 6.98 3.315 7.005 3.459 ;
      RECT 6.975 3.309 6.98 3.456 ;
      RECT 6.935 3.303 6.975 3.453 ;
      RECT 6.92 3.296 6.935 3.448 ;
      RECT 6.9 3.292 6.92 3.443 ;
      RECT 6.885 3.287 6.9 3.439 ;
      RECT 6.87 3.282 6.885 3.437 ;
      RECT 6.855 3.278 6.87 3.436 ;
      RECT 6.84 3.276 6.855 3.432 ;
      RECT 6.83 3.274 6.84 3.427 ;
      RECT 6.815 3.271 6.83 3.423 ;
      RECT 6.805 3.269 6.815 3.418 ;
      RECT 6.785 3.266 6.805 3.414 ;
      RECT 6.74 3.265 6.785 3.412 ;
      RECT 6.68 3.267 6.74 3.413 ;
      RECT 6.66 3.269 6.68 3.415 ;
      RECT 6.63 3.272 6.66 3.416 ;
      RECT 6.58 3.277 6.63 3.418 ;
      RECT 6.575 3.28 6.58 3.42 ;
      RECT 6.565 3.282 6.575 3.423 ;
      RECT 6.56 3.284 6.565 3.426 ;
      RECT 6.51 3.287 6.56 3.433 ;
      RECT 6.49 3.291 6.51 3.445 ;
      RECT 6.48 3.294 6.49 3.451 ;
      RECT 6.47 3.295 6.48 3.454 ;
      RECT 6.431 3.298 6.47 3.456 ;
      RECT 6.345 3.305 6.431 3.459 ;
      RECT 6.271 3.315 6.345 3.463 ;
      RECT 6.185 3.326 6.271 3.468 ;
      RECT 6.17 3.333 6.185 3.47 ;
      RECT 6.115 3.337 6.17 3.471 ;
      RECT 6.101 3.34 6.115 3.473 ;
      RECT 6.015 3.34 6.101 3.475 ;
      RECT 5.975 3.337 6.015 3.478 ;
      RECT 5.951 3.333 5.975 3.48 ;
      RECT 5.865 3.323 5.951 3.483 ;
      RECT 5.835 3.312 5.865 3.484 ;
      RECT 5.816 3.308 5.835 3.483 ;
      RECT 5.73 3.301 5.816 3.48 ;
      RECT 5.67 3.29 5.73 3.477 ;
      RECT 5.65 3.282 5.67 3.475 ;
      RECT 5.615 3.277 5.65 3.474 ;
      RECT 5.59 3.272 5.615 3.473 ;
      RECT 5.56 3.267 5.59 3.472 ;
      RECT 5.535 3.21 5.56 3.471 ;
      RECT 5.52 3.21 5.535 3.495 ;
      RECT 5.325 3.21 5.335 3.495 ;
      RECT 7.1 4.23 7.105 4.37 ;
      RECT 6.76 4.23 6.795 4.368 ;
      RECT 6.335 4.215 6.35 4.36 ;
      RECT 8.165 3.995 8.255 4.255 ;
      RECT 7.995 3.86 8.095 4.255 ;
      RECT 5.03 3.835 5.11 4.045 ;
      RECT 8.12 3.972 8.165 4.255 ;
      RECT 8.11 3.942 8.12 4.255 ;
      RECT 8.095 3.865 8.11 4.255 ;
      RECT 7.91 3.86 7.995 4.22 ;
      RECT 7.905 3.862 7.91 4.215 ;
      RECT 7.9 3.867 7.905 4.215 ;
      RECT 7.865 3.967 7.9 4.215 ;
      RECT 7.855 3.995 7.865 4.215 ;
      RECT 7.845 4.01 7.855 4.215 ;
      RECT 7.835 4.022 7.845 4.215 ;
      RECT 7.83 4.032 7.835 4.215 ;
      RECT 7.815 4.042 7.83 4.217 ;
      RECT 7.81 4.057 7.815 4.219 ;
      RECT 7.795 4.07 7.81 4.221 ;
      RECT 7.79 4.085 7.795 4.224 ;
      RECT 7.77 4.095 7.79 4.228 ;
      RECT 7.755 4.105 7.77 4.231 ;
      RECT 7.72 4.112 7.755 4.236 ;
      RECT 7.676 4.119 7.72 4.244 ;
      RECT 7.59 4.131 7.676 4.257 ;
      RECT 7.565 4.142 7.59 4.268 ;
      RECT 7.535 4.147 7.565 4.273 ;
      RECT 7.5 4.152 7.535 4.281 ;
      RECT 7.47 4.157 7.5 4.288 ;
      RECT 7.445 4.162 7.47 4.293 ;
      RECT 7.38 4.169 7.445 4.302 ;
      RECT 7.31 4.182 7.38 4.318 ;
      RECT 7.28 4.192 7.31 4.33 ;
      RECT 7.255 4.197 7.28 4.337 ;
      RECT 7.2 4.204 7.255 4.345 ;
      RECT 7.195 4.211 7.2 4.35 ;
      RECT 7.19 4.213 7.195 4.351 ;
      RECT 7.175 4.215 7.19 4.353 ;
      RECT 7.17 4.215 7.175 4.356 ;
      RECT 7.105 4.222 7.17 4.363 ;
      RECT 7.07 4.232 7.1 4.373 ;
      RECT 7.053 4.235 7.07 4.375 ;
      RECT 6.967 4.234 7.053 4.374 ;
      RECT 6.881 4.232 6.967 4.371 ;
      RECT 6.795 4.231 6.881 4.369 ;
      RECT 6.694 4.229 6.76 4.368 ;
      RECT 6.608 4.226 6.694 4.366 ;
      RECT 6.522 4.222 6.608 4.364 ;
      RECT 6.436 4.219 6.522 4.363 ;
      RECT 6.35 4.216 6.436 4.361 ;
      RECT 6.25 4.215 6.335 4.358 ;
      RECT 6.2 4.213 6.25 4.356 ;
      RECT 6.18 4.21 6.2 4.354 ;
      RECT 6.16 4.208 6.18 4.351 ;
      RECT 6.135 4.204 6.16 4.348 ;
      RECT 6.09 4.198 6.135 4.343 ;
      RECT 6.05 4.192 6.09 4.335 ;
      RECT 6.025 4.187 6.05 4.328 ;
      RECT 5.97 4.18 6.025 4.32 ;
      RECT 5.946 4.173 5.97 4.313 ;
      RECT 5.86 4.164 5.946 4.303 ;
      RECT 5.83 4.156 5.86 4.293 ;
      RECT 5.8 4.152 5.83 4.288 ;
      RECT 5.795 4.149 5.8 4.285 ;
      RECT 5.79 4.148 5.795 4.285 ;
      RECT 5.715 4.141 5.79 4.278 ;
      RECT 5.676 4.132 5.715 4.267 ;
      RECT 5.59 4.122 5.676 4.255 ;
      RECT 5.55 4.112 5.59 4.243 ;
      RECT 5.511 4.107 5.55 4.236 ;
      RECT 5.425 4.097 5.511 4.225 ;
      RECT 5.385 4.085 5.425 4.214 ;
      RECT 5.35 4.07 5.385 4.207 ;
      RECT 5.34 4.06 5.35 4.204 ;
      RECT 5.32 4.045 5.34 4.202 ;
      RECT 5.29 4.015 5.32 4.198 ;
      RECT 5.28 3.995 5.29 4.193 ;
      RECT 5.275 3.987 5.28 4.19 ;
      RECT 5.27 3.98 5.275 4.188 ;
      RECT 5.255 3.967 5.27 4.181 ;
      RECT 5.25 3.957 5.255 4.173 ;
      RECT 5.245 3.95 5.25 4.168 ;
      RECT 5.24 3.945 5.245 4.164 ;
      RECT 5.225 3.932 5.24 4.156 ;
      RECT 5.22 3.842 5.225 4.145 ;
      RECT 5.215 3.837 5.22 4.138 ;
      RECT 5.14 3.835 5.215 4.098 ;
      RECT 5.11 3.835 5.14 4.053 ;
      RECT 5.015 3.84 5.03 4.04 ;
      RECT 7.5 3.545 7.76 3.805 ;
      RECT 7.485 3.533 7.665 3.77 ;
      RECT 7.48 3.534 7.665 3.768 ;
      RECT 7.465 3.538 7.675 3.758 ;
      RECT 7.46 3.543 7.68 3.728 ;
      RECT 7.465 3.54 7.68 3.758 ;
      RECT 7.48 3.535 7.675 3.768 ;
      RECT 7.5 3.532 7.665 3.805 ;
      RECT 7.5 3.531 7.655 3.805 ;
      RECT 7.525 3.53 7.655 3.805 ;
      RECT 7.085 3.775 7.345 4.035 ;
      RECT 6.96 3.82 7.345 4.03 ;
      RECT 6.95 3.825 7.345 4.025 ;
      RECT 6.965 4.765 6.98 5.075 ;
      RECT 5.56 4.535 5.57 4.665 ;
      RECT 5.34 4.53 5.445 4.665 ;
      RECT 5.255 4.535 5.305 4.665 ;
      RECT 3.805 3.27 3.81 4.375 ;
      RECT 7.06 4.857 7.065 4.993 ;
      RECT 7.055 4.852 7.06 5.053 ;
      RECT 7.05 4.85 7.055 5.066 ;
      RECT 7.035 4.847 7.05 5.068 ;
      RECT 7.03 4.842 7.035 5.07 ;
      RECT 7.025 4.838 7.03 5.073 ;
      RECT 7.01 4.833 7.025 5.075 ;
      RECT 6.98 4.825 7.01 5.075 ;
      RECT 6.941 4.765 6.965 5.075 ;
      RECT 6.855 4.765 6.941 5.072 ;
      RECT 6.825 4.765 6.855 5.065 ;
      RECT 6.8 4.765 6.825 5.058 ;
      RECT 6.775 4.765 6.8 5.05 ;
      RECT 6.76 4.765 6.775 5.043 ;
      RECT 6.735 4.765 6.76 5.035 ;
      RECT 6.72 4.765 6.735 5.028 ;
      RECT 6.68 4.775 6.72 5.017 ;
      RECT 6.67 4.77 6.68 5.007 ;
      RECT 6.666 4.769 6.67 5.004 ;
      RECT 6.58 4.761 6.666 4.987 ;
      RECT 6.547 4.75 6.58 4.964 ;
      RECT 6.461 4.739 6.547 4.942 ;
      RECT 6.375 4.723 6.461 4.911 ;
      RECT 6.305 4.708 6.375 4.883 ;
      RECT 6.295 4.701 6.305 4.87 ;
      RECT 6.265 4.698 6.295 4.86 ;
      RECT 6.24 4.694 6.265 4.853 ;
      RECT 6.225 4.691 6.24 4.848 ;
      RECT 6.22 4.69 6.225 4.843 ;
      RECT 6.19 4.685 6.22 4.836 ;
      RECT 6.185 4.68 6.19 4.831 ;
      RECT 6.17 4.677 6.185 4.826 ;
      RECT 6.165 4.672 6.17 4.821 ;
      RECT 6.145 4.667 6.165 4.818 ;
      RECT 6.13 4.662 6.145 4.81 ;
      RECT 6.115 4.656 6.13 4.805 ;
      RECT 6.085 4.647 6.115 4.798 ;
      RECT 6.08 4.64 6.085 4.79 ;
      RECT 6.075 4.638 6.08 4.788 ;
      RECT 6.07 4.637 6.075 4.785 ;
      RECT 6.03 4.63 6.07 4.778 ;
      RECT 6.016 4.62 6.03 4.768 ;
      RECT 5.965 4.609 6.016 4.756 ;
      RECT 5.94 4.595 5.965 4.742 ;
      RECT 5.915 4.584 5.94 4.734 ;
      RECT 5.895 4.573 5.915 4.728 ;
      RECT 5.885 4.567 5.895 4.723 ;
      RECT 5.88 4.565 5.885 4.719 ;
      RECT 5.86 4.56 5.88 4.714 ;
      RECT 5.83 4.55 5.86 4.704 ;
      RECT 5.825 4.542 5.83 4.697 ;
      RECT 5.81 4.54 5.825 4.693 ;
      RECT 5.79 4.54 5.81 4.688 ;
      RECT 5.785 4.539 5.79 4.686 ;
      RECT 5.78 4.539 5.785 4.683 ;
      RECT 5.74 4.538 5.78 4.678 ;
      RECT 5.715 4.537 5.74 4.673 ;
      RECT 5.655 4.536 5.715 4.67 ;
      RECT 5.57 4.535 5.655 4.668 ;
      RECT 5.531 4.534 5.56 4.665 ;
      RECT 5.445 4.532 5.531 4.665 ;
      RECT 5.305 4.532 5.34 4.665 ;
      RECT 5.215 4.536 5.255 4.668 ;
      RECT 5.2 4.539 5.215 4.675 ;
      RECT 5.19 4.54 5.2 4.682 ;
      RECT 5.165 4.543 5.19 4.687 ;
      RECT 5.16 4.545 5.165 4.69 ;
      RECT 5.11 4.547 5.16 4.691 ;
      RECT 5.071 4.551 5.11 4.693 ;
      RECT 4.985 4.553 5.071 4.696 ;
      RECT 4.967 4.555 4.985 4.698 ;
      RECT 4.881 4.558 4.967 4.7 ;
      RECT 4.795 4.562 4.881 4.703 ;
      RECT 4.758 4.566 4.795 4.706 ;
      RECT 4.672 4.569 4.758 4.709 ;
      RECT 4.586 4.573 4.672 4.712 ;
      RECT 4.5 4.578 4.586 4.716 ;
      RECT 4.48 4.58 4.5 4.719 ;
      RECT 4.46 4.579 4.48 4.72 ;
      RECT 4.411 4.576 4.46 4.721 ;
      RECT 4.325 4.571 4.411 4.724 ;
      RECT 4.275 4.566 4.325 4.726 ;
      RECT 4.251 4.564 4.275 4.727 ;
      RECT 4.165 4.559 4.251 4.729 ;
      RECT 4.14 4.555 4.165 4.728 ;
      RECT 4.13 4.552 4.14 4.726 ;
      RECT 4.12 4.545 4.13 4.723 ;
      RECT 4.115 4.525 4.12 4.718 ;
      RECT 4.105 4.495 4.115 4.713 ;
      RECT 4.09 4.365 4.105 4.704 ;
      RECT 4.085 4.357 4.09 4.697 ;
      RECT 4.065 4.35 4.085 4.689 ;
      RECT 4.06 4.332 4.065 4.681 ;
      RECT 4.05 4.312 4.06 4.676 ;
      RECT 4.045 4.285 4.05 4.672 ;
      RECT 4.04 4.262 4.045 4.669 ;
      RECT 4.02 4.22 4.04 4.661 ;
      RECT 3.985 4.135 4.02 4.645 ;
      RECT 3.98 4.067 3.985 4.633 ;
      RECT 3.965 4.037 3.98 4.627 ;
      RECT 3.96 3.282 3.965 3.528 ;
      RECT 3.95 4.007 3.965 4.618 ;
      RECT 3.955 3.277 3.96 3.56 ;
      RECT 3.95 3.272 3.955 3.603 ;
      RECT 3.945 3.27 3.95 3.638 ;
      RECT 3.93 3.97 3.95 4.608 ;
      RECT 3.94 3.27 3.945 3.675 ;
      RECT 3.925 3.27 3.94 3.773 ;
      RECT 3.925 3.943 3.93 4.601 ;
      RECT 3.92 3.27 3.925 3.848 ;
      RECT 3.92 3.931 3.925 4.598 ;
      RECT 3.915 3.27 3.92 3.88 ;
      RECT 3.915 3.91 3.92 4.595 ;
      RECT 3.91 3.27 3.915 4.592 ;
      RECT 3.875 3.27 3.91 4.578 ;
      RECT 3.86 3.27 3.875 4.56 ;
      RECT 3.84 3.27 3.86 4.55 ;
      RECT 3.815 3.27 3.84 4.533 ;
      RECT 3.81 3.27 3.815 4.483 ;
      RECT 3.8 3.27 3.805 4.313 ;
      RECT 3.795 3.27 3.8 4.22 ;
      RECT 3.79 3.27 3.795 4.133 ;
      RECT 3.785 3.27 3.79 4.065 ;
      RECT 3.78 3.27 3.785 4.008 ;
      RECT 3.77 3.27 3.78 3.903 ;
      RECT 3.765 3.27 3.77 3.775 ;
      RECT 3.76 3.27 3.765 3.693 ;
      RECT 3.755 3.272 3.76 3.61 ;
      RECT 3.75 3.277 3.755 3.543 ;
      RECT 3.745 3.282 3.75 3.47 ;
      RECT 6.56 3.6 6.82 3.86 ;
      RECT 6.58 3.567 6.79 3.86 ;
      RECT 6.58 3.565 6.78 3.86 ;
      RECT 6.59 3.552 6.78 3.86 ;
      RECT 6.59 3.55 6.705 3.86 ;
      RECT 6.065 3.675 6.24 3.955 ;
      RECT 6.06 3.675 6.24 3.953 ;
      RECT 6.06 3.675 6.255 3.95 ;
      RECT 6.05 3.675 6.255 3.948 ;
      RECT 5.995 3.675 6.255 3.935 ;
      RECT 5.995 3.75 6.26 3.913 ;
      RECT 5.54 3.687 5.56 3.93 ;
      RECT 5.54 3.687 5.6 3.929 ;
      RECT 5.535 3.689 5.6 3.928 ;
      RECT 5.535 3.689 5.686 3.927 ;
      RECT 5.535 3.689 5.755 3.926 ;
      RECT 5.535 3.689 5.775 3.918 ;
      RECT 5.515 3.692 5.775 3.916 ;
      RECT 5.5 3.702 5.775 3.901 ;
      RECT 5.5 3.702 5.79 3.9 ;
      RECT 5.495 3.711 5.79 3.892 ;
      RECT 5.495 3.711 5.795 3.888 ;
      RECT 5.6 3.625 5.86 3.885 ;
      RECT 5.49 3.713 5.86 3.77 ;
      RECT 5.56 3.68 5.86 3.885 ;
      RECT 5.525 4.873 5.53 5.08 ;
      RECT 5.475 4.867 5.525 5.079 ;
      RECT 5.442 4.881 5.535 5.078 ;
      RECT 5.356 4.881 5.535 5.077 ;
      RECT 5.27 4.881 5.535 5.076 ;
      RECT 5.27 4.98 5.54 5.073 ;
      RECT 5.265 4.98 5.54 5.068 ;
      RECT 5.26 4.98 5.54 5.05 ;
      RECT 5.255 4.98 5.54 5.033 ;
      RECT 5.215 4.765 5.475 5.025 ;
      RECT 4.675 3.915 4.761 4.329 ;
      RECT 4.675 3.915 4.8 4.326 ;
      RECT 4.675 3.915 4.82 4.316 ;
      RECT 4.63 3.915 4.82 4.313 ;
      RECT 4.63 4.067 4.83 4.303 ;
      RECT 4.63 4.088 4.835 4.297 ;
      RECT 4.63 4.106 4.84 4.293 ;
      RECT 4.63 4.126 4.85 4.288 ;
      RECT 4.605 4.126 4.85 4.285 ;
      RECT 4.595 4.126 4.85 4.263 ;
      RECT 4.595 4.142 4.855 4.233 ;
      RECT 4.56 3.915 4.82 4.22 ;
      RECT 4.56 4.154 4.86 4.175 ;
      RECT 1.57 10.055 1.86 10.285 ;
      RECT 1.63 9.315 1.8 10.285 ;
      RECT 1.54 9.315 1.89 9.605 ;
      RECT 1.165 8.575 1.515 8.865 ;
      RECT 1.025 8.605 1.515 8.775 ;
      RECT 68.185 4.56 68.445 4.82 ;
      RECT 52.925 4.56 53.185 4.82 ;
      RECT 37.665 4.56 37.925 4.82 ;
      RECT 22.405 4.56 22.665 4.82 ;
      RECT 7.145 4.56 7.405 4.82 ;
    LAYER mcon ;
      RECT 78.58 8.61 78.75 8.78 ;
      RECT 78.58 10.09 78.75 10.26 ;
      RECT 78.23 1.395 78.4 1.565 ;
      RECT 78.21 4.055 78.38 4.225 ;
      RECT 78.21 8.24 78.38 8.41 ;
      RECT 77.59 2.205 77.76 2.375 ;
      RECT 77.59 3.685 77.76 3.855 ;
      RECT 77.59 8.61 77.76 8.78 ;
      RECT 77.59 10.09 77.76 10.26 ;
      RECT 77.24 1.395 77.41 1.565 ;
      RECT 77.22 4.055 77.39 4.225 ;
      RECT 77.22 8.24 77.39 8.41 ;
      RECT 76.54 1.4 76.71 1.57 ;
      RECT 76.23 3.32 76.4 3.49 ;
      RECT 76.23 8.975 76.4 9.145 ;
      RECT 75.86 1.4 76.03 1.57 ;
      RECT 75.8 2.21 75.97 2.38 ;
      RECT 75.8 2.95 75.97 3.12 ;
      RECT 75.8 9.345 75.97 9.515 ;
      RECT 75.8 10.085 75.97 10.255 ;
      RECT 75.425 3.69 75.595 3.86 ;
      RECT 75.425 8.605 75.595 8.775 ;
      RECT 75.18 1.4 75.35 1.57 ;
      RECT 74.5 1.4 74.67 1.57 ;
      RECT 73.04 2.71 73.21 2.88 ;
      RECT 72.6 3.575 72.77 3.745 ;
      RECT 72.58 2.71 72.75 2.88 ;
      RECT 72.205 4.32 72.375 4.49 ;
      RECT 72.12 2.71 72.29 2.88 ;
      RECT 72.095 3.595 72.265 3.765 ;
      RECT 71.66 2.71 71.83 2.88 ;
      RECT 71.275 3.285 71.445 3.455 ;
      RECT 71.2 2.71 71.37 2.88 ;
      RECT 70.96 4.325 71.13 4.495 ;
      RECT 70.915 3.815 71.085 3.985 ;
      RECT 70.74 2.71 70.91 2.88 ;
      RECT 70.595 8.975 70.765 9.145 ;
      RECT 70.49 4.025 70.66 4.195 ;
      RECT 70.3 3.245 70.47 3.415 ;
      RECT 70.28 2.71 70.45 2.88 ;
      RECT 70.25 4.855 70.42 5.025 ;
      RECT 70.165 9.345 70.335 9.515 ;
      RECT 70.165 10.085 70.335 10.255 ;
      RECT 69.915 4.295 70.085 4.465 ;
      RECT 69.82 2.71 69.99 2.88 ;
      RECT 69.82 3.455 69.99 3.625 ;
      RECT 69.36 2.71 69.53 2.88 ;
      RECT 69.02 4.68 69.19 4.85 ;
      RECT 68.96 3.88 69.13 4.05 ;
      RECT 68.9 2.71 69.07 2.88 ;
      RECT 68.52 3.55 68.69 3.72 ;
      RECT 68.44 2.71 68.61 2.88 ;
      RECT 68.255 4.6 68.425 4.77 ;
      RECT 68.01 3.84 68.18 4.01 ;
      RECT 67.98 2.71 68.15 2.88 ;
      RECT 67.915 4.87 68.085 5.04 ;
      RECT 67.64 3.565 67.81 3.735 ;
      RECT 67.52 2.71 67.69 2.88 ;
      RECT 67.11 3.765 67.28 3.935 ;
      RECT 67.06 2.71 67.23 2.88 ;
      RECT 66.6 2.71 66.77 2.88 ;
      RECT 66.59 3.71 66.76 3.88 ;
      RECT 66.385 3.31 66.555 3.48 ;
      RECT 66.385 4.89 66.555 5.06 ;
      RECT 66.14 2.71 66.31 2.88 ;
      RECT 66.075 3.855 66.245 4.025 ;
      RECT 65.68 2.71 65.85 2.88 ;
      RECT 65.665 4.08 65.835 4.25 ;
      RECT 65.22 2.71 65.39 2.88 ;
      RECT 64.955 4.38 65.125 4.55 ;
      RECT 64.81 3.29 64.98 3.46 ;
      RECT 64.76 2.71 64.93 2.88 ;
      RECT 63.32 8.61 63.49 8.78 ;
      RECT 63.32 10.09 63.49 10.26 ;
      RECT 62.97 1.395 63.14 1.565 ;
      RECT 62.95 4.055 63.12 4.225 ;
      RECT 62.95 8.24 63.12 8.41 ;
      RECT 62.33 2.205 62.5 2.375 ;
      RECT 62.33 3.685 62.5 3.855 ;
      RECT 62.33 8.61 62.5 8.78 ;
      RECT 62.33 10.09 62.5 10.26 ;
      RECT 61.98 1.395 62.15 1.565 ;
      RECT 61.96 4.055 62.13 4.225 ;
      RECT 61.96 8.24 62.13 8.41 ;
      RECT 61.28 1.4 61.45 1.57 ;
      RECT 60.97 3.32 61.14 3.49 ;
      RECT 60.97 8.975 61.14 9.145 ;
      RECT 60.6 1.4 60.77 1.57 ;
      RECT 60.54 2.21 60.71 2.38 ;
      RECT 60.54 2.95 60.71 3.12 ;
      RECT 60.54 9.345 60.71 9.515 ;
      RECT 60.54 10.085 60.71 10.255 ;
      RECT 60.165 3.69 60.335 3.86 ;
      RECT 60.165 8.605 60.335 8.775 ;
      RECT 59.92 1.4 60.09 1.57 ;
      RECT 59.24 1.4 59.41 1.57 ;
      RECT 57.78 2.71 57.95 2.88 ;
      RECT 57.34 3.575 57.51 3.745 ;
      RECT 57.32 2.71 57.49 2.88 ;
      RECT 56.945 4.32 57.115 4.49 ;
      RECT 56.86 2.71 57.03 2.88 ;
      RECT 56.835 3.595 57.005 3.765 ;
      RECT 56.4 2.71 56.57 2.88 ;
      RECT 56.015 3.285 56.185 3.455 ;
      RECT 55.94 2.71 56.11 2.88 ;
      RECT 55.7 4.325 55.87 4.495 ;
      RECT 55.655 3.815 55.825 3.985 ;
      RECT 55.48 2.71 55.65 2.88 ;
      RECT 55.335 8.975 55.505 9.145 ;
      RECT 55.23 4.025 55.4 4.195 ;
      RECT 55.04 3.245 55.21 3.415 ;
      RECT 55.02 2.71 55.19 2.88 ;
      RECT 54.99 4.855 55.16 5.025 ;
      RECT 54.905 9.345 55.075 9.515 ;
      RECT 54.905 10.085 55.075 10.255 ;
      RECT 54.655 4.295 54.825 4.465 ;
      RECT 54.56 2.71 54.73 2.88 ;
      RECT 54.56 3.455 54.73 3.625 ;
      RECT 54.1 2.71 54.27 2.88 ;
      RECT 53.76 4.68 53.93 4.85 ;
      RECT 53.7 3.88 53.87 4.05 ;
      RECT 53.64 2.71 53.81 2.88 ;
      RECT 53.26 3.55 53.43 3.72 ;
      RECT 53.18 2.71 53.35 2.88 ;
      RECT 52.995 4.6 53.165 4.77 ;
      RECT 52.75 3.84 52.92 4.01 ;
      RECT 52.72 2.71 52.89 2.88 ;
      RECT 52.655 4.87 52.825 5.04 ;
      RECT 52.38 3.565 52.55 3.735 ;
      RECT 52.26 2.71 52.43 2.88 ;
      RECT 51.85 3.765 52.02 3.935 ;
      RECT 51.8 2.71 51.97 2.88 ;
      RECT 51.34 2.71 51.51 2.88 ;
      RECT 51.33 3.71 51.5 3.88 ;
      RECT 51.125 3.31 51.295 3.48 ;
      RECT 51.125 4.89 51.295 5.06 ;
      RECT 50.88 2.71 51.05 2.88 ;
      RECT 50.815 3.855 50.985 4.025 ;
      RECT 50.42 2.71 50.59 2.88 ;
      RECT 50.405 4.08 50.575 4.25 ;
      RECT 49.96 2.71 50.13 2.88 ;
      RECT 49.695 4.38 49.865 4.55 ;
      RECT 49.55 3.29 49.72 3.46 ;
      RECT 49.5 2.71 49.67 2.88 ;
      RECT 48.06 8.61 48.23 8.78 ;
      RECT 48.06 10.09 48.23 10.26 ;
      RECT 47.71 1.395 47.88 1.565 ;
      RECT 47.69 4.055 47.86 4.225 ;
      RECT 47.69 8.24 47.86 8.41 ;
      RECT 47.07 2.205 47.24 2.375 ;
      RECT 47.07 3.685 47.24 3.855 ;
      RECT 47.07 8.61 47.24 8.78 ;
      RECT 47.07 10.09 47.24 10.26 ;
      RECT 46.72 1.395 46.89 1.565 ;
      RECT 46.7 4.055 46.87 4.225 ;
      RECT 46.7 8.24 46.87 8.41 ;
      RECT 46.02 1.4 46.19 1.57 ;
      RECT 45.71 3.32 45.88 3.49 ;
      RECT 45.71 8.975 45.88 9.145 ;
      RECT 45.34 1.4 45.51 1.57 ;
      RECT 45.28 2.21 45.45 2.38 ;
      RECT 45.28 2.95 45.45 3.12 ;
      RECT 45.28 9.345 45.45 9.515 ;
      RECT 45.28 10.085 45.45 10.255 ;
      RECT 44.905 3.69 45.075 3.86 ;
      RECT 44.905 8.605 45.075 8.775 ;
      RECT 44.66 1.4 44.83 1.57 ;
      RECT 43.98 1.4 44.15 1.57 ;
      RECT 42.52 2.71 42.69 2.88 ;
      RECT 42.08 3.575 42.25 3.745 ;
      RECT 42.06 2.71 42.23 2.88 ;
      RECT 41.685 4.32 41.855 4.49 ;
      RECT 41.6 2.71 41.77 2.88 ;
      RECT 41.575 3.595 41.745 3.765 ;
      RECT 41.14 2.71 41.31 2.88 ;
      RECT 40.755 3.285 40.925 3.455 ;
      RECT 40.68 2.71 40.85 2.88 ;
      RECT 40.44 4.325 40.61 4.495 ;
      RECT 40.395 3.815 40.565 3.985 ;
      RECT 40.22 2.71 40.39 2.88 ;
      RECT 40.075 8.975 40.245 9.145 ;
      RECT 39.97 4.025 40.14 4.195 ;
      RECT 39.78 3.245 39.95 3.415 ;
      RECT 39.76 2.71 39.93 2.88 ;
      RECT 39.73 4.855 39.9 5.025 ;
      RECT 39.645 9.345 39.815 9.515 ;
      RECT 39.645 10.085 39.815 10.255 ;
      RECT 39.395 4.295 39.565 4.465 ;
      RECT 39.3 2.71 39.47 2.88 ;
      RECT 39.3 3.455 39.47 3.625 ;
      RECT 38.84 2.71 39.01 2.88 ;
      RECT 38.5 4.68 38.67 4.85 ;
      RECT 38.44 3.88 38.61 4.05 ;
      RECT 38.38 2.71 38.55 2.88 ;
      RECT 38 3.55 38.17 3.72 ;
      RECT 37.92 2.71 38.09 2.88 ;
      RECT 37.735 4.6 37.905 4.77 ;
      RECT 37.49 3.84 37.66 4.01 ;
      RECT 37.46 2.71 37.63 2.88 ;
      RECT 37.395 4.87 37.565 5.04 ;
      RECT 37.12 3.565 37.29 3.735 ;
      RECT 37 2.71 37.17 2.88 ;
      RECT 36.59 3.765 36.76 3.935 ;
      RECT 36.54 2.71 36.71 2.88 ;
      RECT 36.08 2.71 36.25 2.88 ;
      RECT 36.07 3.71 36.24 3.88 ;
      RECT 35.865 3.31 36.035 3.48 ;
      RECT 35.865 4.89 36.035 5.06 ;
      RECT 35.62 2.71 35.79 2.88 ;
      RECT 35.555 3.855 35.725 4.025 ;
      RECT 35.16 2.71 35.33 2.88 ;
      RECT 35.145 4.08 35.315 4.25 ;
      RECT 34.7 2.71 34.87 2.88 ;
      RECT 34.435 4.38 34.605 4.55 ;
      RECT 34.29 3.29 34.46 3.46 ;
      RECT 34.24 2.71 34.41 2.88 ;
      RECT 32.8 8.61 32.97 8.78 ;
      RECT 32.8 10.09 32.97 10.26 ;
      RECT 32.45 1.395 32.62 1.565 ;
      RECT 32.43 4.055 32.6 4.225 ;
      RECT 32.43 8.24 32.6 8.41 ;
      RECT 31.81 2.205 31.98 2.375 ;
      RECT 31.81 3.685 31.98 3.855 ;
      RECT 31.81 8.61 31.98 8.78 ;
      RECT 31.81 10.09 31.98 10.26 ;
      RECT 31.46 1.395 31.63 1.565 ;
      RECT 31.44 4.055 31.61 4.225 ;
      RECT 31.44 8.24 31.61 8.41 ;
      RECT 30.76 1.4 30.93 1.57 ;
      RECT 30.45 3.32 30.62 3.49 ;
      RECT 30.45 8.975 30.62 9.145 ;
      RECT 30.08 1.4 30.25 1.57 ;
      RECT 30.02 2.21 30.19 2.38 ;
      RECT 30.02 2.95 30.19 3.12 ;
      RECT 30.02 9.345 30.19 9.515 ;
      RECT 30.02 10.085 30.19 10.255 ;
      RECT 29.645 3.69 29.815 3.86 ;
      RECT 29.645 8.605 29.815 8.775 ;
      RECT 29.4 1.4 29.57 1.57 ;
      RECT 28.72 1.4 28.89 1.57 ;
      RECT 27.26 2.71 27.43 2.88 ;
      RECT 26.82 3.575 26.99 3.745 ;
      RECT 26.8 2.71 26.97 2.88 ;
      RECT 26.425 4.32 26.595 4.49 ;
      RECT 26.34 2.71 26.51 2.88 ;
      RECT 26.315 3.595 26.485 3.765 ;
      RECT 25.88 2.71 26.05 2.88 ;
      RECT 25.495 3.285 25.665 3.455 ;
      RECT 25.42 2.71 25.59 2.88 ;
      RECT 25.18 4.325 25.35 4.495 ;
      RECT 25.135 3.815 25.305 3.985 ;
      RECT 24.96 2.71 25.13 2.88 ;
      RECT 24.815 8.975 24.985 9.145 ;
      RECT 24.71 4.025 24.88 4.195 ;
      RECT 24.52 3.245 24.69 3.415 ;
      RECT 24.5 2.71 24.67 2.88 ;
      RECT 24.47 4.855 24.64 5.025 ;
      RECT 24.385 9.345 24.555 9.515 ;
      RECT 24.385 10.085 24.555 10.255 ;
      RECT 24.135 4.295 24.305 4.465 ;
      RECT 24.04 2.71 24.21 2.88 ;
      RECT 24.04 3.455 24.21 3.625 ;
      RECT 23.58 2.71 23.75 2.88 ;
      RECT 23.24 4.68 23.41 4.85 ;
      RECT 23.18 3.88 23.35 4.05 ;
      RECT 23.12 2.71 23.29 2.88 ;
      RECT 22.74 3.55 22.91 3.72 ;
      RECT 22.66 2.71 22.83 2.88 ;
      RECT 22.475 4.6 22.645 4.77 ;
      RECT 22.23 3.84 22.4 4.01 ;
      RECT 22.2 2.71 22.37 2.88 ;
      RECT 22.135 4.87 22.305 5.04 ;
      RECT 21.86 3.565 22.03 3.735 ;
      RECT 21.74 2.71 21.91 2.88 ;
      RECT 21.33 3.765 21.5 3.935 ;
      RECT 21.28 2.71 21.45 2.88 ;
      RECT 20.82 2.71 20.99 2.88 ;
      RECT 20.81 3.71 20.98 3.88 ;
      RECT 20.605 3.31 20.775 3.48 ;
      RECT 20.605 4.89 20.775 5.06 ;
      RECT 20.36 2.71 20.53 2.88 ;
      RECT 20.295 3.855 20.465 4.025 ;
      RECT 19.9 2.71 20.07 2.88 ;
      RECT 19.885 4.08 20.055 4.25 ;
      RECT 19.44 2.71 19.61 2.88 ;
      RECT 19.175 4.38 19.345 4.55 ;
      RECT 19.03 3.29 19.2 3.46 ;
      RECT 18.98 2.71 19.15 2.88 ;
      RECT 17.54 8.61 17.71 8.78 ;
      RECT 17.54 10.09 17.71 10.26 ;
      RECT 17.19 1.395 17.36 1.565 ;
      RECT 17.17 4.055 17.34 4.225 ;
      RECT 17.17 8.24 17.34 8.41 ;
      RECT 16.55 2.205 16.72 2.375 ;
      RECT 16.55 3.685 16.72 3.855 ;
      RECT 16.55 8.61 16.72 8.78 ;
      RECT 16.55 10.09 16.72 10.26 ;
      RECT 16.2 1.395 16.37 1.565 ;
      RECT 16.18 4.055 16.35 4.225 ;
      RECT 16.18 8.24 16.35 8.41 ;
      RECT 15.5 1.4 15.67 1.57 ;
      RECT 15.19 3.32 15.36 3.49 ;
      RECT 15.19 8.975 15.36 9.145 ;
      RECT 14.82 1.4 14.99 1.57 ;
      RECT 14.76 2.21 14.93 2.38 ;
      RECT 14.76 2.95 14.93 3.12 ;
      RECT 14.76 9.345 14.93 9.515 ;
      RECT 14.76 10.085 14.93 10.255 ;
      RECT 14.385 3.69 14.555 3.86 ;
      RECT 14.385 8.605 14.555 8.775 ;
      RECT 14.14 1.4 14.31 1.57 ;
      RECT 13.46 1.4 13.63 1.57 ;
      RECT 12 2.71 12.17 2.88 ;
      RECT 11.56 3.575 11.73 3.745 ;
      RECT 11.54 2.71 11.71 2.88 ;
      RECT 11.165 4.32 11.335 4.49 ;
      RECT 11.08 2.71 11.25 2.88 ;
      RECT 11.055 3.595 11.225 3.765 ;
      RECT 10.62 2.71 10.79 2.88 ;
      RECT 10.235 3.285 10.405 3.455 ;
      RECT 10.16 2.71 10.33 2.88 ;
      RECT 9.92 4.325 10.09 4.495 ;
      RECT 9.875 3.815 10.045 3.985 ;
      RECT 9.7 2.71 9.87 2.88 ;
      RECT 9.555 8.975 9.725 9.145 ;
      RECT 9.45 4.025 9.62 4.195 ;
      RECT 9.26 3.245 9.43 3.415 ;
      RECT 9.24 2.71 9.41 2.88 ;
      RECT 9.21 4.855 9.38 5.025 ;
      RECT 9.125 9.345 9.295 9.515 ;
      RECT 9.125 10.085 9.295 10.255 ;
      RECT 8.875 4.295 9.045 4.465 ;
      RECT 8.78 2.71 8.95 2.88 ;
      RECT 8.78 3.455 8.95 3.625 ;
      RECT 8.32 2.71 8.49 2.88 ;
      RECT 7.98 4.68 8.15 4.85 ;
      RECT 7.92 3.88 8.09 4.05 ;
      RECT 7.86 2.71 8.03 2.88 ;
      RECT 7.48 3.55 7.65 3.72 ;
      RECT 7.4 2.71 7.57 2.88 ;
      RECT 7.215 4.6 7.385 4.77 ;
      RECT 6.97 3.84 7.14 4.01 ;
      RECT 6.94 2.71 7.11 2.88 ;
      RECT 6.875 4.87 7.045 5.04 ;
      RECT 6.6 3.565 6.77 3.735 ;
      RECT 6.48 2.71 6.65 2.88 ;
      RECT 6.07 3.765 6.24 3.935 ;
      RECT 6.02 2.71 6.19 2.88 ;
      RECT 5.56 2.71 5.73 2.88 ;
      RECT 5.55 3.71 5.72 3.88 ;
      RECT 5.345 3.31 5.515 3.48 ;
      RECT 5.345 4.89 5.515 5.06 ;
      RECT 5.1 2.71 5.27 2.88 ;
      RECT 5.035 3.855 5.205 4.025 ;
      RECT 4.64 2.71 4.81 2.88 ;
      RECT 4.625 4.08 4.795 4.25 ;
      RECT 4.18 2.71 4.35 2.88 ;
      RECT 3.915 4.38 4.085 4.55 ;
      RECT 3.77 3.29 3.94 3.46 ;
      RECT 3.72 2.71 3.89 2.88 ;
      RECT 1.63 9.345 1.8 9.515 ;
      RECT 1.63 10.085 1.8 10.255 ;
      RECT 1.255 8.605 1.425 8.775 ;
    LAYER li1 ;
      RECT 72.585 0 72.755 3.38 ;
      RECT 71.645 0 71.815 3.38 ;
      RECT 70.685 0 70.855 3.38 ;
      RECT 68.765 0 68.935 3.38 ;
      RECT 67.805 0 67.975 3.38 ;
      RECT 65.885 0 66.055 3.38 ;
      RECT 57.325 0 57.495 3.38 ;
      RECT 56.385 0 56.555 3.38 ;
      RECT 55.425 0 55.595 3.38 ;
      RECT 53.505 0 53.675 3.38 ;
      RECT 52.545 0 52.715 3.38 ;
      RECT 50.625 0 50.795 3.38 ;
      RECT 42.065 0 42.235 3.38 ;
      RECT 41.125 0 41.295 3.38 ;
      RECT 40.165 0 40.335 3.38 ;
      RECT 38.245 0 38.415 3.38 ;
      RECT 37.285 0 37.455 3.38 ;
      RECT 35.365 0 35.535 3.38 ;
      RECT 26.805 0 26.975 3.38 ;
      RECT 25.865 0 26.035 3.38 ;
      RECT 24.905 0 25.075 3.38 ;
      RECT 22.985 0 23.155 3.38 ;
      RECT 22.025 0 22.195 3.38 ;
      RECT 20.105 0 20.275 3.38 ;
      RECT 11.545 0 11.715 3.38 ;
      RECT 10.605 0 10.775 3.38 ;
      RECT 9.645 0 9.815 3.38 ;
      RECT 7.725 0 7.895 3.38 ;
      RECT 6.765 0 6.935 3.38 ;
      RECT 4.845 0 5.015 3.38 ;
      RECT 69.64 0 69.835 2.89 ;
      RECT 65.885 0 66.16 2.89 ;
      RECT 54.38 0 54.575 2.89 ;
      RECT 50.625 0 50.9 2.89 ;
      RECT 39.12 0 39.315 2.89 ;
      RECT 35.365 0 35.64 2.89 ;
      RECT 23.86 0 24.055 2.89 ;
      RECT 20.105 0 20.38 2.89 ;
      RECT 8.6 0 8.795 2.89 ;
      RECT 4.845 0 5.12 2.89 ;
      RECT 64.615 0 73.355 2.88 ;
      RECT 49.355 0 58.095 2.88 ;
      RECT 34.095 0 42.835 2.88 ;
      RECT 18.835 0 27.575 2.88 ;
      RECT 3.575 0 12.315 2.88 ;
      RECT 74.42 0 74.59 2.23 ;
      RECT 59.16 0 59.33 2.23 ;
      RECT 43.9 0 44.07 2.23 ;
      RECT 28.64 0 28.81 2.23 ;
      RECT 13.38 0 13.55 2.23 ;
      RECT 78.15 0 78.32 2.225 ;
      RECT 77.16 0 77.33 2.225 ;
      RECT 62.89 0 63.06 2.225 ;
      RECT 61.9 0 62.07 2.225 ;
      RECT 47.63 0 47.8 2.225 ;
      RECT 46.64 0 46.81 2.225 ;
      RECT 32.37 0 32.54 2.225 ;
      RECT 31.38 0 31.55 2.225 ;
      RECT 17.11 0 17.28 2.225 ;
      RECT 16.12 0 16.29 2.225 ;
      RECT 0.03 0 79.125 1.6 ;
      RECT 78.21 3.035 78.38 4.225 ;
      RECT 78.21 3.035 78.68 3.205 ;
      RECT 78.21 9.26 78.68 9.43 ;
      RECT 78.21 8.24 78.38 9.43 ;
      RECT 77.22 3.035 77.39 4.225 ;
      RECT 77.22 3.035 77.69 3.205 ;
      RECT 77.22 9.26 77.69 9.43 ;
      RECT 77.22 8.24 77.39 9.43 ;
      RECT 75.37 3.93 75.54 5.16 ;
      RECT 75.425 2.15 75.595 4.1 ;
      RECT 75.37 1.87 75.54 2.32 ;
      RECT 75.37 10.145 75.54 10.595 ;
      RECT 75.425 8.365 75.595 10.315 ;
      RECT 75.37 7.305 75.54 8.535 ;
      RECT 74.85 1.87 75.02 5.16 ;
      RECT 74.85 3.37 75.255 3.7 ;
      RECT 74.85 2.53 75.255 2.86 ;
      RECT 74.85 7.305 75.02 10.595 ;
      RECT 74.85 9.605 75.255 9.935 ;
      RECT 74.85 8.765 75.255 9.095 ;
      RECT 72.775 4.421 72.78 4.593 ;
      RECT 72.77 4.414 72.775 4.683 ;
      RECT 72.765 4.408 72.77 4.702 ;
      RECT 72.745 4.402 72.765 4.712 ;
      RECT 72.73 4.397 72.745 4.72 ;
      RECT 72.693 4.391 72.73 4.718 ;
      RECT 72.607 4.377 72.693 4.714 ;
      RECT 72.521 4.359 72.607 4.709 ;
      RECT 72.435 4.34 72.521 4.703 ;
      RECT 72.405 4.328 72.435 4.699 ;
      RECT 72.385 4.322 72.405 4.698 ;
      RECT 72.32 4.32 72.385 4.696 ;
      RECT 72.305 4.32 72.32 4.688 ;
      RECT 72.29 4.32 72.305 4.675 ;
      RECT 72.285 4.32 72.29 4.665 ;
      RECT 72.27 4.32 72.285 4.643 ;
      RECT 72.255 4.32 72.27 4.61 ;
      RECT 72.25 4.32 72.255 4.588 ;
      RECT 72.24 4.32 72.25 4.57 ;
      RECT 72.225 4.32 72.24 4.548 ;
      RECT 72.205 4.32 72.225 4.51 ;
      RECT 72.555 3.605 72.59 4.044 ;
      RECT 72.555 3.605 72.595 4.043 ;
      RECT 72.5 3.665 72.595 4.042 ;
      RECT 72.365 3.837 72.595 4.041 ;
      RECT 72.475 3.715 72.595 4.041 ;
      RECT 72.365 3.837 72.62 4.031 ;
      RECT 72.42 3.782 72.7 3.948 ;
      RECT 72.595 3.576 72.6 4.039 ;
      RECT 72.45 3.752 72.74 3.825 ;
      RECT 72.465 3.735 72.595 4.041 ;
      RECT 72.6 3.575 72.77 3.763 ;
      RECT 72.59 3.578 72.77 3.763 ;
      RECT 72.095 3.455 72.265 3.765 ;
      RECT 72.095 3.455 72.27 3.738 ;
      RECT 72.095 3.455 72.275 3.715 ;
      RECT 72.095 3.455 72.285 3.665 ;
      RECT 72.09 3.56 72.285 3.635 ;
      RECT 72.125 3.13 72.295 3.608 ;
      RECT 72.125 3.13 72.31 3.529 ;
      RECT 72.115 3.34 72.31 3.529 ;
      RECT 72.125 3.14 72.32 3.444 ;
      RECT 72.055 3.882 72.06 4.085 ;
      RECT 72.045 3.87 72.055 4.195 ;
      RECT 72.02 3.87 72.045 4.235 ;
      RECT 71.94 3.87 72.02 4.32 ;
      RECT 71.93 3.87 71.94 4.39 ;
      RECT 71.905 3.87 71.93 4.413 ;
      RECT 71.885 3.87 71.905 4.448 ;
      RECT 71.84 3.88 71.885 4.491 ;
      RECT 71.83 3.892 71.84 4.528 ;
      RECT 71.81 3.906 71.83 4.548 ;
      RECT 71.8 3.924 71.81 4.564 ;
      RECT 71.785 3.95 71.8 4.574 ;
      RECT 71.77 3.991 71.785 4.588 ;
      RECT 71.76 4.026 71.77 4.598 ;
      RECT 71.755 4.042 71.76 4.603 ;
      RECT 71.745 4.057 71.755 4.608 ;
      RECT 71.725 4.1 71.745 4.618 ;
      RECT 71.705 4.137 71.725 4.631 ;
      RECT 71.67 4.16 71.705 4.649 ;
      RECT 71.66 4.174 71.67 4.665 ;
      RECT 71.64 4.184 71.66 4.675 ;
      RECT 71.635 4.193 71.64 4.683 ;
      RECT 71.625 4.2 71.635 4.69 ;
      RECT 71.615 4.207 71.625 4.698 ;
      RECT 71.6 4.217 71.615 4.706 ;
      RECT 71.59 4.231 71.6 4.716 ;
      RECT 71.58 4.243 71.59 4.728 ;
      RECT 71.565 4.265 71.58 4.741 ;
      RECT 71.555 4.287 71.565 4.752 ;
      RECT 71.545 4.307 71.555 4.761 ;
      RECT 71.54 4.322 71.545 4.768 ;
      RECT 71.51 4.355 71.54 4.782 ;
      RECT 71.5 4.39 71.51 4.797 ;
      RECT 71.495 4.397 71.5 4.803 ;
      RECT 71.475 4.412 71.495 4.81 ;
      RECT 71.47 4.427 71.475 4.818 ;
      RECT 71.465 4.436 71.47 4.823 ;
      RECT 71.45 4.442 71.465 4.83 ;
      RECT 71.445 4.448 71.45 4.838 ;
      RECT 71.44 4.452 71.445 4.845 ;
      RECT 71.435 4.456 71.44 4.855 ;
      RECT 71.425 4.461 71.435 4.865 ;
      RECT 71.405 4.472 71.425 4.893 ;
      RECT 71.39 4.484 71.405 4.92 ;
      RECT 71.37 4.497 71.39 4.945 ;
      RECT 71.35 4.512 71.37 4.969 ;
      RECT 71.335 4.527 71.35 4.984 ;
      RECT 71.33 4.538 71.335 4.993 ;
      RECT 71.265 4.583 71.33 5.003 ;
      RECT 71.23 4.642 71.265 5.016 ;
      RECT 71.225 4.665 71.23 5.022 ;
      RECT 71.22 4.672 71.225 5.024 ;
      RECT 71.205 4.682 71.22 5.027 ;
      RECT 71.175 4.707 71.205 5.031 ;
      RECT 71.17 4.725 71.175 5.035 ;
      RECT 71.165 4.732 71.17 5.036 ;
      RECT 71.145 4.74 71.165 5.04 ;
      RECT 71.135 4.747 71.145 5.044 ;
      RECT 71.091 4.758 71.135 5.051 ;
      RECT 71.005 4.786 71.091 5.067 ;
      RECT 70.945 4.81 71.005 5.085 ;
      RECT 70.9 4.82 70.945 5.099 ;
      RECT 70.841 4.828 70.9 5.113 ;
      RECT 70.755 4.835 70.841 5.132 ;
      RECT 70.73 4.84 70.755 5.147 ;
      RECT 70.65 4.843 70.73 5.15 ;
      RECT 70.57 4.847 70.65 5.137 ;
      RECT 70.561 4.85 70.57 5.122 ;
      RECT 70.475 4.85 70.561 5.107 ;
      RECT 70.415 4.852 70.475 5.084 ;
      RECT 70.411 4.855 70.415 5.074 ;
      RECT 70.325 4.855 70.411 5.059 ;
      RECT 70.25 4.855 70.325 5.035 ;
      RECT 71.565 3.864 71.575 4.04 ;
      RECT 71.52 3.831 71.565 4.04 ;
      RECT 71.475 3.782 71.52 4.04 ;
      RECT 71.445 3.752 71.475 4.041 ;
      RECT 71.44 3.735 71.445 4.042 ;
      RECT 71.415 3.715 71.44 4.043 ;
      RECT 71.4 3.69 71.415 4.044 ;
      RECT 71.395 3.677 71.4 4.045 ;
      RECT 71.39 3.671 71.395 4.043 ;
      RECT 71.385 3.663 71.39 4.037 ;
      RECT 71.36 3.655 71.385 4.017 ;
      RECT 71.34 3.644 71.36 3.988 ;
      RECT 71.31 3.629 71.34 3.959 ;
      RECT 71.29 3.615 71.31 3.931 ;
      RECT 71.28 3.609 71.29 3.91 ;
      RECT 71.275 3.606 71.28 3.893 ;
      RECT 71.27 3.603 71.275 3.878 ;
      RECT 71.255 3.598 71.27 3.843 ;
      RECT 71.25 3.594 71.255 3.81 ;
      RECT 71.23 3.589 71.25 3.786 ;
      RECT 71.2 3.581 71.23 3.751 ;
      RECT 71.185 3.575 71.2 3.728 ;
      RECT 71.145 3.568 71.185 3.713 ;
      RECT 71.12 3.56 71.145 3.693 ;
      RECT 71.1 3.555 71.12 3.683 ;
      RECT 71.065 3.549 71.1 3.678 ;
      RECT 71.02 3.54 71.065 3.677 ;
      RECT 70.99 3.536 71.02 3.679 ;
      RECT 70.905 3.544 70.99 3.683 ;
      RECT 70.835 3.555 70.905 3.705 ;
      RECT 70.822 3.561 70.835 3.728 ;
      RECT 70.736 3.568 70.822 3.75 ;
      RECT 70.65 3.58 70.736 3.787 ;
      RECT 70.65 3.957 70.66 4.195 ;
      RECT 70.645 3.586 70.65 3.81 ;
      RECT 70.64 3.842 70.65 4.195 ;
      RECT 70.64 3.587 70.645 3.815 ;
      RECT 70.635 3.588 70.64 4.195 ;
      RECT 70.611 3.59 70.635 4.196 ;
      RECT 70.525 3.598 70.611 4.198 ;
      RECT 70.505 3.612 70.525 4.201 ;
      RECT 70.5 3.64 70.505 4.202 ;
      RECT 70.495 3.652 70.5 4.203 ;
      RECT 70.49 3.667 70.495 4.204 ;
      RECT 70.48 3.697 70.49 4.205 ;
      RECT 70.475 3.735 70.48 4.203 ;
      RECT 70.47 3.755 70.475 4.198 ;
      RECT 70.455 3.79 70.47 4.183 ;
      RECT 70.445 3.842 70.455 4.163 ;
      RECT 70.44 3.872 70.445 4.151 ;
      RECT 70.425 3.885 70.44 4.134 ;
      RECT 70.4 3.889 70.425 4.101 ;
      RECT 70.385 3.887 70.4 4.078 ;
      RECT 70.37 3.886 70.385 4.075 ;
      RECT 70.31 3.884 70.37 4.073 ;
      RECT 70.3 3.882 70.31 4.068 ;
      RECT 70.26 3.881 70.3 4.065 ;
      RECT 70.19 3.878 70.26 4.063 ;
      RECT 70.135 3.876 70.19 4.058 ;
      RECT 70.065 3.87 70.135 4.053 ;
      RECT 70.056 3.87 70.065 4.05 ;
      RECT 69.97 3.87 70.056 4.045 ;
      RECT 69.965 3.87 69.97 4.04 ;
      RECT 71.27 3.105 71.445 3.455 ;
      RECT 71.27 3.12 71.455 3.453 ;
      RECT 71.245 3.07 71.39 3.45 ;
      RECT 71.225 3.071 71.39 3.443 ;
      RECT 71.215 3.072 71.4 3.438 ;
      RECT 71.185 3.073 71.4 3.425 ;
      RECT 71.135 3.074 71.4 3.401 ;
      RECT 71.13 3.076 71.4 3.386 ;
      RECT 71.13 3.142 71.46 3.38 ;
      RECT 71.11 3.083 71.415 3.36 ;
      RECT 71.1 3.092 71.425 3.215 ;
      RECT 71.11 3.087 71.425 3.36 ;
      RECT 71.13 3.077 71.415 3.386 ;
      RECT 70.715 4.402 70.885 4.69 ;
      RECT 70.71 4.42 70.895 4.685 ;
      RECT 70.675 4.428 70.96 4.605 ;
      RECT 70.675 4.428 71.046 4.595 ;
      RECT 70.675 4.428 71.1 4.541 ;
      RECT 70.96 4.325 71.13 4.509 ;
      RECT 70.675 4.48 71.135 4.497 ;
      RECT 70.66 4.45 71.13 4.493 ;
      RECT 70.92 4.332 70.96 4.644 ;
      RECT 70.8 4.369 71.13 4.509 ;
      RECT 70.895 4.344 70.92 4.67 ;
      RECT 70.885 4.351 71.13 4.509 ;
      RECT 71.016 3.815 71.085 4.074 ;
      RECT 71.016 3.87 71.09 4.073 ;
      RECT 70.93 3.87 71.09 4.072 ;
      RECT 70.925 3.87 71.095 4.065 ;
      RECT 70.915 3.815 71.085 4.06 ;
      RECT 70.295 3.114 70.47 3.415 ;
      RECT 70.28 3.102 70.295 3.4 ;
      RECT 70.25 3.101 70.28 3.353 ;
      RECT 70.25 3.119 70.475 3.348 ;
      RECT 70.235 3.103 70.295 3.313 ;
      RECT 70.23 3.125 70.485 3.213 ;
      RECT 70.23 3.108 70.381 3.213 ;
      RECT 70.23 3.11 70.385 3.213 ;
      RECT 70.235 3.106 70.381 3.313 ;
      RECT 70.34 4.342 70.345 4.69 ;
      RECT 70.33 4.332 70.34 4.696 ;
      RECT 70.295 4.322 70.33 4.698 ;
      RECT 70.257 4.317 70.295 4.702 ;
      RECT 70.171 4.31 70.257 4.709 ;
      RECT 70.085 4.3 70.171 4.719 ;
      RECT 70.04 4.295 70.085 4.727 ;
      RECT 70.036 4.295 70.04 4.731 ;
      RECT 69.95 4.295 70.036 4.738 ;
      RECT 69.935 4.295 69.95 4.738 ;
      RECT 69.925 4.293 69.935 4.71 ;
      RECT 69.915 4.289 69.925 4.653 ;
      RECT 69.895 4.283 69.915 4.585 ;
      RECT 69.89 4.279 69.895 4.533 ;
      RECT 69.88 4.278 69.89 4.5 ;
      RECT 69.83 4.276 69.88 4.485 ;
      RECT 69.805 4.274 69.83 4.48 ;
      RECT 69.762 4.272 69.805 4.476 ;
      RECT 69.676 4.268 69.762 4.464 ;
      RECT 69.59 4.263 69.676 4.448 ;
      RECT 69.56 4.26 69.59 4.435 ;
      RECT 69.535 4.259 69.56 4.423 ;
      RECT 69.53 4.259 69.535 4.413 ;
      RECT 69.49 4.258 69.53 4.405 ;
      RECT 69.475 4.257 69.49 4.398 ;
      RECT 69.425 4.256 69.475 4.39 ;
      RECT 69.423 4.255 69.425 4.385 ;
      RECT 69.337 4.253 69.423 4.385 ;
      RECT 69.251 4.248 69.337 4.385 ;
      RECT 69.165 4.244 69.251 4.385 ;
      RECT 69.116 4.24 69.165 4.383 ;
      RECT 69.03 4.237 69.116 4.378 ;
      RECT 69.007 4.234 69.03 4.374 ;
      RECT 68.921 4.231 69.007 4.369 ;
      RECT 68.835 4.227 68.921 4.36 ;
      RECT 68.81 4.22 68.835 4.355 ;
      RECT 68.75 4.185 68.81 4.352 ;
      RECT 68.73 4.11 68.75 4.349 ;
      RECT 68.725 4.052 68.73 4.348 ;
      RECT 68.7 3.992 68.725 4.347 ;
      RECT 68.625 3.87 68.7 4.343 ;
      RECT 68.615 3.87 68.625 4.335 ;
      RECT 68.6 3.87 68.615 4.325 ;
      RECT 68.585 3.87 68.6 4.295 ;
      RECT 68.57 3.87 68.585 4.24 ;
      RECT 68.555 3.87 68.57 4.178 ;
      RECT 68.53 3.87 68.555 4.103 ;
      RECT 68.525 3.87 68.53 4.053 ;
      RECT 69.87 3.415 69.89 3.724 ;
      RECT 69.856 3.417 69.905 3.721 ;
      RECT 69.856 3.422 69.925 3.712 ;
      RECT 69.77 3.42 69.905 3.706 ;
      RECT 69.77 3.428 69.96 3.689 ;
      RECT 69.735 3.43 69.96 3.688 ;
      RECT 69.705 3.438 69.96 3.679 ;
      RECT 69.695 3.443 69.98 3.665 ;
      RECT 69.735 3.433 69.98 3.665 ;
      RECT 69.735 3.436 69.99 3.653 ;
      RECT 69.705 3.438 70 3.64 ;
      RECT 69.705 3.442 70.01 3.583 ;
      RECT 69.695 3.447 70.015 3.498 ;
      RECT 69.856 3.415 69.89 3.721 ;
      RECT 69.295 3.518 69.3 3.73 ;
      RECT 69.17 3.515 69.185 3.73 ;
      RECT 68.635 3.545 68.705 3.73 ;
      RECT 68.52 3.545 68.555 3.725 ;
      RECT 69.641 3.847 69.66 4.041 ;
      RECT 69.555 3.802 69.641 4.042 ;
      RECT 69.545 3.755 69.555 4.044 ;
      RECT 69.54 3.735 69.545 4.045 ;
      RECT 69.52 3.7 69.54 4.046 ;
      RECT 69.505 3.65 69.52 4.047 ;
      RECT 69.485 3.587 69.505 4.048 ;
      RECT 69.475 3.55 69.485 4.049 ;
      RECT 69.46 3.539 69.475 4.05 ;
      RECT 69.455 3.531 69.46 4.048 ;
      RECT 69.445 3.53 69.455 4.04 ;
      RECT 69.415 3.527 69.445 4.019 ;
      RECT 69.34 3.522 69.415 3.964 ;
      RECT 69.325 3.518 69.34 3.91 ;
      RECT 69.315 3.518 69.325 3.805 ;
      RECT 69.3 3.518 69.315 3.738 ;
      RECT 69.285 3.518 69.295 3.728 ;
      RECT 69.23 3.517 69.285 3.725 ;
      RECT 69.185 3.515 69.23 3.728 ;
      RECT 69.157 3.515 69.17 3.731 ;
      RECT 69.071 3.519 69.157 3.733 ;
      RECT 68.985 3.525 69.071 3.738 ;
      RECT 68.965 3.529 68.985 3.74 ;
      RECT 68.963 3.53 68.965 3.739 ;
      RECT 68.877 3.532 68.963 3.738 ;
      RECT 68.791 3.537 68.877 3.735 ;
      RECT 68.705 3.542 68.791 3.732 ;
      RECT 68.555 3.545 68.635 3.728 ;
      RECT 69.215 7.305 69.385 10.595 ;
      RECT 69.215 9.605 69.62 9.935 ;
      RECT 69.215 8.765 69.62 9.095 ;
      RECT 69.331 4.52 69.38 4.854 ;
      RECT 69.331 4.52 69.385 4.853 ;
      RECT 69.245 4.52 69.385 4.852 ;
      RECT 69.02 4.628 69.39 4.85 ;
      RECT 69.245 4.52 69.415 4.843 ;
      RECT 69.215 4.532 69.42 4.834 ;
      RECT 69.2 4.55 69.425 4.831 ;
      RECT 69.015 4.634 69.425 4.758 ;
      RECT 69.01 4.641 69.425 4.718 ;
      RECT 69.025 4.607 69.425 4.831 ;
      RECT 69.186 4.553 69.39 4.85 ;
      RECT 69.1 4.573 69.425 4.831 ;
      RECT 69.2 4.547 69.42 4.834 ;
      RECT 68.97 3.871 69.16 4.065 ;
      RECT 68.965 3.873 69.16 4.064 ;
      RECT 68.96 3.877 69.175 4.061 ;
      RECT 68.975 3.87 69.175 4.061 ;
      RECT 68.96 3.98 69.18 4.056 ;
      RECT 68.255 4.48 68.346 4.778 ;
      RECT 68.25 4.482 68.425 4.773 ;
      RECT 68.255 4.48 68.425 4.773 ;
      RECT 68.25 4.486 68.445 4.771 ;
      RECT 68.25 4.541 68.485 4.77 ;
      RECT 68.25 4.576 68.5 4.764 ;
      RECT 68.25 4.61 68.51 4.754 ;
      RECT 68.24 4.49 68.445 4.605 ;
      RECT 68.24 4.51 68.46 4.605 ;
      RECT 68.24 4.493 68.45 4.605 ;
      RECT 68.465 3.261 68.47 3.323 ;
      RECT 68.46 3.183 68.465 3.346 ;
      RECT 68.455 3.14 68.46 3.357 ;
      RECT 68.45 3.13 68.455 3.369 ;
      RECT 68.445 3.13 68.45 3.378 ;
      RECT 68.42 3.13 68.445 3.41 ;
      RECT 68.415 3.13 68.42 3.443 ;
      RECT 68.4 3.13 68.415 3.468 ;
      RECT 68.39 3.13 68.4 3.495 ;
      RECT 68.385 3.13 68.39 3.508 ;
      RECT 68.38 3.13 68.385 3.523 ;
      RECT 68.37 3.13 68.38 3.538 ;
      RECT 68.365 3.13 68.37 3.558 ;
      RECT 68.34 3.13 68.365 3.593 ;
      RECT 68.295 3.13 68.34 3.638 ;
      RECT 68.285 3.13 68.295 3.651 ;
      RECT 68.2 3.215 68.285 3.658 ;
      RECT 68.165 3.337 68.2 3.667 ;
      RECT 68.16 3.377 68.165 3.671 ;
      RECT 68.14 3.4 68.16 3.673 ;
      RECT 68.135 3.43 68.14 3.676 ;
      RECT 68.125 3.442 68.135 3.677 ;
      RECT 68.08 3.465 68.125 3.682 ;
      RECT 68.04 3.495 68.08 3.69 ;
      RECT 68.005 3.507 68.04 3.696 ;
      RECT 68 3.512 68.005 3.7 ;
      RECT 67.93 3.522 68 3.707 ;
      RECT 67.89 3.532 67.93 3.717 ;
      RECT 67.87 3.537 67.89 3.723 ;
      RECT 67.86 3.541 67.87 3.728 ;
      RECT 67.855 3.544 67.86 3.731 ;
      RECT 67.845 3.545 67.855 3.732 ;
      RECT 67.82 3.547 67.845 3.736 ;
      RECT 67.81 3.552 67.82 3.739 ;
      RECT 67.765 3.56 67.81 3.74 ;
      RECT 67.64 3.565 67.765 3.74 ;
      RECT 68.195 3.862 68.215 4.044 ;
      RECT 68.146 3.847 68.195 4.043 ;
      RECT 68.06 3.862 68.215 4.041 ;
      RECT 68.045 3.862 68.215 4.04 ;
      RECT 68.01 3.84 68.18 4.025 ;
      RECT 68.08 4.86 68.095 5.069 ;
      RECT 68.08 4.868 68.1 5.068 ;
      RECT 68.025 4.868 68.1 5.067 ;
      RECT 68.005 4.872 68.105 5.065 ;
      RECT 67.985 4.822 68.025 5.064 ;
      RECT 67.93 4.88 68.11 5.062 ;
      RECT 67.895 4.837 68.025 5.06 ;
      RECT 67.891 4.84 68.08 5.059 ;
      RECT 67.805 4.848 68.08 5.057 ;
      RECT 67.805 4.892 68.115 5.05 ;
      RECT 67.795 4.985 68.115 5.048 ;
      RECT 67.805 4.904 68.12 5.033 ;
      RECT 67.805 4.925 68.135 5.003 ;
      RECT 67.805 4.952 68.14 4.973 ;
      RECT 67.93 4.83 68.025 5.062 ;
      RECT 67.56 3.875 67.565 4.413 ;
      RECT 67.365 4.205 67.37 4.4 ;
      RECT 65.665 3.87 65.68 4.25 ;
      RECT 67.73 3.87 67.735 4.04 ;
      RECT 67.725 3.87 67.73 4.05 ;
      RECT 67.72 3.87 67.725 4.063 ;
      RECT 67.695 3.87 67.72 4.105 ;
      RECT 67.67 3.87 67.695 4.178 ;
      RECT 67.655 3.87 67.67 4.23 ;
      RECT 67.65 3.87 67.655 4.26 ;
      RECT 67.625 3.87 67.65 4.3 ;
      RECT 67.61 3.87 67.625 4.355 ;
      RECT 67.605 3.87 67.61 4.388 ;
      RECT 67.58 3.87 67.605 4.408 ;
      RECT 67.565 3.87 67.58 4.414 ;
      RECT 67.495 3.905 67.56 4.41 ;
      RECT 67.445 3.96 67.495 4.405 ;
      RECT 67.435 3.992 67.445 4.403 ;
      RECT 67.43 4.017 67.435 4.403 ;
      RECT 67.41 4.09 67.43 4.403 ;
      RECT 67.4 4.17 67.41 4.402 ;
      RECT 67.385 4.2 67.4 4.402 ;
      RECT 67.37 4.205 67.385 4.401 ;
      RECT 67.31 4.207 67.365 4.398 ;
      RECT 67.28 4.212 67.31 4.394 ;
      RECT 67.278 4.215 67.28 4.393 ;
      RECT 67.192 4.217 67.278 4.39 ;
      RECT 67.106 4.223 67.192 4.384 ;
      RECT 67.02 4.228 67.106 4.378 ;
      RECT 66.947 4.233 67.02 4.379 ;
      RECT 66.861 4.239 66.947 4.387 ;
      RECT 66.775 4.245 66.861 4.396 ;
      RECT 66.755 4.249 66.775 4.401 ;
      RECT 66.708 4.251 66.755 4.404 ;
      RECT 66.622 4.256 66.708 4.41 ;
      RECT 66.536 4.261 66.622 4.419 ;
      RECT 66.45 4.267 66.536 4.427 ;
      RECT 66.365 4.265 66.45 4.436 ;
      RECT 66.361 4.26 66.365 4.44 ;
      RECT 66.275 4.255 66.361 4.432 ;
      RECT 66.211 4.246 66.275 4.42 ;
      RECT 66.125 4.237 66.211 4.407 ;
      RECT 66.101 4.23 66.125 4.398 ;
      RECT 66.015 4.224 66.101 4.385 ;
      RECT 65.975 4.217 66.015 4.371 ;
      RECT 65.97 4.207 65.975 4.367 ;
      RECT 65.96 4.195 65.97 4.366 ;
      RECT 65.94 4.165 65.96 4.363 ;
      RECT 65.885 4.085 65.94 4.357 ;
      RECT 65.865 4.004 65.885 4.352 ;
      RECT 65.845 3.962 65.865 4.348 ;
      RECT 65.82 3.915 65.845 4.342 ;
      RECT 65.815 3.89 65.82 4.339 ;
      RECT 65.78 3.87 65.815 4.334 ;
      RECT 65.771 3.87 65.78 4.327 ;
      RECT 65.685 3.87 65.771 4.297 ;
      RECT 65.68 3.87 65.685 4.26 ;
      RECT 65.645 3.87 65.665 4.182 ;
      RECT 65.64 3.912 65.645 4.147 ;
      RECT 65.635 3.987 65.64 4.103 ;
      RECT 67.085 3.792 67.26 4.04 ;
      RECT 67.085 3.792 67.265 4.038 ;
      RECT 67.08 3.824 67.265 3.998 ;
      RECT 67.11 3.765 67.28 3.985 ;
      RECT 67.075 3.842 67.28 3.918 ;
      RECT 66.385 3.305 66.555 3.48 ;
      RECT 66.385 3.305 66.727 3.472 ;
      RECT 66.385 3.305 66.81 3.466 ;
      RECT 66.385 3.305 66.845 3.462 ;
      RECT 66.385 3.305 66.865 3.461 ;
      RECT 66.385 3.305 66.951 3.457 ;
      RECT 66.845 3.13 67.015 3.452 ;
      RECT 66.42 3.237 67.045 3.45 ;
      RECT 66.41 3.292 67.05 3.448 ;
      RECT 66.385 3.328 67.06 3.443 ;
      RECT 66.385 3.355 67.065 3.373 ;
      RECT 66.45 3.18 67.025 3.45 ;
      RECT 66.641 3.165 67.025 3.45 ;
      RECT 66.475 3.168 67.025 3.45 ;
      RECT 66.555 3.166 66.641 3.477 ;
      RECT 66.641 3.163 67.02 3.45 ;
      RECT 66.825 3.14 67.02 3.45 ;
      RECT 66.727 3.161 67.02 3.45 ;
      RECT 66.81 3.155 66.825 3.463 ;
      RECT 66.96 4.52 66.965 4.72 ;
      RECT 66.425 4.585 66.47 4.72 ;
      RECT 66.995 4.52 67.015 4.693 ;
      RECT 66.965 4.52 66.995 4.708 ;
      RECT 66.9 4.52 66.96 4.745 ;
      RECT 66.885 4.52 66.9 4.775 ;
      RECT 66.87 4.52 66.885 4.788 ;
      RECT 66.85 4.52 66.87 4.803 ;
      RECT 66.845 4.52 66.85 4.812 ;
      RECT 66.835 4.524 66.845 4.817 ;
      RECT 66.82 4.534 66.835 4.828 ;
      RECT 66.795 4.55 66.82 4.838 ;
      RECT 66.785 4.564 66.795 4.84 ;
      RECT 66.765 4.576 66.785 4.837 ;
      RECT 66.735 4.597 66.765 4.831 ;
      RECT 66.725 4.609 66.735 4.826 ;
      RECT 66.715 4.607 66.725 4.823 ;
      RECT 66.7 4.606 66.715 4.818 ;
      RECT 66.695 4.605 66.7 4.813 ;
      RECT 66.66 4.603 66.695 4.803 ;
      RECT 66.64 4.6 66.66 4.785 ;
      RECT 66.63 4.598 66.64 4.78 ;
      RECT 66.62 4.597 66.63 4.775 ;
      RECT 66.585 4.595 66.62 4.763 ;
      RECT 66.53 4.591 66.585 4.743 ;
      RECT 66.52 4.589 66.53 4.728 ;
      RECT 66.515 4.589 66.52 4.723 ;
      RECT 66.47 4.587 66.515 4.72 ;
      RECT 66.375 4.585 66.425 4.724 ;
      RECT 66.365 4.586 66.375 4.729 ;
      RECT 66.305 4.593 66.365 4.743 ;
      RECT 66.28 4.601 66.305 4.763 ;
      RECT 66.27 4.605 66.28 4.775 ;
      RECT 66.265 4.606 66.27 4.78 ;
      RECT 66.25 4.608 66.265 4.783 ;
      RECT 66.235 4.61 66.25 4.788 ;
      RECT 66.23 4.61 66.235 4.791 ;
      RECT 66.185 4.615 66.23 4.802 ;
      RECT 66.18 4.619 66.185 4.814 ;
      RECT 66.155 4.615 66.18 4.818 ;
      RECT 66.145 4.611 66.155 4.822 ;
      RECT 66.135 4.61 66.145 4.826 ;
      RECT 66.12 4.6 66.135 4.832 ;
      RECT 66.115 4.588 66.12 4.836 ;
      RECT 66.11 4.585 66.115 4.837 ;
      RECT 66.105 4.582 66.11 4.839 ;
      RECT 66.09 4.57 66.105 4.838 ;
      RECT 66.075 4.552 66.09 4.835 ;
      RECT 66.055 4.531 66.075 4.828 ;
      RECT 65.99 4.52 66.055 4.8 ;
      RECT 65.986 4.52 65.99 4.779 ;
      RECT 65.9 4.52 65.986 4.749 ;
      RECT 65.885 4.52 65.9 4.705 ;
      RECT 66.46 3.62 66.465 3.855 ;
      RECT 65.59 3.536 65.595 3.74 ;
      RECT 66.17 3.565 66.175 3.72 ;
      RECT 66.09 3.545 66.095 3.72 ;
      RECT 66.76 3.687 66.775 4.04 ;
      RECT 66.686 3.672 66.76 4.04 ;
      RECT 66.6 3.655 66.686 4.04 ;
      RECT 66.59 3.645 66.6 4.038 ;
      RECT 66.585 3.643 66.59 4.033 ;
      RECT 66.57 3.641 66.585 4.019 ;
      RECT 66.5 3.633 66.57 3.959 ;
      RECT 66.48 3.624 66.5 3.893 ;
      RECT 66.475 3.621 66.48 3.873 ;
      RECT 66.465 3.62 66.475 3.863 ;
      RECT 66.455 3.62 66.46 3.847 ;
      RECT 66.445 3.619 66.455 3.837 ;
      RECT 66.435 3.617 66.445 3.825 ;
      RECT 66.42 3.614 66.435 3.805 ;
      RECT 66.41 3.612 66.42 3.79 ;
      RECT 66.39 3.609 66.41 3.778 ;
      RECT 66.385 3.607 66.39 3.768 ;
      RECT 66.36 3.605 66.385 3.755 ;
      RECT 66.33 3.6 66.36 3.74 ;
      RECT 66.25 3.591 66.33 3.731 ;
      RECT 66.205 3.58 66.25 3.724 ;
      RECT 66.185 3.571 66.205 3.721 ;
      RECT 66.175 3.566 66.185 3.72 ;
      RECT 66.13 3.56 66.17 3.72 ;
      RECT 66.115 3.552 66.13 3.72 ;
      RECT 66.095 3.547 66.115 3.72 ;
      RECT 66.075 3.544 66.09 3.72 ;
      RECT 65.992 3.543 66.075 3.719 ;
      RECT 65.906 3.542 65.992 3.715 ;
      RECT 65.82 3.54 65.906 3.712 ;
      RECT 65.767 3.539 65.82 3.714 ;
      RECT 65.681 3.538 65.767 3.723 ;
      RECT 65.595 3.537 65.681 3.735 ;
      RECT 65.575 3.536 65.59 3.743 ;
      RECT 65.495 3.535 65.575 3.755 ;
      RECT 65.47 3.535 65.495 3.768 ;
      RECT 65.445 3.535 65.47 3.783 ;
      RECT 65.44 3.535 65.445 3.805 ;
      RECT 65.435 3.535 65.44 3.823 ;
      RECT 65.43 3.535 65.435 3.84 ;
      RECT 65.425 3.535 65.43 3.853 ;
      RECT 65.42 3.535 65.425 3.863 ;
      RECT 65.38 3.535 65.42 3.948 ;
      RECT 65.365 3.535 65.38 4.033 ;
      RECT 65.355 3.536 65.365 4.045 ;
      RECT 65.32 3.541 65.355 4.05 ;
      RECT 65.28 3.55 65.32 4.05 ;
      RECT 65.265 3.56 65.28 4.05 ;
      RECT 65.26 3.57 65.265 4.05 ;
      RECT 65.24 3.597 65.26 4.05 ;
      RECT 65.19 3.68 65.24 4.05 ;
      RECT 65.185 3.742 65.19 4.05 ;
      RECT 65.175 3.755 65.185 4.05 ;
      RECT 65.165 3.777 65.175 4.05 ;
      RECT 65.155 3.802 65.165 4.045 ;
      RECT 65.15 3.84 65.155 4.038 ;
      RECT 65.14 3.95 65.15 4.033 ;
      RECT 66.535 4.871 66.55 5.13 ;
      RECT 66.535 4.886 66.555 5.129 ;
      RECT 66.451 4.886 66.555 5.127 ;
      RECT 66.451 4.9 66.56 5.126 ;
      RECT 66.365 4.942 66.565 5.123 ;
      RECT 66.36 4.885 66.55 5.118 ;
      RECT 66.36 4.956 66.57 5.115 ;
      RECT 66.355 4.987 66.57 5.113 ;
      RECT 66.36 4.984 66.585 5.103 ;
      RECT 66.355 5.03 66.6 5.088 ;
      RECT 66.355 5.058 66.605 5.073 ;
      RECT 66.365 4.86 66.535 5.123 ;
      RECT 66.125 3.87 66.295 4.04 ;
      RECT 66.09 3.87 66.295 4.035 ;
      RECT 66.08 3.87 66.295 4.028 ;
      RECT 66.075 3.855 66.245 4.025 ;
      RECT 64.905 4.392 65.17 4.835 ;
      RECT 64.9 4.363 65.115 4.833 ;
      RECT 64.895 4.517 65.175 4.828 ;
      RECT 64.9 4.412 65.175 4.828 ;
      RECT 64.9 4.423 65.185 4.815 ;
      RECT 64.9 4.37 65.145 4.833 ;
      RECT 64.905 4.357 65.115 4.835 ;
      RECT 64.905 4.355 65.065 4.835 ;
      RECT 65.006 4.347 65.065 4.835 ;
      RECT 64.92 4.348 65.065 4.835 ;
      RECT 65.006 4.346 65.055 4.835 ;
      RECT 64.81 3.161 64.985 3.46 ;
      RECT 64.86 3.123 64.985 3.46 ;
      RECT 64.845 3.125 65.071 3.452 ;
      RECT 64.845 3.128 65.11 3.439 ;
      RECT 64.845 3.129 65.12 3.425 ;
      RECT 64.8 3.18 65.12 3.415 ;
      RECT 64.845 3.13 65.125 3.41 ;
      RECT 64.8 3.34 65.13 3.4 ;
      RECT 64.785 3.2 65.125 3.34 ;
      RECT 64.78 3.216 65.125 3.28 ;
      RECT 64.825 3.14 65.125 3.41 ;
      RECT 64.86 3.121 64.946 3.46 ;
      RECT 62.95 3.035 63.12 4.225 ;
      RECT 62.95 3.035 63.42 3.205 ;
      RECT 62.95 9.26 63.42 9.43 ;
      RECT 62.95 8.24 63.12 9.43 ;
      RECT 61.96 3.035 62.13 4.225 ;
      RECT 61.96 3.035 62.43 3.205 ;
      RECT 61.96 9.26 62.43 9.43 ;
      RECT 61.96 8.24 62.13 9.43 ;
      RECT 60.11 3.93 60.28 5.16 ;
      RECT 60.165 2.15 60.335 4.1 ;
      RECT 60.11 1.87 60.28 2.32 ;
      RECT 60.11 10.145 60.28 10.595 ;
      RECT 60.165 8.365 60.335 10.315 ;
      RECT 60.11 7.305 60.28 8.535 ;
      RECT 59.59 1.87 59.76 5.16 ;
      RECT 59.59 3.37 59.995 3.7 ;
      RECT 59.59 2.53 59.995 2.86 ;
      RECT 59.59 7.305 59.76 10.595 ;
      RECT 59.59 9.605 59.995 9.935 ;
      RECT 59.59 8.765 59.995 9.095 ;
      RECT 57.515 4.421 57.52 4.593 ;
      RECT 57.51 4.414 57.515 4.683 ;
      RECT 57.505 4.408 57.51 4.702 ;
      RECT 57.485 4.402 57.505 4.712 ;
      RECT 57.47 4.397 57.485 4.72 ;
      RECT 57.433 4.391 57.47 4.718 ;
      RECT 57.347 4.377 57.433 4.714 ;
      RECT 57.261 4.359 57.347 4.709 ;
      RECT 57.175 4.34 57.261 4.703 ;
      RECT 57.145 4.328 57.175 4.699 ;
      RECT 57.125 4.322 57.145 4.698 ;
      RECT 57.06 4.32 57.125 4.696 ;
      RECT 57.045 4.32 57.06 4.688 ;
      RECT 57.03 4.32 57.045 4.675 ;
      RECT 57.025 4.32 57.03 4.665 ;
      RECT 57.01 4.32 57.025 4.643 ;
      RECT 56.995 4.32 57.01 4.61 ;
      RECT 56.99 4.32 56.995 4.588 ;
      RECT 56.98 4.32 56.99 4.57 ;
      RECT 56.965 4.32 56.98 4.548 ;
      RECT 56.945 4.32 56.965 4.51 ;
      RECT 57.295 3.605 57.33 4.044 ;
      RECT 57.295 3.605 57.335 4.043 ;
      RECT 57.24 3.665 57.335 4.042 ;
      RECT 57.105 3.837 57.335 4.041 ;
      RECT 57.215 3.715 57.335 4.041 ;
      RECT 57.105 3.837 57.36 4.031 ;
      RECT 57.16 3.782 57.44 3.948 ;
      RECT 57.335 3.576 57.34 4.039 ;
      RECT 57.19 3.752 57.48 3.825 ;
      RECT 57.205 3.735 57.335 4.041 ;
      RECT 57.34 3.575 57.51 3.763 ;
      RECT 57.33 3.578 57.51 3.763 ;
      RECT 56.835 3.455 57.005 3.765 ;
      RECT 56.835 3.455 57.01 3.738 ;
      RECT 56.835 3.455 57.015 3.715 ;
      RECT 56.835 3.455 57.025 3.665 ;
      RECT 56.83 3.56 57.025 3.635 ;
      RECT 56.865 3.13 57.035 3.608 ;
      RECT 56.865 3.13 57.05 3.529 ;
      RECT 56.855 3.34 57.05 3.529 ;
      RECT 56.865 3.14 57.06 3.444 ;
      RECT 56.795 3.882 56.8 4.085 ;
      RECT 56.785 3.87 56.795 4.195 ;
      RECT 56.76 3.87 56.785 4.235 ;
      RECT 56.68 3.87 56.76 4.32 ;
      RECT 56.67 3.87 56.68 4.39 ;
      RECT 56.645 3.87 56.67 4.413 ;
      RECT 56.625 3.87 56.645 4.448 ;
      RECT 56.58 3.88 56.625 4.491 ;
      RECT 56.57 3.892 56.58 4.528 ;
      RECT 56.55 3.906 56.57 4.548 ;
      RECT 56.54 3.924 56.55 4.564 ;
      RECT 56.525 3.95 56.54 4.574 ;
      RECT 56.51 3.991 56.525 4.588 ;
      RECT 56.5 4.026 56.51 4.598 ;
      RECT 56.495 4.042 56.5 4.603 ;
      RECT 56.485 4.057 56.495 4.608 ;
      RECT 56.465 4.1 56.485 4.618 ;
      RECT 56.445 4.137 56.465 4.631 ;
      RECT 56.41 4.16 56.445 4.649 ;
      RECT 56.4 4.174 56.41 4.665 ;
      RECT 56.38 4.184 56.4 4.675 ;
      RECT 56.375 4.193 56.38 4.683 ;
      RECT 56.365 4.2 56.375 4.69 ;
      RECT 56.355 4.207 56.365 4.698 ;
      RECT 56.34 4.217 56.355 4.706 ;
      RECT 56.33 4.231 56.34 4.716 ;
      RECT 56.32 4.243 56.33 4.728 ;
      RECT 56.305 4.265 56.32 4.741 ;
      RECT 56.295 4.287 56.305 4.752 ;
      RECT 56.285 4.307 56.295 4.761 ;
      RECT 56.28 4.322 56.285 4.768 ;
      RECT 56.25 4.355 56.28 4.782 ;
      RECT 56.24 4.39 56.25 4.797 ;
      RECT 56.235 4.397 56.24 4.803 ;
      RECT 56.215 4.412 56.235 4.81 ;
      RECT 56.21 4.427 56.215 4.818 ;
      RECT 56.205 4.436 56.21 4.823 ;
      RECT 56.19 4.442 56.205 4.83 ;
      RECT 56.185 4.448 56.19 4.838 ;
      RECT 56.18 4.452 56.185 4.845 ;
      RECT 56.175 4.456 56.18 4.855 ;
      RECT 56.165 4.461 56.175 4.865 ;
      RECT 56.145 4.472 56.165 4.893 ;
      RECT 56.13 4.484 56.145 4.92 ;
      RECT 56.11 4.497 56.13 4.945 ;
      RECT 56.09 4.512 56.11 4.969 ;
      RECT 56.075 4.527 56.09 4.984 ;
      RECT 56.07 4.538 56.075 4.993 ;
      RECT 56.005 4.583 56.07 5.003 ;
      RECT 55.97 4.642 56.005 5.016 ;
      RECT 55.965 4.665 55.97 5.022 ;
      RECT 55.96 4.672 55.965 5.024 ;
      RECT 55.945 4.682 55.96 5.027 ;
      RECT 55.915 4.707 55.945 5.031 ;
      RECT 55.91 4.725 55.915 5.035 ;
      RECT 55.905 4.732 55.91 5.036 ;
      RECT 55.885 4.74 55.905 5.04 ;
      RECT 55.875 4.747 55.885 5.044 ;
      RECT 55.831 4.758 55.875 5.051 ;
      RECT 55.745 4.786 55.831 5.067 ;
      RECT 55.685 4.81 55.745 5.085 ;
      RECT 55.64 4.82 55.685 5.099 ;
      RECT 55.581 4.828 55.64 5.113 ;
      RECT 55.495 4.835 55.581 5.132 ;
      RECT 55.47 4.84 55.495 5.147 ;
      RECT 55.39 4.843 55.47 5.15 ;
      RECT 55.31 4.847 55.39 5.137 ;
      RECT 55.301 4.85 55.31 5.122 ;
      RECT 55.215 4.85 55.301 5.107 ;
      RECT 55.155 4.852 55.215 5.084 ;
      RECT 55.151 4.855 55.155 5.074 ;
      RECT 55.065 4.855 55.151 5.059 ;
      RECT 54.99 4.855 55.065 5.035 ;
      RECT 56.305 3.864 56.315 4.04 ;
      RECT 56.26 3.831 56.305 4.04 ;
      RECT 56.215 3.782 56.26 4.04 ;
      RECT 56.185 3.752 56.215 4.041 ;
      RECT 56.18 3.735 56.185 4.042 ;
      RECT 56.155 3.715 56.18 4.043 ;
      RECT 56.14 3.69 56.155 4.044 ;
      RECT 56.135 3.677 56.14 4.045 ;
      RECT 56.13 3.671 56.135 4.043 ;
      RECT 56.125 3.663 56.13 4.037 ;
      RECT 56.1 3.655 56.125 4.017 ;
      RECT 56.08 3.644 56.1 3.988 ;
      RECT 56.05 3.629 56.08 3.959 ;
      RECT 56.03 3.615 56.05 3.931 ;
      RECT 56.02 3.609 56.03 3.91 ;
      RECT 56.015 3.606 56.02 3.893 ;
      RECT 56.01 3.603 56.015 3.878 ;
      RECT 55.995 3.598 56.01 3.843 ;
      RECT 55.99 3.594 55.995 3.81 ;
      RECT 55.97 3.589 55.99 3.786 ;
      RECT 55.94 3.581 55.97 3.751 ;
      RECT 55.925 3.575 55.94 3.728 ;
      RECT 55.885 3.568 55.925 3.713 ;
      RECT 55.86 3.56 55.885 3.693 ;
      RECT 55.84 3.555 55.86 3.683 ;
      RECT 55.805 3.549 55.84 3.678 ;
      RECT 55.76 3.54 55.805 3.677 ;
      RECT 55.73 3.536 55.76 3.679 ;
      RECT 55.645 3.544 55.73 3.683 ;
      RECT 55.575 3.555 55.645 3.705 ;
      RECT 55.562 3.561 55.575 3.728 ;
      RECT 55.476 3.568 55.562 3.75 ;
      RECT 55.39 3.58 55.476 3.787 ;
      RECT 55.39 3.957 55.4 4.195 ;
      RECT 55.385 3.586 55.39 3.81 ;
      RECT 55.38 3.842 55.39 4.195 ;
      RECT 55.38 3.587 55.385 3.815 ;
      RECT 55.375 3.588 55.38 4.195 ;
      RECT 55.351 3.59 55.375 4.196 ;
      RECT 55.265 3.598 55.351 4.198 ;
      RECT 55.245 3.612 55.265 4.201 ;
      RECT 55.24 3.64 55.245 4.202 ;
      RECT 55.235 3.652 55.24 4.203 ;
      RECT 55.23 3.667 55.235 4.204 ;
      RECT 55.22 3.697 55.23 4.205 ;
      RECT 55.215 3.735 55.22 4.203 ;
      RECT 55.21 3.755 55.215 4.198 ;
      RECT 55.195 3.79 55.21 4.183 ;
      RECT 55.185 3.842 55.195 4.163 ;
      RECT 55.18 3.872 55.185 4.151 ;
      RECT 55.165 3.885 55.18 4.134 ;
      RECT 55.14 3.889 55.165 4.101 ;
      RECT 55.125 3.887 55.14 4.078 ;
      RECT 55.11 3.886 55.125 4.075 ;
      RECT 55.05 3.884 55.11 4.073 ;
      RECT 55.04 3.882 55.05 4.068 ;
      RECT 55 3.881 55.04 4.065 ;
      RECT 54.93 3.878 55 4.063 ;
      RECT 54.875 3.876 54.93 4.058 ;
      RECT 54.805 3.87 54.875 4.053 ;
      RECT 54.796 3.87 54.805 4.05 ;
      RECT 54.71 3.87 54.796 4.045 ;
      RECT 54.705 3.87 54.71 4.04 ;
      RECT 56.01 3.105 56.185 3.455 ;
      RECT 56.01 3.12 56.195 3.453 ;
      RECT 55.985 3.07 56.13 3.45 ;
      RECT 55.965 3.071 56.13 3.443 ;
      RECT 55.955 3.072 56.14 3.438 ;
      RECT 55.925 3.073 56.14 3.425 ;
      RECT 55.875 3.074 56.14 3.401 ;
      RECT 55.87 3.076 56.14 3.386 ;
      RECT 55.87 3.142 56.2 3.38 ;
      RECT 55.85 3.083 56.155 3.36 ;
      RECT 55.84 3.092 56.165 3.215 ;
      RECT 55.85 3.087 56.165 3.36 ;
      RECT 55.87 3.077 56.155 3.386 ;
      RECT 55.455 4.402 55.625 4.69 ;
      RECT 55.45 4.42 55.635 4.685 ;
      RECT 55.415 4.428 55.7 4.605 ;
      RECT 55.415 4.428 55.786 4.595 ;
      RECT 55.415 4.428 55.84 4.541 ;
      RECT 55.7 4.325 55.87 4.509 ;
      RECT 55.415 4.48 55.875 4.497 ;
      RECT 55.4 4.45 55.87 4.493 ;
      RECT 55.66 4.332 55.7 4.644 ;
      RECT 55.54 4.369 55.87 4.509 ;
      RECT 55.635 4.344 55.66 4.67 ;
      RECT 55.625 4.351 55.87 4.509 ;
      RECT 55.756 3.815 55.825 4.074 ;
      RECT 55.756 3.87 55.83 4.073 ;
      RECT 55.67 3.87 55.83 4.072 ;
      RECT 55.665 3.87 55.835 4.065 ;
      RECT 55.655 3.815 55.825 4.06 ;
      RECT 55.035 3.114 55.21 3.415 ;
      RECT 55.02 3.102 55.035 3.4 ;
      RECT 54.99 3.101 55.02 3.353 ;
      RECT 54.99 3.119 55.215 3.348 ;
      RECT 54.975 3.103 55.035 3.313 ;
      RECT 54.97 3.125 55.225 3.213 ;
      RECT 54.97 3.108 55.121 3.213 ;
      RECT 54.97 3.11 55.125 3.213 ;
      RECT 54.975 3.106 55.121 3.313 ;
      RECT 55.08 4.342 55.085 4.69 ;
      RECT 55.07 4.332 55.08 4.696 ;
      RECT 55.035 4.322 55.07 4.698 ;
      RECT 54.997 4.317 55.035 4.702 ;
      RECT 54.911 4.31 54.997 4.709 ;
      RECT 54.825 4.3 54.911 4.719 ;
      RECT 54.78 4.295 54.825 4.727 ;
      RECT 54.776 4.295 54.78 4.731 ;
      RECT 54.69 4.295 54.776 4.738 ;
      RECT 54.675 4.295 54.69 4.738 ;
      RECT 54.665 4.293 54.675 4.71 ;
      RECT 54.655 4.289 54.665 4.653 ;
      RECT 54.635 4.283 54.655 4.585 ;
      RECT 54.63 4.279 54.635 4.533 ;
      RECT 54.62 4.278 54.63 4.5 ;
      RECT 54.57 4.276 54.62 4.485 ;
      RECT 54.545 4.274 54.57 4.48 ;
      RECT 54.502 4.272 54.545 4.476 ;
      RECT 54.416 4.268 54.502 4.464 ;
      RECT 54.33 4.263 54.416 4.448 ;
      RECT 54.3 4.26 54.33 4.435 ;
      RECT 54.275 4.259 54.3 4.423 ;
      RECT 54.27 4.259 54.275 4.413 ;
      RECT 54.23 4.258 54.27 4.405 ;
      RECT 54.215 4.257 54.23 4.398 ;
      RECT 54.165 4.256 54.215 4.39 ;
      RECT 54.163 4.255 54.165 4.385 ;
      RECT 54.077 4.253 54.163 4.385 ;
      RECT 53.991 4.248 54.077 4.385 ;
      RECT 53.905 4.244 53.991 4.385 ;
      RECT 53.856 4.24 53.905 4.383 ;
      RECT 53.77 4.237 53.856 4.378 ;
      RECT 53.747 4.234 53.77 4.374 ;
      RECT 53.661 4.231 53.747 4.369 ;
      RECT 53.575 4.227 53.661 4.36 ;
      RECT 53.55 4.22 53.575 4.355 ;
      RECT 53.49 4.185 53.55 4.352 ;
      RECT 53.47 4.11 53.49 4.349 ;
      RECT 53.465 4.052 53.47 4.348 ;
      RECT 53.44 3.992 53.465 4.347 ;
      RECT 53.365 3.87 53.44 4.343 ;
      RECT 53.355 3.87 53.365 4.335 ;
      RECT 53.34 3.87 53.355 4.325 ;
      RECT 53.325 3.87 53.34 4.295 ;
      RECT 53.31 3.87 53.325 4.24 ;
      RECT 53.295 3.87 53.31 4.178 ;
      RECT 53.27 3.87 53.295 4.103 ;
      RECT 53.265 3.87 53.27 4.053 ;
      RECT 54.61 3.415 54.63 3.724 ;
      RECT 54.596 3.417 54.645 3.721 ;
      RECT 54.596 3.422 54.665 3.712 ;
      RECT 54.51 3.42 54.645 3.706 ;
      RECT 54.51 3.428 54.7 3.689 ;
      RECT 54.475 3.43 54.7 3.688 ;
      RECT 54.445 3.438 54.7 3.679 ;
      RECT 54.435 3.443 54.72 3.665 ;
      RECT 54.475 3.433 54.72 3.665 ;
      RECT 54.475 3.436 54.73 3.653 ;
      RECT 54.445 3.438 54.74 3.64 ;
      RECT 54.445 3.442 54.75 3.583 ;
      RECT 54.435 3.447 54.755 3.498 ;
      RECT 54.596 3.415 54.63 3.721 ;
      RECT 54.035 3.518 54.04 3.73 ;
      RECT 53.91 3.515 53.925 3.73 ;
      RECT 53.375 3.545 53.445 3.73 ;
      RECT 53.26 3.545 53.295 3.725 ;
      RECT 54.381 3.847 54.4 4.041 ;
      RECT 54.295 3.802 54.381 4.042 ;
      RECT 54.285 3.755 54.295 4.044 ;
      RECT 54.28 3.735 54.285 4.045 ;
      RECT 54.26 3.7 54.28 4.046 ;
      RECT 54.245 3.65 54.26 4.047 ;
      RECT 54.225 3.587 54.245 4.048 ;
      RECT 54.215 3.55 54.225 4.049 ;
      RECT 54.2 3.539 54.215 4.05 ;
      RECT 54.195 3.531 54.2 4.048 ;
      RECT 54.185 3.53 54.195 4.04 ;
      RECT 54.155 3.527 54.185 4.019 ;
      RECT 54.08 3.522 54.155 3.964 ;
      RECT 54.065 3.518 54.08 3.91 ;
      RECT 54.055 3.518 54.065 3.805 ;
      RECT 54.04 3.518 54.055 3.738 ;
      RECT 54.025 3.518 54.035 3.728 ;
      RECT 53.97 3.517 54.025 3.725 ;
      RECT 53.925 3.515 53.97 3.728 ;
      RECT 53.897 3.515 53.91 3.731 ;
      RECT 53.811 3.519 53.897 3.733 ;
      RECT 53.725 3.525 53.811 3.738 ;
      RECT 53.705 3.529 53.725 3.74 ;
      RECT 53.703 3.53 53.705 3.739 ;
      RECT 53.617 3.532 53.703 3.738 ;
      RECT 53.531 3.537 53.617 3.735 ;
      RECT 53.445 3.542 53.531 3.732 ;
      RECT 53.295 3.545 53.375 3.728 ;
      RECT 53.955 7.305 54.125 10.595 ;
      RECT 53.955 9.605 54.36 9.935 ;
      RECT 53.955 8.765 54.36 9.095 ;
      RECT 54.071 4.52 54.12 4.854 ;
      RECT 54.071 4.52 54.125 4.853 ;
      RECT 53.985 4.52 54.125 4.852 ;
      RECT 53.76 4.628 54.13 4.85 ;
      RECT 53.985 4.52 54.155 4.843 ;
      RECT 53.955 4.532 54.16 4.834 ;
      RECT 53.94 4.55 54.165 4.831 ;
      RECT 53.755 4.634 54.165 4.758 ;
      RECT 53.75 4.641 54.165 4.718 ;
      RECT 53.765 4.607 54.165 4.831 ;
      RECT 53.926 4.553 54.13 4.85 ;
      RECT 53.84 4.573 54.165 4.831 ;
      RECT 53.94 4.547 54.16 4.834 ;
      RECT 53.71 3.871 53.9 4.065 ;
      RECT 53.705 3.873 53.9 4.064 ;
      RECT 53.7 3.877 53.915 4.061 ;
      RECT 53.715 3.87 53.915 4.061 ;
      RECT 53.7 3.98 53.92 4.056 ;
      RECT 52.995 4.48 53.086 4.778 ;
      RECT 52.99 4.482 53.165 4.773 ;
      RECT 52.995 4.48 53.165 4.773 ;
      RECT 52.99 4.486 53.185 4.771 ;
      RECT 52.99 4.541 53.225 4.77 ;
      RECT 52.99 4.576 53.24 4.764 ;
      RECT 52.99 4.61 53.25 4.754 ;
      RECT 52.98 4.49 53.185 4.605 ;
      RECT 52.98 4.51 53.2 4.605 ;
      RECT 52.98 4.493 53.19 4.605 ;
      RECT 53.205 3.261 53.21 3.323 ;
      RECT 53.2 3.183 53.205 3.346 ;
      RECT 53.195 3.14 53.2 3.357 ;
      RECT 53.19 3.13 53.195 3.369 ;
      RECT 53.185 3.13 53.19 3.378 ;
      RECT 53.16 3.13 53.185 3.41 ;
      RECT 53.155 3.13 53.16 3.443 ;
      RECT 53.14 3.13 53.155 3.468 ;
      RECT 53.13 3.13 53.14 3.495 ;
      RECT 53.125 3.13 53.13 3.508 ;
      RECT 53.12 3.13 53.125 3.523 ;
      RECT 53.11 3.13 53.12 3.538 ;
      RECT 53.105 3.13 53.11 3.558 ;
      RECT 53.08 3.13 53.105 3.593 ;
      RECT 53.035 3.13 53.08 3.638 ;
      RECT 53.025 3.13 53.035 3.651 ;
      RECT 52.94 3.215 53.025 3.658 ;
      RECT 52.905 3.337 52.94 3.667 ;
      RECT 52.9 3.377 52.905 3.671 ;
      RECT 52.88 3.4 52.9 3.673 ;
      RECT 52.875 3.43 52.88 3.676 ;
      RECT 52.865 3.442 52.875 3.677 ;
      RECT 52.82 3.465 52.865 3.682 ;
      RECT 52.78 3.495 52.82 3.69 ;
      RECT 52.745 3.507 52.78 3.696 ;
      RECT 52.74 3.512 52.745 3.7 ;
      RECT 52.67 3.522 52.74 3.707 ;
      RECT 52.63 3.532 52.67 3.717 ;
      RECT 52.61 3.537 52.63 3.723 ;
      RECT 52.6 3.541 52.61 3.728 ;
      RECT 52.595 3.544 52.6 3.731 ;
      RECT 52.585 3.545 52.595 3.732 ;
      RECT 52.56 3.547 52.585 3.736 ;
      RECT 52.55 3.552 52.56 3.739 ;
      RECT 52.505 3.56 52.55 3.74 ;
      RECT 52.38 3.565 52.505 3.74 ;
      RECT 52.935 3.862 52.955 4.044 ;
      RECT 52.886 3.847 52.935 4.043 ;
      RECT 52.8 3.862 52.955 4.041 ;
      RECT 52.785 3.862 52.955 4.04 ;
      RECT 52.75 3.84 52.92 4.025 ;
      RECT 52.82 4.86 52.835 5.069 ;
      RECT 52.82 4.868 52.84 5.068 ;
      RECT 52.765 4.868 52.84 5.067 ;
      RECT 52.745 4.872 52.845 5.065 ;
      RECT 52.725 4.822 52.765 5.064 ;
      RECT 52.67 4.88 52.85 5.062 ;
      RECT 52.635 4.837 52.765 5.06 ;
      RECT 52.631 4.84 52.82 5.059 ;
      RECT 52.545 4.848 52.82 5.057 ;
      RECT 52.545 4.892 52.855 5.05 ;
      RECT 52.535 4.985 52.855 5.048 ;
      RECT 52.545 4.904 52.86 5.033 ;
      RECT 52.545 4.925 52.875 5.003 ;
      RECT 52.545 4.952 52.88 4.973 ;
      RECT 52.67 4.83 52.765 5.062 ;
      RECT 52.3 3.875 52.305 4.413 ;
      RECT 52.105 4.205 52.11 4.4 ;
      RECT 50.405 3.87 50.42 4.25 ;
      RECT 52.47 3.87 52.475 4.04 ;
      RECT 52.465 3.87 52.47 4.05 ;
      RECT 52.46 3.87 52.465 4.063 ;
      RECT 52.435 3.87 52.46 4.105 ;
      RECT 52.41 3.87 52.435 4.178 ;
      RECT 52.395 3.87 52.41 4.23 ;
      RECT 52.39 3.87 52.395 4.26 ;
      RECT 52.365 3.87 52.39 4.3 ;
      RECT 52.35 3.87 52.365 4.355 ;
      RECT 52.345 3.87 52.35 4.388 ;
      RECT 52.32 3.87 52.345 4.408 ;
      RECT 52.305 3.87 52.32 4.414 ;
      RECT 52.235 3.905 52.3 4.41 ;
      RECT 52.185 3.96 52.235 4.405 ;
      RECT 52.175 3.992 52.185 4.403 ;
      RECT 52.17 4.017 52.175 4.403 ;
      RECT 52.15 4.09 52.17 4.403 ;
      RECT 52.14 4.17 52.15 4.402 ;
      RECT 52.125 4.2 52.14 4.402 ;
      RECT 52.11 4.205 52.125 4.401 ;
      RECT 52.05 4.207 52.105 4.398 ;
      RECT 52.02 4.212 52.05 4.394 ;
      RECT 52.018 4.215 52.02 4.393 ;
      RECT 51.932 4.217 52.018 4.39 ;
      RECT 51.846 4.223 51.932 4.384 ;
      RECT 51.76 4.228 51.846 4.378 ;
      RECT 51.687 4.233 51.76 4.379 ;
      RECT 51.601 4.239 51.687 4.387 ;
      RECT 51.515 4.245 51.601 4.396 ;
      RECT 51.495 4.249 51.515 4.401 ;
      RECT 51.448 4.251 51.495 4.404 ;
      RECT 51.362 4.256 51.448 4.41 ;
      RECT 51.276 4.261 51.362 4.419 ;
      RECT 51.19 4.267 51.276 4.427 ;
      RECT 51.105 4.265 51.19 4.436 ;
      RECT 51.101 4.26 51.105 4.44 ;
      RECT 51.015 4.255 51.101 4.432 ;
      RECT 50.951 4.246 51.015 4.42 ;
      RECT 50.865 4.237 50.951 4.407 ;
      RECT 50.841 4.23 50.865 4.398 ;
      RECT 50.755 4.224 50.841 4.385 ;
      RECT 50.715 4.217 50.755 4.371 ;
      RECT 50.71 4.207 50.715 4.367 ;
      RECT 50.7 4.195 50.71 4.366 ;
      RECT 50.68 4.165 50.7 4.363 ;
      RECT 50.625 4.085 50.68 4.357 ;
      RECT 50.605 4.004 50.625 4.352 ;
      RECT 50.585 3.962 50.605 4.348 ;
      RECT 50.56 3.915 50.585 4.342 ;
      RECT 50.555 3.89 50.56 4.339 ;
      RECT 50.52 3.87 50.555 4.334 ;
      RECT 50.511 3.87 50.52 4.327 ;
      RECT 50.425 3.87 50.511 4.297 ;
      RECT 50.42 3.87 50.425 4.26 ;
      RECT 50.385 3.87 50.405 4.182 ;
      RECT 50.38 3.912 50.385 4.147 ;
      RECT 50.375 3.987 50.38 4.103 ;
      RECT 51.825 3.792 52 4.04 ;
      RECT 51.825 3.792 52.005 4.038 ;
      RECT 51.82 3.824 52.005 3.998 ;
      RECT 51.85 3.765 52.02 3.985 ;
      RECT 51.815 3.842 52.02 3.918 ;
      RECT 51.125 3.305 51.295 3.48 ;
      RECT 51.125 3.305 51.467 3.472 ;
      RECT 51.125 3.305 51.55 3.466 ;
      RECT 51.125 3.305 51.585 3.462 ;
      RECT 51.125 3.305 51.605 3.461 ;
      RECT 51.125 3.305 51.691 3.457 ;
      RECT 51.585 3.13 51.755 3.452 ;
      RECT 51.16 3.237 51.785 3.45 ;
      RECT 51.15 3.292 51.79 3.448 ;
      RECT 51.125 3.328 51.8 3.443 ;
      RECT 51.125 3.355 51.805 3.373 ;
      RECT 51.19 3.18 51.765 3.45 ;
      RECT 51.381 3.165 51.765 3.45 ;
      RECT 51.215 3.168 51.765 3.45 ;
      RECT 51.295 3.166 51.381 3.477 ;
      RECT 51.381 3.163 51.76 3.45 ;
      RECT 51.565 3.14 51.76 3.45 ;
      RECT 51.467 3.161 51.76 3.45 ;
      RECT 51.55 3.155 51.565 3.463 ;
      RECT 51.7 4.52 51.705 4.72 ;
      RECT 51.165 4.585 51.21 4.72 ;
      RECT 51.735 4.52 51.755 4.693 ;
      RECT 51.705 4.52 51.735 4.708 ;
      RECT 51.64 4.52 51.7 4.745 ;
      RECT 51.625 4.52 51.64 4.775 ;
      RECT 51.61 4.52 51.625 4.788 ;
      RECT 51.59 4.52 51.61 4.803 ;
      RECT 51.585 4.52 51.59 4.812 ;
      RECT 51.575 4.524 51.585 4.817 ;
      RECT 51.56 4.534 51.575 4.828 ;
      RECT 51.535 4.55 51.56 4.838 ;
      RECT 51.525 4.564 51.535 4.84 ;
      RECT 51.505 4.576 51.525 4.837 ;
      RECT 51.475 4.597 51.505 4.831 ;
      RECT 51.465 4.609 51.475 4.826 ;
      RECT 51.455 4.607 51.465 4.823 ;
      RECT 51.44 4.606 51.455 4.818 ;
      RECT 51.435 4.605 51.44 4.813 ;
      RECT 51.4 4.603 51.435 4.803 ;
      RECT 51.38 4.6 51.4 4.785 ;
      RECT 51.37 4.598 51.38 4.78 ;
      RECT 51.36 4.597 51.37 4.775 ;
      RECT 51.325 4.595 51.36 4.763 ;
      RECT 51.27 4.591 51.325 4.743 ;
      RECT 51.26 4.589 51.27 4.728 ;
      RECT 51.255 4.589 51.26 4.723 ;
      RECT 51.21 4.587 51.255 4.72 ;
      RECT 51.115 4.585 51.165 4.724 ;
      RECT 51.105 4.586 51.115 4.729 ;
      RECT 51.045 4.593 51.105 4.743 ;
      RECT 51.02 4.601 51.045 4.763 ;
      RECT 51.01 4.605 51.02 4.775 ;
      RECT 51.005 4.606 51.01 4.78 ;
      RECT 50.99 4.608 51.005 4.783 ;
      RECT 50.975 4.61 50.99 4.788 ;
      RECT 50.97 4.61 50.975 4.791 ;
      RECT 50.925 4.615 50.97 4.802 ;
      RECT 50.92 4.619 50.925 4.814 ;
      RECT 50.895 4.615 50.92 4.818 ;
      RECT 50.885 4.611 50.895 4.822 ;
      RECT 50.875 4.61 50.885 4.826 ;
      RECT 50.86 4.6 50.875 4.832 ;
      RECT 50.855 4.588 50.86 4.836 ;
      RECT 50.85 4.585 50.855 4.837 ;
      RECT 50.845 4.582 50.85 4.839 ;
      RECT 50.83 4.57 50.845 4.838 ;
      RECT 50.815 4.552 50.83 4.835 ;
      RECT 50.795 4.531 50.815 4.828 ;
      RECT 50.73 4.52 50.795 4.8 ;
      RECT 50.726 4.52 50.73 4.779 ;
      RECT 50.64 4.52 50.726 4.749 ;
      RECT 50.625 4.52 50.64 4.705 ;
      RECT 51.2 3.62 51.205 3.855 ;
      RECT 50.33 3.536 50.335 3.74 ;
      RECT 50.91 3.565 50.915 3.72 ;
      RECT 50.83 3.545 50.835 3.72 ;
      RECT 51.5 3.687 51.515 4.04 ;
      RECT 51.426 3.672 51.5 4.04 ;
      RECT 51.34 3.655 51.426 4.04 ;
      RECT 51.33 3.645 51.34 4.038 ;
      RECT 51.325 3.643 51.33 4.033 ;
      RECT 51.31 3.641 51.325 4.019 ;
      RECT 51.24 3.633 51.31 3.959 ;
      RECT 51.22 3.624 51.24 3.893 ;
      RECT 51.215 3.621 51.22 3.873 ;
      RECT 51.205 3.62 51.215 3.863 ;
      RECT 51.195 3.62 51.2 3.847 ;
      RECT 51.185 3.619 51.195 3.837 ;
      RECT 51.175 3.617 51.185 3.825 ;
      RECT 51.16 3.614 51.175 3.805 ;
      RECT 51.15 3.612 51.16 3.79 ;
      RECT 51.13 3.609 51.15 3.778 ;
      RECT 51.125 3.607 51.13 3.768 ;
      RECT 51.1 3.605 51.125 3.755 ;
      RECT 51.07 3.6 51.1 3.74 ;
      RECT 50.99 3.591 51.07 3.731 ;
      RECT 50.945 3.58 50.99 3.724 ;
      RECT 50.925 3.571 50.945 3.721 ;
      RECT 50.915 3.566 50.925 3.72 ;
      RECT 50.87 3.56 50.91 3.72 ;
      RECT 50.855 3.552 50.87 3.72 ;
      RECT 50.835 3.547 50.855 3.72 ;
      RECT 50.815 3.544 50.83 3.72 ;
      RECT 50.732 3.543 50.815 3.719 ;
      RECT 50.646 3.542 50.732 3.715 ;
      RECT 50.56 3.54 50.646 3.712 ;
      RECT 50.507 3.539 50.56 3.714 ;
      RECT 50.421 3.538 50.507 3.723 ;
      RECT 50.335 3.537 50.421 3.735 ;
      RECT 50.315 3.536 50.33 3.743 ;
      RECT 50.235 3.535 50.315 3.755 ;
      RECT 50.21 3.535 50.235 3.768 ;
      RECT 50.185 3.535 50.21 3.783 ;
      RECT 50.18 3.535 50.185 3.805 ;
      RECT 50.175 3.535 50.18 3.823 ;
      RECT 50.17 3.535 50.175 3.84 ;
      RECT 50.165 3.535 50.17 3.853 ;
      RECT 50.16 3.535 50.165 3.863 ;
      RECT 50.12 3.535 50.16 3.948 ;
      RECT 50.105 3.535 50.12 4.033 ;
      RECT 50.095 3.536 50.105 4.045 ;
      RECT 50.06 3.541 50.095 4.05 ;
      RECT 50.02 3.55 50.06 4.05 ;
      RECT 50.005 3.56 50.02 4.05 ;
      RECT 50 3.57 50.005 4.05 ;
      RECT 49.98 3.597 50 4.05 ;
      RECT 49.93 3.68 49.98 4.05 ;
      RECT 49.925 3.742 49.93 4.05 ;
      RECT 49.915 3.755 49.925 4.05 ;
      RECT 49.905 3.777 49.915 4.05 ;
      RECT 49.895 3.802 49.905 4.045 ;
      RECT 49.89 3.84 49.895 4.038 ;
      RECT 49.88 3.95 49.89 4.033 ;
      RECT 51.275 4.871 51.29 5.13 ;
      RECT 51.275 4.886 51.295 5.129 ;
      RECT 51.191 4.886 51.295 5.127 ;
      RECT 51.191 4.9 51.3 5.126 ;
      RECT 51.105 4.942 51.305 5.123 ;
      RECT 51.1 4.885 51.29 5.118 ;
      RECT 51.1 4.956 51.31 5.115 ;
      RECT 51.095 4.987 51.31 5.113 ;
      RECT 51.1 4.984 51.325 5.103 ;
      RECT 51.095 5.03 51.34 5.088 ;
      RECT 51.095 5.058 51.345 5.073 ;
      RECT 51.105 4.86 51.275 5.123 ;
      RECT 50.865 3.87 51.035 4.04 ;
      RECT 50.83 3.87 51.035 4.035 ;
      RECT 50.82 3.87 51.035 4.028 ;
      RECT 50.815 3.855 50.985 4.025 ;
      RECT 49.645 4.392 49.91 4.835 ;
      RECT 49.64 4.363 49.855 4.833 ;
      RECT 49.635 4.517 49.915 4.828 ;
      RECT 49.64 4.412 49.915 4.828 ;
      RECT 49.64 4.423 49.925 4.815 ;
      RECT 49.64 4.37 49.885 4.833 ;
      RECT 49.645 4.357 49.855 4.835 ;
      RECT 49.645 4.355 49.805 4.835 ;
      RECT 49.746 4.347 49.805 4.835 ;
      RECT 49.66 4.348 49.805 4.835 ;
      RECT 49.746 4.346 49.795 4.835 ;
      RECT 49.55 3.161 49.725 3.46 ;
      RECT 49.6 3.123 49.725 3.46 ;
      RECT 49.585 3.125 49.811 3.452 ;
      RECT 49.585 3.128 49.85 3.439 ;
      RECT 49.585 3.129 49.86 3.425 ;
      RECT 49.54 3.18 49.86 3.415 ;
      RECT 49.585 3.13 49.865 3.41 ;
      RECT 49.54 3.34 49.87 3.4 ;
      RECT 49.525 3.2 49.865 3.34 ;
      RECT 49.52 3.216 49.865 3.28 ;
      RECT 49.565 3.14 49.865 3.41 ;
      RECT 49.6 3.121 49.686 3.46 ;
      RECT 47.69 3.035 47.86 4.225 ;
      RECT 47.69 3.035 48.16 3.205 ;
      RECT 47.69 9.26 48.16 9.43 ;
      RECT 47.69 8.24 47.86 9.43 ;
      RECT 46.7 3.035 46.87 4.225 ;
      RECT 46.7 3.035 47.17 3.205 ;
      RECT 46.7 9.26 47.17 9.43 ;
      RECT 46.7 8.24 46.87 9.43 ;
      RECT 44.85 3.93 45.02 5.16 ;
      RECT 44.905 2.15 45.075 4.1 ;
      RECT 44.85 1.87 45.02 2.32 ;
      RECT 44.85 10.145 45.02 10.595 ;
      RECT 44.905 8.365 45.075 10.315 ;
      RECT 44.85 7.305 45.02 8.535 ;
      RECT 44.33 1.87 44.5 5.16 ;
      RECT 44.33 3.37 44.735 3.7 ;
      RECT 44.33 2.53 44.735 2.86 ;
      RECT 44.33 7.305 44.5 10.595 ;
      RECT 44.33 9.605 44.735 9.935 ;
      RECT 44.33 8.765 44.735 9.095 ;
      RECT 42.255 4.421 42.26 4.593 ;
      RECT 42.25 4.414 42.255 4.683 ;
      RECT 42.245 4.408 42.25 4.702 ;
      RECT 42.225 4.402 42.245 4.712 ;
      RECT 42.21 4.397 42.225 4.72 ;
      RECT 42.173 4.391 42.21 4.718 ;
      RECT 42.087 4.377 42.173 4.714 ;
      RECT 42.001 4.359 42.087 4.709 ;
      RECT 41.915 4.34 42.001 4.703 ;
      RECT 41.885 4.328 41.915 4.699 ;
      RECT 41.865 4.322 41.885 4.698 ;
      RECT 41.8 4.32 41.865 4.696 ;
      RECT 41.785 4.32 41.8 4.688 ;
      RECT 41.77 4.32 41.785 4.675 ;
      RECT 41.765 4.32 41.77 4.665 ;
      RECT 41.75 4.32 41.765 4.643 ;
      RECT 41.735 4.32 41.75 4.61 ;
      RECT 41.73 4.32 41.735 4.588 ;
      RECT 41.72 4.32 41.73 4.57 ;
      RECT 41.705 4.32 41.72 4.548 ;
      RECT 41.685 4.32 41.705 4.51 ;
      RECT 42.035 3.605 42.07 4.044 ;
      RECT 42.035 3.605 42.075 4.043 ;
      RECT 41.98 3.665 42.075 4.042 ;
      RECT 41.845 3.837 42.075 4.041 ;
      RECT 41.955 3.715 42.075 4.041 ;
      RECT 41.845 3.837 42.1 4.031 ;
      RECT 41.9 3.782 42.18 3.948 ;
      RECT 42.075 3.576 42.08 4.039 ;
      RECT 41.93 3.752 42.22 3.825 ;
      RECT 41.945 3.735 42.075 4.041 ;
      RECT 42.08 3.575 42.25 3.763 ;
      RECT 42.07 3.578 42.25 3.763 ;
      RECT 41.575 3.455 41.745 3.765 ;
      RECT 41.575 3.455 41.75 3.738 ;
      RECT 41.575 3.455 41.755 3.715 ;
      RECT 41.575 3.455 41.765 3.665 ;
      RECT 41.57 3.56 41.765 3.635 ;
      RECT 41.605 3.13 41.775 3.608 ;
      RECT 41.605 3.13 41.79 3.529 ;
      RECT 41.595 3.34 41.79 3.529 ;
      RECT 41.605 3.14 41.8 3.444 ;
      RECT 41.535 3.882 41.54 4.085 ;
      RECT 41.525 3.87 41.535 4.195 ;
      RECT 41.5 3.87 41.525 4.235 ;
      RECT 41.42 3.87 41.5 4.32 ;
      RECT 41.41 3.87 41.42 4.39 ;
      RECT 41.385 3.87 41.41 4.413 ;
      RECT 41.365 3.87 41.385 4.448 ;
      RECT 41.32 3.88 41.365 4.491 ;
      RECT 41.31 3.892 41.32 4.528 ;
      RECT 41.29 3.906 41.31 4.548 ;
      RECT 41.28 3.924 41.29 4.564 ;
      RECT 41.265 3.95 41.28 4.574 ;
      RECT 41.25 3.991 41.265 4.588 ;
      RECT 41.24 4.026 41.25 4.598 ;
      RECT 41.235 4.042 41.24 4.603 ;
      RECT 41.225 4.057 41.235 4.608 ;
      RECT 41.205 4.1 41.225 4.618 ;
      RECT 41.185 4.137 41.205 4.631 ;
      RECT 41.15 4.16 41.185 4.649 ;
      RECT 41.14 4.174 41.15 4.665 ;
      RECT 41.12 4.184 41.14 4.675 ;
      RECT 41.115 4.193 41.12 4.683 ;
      RECT 41.105 4.2 41.115 4.69 ;
      RECT 41.095 4.207 41.105 4.698 ;
      RECT 41.08 4.217 41.095 4.706 ;
      RECT 41.07 4.231 41.08 4.716 ;
      RECT 41.06 4.243 41.07 4.728 ;
      RECT 41.045 4.265 41.06 4.741 ;
      RECT 41.035 4.287 41.045 4.752 ;
      RECT 41.025 4.307 41.035 4.761 ;
      RECT 41.02 4.322 41.025 4.768 ;
      RECT 40.99 4.355 41.02 4.782 ;
      RECT 40.98 4.39 40.99 4.797 ;
      RECT 40.975 4.397 40.98 4.803 ;
      RECT 40.955 4.412 40.975 4.81 ;
      RECT 40.95 4.427 40.955 4.818 ;
      RECT 40.945 4.436 40.95 4.823 ;
      RECT 40.93 4.442 40.945 4.83 ;
      RECT 40.925 4.448 40.93 4.838 ;
      RECT 40.92 4.452 40.925 4.845 ;
      RECT 40.915 4.456 40.92 4.855 ;
      RECT 40.905 4.461 40.915 4.865 ;
      RECT 40.885 4.472 40.905 4.893 ;
      RECT 40.87 4.484 40.885 4.92 ;
      RECT 40.85 4.497 40.87 4.945 ;
      RECT 40.83 4.512 40.85 4.969 ;
      RECT 40.815 4.527 40.83 4.984 ;
      RECT 40.81 4.538 40.815 4.993 ;
      RECT 40.745 4.583 40.81 5.003 ;
      RECT 40.71 4.642 40.745 5.016 ;
      RECT 40.705 4.665 40.71 5.022 ;
      RECT 40.7 4.672 40.705 5.024 ;
      RECT 40.685 4.682 40.7 5.027 ;
      RECT 40.655 4.707 40.685 5.031 ;
      RECT 40.65 4.725 40.655 5.035 ;
      RECT 40.645 4.732 40.65 5.036 ;
      RECT 40.625 4.74 40.645 5.04 ;
      RECT 40.615 4.747 40.625 5.044 ;
      RECT 40.571 4.758 40.615 5.051 ;
      RECT 40.485 4.786 40.571 5.067 ;
      RECT 40.425 4.81 40.485 5.085 ;
      RECT 40.38 4.82 40.425 5.099 ;
      RECT 40.321 4.828 40.38 5.113 ;
      RECT 40.235 4.835 40.321 5.132 ;
      RECT 40.21 4.84 40.235 5.147 ;
      RECT 40.13 4.843 40.21 5.15 ;
      RECT 40.05 4.847 40.13 5.137 ;
      RECT 40.041 4.85 40.05 5.122 ;
      RECT 39.955 4.85 40.041 5.107 ;
      RECT 39.895 4.852 39.955 5.084 ;
      RECT 39.891 4.855 39.895 5.074 ;
      RECT 39.805 4.855 39.891 5.059 ;
      RECT 39.73 4.855 39.805 5.035 ;
      RECT 41.045 3.864 41.055 4.04 ;
      RECT 41 3.831 41.045 4.04 ;
      RECT 40.955 3.782 41 4.04 ;
      RECT 40.925 3.752 40.955 4.041 ;
      RECT 40.92 3.735 40.925 4.042 ;
      RECT 40.895 3.715 40.92 4.043 ;
      RECT 40.88 3.69 40.895 4.044 ;
      RECT 40.875 3.677 40.88 4.045 ;
      RECT 40.87 3.671 40.875 4.043 ;
      RECT 40.865 3.663 40.87 4.037 ;
      RECT 40.84 3.655 40.865 4.017 ;
      RECT 40.82 3.644 40.84 3.988 ;
      RECT 40.79 3.629 40.82 3.959 ;
      RECT 40.77 3.615 40.79 3.931 ;
      RECT 40.76 3.609 40.77 3.91 ;
      RECT 40.755 3.606 40.76 3.893 ;
      RECT 40.75 3.603 40.755 3.878 ;
      RECT 40.735 3.598 40.75 3.843 ;
      RECT 40.73 3.594 40.735 3.81 ;
      RECT 40.71 3.589 40.73 3.786 ;
      RECT 40.68 3.581 40.71 3.751 ;
      RECT 40.665 3.575 40.68 3.728 ;
      RECT 40.625 3.568 40.665 3.713 ;
      RECT 40.6 3.56 40.625 3.693 ;
      RECT 40.58 3.555 40.6 3.683 ;
      RECT 40.545 3.549 40.58 3.678 ;
      RECT 40.5 3.54 40.545 3.677 ;
      RECT 40.47 3.536 40.5 3.679 ;
      RECT 40.385 3.544 40.47 3.683 ;
      RECT 40.315 3.555 40.385 3.705 ;
      RECT 40.302 3.561 40.315 3.728 ;
      RECT 40.216 3.568 40.302 3.75 ;
      RECT 40.13 3.58 40.216 3.787 ;
      RECT 40.13 3.957 40.14 4.195 ;
      RECT 40.125 3.586 40.13 3.81 ;
      RECT 40.12 3.842 40.13 4.195 ;
      RECT 40.12 3.587 40.125 3.815 ;
      RECT 40.115 3.588 40.12 4.195 ;
      RECT 40.091 3.59 40.115 4.196 ;
      RECT 40.005 3.598 40.091 4.198 ;
      RECT 39.985 3.612 40.005 4.201 ;
      RECT 39.98 3.64 39.985 4.202 ;
      RECT 39.975 3.652 39.98 4.203 ;
      RECT 39.97 3.667 39.975 4.204 ;
      RECT 39.96 3.697 39.97 4.205 ;
      RECT 39.955 3.735 39.96 4.203 ;
      RECT 39.95 3.755 39.955 4.198 ;
      RECT 39.935 3.79 39.95 4.183 ;
      RECT 39.925 3.842 39.935 4.163 ;
      RECT 39.92 3.872 39.925 4.151 ;
      RECT 39.905 3.885 39.92 4.134 ;
      RECT 39.88 3.889 39.905 4.101 ;
      RECT 39.865 3.887 39.88 4.078 ;
      RECT 39.85 3.886 39.865 4.075 ;
      RECT 39.79 3.884 39.85 4.073 ;
      RECT 39.78 3.882 39.79 4.068 ;
      RECT 39.74 3.881 39.78 4.065 ;
      RECT 39.67 3.878 39.74 4.063 ;
      RECT 39.615 3.876 39.67 4.058 ;
      RECT 39.545 3.87 39.615 4.053 ;
      RECT 39.536 3.87 39.545 4.05 ;
      RECT 39.45 3.87 39.536 4.045 ;
      RECT 39.445 3.87 39.45 4.04 ;
      RECT 40.75 3.105 40.925 3.455 ;
      RECT 40.75 3.12 40.935 3.453 ;
      RECT 40.725 3.07 40.87 3.45 ;
      RECT 40.705 3.071 40.87 3.443 ;
      RECT 40.695 3.072 40.88 3.438 ;
      RECT 40.665 3.073 40.88 3.425 ;
      RECT 40.615 3.074 40.88 3.401 ;
      RECT 40.61 3.076 40.88 3.386 ;
      RECT 40.61 3.142 40.94 3.38 ;
      RECT 40.59 3.083 40.895 3.36 ;
      RECT 40.58 3.092 40.905 3.215 ;
      RECT 40.59 3.087 40.905 3.36 ;
      RECT 40.61 3.077 40.895 3.386 ;
      RECT 40.195 4.402 40.365 4.69 ;
      RECT 40.19 4.42 40.375 4.685 ;
      RECT 40.155 4.428 40.44 4.605 ;
      RECT 40.155 4.428 40.526 4.595 ;
      RECT 40.155 4.428 40.58 4.541 ;
      RECT 40.44 4.325 40.61 4.509 ;
      RECT 40.155 4.48 40.615 4.497 ;
      RECT 40.14 4.45 40.61 4.493 ;
      RECT 40.4 4.332 40.44 4.644 ;
      RECT 40.28 4.369 40.61 4.509 ;
      RECT 40.375 4.344 40.4 4.67 ;
      RECT 40.365 4.351 40.61 4.509 ;
      RECT 40.496 3.815 40.565 4.074 ;
      RECT 40.496 3.87 40.57 4.073 ;
      RECT 40.41 3.87 40.57 4.072 ;
      RECT 40.405 3.87 40.575 4.065 ;
      RECT 40.395 3.815 40.565 4.06 ;
      RECT 39.775 3.114 39.95 3.415 ;
      RECT 39.76 3.102 39.775 3.4 ;
      RECT 39.73 3.101 39.76 3.353 ;
      RECT 39.73 3.119 39.955 3.348 ;
      RECT 39.715 3.103 39.775 3.313 ;
      RECT 39.71 3.125 39.965 3.213 ;
      RECT 39.71 3.108 39.861 3.213 ;
      RECT 39.71 3.11 39.865 3.213 ;
      RECT 39.715 3.106 39.861 3.313 ;
      RECT 39.82 4.342 39.825 4.69 ;
      RECT 39.81 4.332 39.82 4.696 ;
      RECT 39.775 4.322 39.81 4.698 ;
      RECT 39.737 4.317 39.775 4.702 ;
      RECT 39.651 4.31 39.737 4.709 ;
      RECT 39.565 4.3 39.651 4.719 ;
      RECT 39.52 4.295 39.565 4.727 ;
      RECT 39.516 4.295 39.52 4.731 ;
      RECT 39.43 4.295 39.516 4.738 ;
      RECT 39.415 4.295 39.43 4.738 ;
      RECT 39.405 4.293 39.415 4.71 ;
      RECT 39.395 4.289 39.405 4.653 ;
      RECT 39.375 4.283 39.395 4.585 ;
      RECT 39.37 4.279 39.375 4.533 ;
      RECT 39.36 4.278 39.37 4.5 ;
      RECT 39.31 4.276 39.36 4.485 ;
      RECT 39.285 4.274 39.31 4.48 ;
      RECT 39.242 4.272 39.285 4.476 ;
      RECT 39.156 4.268 39.242 4.464 ;
      RECT 39.07 4.263 39.156 4.448 ;
      RECT 39.04 4.26 39.07 4.435 ;
      RECT 39.015 4.259 39.04 4.423 ;
      RECT 39.01 4.259 39.015 4.413 ;
      RECT 38.97 4.258 39.01 4.405 ;
      RECT 38.955 4.257 38.97 4.398 ;
      RECT 38.905 4.256 38.955 4.39 ;
      RECT 38.903 4.255 38.905 4.385 ;
      RECT 38.817 4.253 38.903 4.385 ;
      RECT 38.731 4.248 38.817 4.385 ;
      RECT 38.645 4.244 38.731 4.385 ;
      RECT 38.596 4.24 38.645 4.383 ;
      RECT 38.51 4.237 38.596 4.378 ;
      RECT 38.487 4.234 38.51 4.374 ;
      RECT 38.401 4.231 38.487 4.369 ;
      RECT 38.315 4.227 38.401 4.36 ;
      RECT 38.29 4.22 38.315 4.355 ;
      RECT 38.23 4.185 38.29 4.352 ;
      RECT 38.21 4.11 38.23 4.349 ;
      RECT 38.205 4.052 38.21 4.348 ;
      RECT 38.18 3.992 38.205 4.347 ;
      RECT 38.105 3.87 38.18 4.343 ;
      RECT 38.095 3.87 38.105 4.335 ;
      RECT 38.08 3.87 38.095 4.325 ;
      RECT 38.065 3.87 38.08 4.295 ;
      RECT 38.05 3.87 38.065 4.24 ;
      RECT 38.035 3.87 38.05 4.178 ;
      RECT 38.01 3.87 38.035 4.103 ;
      RECT 38.005 3.87 38.01 4.053 ;
      RECT 39.35 3.415 39.37 3.724 ;
      RECT 39.336 3.417 39.385 3.721 ;
      RECT 39.336 3.422 39.405 3.712 ;
      RECT 39.25 3.42 39.385 3.706 ;
      RECT 39.25 3.428 39.44 3.689 ;
      RECT 39.215 3.43 39.44 3.688 ;
      RECT 39.185 3.438 39.44 3.679 ;
      RECT 39.175 3.443 39.46 3.665 ;
      RECT 39.215 3.433 39.46 3.665 ;
      RECT 39.215 3.436 39.47 3.653 ;
      RECT 39.185 3.438 39.48 3.64 ;
      RECT 39.185 3.442 39.49 3.583 ;
      RECT 39.175 3.447 39.495 3.498 ;
      RECT 39.336 3.415 39.37 3.721 ;
      RECT 38.775 3.518 38.78 3.73 ;
      RECT 38.65 3.515 38.665 3.73 ;
      RECT 38.115 3.545 38.185 3.73 ;
      RECT 38 3.545 38.035 3.725 ;
      RECT 39.121 3.847 39.14 4.041 ;
      RECT 39.035 3.802 39.121 4.042 ;
      RECT 39.025 3.755 39.035 4.044 ;
      RECT 39.02 3.735 39.025 4.045 ;
      RECT 39 3.7 39.02 4.046 ;
      RECT 38.985 3.65 39 4.047 ;
      RECT 38.965 3.587 38.985 4.048 ;
      RECT 38.955 3.55 38.965 4.049 ;
      RECT 38.94 3.539 38.955 4.05 ;
      RECT 38.935 3.531 38.94 4.048 ;
      RECT 38.925 3.53 38.935 4.04 ;
      RECT 38.895 3.527 38.925 4.019 ;
      RECT 38.82 3.522 38.895 3.964 ;
      RECT 38.805 3.518 38.82 3.91 ;
      RECT 38.795 3.518 38.805 3.805 ;
      RECT 38.78 3.518 38.795 3.738 ;
      RECT 38.765 3.518 38.775 3.728 ;
      RECT 38.71 3.517 38.765 3.725 ;
      RECT 38.665 3.515 38.71 3.728 ;
      RECT 38.637 3.515 38.65 3.731 ;
      RECT 38.551 3.519 38.637 3.733 ;
      RECT 38.465 3.525 38.551 3.738 ;
      RECT 38.445 3.529 38.465 3.74 ;
      RECT 38.443 3.53 38.445 3.739 ;
      RECT 38.357 3.532 38.443 3.738 ;
      RECT 38.271 3.537 38.357 3.735 ;
      RECT 38.185 3.542 38.271 3.732 ;
      RECT 38.035 3.545 38.115 3.728 ;
      RECT 38.695 7.305 38.865 10.595 ;
      RECT 38.695 9.605 39.1 9.935 ;
      RECT 38.695 8.765 39.1 9.095 ;
      RECT 38.811 4.52 38.86 4.854 ;
      RECT 38.811 4.52 38.865 4.853 ;
      RECT 38.725 4.52 38.865 4.852 ;
      RECT 38.5 4.628 38.87 4.85 ;
      RECT 38.725 4.52 38.895 4.843 ;
      RECT 38.695 4.532 38.9 4.834 ;
      RECT 38.68 4.55 38.905 4.831 ;
      RECT 38.495 4.634 38.905 4.758 ;
      RECT 38.49 4.641 38.905 4.718 ;
      RECT 38.505 4.607 38.905 4.831 ;
      RECT 38.666 4.553 38.87 4.85 ;
      RECT 38.58 4.573 38.905 4.831 ;
      RECT 38.68 4.547 38.9 4.834 ;
      RECT 38.45 3.871 38.64 4.065 ;
      RECT 38.445 3.873 38.64 4.064 ;
      RECT 38.44 3.877 38.655 4.061 ;
      RECT 38.455 3.87 38.655 4.061 ;
      RECT 38.44 3.98 38.66 4.056 ;
      RECT 37.735 4.48 37.826 4.778 ;
      RECT 37.73 4.482 37.905 4.773 ;
      RECT 37.735 4.48 37.905 4.773 ;
      RECT 37.73 4.486 37.925 4.771 ;
      RECT 37.73 4.541 37.965 4.77 ;
      RECT 37.73 4.576 37.98 4.764 ;
      RECT 37.73 4.61 37.99 4.754 ;
      RECT 37.72 4.49 37.925 4.605 ;
      RECT 37.72 4.51 37.94 4.605 ;
      RECT 37.72 4.493 37.93 4.605 ;
      RECT 37.945 3.261 37.95 3.323 ;
      RECT 37.94 3.183 37.945 3.346 ;
      RECT 37.935 3.14 37.94 3.357 ;
      RECT 37.93 3.13 37.935 3.369 ;
      RECT 37.925 3.13 37.93 3.378 ;
      RECT 37.9 3.13 37.925 3.41 ;
      RECT 37.895 3.13 37.9 3.443 ;
      RECT 37.88 3.13 37.895 3.468 ;
      RECT 37.87 3.13 37.88 3.495 ;
      RECT 37.865 3.13 37.87 3.508 ;
      RECT 37.86 3.13 37.865 3.523 ;
      RECT 37.85 3.13 37.86 3.538 ;
      RECT 37.845 3.13 37.85 3.558 ;
      RECT 37.82 3.13 37.845 3.593 ;
      RECT 37.775 3.13 37.82 3.638 ;
      RECT 37.765 3.13 37.775 3.651 ;
      RECT 37.68 3.215 37.765 3.658 ;
      RECT 37.645 3.337 37.68 3.667 ;
      RECT 37.64 3.377 37.645 3.671 ;
      RECT 37.62 3.4 37.64 3.673 ;
      RECT 37.615 3.43 37.62 3.676 ;
      RECT 37.605 3.442 37.615 3.677 ;
      RECT 37.56 3.465 37.605 3.682 ;
      RECT 37.52 3.495 37.56 3.69 ;
      RECT 37.485 3.507 37.52 3.696 ;
      RECT 37.48 3.512 37.485 3.7 ;
      RECT 37.41 3.522 37.48 3.707 ;
      RECT 37.37 3.532 37.41 3.717 ;
      RECT 37.35 3.537 37.37 3.723 ;
      RECT 37.34 3.541 37.35 3.728 ;
      RECT 37.335 3.544 37.34 3.731 ;
      RECT 37.325 3.545 37.335 3.732 ;
      RECT 37.3 3.547 37.325 3.736 ;
      RECT 37.29 3.552 37.3 3.739 ;
      RECT 37.245 3.56 37.29 3.74 ;
      RECT 37.12 3.565 37.245 3.74 ;
      RECT 37.675 3.862 37.695 4.044 ;
      RECT 37.626 3.847 37.675 4.043 ;
      RECT 37.54 3.862 37.695 4.041 ;
      RECT 37.525 3.862 37.695 4.04 ;
      RECT 37.49 3.84 37.66 4.025 ;
      RECT 37.56 4.86 37.575 5.069 ;
      RECT 37.56 4.868 37.58 5.068 ;
      RECT 37.505 4.868 37.58 5.067 ;
      RECT 37.485 4.872 37.585 5.065 ;
      RECT 37.465 4.822 37.505 5.064 ;
      RECT 37.41 4.88 37.59 5.062 ;
      RECT 37.375 4.837 37.505 5.06 ;
      RECT 37.371 4.84 37.56 5.059 ;
      RECT 37.285 4.848 37.56 5.057 ;
      RECT 37.285 4.892 37.595 5.05 ;
      RECT 37.275 4.985 37.595 5.048 ;
      RECT 37.285 4.904 37.6 5.033 ;
      RECT 37.285 4.925 37.615 5.003 ;
      RECT 37.285 4.952 37.62 4.973 ;
      RECT 37.41 4.83 37.505 5.062 ;
      RECT 37.04 3.875 37.045 4.413 ;
      RECT 36.845 4.205 36.85 4.4 ;
      RECT 35.145 3.87 35.16 4.25 ;
      RECT 37.21 3.87 37.215 4.04 ;
      RECT 37.205 3.87 37.21 4.05 ;
      RECT 37.2 3.87 37.205 4.063 ;
      RECT 37.175 3.87 37.2 4.105 ;
      RECT 37.15 3.87 37.175 4.178 ;
      RECT 37.135 3.87 37.15 4.23 ;
      RECT 37.13 3.87 37.135 4.26 ;
      RECT 37.105 3.87 37.13 4.3 ;
      RECT 37.09 3.87 37.105 4.355 ;
      RECT 37.085 3.87 37.09 4.388 ;
      RECT 37.06 3.87 37.085 4.408 ;
      RECT 37.045 3.87 37.06 4.414 ;
      RECT 36.975 3.905 37.04 4.41 ;
      RECT 36.925 3.96 36.975 4.405 ;
      RECT 36.915 3.992 36.925 4.403 ;
      RECT 36.91 4.017 36.915 4.403 ;
      RECT 36.89 4.09 36.91 4.403 ;
      RECT 36.88 4.17 36.89 4.402 ;
      RECT 36.865 4.2 36.88 4.402 ;
      RECT 36.85 4.205 36.865 4.401 ;
      RECT 36.79 4.207 36.845 4.398 ;
      RECT 36.76 4.212 36.79 4.394 ;
      RECT 36.758 4.215 36.76 4.393 ;
      RECT 36.672 4.217 36.758 4.39 ;
      RECT 36.586 4.223 36.672 4.384 ;
      RECT 36.5 4.228 36.586 4.378 ;
      RECT 36.427 4.233 36.5 4.379 ;
      RECT 36.341 4.239 36.427 4.387 ;
      RECT 36.255 4.245 36.341 4.396 ;
      RECT 36.235 4.249 36.255 4.401 ;
      RECT 36.188 4.251 36.235 4.404 ;
      RECT 36.102 4.256 36.188 4.41 ;
      RECT 36.016 4.261 36.102 4.419 ;
      RECT 35.93 4.267 36.016 4.427 ;
      RECT 35.845 4.265 35.93 4.436 ;
      RECT 35.841 4.26 35.845 4.44 ;
      RECT 35.755 4.255 35.841 4.432 ;
      RECT 35.691 4.246 35.755 4.42 ;
      RECT 35.605 4.237 35.691 4.407 ;
      RECT 35.581 4.23 35.605 4.398 ;
      RECT 35.495 4.224 35.581 4.385 ;
      RECT 35.455 4.217 35.495 4.371 ;
      RECT 35.45 4.207 35.455 4.367 ;
      RECT 35.44 4.195 35.45 4.366 ;
      RECT 35.42 4.165 35.44 4.363 ;
      RECT 35.365 4.085 35.42 4.357 ;
      RECT 35.345 4.004 35.365 4.352 ;
      RECT 35.325 3.962 35.345 4.348 ;
      RECT 35.3 3.915 35.325 4.342 ;
      RECT 35.295 3.89 35.3 4.339 ;
      RECT 35.26 3.87 35.295 4.334 ;
      RECT 35.251 3.87 35.26 4.327 ;
      RECT 35.165 3.87 35.251 4.297 ;
      RECT 35.16 3.87 35.165 4.26 ;
      RECT 35.125 3.87 35.145 4.182 ;
      RECT 35.12 3.912 35.125 4.147 ;
      RECT 35.115 3.987 35.12 4.103 ;
      RECT 36.565 3.792 36.74 4.04 ;
      RECT 36.565 3.792 36.745 4.038 ;
      RECT 36.56 3.824 36.745 3.998 ;
      RECT 36.59 3.765 36.76 3.985 ;
      RECT 36.555 3.842 36.76 3.918 ;
      RECT 35.865 3.305 36.035 3.48 ;
      RECT 35.865 3.305 36.207 3.472 ;
      RECT 35.865 3.305 36.29 3.466 ;
      RECT 35.865 3.305 36.325 3.462 ;
      RECT 35.865 3.305 36.345 3.461 ;
      RECT 35.865 3.305 36.431 3.457 ;
      RECT 36.325 3.13 36.495 3.452 ;
      RECT 35.9 3.237 36.525 3.45 ;
      RECT 35.89 3.292 36.53 3.448 ;
      RECT 35.865 3.328 36.54 3.443 ;
      RECT 35.865 3.355 36.545 3.373 ;
      RECT 35.93 3.18 36.505 3.45 ;
      RECT 36.121 3.165 36.505 3.45 ;
      RECT 35.955 3.168 36.505 3.45 ;
      RECT 36.035 3.166 36.121 3.477 ;
      RECT 36.121 3.163 36.5 3.45 ;
      RECT 36.305 3.14 36.5 3.45 ;
      RECT 36.207 3.161 36.5 3.45 ;
      RECT 36.29 3.155 36.305 3.463 ;
      RECT 36.44 4.52 36.445 4.72 ;
      RECT 35.905 4.585 35.95 4.72 ;
      RECT 36.475 4.52 36.495 4.693 ;
      RECT 36.445 4.52 36.475 4.708 ;
      RECT 36.38 4.52 36.44 4.745 ;
      RECT 36.365 4.52 36.38 4.775 ;
      RECT 36.35 4.52 36.365 4.788 ;
      RECT 36.33 4.52 36.35 4.803 ;
      RECT 36.325 4.52 36.33 4.812 ;
      RECT 36.315 4.524 36.325 4.817 ;
      RECT 36.3 4.534 36.315 4.828 ;
      RECT 36.275 4.55 36.3 4.838 ;
      RECT 36.265 4.564 36.275 4.84 ;
      RECT 36.245 4.576 36.265 4.837 ;
      RECT 36.215 4.597 36.245 4.831 ;
      RECT 36.205 4.609 36.215 4.826 ;
      RECT 36.195 4.607 36.205 4.823 ;
      RECT 36.18 4.606 36.195 4.818 ;
      RECT 36.175 4.605 36.18 4.813 ;
      RECT 36.14 4.603 36.175 4.803 ;
      RECT 36.12 4.6 36.14 4.785 ;
      RECT 36.11 4.598 36.12 4.78 ;
      RECT 36.1 4.597 36.11 4.775 ;
      RECT 36.065 4.595 36.1 4.763 ;
      RECT 36.01 4.591 36.065 4.743 ;
      RECT 36 4.589 36.01 4.728 ;
      RECT 35.995 4.589 36 4.723 ;
      RECT 35.95 4.587 35.995 4.72 ;
      RECT 35.855 4.585 35.905 4.724 ;
      RECT 35.845 4.586 35.855 4.729 ;
      RECT 35.785 4.593 35.845 4.743 ;
      RECT 35.76 4.601 35.785 4.763 ;
      RECT 35.75 4.605 35.76 4.775 ;
      RECT 35.745 4.606 35.75 4.78 ;
      RECT 35.73 4.608 35.745 4.783 ;
      RECT 35.715 4.61 35.73 4.788 ;
      RECT 35.71 4.61 35.715 4.791 ;
      RECT 35.665 4.615 35.71 4.802 ;
      RECT 35.66 4.619 35.665 4.814 ;
      RECT 35.635 4.615 35.66 4.818 ;
      RECT 35.625 4.611 35.635 4.822 ;
      RECT 35.615 4.61 35.625 4.826 ;
      RECT 35.6 4.6 35.615 4.832 ;
      RECT 35.595 4.588 35.6 4.836 ;
      RECT 35.59 4.585 35.595 4.837 ;
      RECT 35.585 4.582 35.59 4.839 ;
      RECT 35.57 4.57 35.585 4.838 ;
      RECT 35.555 4.552 35.57 4.835 ;
      RECT 35.535 4.531 35.555 4.828 ;
      RECT 35.47 4.52 35.535 4.8 ;
      RECT 35.466 4.52 35.47 4.779 ;
      RECT 35.38 4.52 35.466 4.749 ;
      RECT 35.365 4.52 35.38 4.705 ;
      RECT 35.94 3.62 35.945 3.855 ;
      RECT 35.07 3.536 35.075 3.74 ;
      RECT 35.65 3.565 35.655 3.72 ;
      RECT 35.57 3.545 35.575 3.72 ;
      RECT 36.24 3.687 36.255 4.04 ;
      RECT 36.166 3.672 36.24 4.04 ;
      RECT 36.08 3.655 36.166 4.04 ;
      RECT 36.07 3.645 36.08 4.038 ;
      RECT 36.065 3.643 36.07 4.033 ;
      RECT 36.05 3.641 36.065 4.019 ;
      RECT 35.98 3.633 36.05 3.959 ;
      RECT 35.96 3.624 35.98 3.893 ;
      RECT 35.955 3.621 35.96 3.873 ;
      RECT 35.945 3.62 35.955 3.863 ;
      RECT 35.935 3.62 35.94 3.847 ;
      RECT 35.925 3.619 35.935 3.837 ;
      RECT 35.915 3.617 35.925 3.825 ;
      RECT 35.9 3.614 35.915 3.805 ;
      RECT 35.89 3.612 35.9 3.79 ;
      RECT 35.87 3.609 35.89 3.778 ;
      RECT 35.865 3.607 35.87 3.768 ;
      RECT 35.84 3.605 35.865 3.755 ;
      RECT 35.81 3.6 35.84 3.74 ;
      RECT 35.73 3.591 35.81 3.731 ;
      RECT 35.685 3.58 35.73 3.724 ;
      RECT 35.665 3.571 35.685 3.721 ;
      RECT 35.655 3.566 35.665 3.72 ;
      RECT 35.61 3.56 35.65 3.72 ;
      RECT 35.595 3.552 35.61 3.72 ;
      RECT 35.575 3.547 35.595 3.72 ;
      RECT 35.555 3.544 35.57 3.72 ;
      RECT 35.472 3.543 35.555 3.719 ;
      RECT 35.386 3.542 35.472 3.715 ;
      RECT 35.3 3.54 35.386 3.712 ;
      RECT 35.247 3.539 35.3 3.714 ;
      RECT 35.161 3.538 35.247 3.723 ;
      RECT 35.075 3.537 35.161 3.735 ;
      RECT 35.055 3.536 35.07 3.743 ;
      RECT 34.975 3.535 35.055 3.755 ;
      RECT 34.95 3.535 34.975 3.768 ;
      RECT 34.925 3.535 34.95 3.783 ;
      RECT 34.92 3.535 34.925 3.805 ;
      RECT 34.915 3.535 34.92 3.823 ;
      RECT 34.91 3.535 34.915 3.84 ;
      RECT 34.905 3.535 34.91 3.853 ;
      RECT 34.9 3.535 34.905 3.863 ;
      RECT 34.86 3.535 34.9 3.948 ;
      RECT 34.845 3.535 34.86 4.033 ;
      RECT 34.835 3.536 34.845 4.045 ;
      RECT 34.8 3.541 34.835 4.05 ;
      RECT 34.76 3.55 34.8 4.05 ;
      RECT 34.745 3.56 34.76 4.05 ;
      RECT 34.74 3.57 34.745 4.05 ;
      RECT 34.72 3.597 34.74 4.05 ;
      RECT 34.67 3.68 34.72 4.05 ;
      RECT 34.665 3.742 34.67 4.05 ;
      RECT 34.655 3.755 34.665 4.05 ;
      RECT 34.645 3.777 34.655 4.05 ;
      RECT 34.635 3.802 34.645 4.045 ;
      RECT 34.63 3.84 34.635 4.038 ;
      RECT 34.62 3.95 34.63 4.033 ;
      RECT 36.015 4.871 36.03 5.13 ;
      RECT 36.015 4.886 36.035 5.129 ;
      RECT 35.931 4.886 36.035 5.127 ;
      RECT 35.931 4.9 36.04 5.126 ;
      RECT 35.845 4.942 36.045 5.123 ;
      RECT 35.84 4.885 36.03 5.118 ;
      RECT 35.84 4.956 36.05 5.115 ;
      RECT 35.835 4.987 36.05 5.113 ;
      RECT 35.84 4.984 36.065 5.103 ;
      RECT 35.835 5.03 36.08 5.088 ;
      RECT 35.835 5.058 36.085 5.073 ;
      RECT 35.845 4.86 36.015 5.123 ;
      RECT 35.605 3.87 35.775 4.04 ;
      RECT 35.57 3.87 35.775 4.035 ;
      RECT 35.56 3.87 35.775 4.028 ;
      RECT 35.555 3.855 35.725 4.025 ;
      RECT 34.385 4.392 34.65 4.835 ;
      RECT 34.38 4.363 34.595 4.833 ;
      RECT 34.375 4.517 34.655 4.828 ;
      RECT 34.38 4.412 34.655 4.828 ;
      RECT 34.38 4.423 34.665 4.815 ;
      RECT 34.38 4.37 34.625 4.833 ;
      RECT 34.385 4.357 34.595 4.835 ;
      RECT 34.385 4.355 34.545 4.835 ;
      RECT 34.486 4.347 34.545 4.835 ;
      RECT 34.4 4.348 34.545 4.835 ;
      RECT 34.486 4.346 34.535 4.835 ;
      RECT 34.29 3.161 34.465 3.46 ;
      RECT 34.34 3.123 34.465 3.46 ;
      RECT 34.325 3.125 34.551 3.452 ;
      RECT 34.325 3.128 34.59 3.439 ;
      RECT 34.325 3.129 34.6 3.425 ;
      RECT 34.28 3.18 34.6 3.415 ;
      RECT 34.325 3.13 34.605 3.41 ;
      RECT 34.28 3.34 34.61 3.4 ;
      RECT 34.265 3.2 34.605 3.34 ;
      RECT 34.26 3.216 34.605 3.28 ;
      RECT 34.305 3.14 34.605 3.41 ;
      RECT 34.34 3.121 34.426 3.46 ;
      RECT 32.43 3.035 32.6 4.225 ;
      RECT 32.43 3.035 32.9 3.205 ;
      RECT 32.43 9.26 32.9 9.43 ;
      RECT 32.43 8.24 32.6 9.43 ;
      RECT 31.44 3.035 31.61 4.225 ;
      RECT 31.44 3.035 31.91 3.205 ;
      RECT 31.44 9.26 31.91 9.43 ;
      RECT 31.44 8.24 31.61 9.43 ;
      RECT 29.59 3.93 29.76 5.16 ;
      RECT 29.645 2.15 29.815 4.1 ;
      RECT 29.59 1.87 29.76 2.32 ;
      RECT 29.59 10.145 29.76 10.595 ;
      RECT 29.645 8.365 29.815 10.315 ;
      RECT 29.59 7.305 29.76 8.535 ;
      RECT 29.07 1.87 29.24 5.16 ;
      RECT 29.07 3.37 29.475 3.7 ;
      RECT 29.07 2.53 29.475 2.86 ;
      RECT 29.07 7.305 29.24 10.595 ;
      RECT 29.07 9.605 29.475 9.935 ;
      RECT 29.07 8.765 29.475 9.095 ;
      RECT 26.995 4.421 27 4.593 ;
      RECT 26.99 4.414 26.995 4.683 ;
      RECT 26.985 4.408 26.99 4.702 ;
      RECT 26.965 4.402 26.985 4.712 ;
      RECT 26.95 4.397 26.965 4.72 ;
      RECT 26.913 4.391 26.95 4.718 ;
      RECT 26.827 4.377 26.913 4.714 ;
      RECT 26.741 4.359 26.827 4.709 ;
      RECT 26.655 4.34 26.741 4.703 ;
      RECT 26.625 4.328 26.655 4.699 ;
      RECT 26.605 4.322 26.625 4.698 ;
      RECT 26.54 4.32 26.605 4.696 ;
      RECT 26.525 4.32 26.54 4.688 ;
      RECT 26.51 4.32 26.525 4.675 ;
      RECT 26.505 4.32 26.51 4.665 ;
      RECT 26.49 4.32 26.505 4.643 ;
      RECT 26.475 4.32 26.49 4.61 ;
      RECT 26.47 4.32 26.475 4.588 ;
      RECT 26.46 4.32 26.47 4.57 ;
      RECT 26.445 4.32 26.46 4.548 ;
      RECT 26.425 4.32 26.445 4.51 ;
      RECT 26.775 3.605 26.81 4.044 ;
      RECT 26.775 3.605 26.815 4.043 ;
      RECT 26.72 3.665 26.815 4.042 ;
      RECT 26.585 3.837 26.815 4.041 ;
      RECT 26.695 3.715 26.815 4.041 ;
      RECT 26.585 3.837 26.84 4.031 ;
      RECT 26.64 3.782 26.92 3.948 ;
      RECT 26.815 3.576 26.82 4.039 ;
      RECT 26.67 3.752 26.96 3.825 ;
      RECT 26.685 3.735 26.815 4.041 ;
      RECT 26.82 3.575 26.99 3.763 ;
      RECT 26.81 3.578 26.99 3.763 ;
      RECT 26.315 3.455 26.485 3.765 ;
      RECT 26.315 3.455 26.49 3.738 ;
      RECT 26.315 3.455 26.495 3.715 ;
      RECT 26.315 3.455 26.505 3.665 ;
      RECT 26.31 3.56 26.505 3.635 ;
      RECT 26.345 3.13 26.515 3.608 ;
      RECT 26.345 3.13 26.53 3.529 ;
      RECT 26.335 3.34 26.53 3.529 ;
      RECT 26.345 3.14 26.54 3.444 ;
      RECT 26.275 3.882 26.28 4.085 ;
      RECT 26.265 3.87 26.275 4.195 ;
      RECT 26.24 3.87 26.265 4.235 ;
      RECT 26.16 3.87 26.24 4.32 ;
      RECT 26.15 3.87 26.16 4.39 ;
      RECT 26.125 3.87 26.15 4.413 ;
      RECT 26.105 3.87 26.125 4.448 ;
      RECT 26.06 3.88 26.105 4.491 ;
      RECT 26.05 3.892 26.06 4.528 ;
      RECT 26.03 3.906 26.05 4.548 ;
      RECT 26.02 3.924 26.03 4.564 ;
      RECT 26.005 3.95 26.02 4.574 ;
      RECT 25.99 3.991 26.005 4.588 ;
      RECT 25.98 4.026 25.99 4.598 ;
      RECT 25.975 4.042 25.98 4.603 ;
      RECT 25.965 4.057 25.975 4.608 ;
      RECT 25.945 4.1 25.965 4.618 ;
      RECT 25.925 4.137 25.945 4.631 ;
      RECT 25.89 4.16 25.925 4.649 ;
      RECT 25.88 4.174 25.89 4.665 ;
      RECT 25.86 4.184 25.88 4.675 ;
      RECT 25.855 4.193 25.86 4.683 ;
      RECT 25.845 4.2 25.855 4.69 ;
      RECT 25.835 4.207 25.845 4.698 ;
      RECT 25.82 4.217 25.835 4.706 ;
      RECT 25.81 4.231 25.82 4.716 ;
      RECT 25.8 4.243 25.81 4.728 ;
      RECT 25.785 4.265 25.8 4.741 ;
      RECT 25.775 4.287 25.785 4.752 ;
      RECT 25.765 4.307 25.775 4.761 ;
      RECT 25.76 4.322 25.765 4.768 ;
      RECT 25.73 4.355 25.76 4.782 ;
      RECT 25.72 4.39 25.73 4.797 ;
      RECT 25.715 4.397 25.72 4.803 ;
      RECT 25.695 4.412 25.715 4.81 ;
      RECT 25.69 4.427 25.695 4.818 ;
      RECT 25.685 4.436 25.69 4.823 ;
      RECT 25.67 4.442 25.685 4.83 ;
      RECT 25.665 4.448 25.67 4.838 ;
      RECT 25.66 4.452 25.665 4.845 ;
      RECT 25.655 4.456 25.66 4.855 ;
      RECT 25.645 4.461 25.655 4.865 ;
      RECT 25.625 4.472 25.645 4.893 ;
      RECT 25.61 4.484 25.625 4.92 ;
      RECT 25.59 4.497 25.61 4.945 ;
      RECT 25.57 4.512 25.59 4.969 ;
      RECT 25.555 4.527 25.57 4.984 ;
      RECT 25.55 4.538 25.555 4.993 ;
      RECT 25.485 4.583 25.55 5.003 ;
      RECT 25.45 4.642 25.485 5.016 ;
      RECT 25.445 4.665 25.45 5.022 ;
      RECT 25.44 4.672 25.445 5.024 ;
      RECT 25.425 4.682 25.44 5.027 ;
      RECT 25.395 4.707 25.425 5.031 ;
      RECT 25.39 4.725 25.395 5.035 ;
      RECT 25.385 4.732 25.39 5.036 ;
      RECT 25.365 4.74 25.385 5.04 ;
      RECT 25.355 4.747 25.365 5.044 ;
      RECT 25.311 4.758 25.355 5.051 ;
      RECT 25.225 4.786 25.311 5.067 ;
      RECT 25.165 4.81 25.225 5.085 ;
      RECT 25.12 4.82 25.165 5.099 ;
      RECT 25.061 4.828 25.12 5.113 ;
      RECT 24.975 4.835 25.061 5.132 ;
      RECT 24.95 4.84 24.975 5.147 ;
      RECT 24.87 4.843 24.95 5.15 ;
      RECT 24.79 4.847 24.87 5.137 ;
      RECT 24.781 4.85 24.79 5.122 ;
      RECT 24.695 4.85 24.781 5.107 ;
      RECT 24.635 4.852 24.695 5.084 ;
      RECT 24.631 4.855 24.635 5.074 ;
      RECT 24.545 4.855 24.631 5.059 ;
      RECT 24.47 4.855 24.545 5.035 ;
      RECT 25.785 3.864 25.795 4.04 ;
      RECT 25.74 3.831 25.785 4.04 ;
      RECT 25.695 3.782 25.74 4.04 ;
      RECT 25.665 3.752 25.695 4.041 ;
      RECT 25.66 3.735 25.665 4.042 ;
      RECT 25.635 3.715 25.66 4.043 ;
      RECT 25.62 3.69 25.635 4.044 ;
      RECT 25.615 3.677 25.62 4.045 ;
      RECT 25.61 3.671 25.615 4.043 ;
      RECT 25.605 3.663 25.61 4.037 ;
      RECT 25.58 3.655 25.605 4.017 ;
      RECT 25.56 3.644 25.58 3.988 ;
      RECT 25.53 3.629 25.56 3.959 ;
      RECT 25.51 3.615 25.53 3.931 ;
      RECT 25.5 3.609 25.51 3.91 ;
      RECT 25.495 3.606 25.5 3.893 ;
      RECT 25.49 3.603 25.495 3.878 ;
      RECT 25.475 3.598 25.49 3.843 ;
      RECT 25.47 3.594 25.475 3.81 ;
      RECT 25.45 3.589 25.47 3.786 ;
      RECT 25.42 3.581 25.45 3.751 ;
      RECT 25.405 3.575 25.42 3.728 ;
      RECT 25.365 3.568 25.405 3.713 ;
      RECT 25.34 3.56 25.365 3.693 ;
      RECT 25.32 3.555 25.34 3.683 ;
      RECT 25.285 3.549 25.32 3.678 ;
      RECT 25.24 3.54 25.285 3.677 ;
      RECT 25.21 3.536 25.24 3.679 ;
      RECT 25.125 3.544 25.21 3.683 ;
      RECT 25.055 3.555 25.125 3.705 ;
      RECT 25.042 3.561 25.055 3.728 ;
      RECT 24.956 3.568 25.042 3.75 ;
      RECT 24.87 3.58 24.956 3.787 ;
      RECT 24.87 3.957 24.88 4.195 ;
      RECT 24.865 3.586 24.87 3.81 ;
      RECT 24.86 3.842 24.87 4.195 ;
      RECT 24.86 3.587 24.865 3.815 ;
      RECT 24.855 3.588 24.86 4.195 ;
      RECT 24.831 3.59 24.855 4.196 ;
      RECT 24.745 3.598 24.831 4.198 ;
      RECT 24.725 3.612 24.745 4.201 ;
      RECT 24.72 3.64 24.725 4.202 ;
      RECT 24.715 3.652 24.72 4.203 ;
      RECT 24.71 3.667 24.715 4.204 ;
      RECT 24.7 3.697 24.71 4.205 ;
      RECT 24.695 3.735 24.7 4.203 ;
      RECT 24.69 3.755 24.695 4.198 ;
      RECT 24.675 3.79 24.69 4.183 ;
      RECT 24.665 3.842 24.675 4.163 ;
      RECT 24.66 3.872 24.665 4.151 ;
      RECT 24.645 3.885 24.66 4.134 ;
      RECT 24.62 3.889 24.645 4.101 ;
      RECT 24.605 3.887 24.62 4.078 ;
      RECT 24.59 3.886 24.605 4.075 ;
      RECT 24.53 3.884 24.59 4.073 ;
      RECT 24.52 3.882 24.53 4.068 ;
      RECT 24.48 3.881 24.52 4.065 ;
      RECT 24.41 3.878 24.48 4.063 ;
      RECT 24.355 3.876 24.41 4.058 ;
      RECT 24.285 3.87 24.355 4.053 ;
      RECT 24.276 3.87 24.285 4.05 ;
      RECT 24.19 3.87 24.276 4.045 ;
      RECT 24.185 3.87 24.19 4.04 ;
      RECT 25.49 3.105 25.665 3.455 ;
      RECT 25.49 3.12 25.675 3.453 ;
      RECT 25.465 3.07 25.61 3.45 ;
      RECT 25.445 3.071 25.61 3.443 ;
      RECT 25.435 3.072 25.62 3.438 ;
      RECT 25.405 3.073 25.62 3.425 ;
      RECT 25.355 3.074 25.62 3.401 ;
      RECT 25.35 3.076 25.62 3.386 ;
      RECT 25.35 3.142 25.68 3.38 ;
      RECT 25.33 3.083 25.635 3.36 ;
      RECT 25.32 3.092 25.645 3.215 ;
      RECT 25.33 3.087 25.645 3.36 ;
      RECT 25.35 3.077 25.635 3.386 ;
      RECT 24.935 4.402 25.105 4.69 ;
      RECT 24.93 4.42 25.115 4.685 ;
      RECT 24.895 4.428 25.18 4.605 ;
      RECT 24.895 4.428 25.266 4.595 ;
      RECT 24.895 4.428 25.32 4.541 ;
      RECT 25.18 4.325 25.35 4.509 ;
      RECT 24.895 4.48 25.355 4.497 ;
      RECT 24.88 4.45 25.35 4.493 ;
      RECT 25.14 4.332 25.18 4.644 ;
      RECT 25.02 4.369 25.35 4.509 ;
      RECT 25.115 4.344 25.14 4.67 ;
      RECT 25.105 4.351 25.35 4.509 ;
      RECT 25.236 3.815 25.305 4.074 ;
      RECT 25.236 3.87 25.31 4.073 ;
      RECT 25.15 3.87 25.31 4.072 ;
      RECT 25.145 3.87 25.315 4.065 ;
      RECT 25.135 3.815 25.305 4.06 ;
      RECT 24.515 3.114 24.69 3.415 ;
      RECT 24.5 3.102 24.515 3.4 ;
      RECT 24.47 3.101 24.5 3.353 ;
      RECT 24.47 3.119 24.695 3.348 ;
      RECT 24.455 3.103 24.515 3.313 ;
      RECT 24.45 3.125 24.705 3.213 ;
      RECT 24.45 3.108 24.601 3.213 ;
      RECT 24.45 3.11 24.605 3.213 ;
      RECT 24.455 3.106 24.601 3.313 ;
      RECT 24.56 4.342 24.565 4.69 ;
      RECT 24.55 4.332 24.56 4.696 ;
      RECT 24.515 4.322 24.55 4.698 ;
      RECT 24.477 4.317 24.515 4.702 ;
      RECT 24.391 4.31 24.477 4.709 ;
      RECT 24.305 4.3 24.391 4.719 ;
      RECT 24.26 4.295 24.305 4.727 ;
      RECT 24.256 4.295 24.26 4.731 ;
      RECT 24.17 4.295 24.256 4.738 ;
      RECT 24.155 4.295 24.17 4.738 ;
      RECT 24.145 4.293 24.155 4.71 ;
      RECT 24.135 4.289 24.145 4.653 ;
      RECT 24.115 4.283 24.135 4.585 ;
      RECT 24.11 4.279 24.115 4.533 ;
      RECT 24.1 4.278 24.11 4.5 ;
      RECT 24.05 4.276 24.1 4.485 ;
      RECT 24.025 4.274 24.05 4.48 ;
      RECT 23.982 4.272 24.025 4.476 ;
      RECT 23.896 4.268 23.982 4.464 ;
      RECT 23.81 4.263 23.896 4.448 ;
      RECT 23.78 4.26 23.81 4.435 ;
      RECT 23.755 4.259 23.78 4.423 ;
      RECT 23.75 4.259 23.755 4.413 ;
      RECT 23.71 4.258 23.75 4.405 ;
      RECT 23.695 4.257 23.71 4.398 ;
      RECT 23.645 4.256 23.695 4.39 ;
      RECT 23.643 4.255 23.645 4.385 ;
      RECT 23.557 4.253 23.643 4.385 ;
      RECT 23.471 4.248 23.557 4.385 ;
      RECT 23.385 4.244 23.471 4.385 ;
      RECT 23.336 4.24 23.385 4.383 ;
      RECT 23.25 4.237 23.336 4.378 ;
      RECT 23.227 4.234 23.25 4.374 ;
      RECT 23.141 4.231 23.227 4.369 ;
      RECT 23.055 4.227 23.141 4.36 ;
      RECT 23.03 4.22 23.055 4.355 ;
      RECT 22.97 4.185 23.03 4.352 ;
      RECT 22.95 4.11 22.97 4.349 ;
      RECT 22.945 4.052 22.95 4.348 ;
      RECT 22.92 3.992 22.945 4.347 ;
      RECT 22.845 3.87 22.92 4.343 ;
      RECT 22.835 3.87 22.845 4.335 ;
      RECT 22.82 3.87 22.835 4.325 ;
      RECT 22.805 3.87 22.82 4.295 ;
      RECT 22.79 3.87 22.805 4.24 ;
      RECT 22.775 3.87 22.79 4.178 ;
      RECT 22.75 3.87 22.775 4.103 ;
      RECT 22.745 3.87 22.75 4.053 ;
      RECT 24.09 3.415 24.11 3.724 ;
      RECT 24.076 3.417 24.125 3.721 ;
      RECT 24.076 3.422 24.145 3.712 ;
      RECT 23.99 3.42 24.125 3.706 ;
      RECT 23.99 3.428 24.18 3.689 ;
      RECT 23.955 3.43 24.18 3.688 ;
      RECT 23.925 3.438 24.18 3.679 ;
      RECT 23.915 3.443 24.2 3.665 ;
      RECT 23.955 3.433 24.2 3.665 ;
      RECT 23.955 3.436 24.21 3.653 ;
      RECT 23.925 3.438 24.22 3.64 ;
      RECT 23.925 3.442 24.23 3.583 ;
      RECT 23.915 3.447 24.235 3.498 ;
      RECT 24.076 3.415 24.11 3.721 ;
      RECT 23.515 3.518 23.52 3.73 ;
      RECT 23.39 3.515 23.405 3.73 ;
      RECT 22.855 3.545 22.925 3.73 ;
      RECT 22.74 3.545 22.775 3.725 ;
      RECT 23.861 3.847 23.88 4.041 ;
      RECT 23.775 3.802 23.861 4.042 ;
      RECT 23.765 3.755 23.775 4.044 ;
      RECT 23.76 3.735 23.765 4.045 ;
      RECT 23.74 3.7 23.76 4.046 ;
      RECT 23.725 3.65 23.74 4.047 ;
      RECT 23.705 3.587 23.725 4.048 ;
      RECT 23.695 3.55 23.705 4.049 ;
      RECT 23.68 3.539 23.695 4.05 ;
      RECT 23.675 3.531 23.68 4.048 ;
      RECT 23.665 3.53 23.675 4.04 ;
      RECT 23.635 3.527 23.665 4.019 ;
      RECT 23.56 3.522 23.635 3.964 ;
      RECT 23.545 3.518 23.56 3.91 ;
      RECT 23.535 3.518 23.545 3.805 ;
      RECT 23.52 3.518 23.535 3.738 ;
      RECT 23.505 3.518 23.515 3.728 ;
      RECT 23.45 3.517 23.505 3.725 ;
      RECT 23.405 3.515 23.45 3.728 ;
      RECT 23.377 3.515 23.39 3.731 ;
      RECT 23.291 3.519 23.377 3.733 ;
      RECT 23.205 3.525 23.291 3.738 ;
      RECT 23.185 3.529 23.205 3.74 ;
      RECT 23.183 3.53 23.185 3.739 ;
      RECT 23.097 3.532 23.183 3.738 ;
      RECT 23.011 3.537 23.097 3.735 ;
      RECT 22.925 3.542 23.011 3.732 ;
      RECT 22.775 3.545 22.855 3.728 ;
      RECT 23.435 7.305 23.605 10.595 ;
      RECT 23.435 9.605 23.84 9.935 ;
      RECT 23.435 8.765 23.84 9.095 ;
      RECT 23.551 4.52 23.6 4.854 ;
      RECT 23.551 4.52 23.605 4.853 ;
      RECT 23.465 4.52 23.605 4.852 ;
      RECT 23.24 4.628 23.61 4.85 ;
      RECT 23.465 4.52 23.635 4.843 ;
      RECT 23.435 4.532 23.64 4.834 ;
      RECT 23.42 4.55 23.645 4.831 ;
      RECT 23.235 4.634 23.645 4.758 ;
      RECT 23.23 4.641 23.645 4.718 ;
      RECT 23.245 4.607 23.645 4.831 ;
      RECT 23.406 4.553 23.61 4.85 ;
      RECT 23.32 4.573 23.645 4.831 ;
      RECT 23.42 4.547 23.64 4.834 ;
      RECT 23.19 3.871 23.38 4.065 ;
      RECT 23.185 3.873 23.38 4.064 ;
      RECT 23.18 3.877 23.395 4.061 ;
      RECT 23.195 3.87 23.395 4.061 ;
      RECT 23.18 3.98 23.4 4.056 ;
      RECT 22.475 4.48 22.566 4.778 ;
      RECT 22.47 4.482 22.645 4.773 ;
      RECT 22.475 4.48 22.645 4.773 ;
      RECT 22.47 4.486 22.665 4.771 ;
      RECT 22.47 4.541 22.705 4.77 ;
      RECT 22.47 4.576 22.72 4.764 ;
      RECT 22.47 4.61 22.73 4.754 ;
      RECT 22.46 4.49 22.665 4.605 ;
      RECT 22.46 4.51 22.68 4.605 ;
      RECT 22.46 4.493 22.67 4.605 ;
      RECT 22.685 3.261 22.69 3.323 ;
      RECT 22.68 3.183 22.685 3.346 ;
      RECT 22.675 3.14 22.68 3.357 ;
      RECT 22.67 3.13 22.675 3.369 ;
      RECT 22.665 3.13 22.67 3.378 ;
      RECT 22.64 3.13 22.665 3.41 ;
      RECT 22.635 3.13 22.64 3.443 ;
      RECT 22.62 3.13 22.635 3.468 ;
      RECT 22.61 3.13 22.62 3.495 ;
      RECT 22.605 3.13 22.61 3.508 ;
      RECT 22.6 3.13 22.605 3.523 ;
      RECT 22.59 3.13 22.6 3.538 ;
      RECT 22.585 3.13 22.59 3.558 ;
      RECT 22.56 3.13 22.585 3.593 ;
      RECT 22.515 3.13 22.56 3.638 ;
      RECT 22.505 3.13 22.515 3.651 ;
      RECT 22.42 3.215 22.505 3.658 ;
      RECT 22.385 3.337 22.42 3.667 ;
      RECT 22.38 3.377 22.385 3.671 ;
      RECT 22.36 3.4 22.38 3.673 ;
      RECT 22.355 3.43 22.36 3.676 ;
      RECT 22.345 3.442 22.355 3.677 ;
      RECT 22.3 3.465 22.345 3.682 ;
      RECT 22.26 3.495 22.3 3.69 ;
      RECT 22.225 3.507 22.26 3.696 ;
      RECT 22.22 3.512 22.225 3.7 ;
      RECT 22.15 3.522 22.22 3.707 ;
      RECT 22.11 3.532 22.15 3.717 ;
      RECT 22.09 3.537 22.11 3.723 ;
      RECT 22.08 3.541 22.09 3.728 ;
      RECT 22.075 3.544 22.08 3.731 ;
      RECT 22.065 3.545 22.075 3.732 ;
      RECT 22.04 3.547 22.065 3.736 ;
      RECT 22.03 3.552 22.04 3.739 ;
      RECT 21.985 3.56 22.03 3.74 ;
      RECT 21.86 3.565 21.985 3.74 ;
      RECT 22.415 3.862 22.435 4.044 ;
      RECT 22.366 3.847 22.415 4.043 ;
      RECT 22.28 3.862 22.435 4.041 ;
      RECT 22.265 3.862 22.435 4.04 ;
      RECT 22.23 3.84 22.4 4.025 ;
      RECT 22.3 4.86 22.315 5.069 ;
      RECT 22.3 4.868 22.32 5.068 ;
      RECT 22.245 4.868 22.32 5.067 ;
      RECT 22.225 4.872 22.325 5.065 ;
      RECT 22.205 4.822 22.245 5.064 ;
      RECT 22.15 4.88 22.33 5.062 ;
      RECT 22.115 4.837 22.245 5.06 ;
      RECT 22.111 4.84 22.3 5.059 ;
      RECT 22.025 4.848 22.3 5.057 ;
      RECT 22.025 4.892 22.335 5.05 ;
      RECT 22.015 4.985 22.335 5.048 ;
      RECT 22.025 4.904 22.34 5.033 ;
      RECT 22.025 4.925 22.355 5.003 ;
      RECT 22.025 4.952 22.36 4.973 ;
      RECT 22.15 4.83 22.245 5.062 ;
      RECT 21.78 3.875 21.785 4.413 ;
      RECT 21.585 4.205 21.59 4.4 ;
      RECT 19.885 3.87 19.9 4.25 ;
      RECT 21.95 3.87 21.955 4.04 ;
      RECT 21.945 3.87 21.95 4.05 ;
      RECT 21.94 3.87 21.945 4.063 ;
      RECT 21.915 3.87 21.94 4.105 ;
      RECT 21.89 3.87 21.915 4.178 ;
      RECT 21.875 3.87 21.89 4.23 ;
      RECT 21.87 3.87 21.875 4.26 ;
      RECT 21.845 3.87 21.87 4.3 ;
      RECT 21.83 3.87 21.845 4.355 ;
      RECT 21.825 3.87 21.83 4.388 ;
      RECT 21.8 3.87 21.825 4.408 ;
      RECT 21.785 3.87 21.8 4.414 ;
      RECT 21.715 3.905 21.78 4.41 ;
      RECT 21.665 3.96 21.715 4.405 ;
      RECT 21.655 3.992 21.665 4.403 ;
      RECT 21.65 4.017 21.655 4.403 ;
      RECT 21.63 4.09 21.65 4.403 ;
      RECT 21.62 4.17 21.63 4.402 ;
      RECT 21.605 4.2 21.62 4.402 ;
      RECT 21.59 4.205 21.605 4.401 ;
      RECT 21.53 4.207 21.585 4.398 ;
      RECT 21.5 4.212 21.53 4.394 ;
      RECT 21.498 4.215 21.5 4.393 ;
      RECT 21.412 4.217 21.498 4.39 ;
      RECT 21.326 4.223 21.412 4.384 ;
      RECT 21.24 4.228 21.326 4.378 ;
      RECT 21.167 4.233 21.24 4.379 ;
      RECT 21.081 4.239 21.167 4.387 ;
      RECT 20.995 4.245 21.081 4.396 ;
      RECT 20.975 4.249 20.995 4.401 ;
      RECT 20.928 4.251 20.975 4.404 ;
      RECT 20.842 4.256 20.928 4.41 ;
      RECT 20.756 4.261 20.842 4.419 ;
      RECT 20.67 4.267 20.756 4.427 ;
      RECT 20.585 4.265 20.67 4.436 ;
      RECT 20.581 4.26 20.585 4.44 ;
      RECT 20.495 4.255 20.581 4.432 ;
      RECT 20.431 4.246 20.495 4.42 ;
      RECT 20.345 4.237 20.431 4.407 ;
      RECT 20.321 4.23 20.345 4.398 ;
      RECT 20.235 4.224 20.321 4.385 ;
      RECT 20.195 4.217 20.235 4.371 ;
      RECT 20.19 4.207 20.195 4.367 ;
      RECT 20.18 4.195 20.19 4.366 ;
      RECT 20.16 4.165 20.18 4.363 ;
      RECT 20.105 4.085 20.16 4.357 ;
      RECT 20.085 4.004 20.105 4.352 ;
      RECT 20.065 3.962 20.085 4.348 ;
      RECT 20.04 3.915 20.065 4.342 ;
      RECT 20.035 3.89 20.04 4.339 ;
      RECT 20 3.87 20.035 4.334 ;
      RECT 19.991 3.87 20 4.327 ;
      RECT 19.905 3.87 19.991 4.297 ;
      RECT 19.9 3.87 19.905 4.26 ;
      RECT 19.865 3.87 19.885 4.182 ;
      RECT 19.86 3.912 19.865 4.147 ;
      RECT 19.855 3.987 19.86 4.103 ;
      RECT 21.305 3.792 21.48 4.04 ;
      RECT 21.305 3.792 21.485 4.038 ;
      RECT 21.3 3.824 21.485 3.998 ;
      RECT 21.33 3.765 21.5 3.985 ;
      RECT 21.295 3.842 21.5 3.918 ;
      RECT 20.605 3.305 20.775 3.48 ;
      RECT 20.605 3.305 20.947 3.472 ;
      RECT 20.605 3.305 21.03 3.466 ;
      RECT 20.605 3.305 21.065 3.462 ;
      RECT 20.605 3.305 21.085 3.461 ;
      RECT 20.605 3.305 21.171 3.457 ;
      RECT 21.065 3.13 21.235 3.452 ;
      RECT 20.64 3.237 21.265 3.45 ;
      RECT 20.63 3.292 21.27 3.448 ;
      RECT 20.605 3.328 21.28 3.443 ;
      RECT 20.605 3.355 21.285 3.373 ;
      RECT 20.67 3.18 21.245 3.45 ;
      RECT 20.861 3.165 21.245 3.45 ;
      RECT 20.695 3.168 21.245 3.45 ;
      RECT 20.775 3.166 20.861 3.477 ;
      RECT 20.861 3.163 21.24 3.45 ;
      RECT 21.045 3.14 21.24 3.45 ;
      RECT 20.947 3.161 21.24 3.45 ;
      RECT 21.03 3.155 21.045 3.463 ;
      RECT 21.18 4.52 21.185 4.72 ;
      RECT 20.645 4.585 20.69 4.72 ;
      RECT 21.215 4.52 21.235 4.693 ;
      RECT 21.185 4.52 21.215 4.708 ;
      RECT 21.12 4.52 21.18 4.745 ;
      RECT 21.105 4.52 21.12 4.775 ;
      RECT 21.09 4.52 21.105 4.788 ;
      RECT 21.07 4.52 21.09 4.803 ;
      RECT 21.065 4.52 21.07 4.812 ;
      RECT 21.055 4.524 21.065 4.817 ;
      RECT 21.04 4.534 21.055 4.828 ;
      RECT 21.015 4.55 21.04 4.838 ;
      RECT 21.005 4.564 21.015 4.84 ;
      RECT 20.985 4.576 21.005 4.837 ;
      RECT 20.955 4.597 20.985 4.831 ;
      RECT 20.945 4.609 20.955 4.826 ;
      RECT 20.935 4.607 20.945 4.823 ;
      RECT 20.92 4.606 20.935 4.818 ;
      RECT 20.915 4.605 20.92 4.813 ;
      RECT 20.88 4.603 20.915 4.803 ;
      RECT 20.86 4.6 20.88 4.785 ;
      RECT 20.85 4.598 20.86 4.78 ;
      RECT 20.84 4.597 20.85 4.775 ;
      RECT 20.805 4.595 20.84 4.763 ;
      RECT 20.75 4.591 20.805 4.743 ;
      RECT 20.74 4.589 20.75 4.728 ;
      RECT 20.735 4.589 20.74 4.723 ;
      RECT 20.69 4.587 20.735 4.72 ;
      RECT 20.595 4.585 20.645 4.724 ;
      RECT 20.585 4.586 20.595 4.729 ;
      RECT 20.525 4.593 20.585 4.743 ;
      RECT 20.5 4.601 20.525 4.763 ;
      RECT 20.49 4.605 20.5 4.775 ;
      RECT 20.485 4.606 20.49 4.78 ;
      RECT 20.47 4.608 20.485 4.783 ;
      RECT 20.455 4.61 20.47 4.788 ;
      RECT 20.45 4.61 20.455 4.791 ;
      RECT 20.405 4.615 20.45 4.802 ;
      RECT 20.4 4.619 20.405 4.814 ;
      RECT 20.375 4.615 20.4 4.818 ;
      RECT 20.365 4.611 20.375 4.822 ;
      RECT 20.355 4.61 20.365 4.826 ;
      RECT 20.34 4.6 20.355 4.832 ;
      RECT 20.335 4.588 20.34 4.836 ;
      RECT 20.33 4.585 20.335 4.837 ;
      RECT 20.325 4.582 20.33 4.839 ;
      RECT 20.31 4.57 20.325 4.838 ;
      RECT 20.295 4.552 20.31 4.835 ;
      RECT 20.275 4.531 20.295 4.828 ;
      RECT 20.21 4.52 20.275 4.8 ;
      RECT 20.206 4.52 20.21 4.779 ;
      RECT 20.12 4.52 20.206 4.749 ;
      RECT 20.105 4.52 20.12 4.705 ;
      RECT 20.68 3.62 20.685 3.855 ;
      RECT 19.81 3.536 19.815 3.74 ;
      RECT 20.39 3.565 20.395 3.72 ;
      RECT 20.31 3.545 20.315 3.72 ;
      RECT 20.98 3.687 20.995 4.04 ;
      RECT 20.906 3.672 20.98 4.04 ;
      RECT 20.82 3.655 20.906 4.04 ;
      RECT 20.81 3.645 20.82 4.038 ;
      RECT 20.805 3.643 20.81 4.033 ;
      RECT 20.79 3.641 20.805 4.019 ;
      RECT 20.72 3.633 20.79 3.959 ;
      RECT 20.7 3.624 20.72 3.893 ;
      RECT 20.695 3.621 20.7 3.873 ;
      RECT 20.685 3.62 20.695 3.863 ;
      RECT 20.675 3.62 20.68 3.847 ;
      RECT 20.665 3.619 20.675 3.837 ;
      RECT 20.655 3.617 20.665 3.825 ;
      RECT 20.64 3.614 20.655 3.805 ;
      RECT 20.63 3.612 20.64 3.79 ;
      RECT 20.61 3.609 20.63 3.778 ;
      RECT 20.605 3.607 20.61 3.768 ;
      RECT 20.58 3.605 20.605 3.755 ;
      RECT 20.55 3.6 20.58 3.74 ;
      RECT 20.47 3.591 20.55 3.731 ;
      RECT 20.425 3.58 20.47 3.724 ;
      RECT 20.405 3.571 20.425 3.721 ;
      RECT 20.395 3.566 20.405 3.72 ;
      RECT 20.35 3.56 20.39 3.72 ;
      RECT 20.335 3.552 20.35 3.72 ;
      RECT 20.315 3.547 20.335 3.72 ;
      RECT 20.295 3.544 20.31 3.72 ;
      RECT 20.212 3.543 20.295 3.719 ;
      RECT 20.126 3.542 20.212 3.715 ;
      RECT 20.04 3.54 20.126 3.712 ;
      RECT 19.987 3.539 20.04 3.714 ;
      RECT 19.901 3.538 19.987 3.723 ;
      RECT 19.815 3.537 19.901 3.735 ;
      RECT 19.795 3.536 19.81 3.743 ;
      RECT 19.715 3.535 19.795 3.755 ;
      RECT 19.69 3.535 19.715 3.768 ;
      RECT 19.665 3.535 19.69 3.783 ;
      RECT 19.66 3.535 19.665 3.805 ;
      RECT 19.655 3.535 19.66 3.823 ;
      RECT 19.65 3.535 19.655 3.84 ;
      RECT 19.645 3.535 19.65 3.853 ;
      RECT 19.64 3.535 19.645 3.863 ;
      RECT 19.6 3.535 19.64 3.948 ;
      RECT 19.585 3.535 19.6 4.033 ;
      RECT 19.575 3.536 19.585 4.045 ;
      RECT 19.54 3.541 19.575 4.05 ;
      RECT 19.5 3.55 19.54 4.05 ;
      RECT 19.485 3.56 19.5 4.05 ;
      RECT 19.48 3.57 19.485 4.05 ;
      RECT 19.46 3.597 19.48 4.05 ;
      RECT 19.41 3.68 19.46 4.05 ;
      RECT 19.405 3.742 19.41 4.05 ;
      RECT 19.395 3.755 19.405 4.05 ;
      RECT 19.385 3.777 19.395 4.05 ;
      RECT 19.375 3.802 19.385 4.045 ;
      RECT 19.37 3.84 19.375 4.038 ;
      RECT 19.36 3.95 19.37 4.033 ;
      RECT 20.755 4.871 20.77 5.13 ;
      RECT 20.755 4.886 20.775 5.129 ;
      RECT 20.671 4.886 20.775 5.127 ;
      RECT 20.671 4.9 20.78 5.126 ;
      RECT 20.585 4.942 20.785 5.123 ;
      RECT 20.58 4.885 20.77 5.118 ;
      RECT 20.58 4.956 20.79 5.115 ;
      RECT 20.575 4.987 20.79 5.113 ;
      RECT 20.58 4.984 20.805 5.103 ;
      RECT 20.575 5.03 20.82 5.088 ;
      RECT 20.575 5.058 20.825 5.073 ;
      RECT 20.585 4.86 20.755 5.123 ;
      RECT 20.345 3.87 20.515 4.04 ;
      RECT 20.31 3.87 20.515 4.035 ;
      RECT 20.3 3.87 20.515 4.028 ;
      RECT 20.295 3.855 20.465 4.025 ;
      RECT 19.125 4.392 19.39 4.835 ;
      RECT 19.12 4.363 19.335 4.833 ;
      RECT 19.115 4.517 19.395 4.828 ;
      RECT 19.12 4.412 19.395 4.828 ;
      RECT 19.12 4.423 19.405 4.815 ;
      RECT 19.12 4.37 19.365 4.833 ;
      RECT 19.125 4.357 19.335 4.835 ;
      RECT 19.125 4.355 19.285 4.835 ;
      RECT 19.226 4.347 19.285 4.835 ;
      RECT 19.14 4.348 19.285 4.835 ;
      RECT 19.226 4.346 19.275 4.835 ;
      RECT 19.03 3.161 19.205 3.46 ;
      RECT 19.08 3.123 19.205 3.46 ;
      RECT 19.065 3.125 19.291 3.452 ;
      RECT 19.065 3.128 19.33 3.439 ;
      RECT 19.065 3.129 19.34 3.425 ;
      RECT 19.02 3.18 19.34 3.415 ;
      RECT 19.065 3.13 19.345 3.41 ;
      RECT 19.02 3.34 19.35 3.4 ;
      RECT 19.005 3.2 19.345 3.34 ;
      RECT 19 3.216 19.345 3.28 ;
      RECT 19.045 3.14 19.345 3.41 ;
      RECT 19.08 3.121 19.166 3.46 ;
      RECT 17.17 3.035 17.34 4.225 ;
      RECT 17.17 3.035 17.64 3.205 ;
      RECT 17.17 9.26 17.64 9.43 ;
      RECT 17.17 8.24 17.34 9.43 ;
      RECT 16.18 3.035 16.35 4.225 ;
      RECT 16.18 3.035 16.65 3.205 ;
      RECT 16.18 9.26 16.65 9.43 ;
      RECT 16.18 8.24 16.35 9.43 ;
      RECT 14.33 3.93 14.5 5.16 ;
      RECT 14.385 2.15 14.555 4.1 ;
      RECT 14.33 1.87 14.5 2.32 ;
      RECT 14.33 10.145 14.5 10.595 ;
      RECT 14.385 8.365 14.555 10.315 ;
      RECT 14.33 7.305 14.5 8.535 ;
      RECT 13.81 1.87 13.98 5.16 ;
      RECT 13.81 3.37 14.215 3.7 ;
      RECT 13.81 2.53 14.215 2.86 ;
      RECT 13.81 7.305 13.98 10.595 ;
      RECT 13.81 9.605 14.215 9.935 ;
      RECT 13.81 8.765 14.215 9.095 ;
      RECT 11.735 4.421 11.74 4.593 ;
      RECT 11.73 4.414 11.735 4.683 ;
      RECT 11.725 4.408 11.73 4.702 ;
      RECT 11.705 4.402 11.725 4.712 ;
      RECT 11.69 4.397 11.705 4.72 ;
      RECT 11.653 4.391 11.69 4.718 ;
      RECT 11.567 4.377 11.653 4.714 ;
      RECT 11.481 4.359 11.567 4.709 ;
      RECT 11.395 4.34 11.481 4.703 ;
      RECT 11.365 4.328 11.395 4.699 ;
      RECT 11.345 4.322 11.365 4.698 ;
      RECT 11.28 4.32 11.345 4.696 ;
      RECT 11.265 4.32 11.28 4.688 ;
      RECT 11.25 4.32 11.265 4.675 ;
      RECT 11.245 4.32 11.25 4.665 ;
      RECT 11.23 4.32 11.245 4.643 ;
      RECT 11.215 4.32 11.23 4.61 ;
      RECT 11.21 4.32 11.215 4.588 ;
      RECT 11.2 4.32 11.21 4.57 ;
      RECT 11.185 4.32 11.2 4.548 ;
      RECT 11.165 4.32 11.185 4.51 ;
      RECT 11.515 3.605 11.55 4.044 ;
      RECT 11.515 3.605 11.555 4.043 ;
      RECT 11.46 3.665 11.555 4.042 ;
      RECT 11.325 3.837 11.555 4.041 ;
      RECT 11.435 3.715 11.555 4.041 ;
      RECT 11.325 3.837 11.58 4.031 ;
      RECT 11.38 3.782 11.66 3.948 ;
      RECT 11.555 3.576 11.56 4.039 ;
      RECT 11.41 3.752 11.7 3.825 ;
      RECT 11.425 3.735 11.555 4.041 ;
      RECT 11.56 3.575 11.73 3.763 ;
      RECT 11.55 3.578 11.73 3.763 ;
      RECT 11.055 3.455 11.225 3.765 ;
      RECT 11.055 3.455 11.23 3.738 ;
      RECT 11.055 3.455 11.235 3.715 ;
      RECT 11.055 3.455 11.245 3.665 ;
      RECT 11.05 3.56 11.245 3.635 ;
      RECT 11.085 3.13 11.255 3.608 ;
      RECT 11.085 3.13 11.27 3.529 ;
      RECT 11.075 3.34 11.27 3.529 ;
      RECT 11.085 3.14 11.28 3.444 ;
      RECT 11.015 3.882 11.02 4.085 ;
      RECT 11.005 3.87 11.015 4.195 ;
      RECT 10.98 3.87 11.005 4.235 ;
      RECT 10.9 3.87 10.98 4.32 ;
      RECT 10.89 3.87 10.9 4.39 ;
      RECT 10.865 3.87 10.89 4.413 ;
      RECT 10.845 3.87 10.865 4.448 ;
      RECT 10.8 3.88 10.845 4.491 ;
      RECT 10.79 3.892 10.8 4.528 ;
      RECT 10.77 3.906 10.79 4.548 ;
      RECT 10.76 3.924 10.77 4.564 ;
      RECT 10.745 3.95 10.76 4.574 ;
      RECT 10.73 3.991 10.745 4.588 ;
      RECT 10.72 4.026 10.73 4.598 ;
      RECT 10.715 4.042 10.72 4.603 ;
      RECT 10.705 4.057 10.715 4.608 ;
      RECT 10.685 4.1 10.705 4.618 ;
      RECT 10.665 4.137 10.685 4.631 ;
      RECT 10.63 4.16 10.665 4.649 ;
      RECT 10.62 4.174 10.63 4.665 ;
      RECT 10.6 4.184 10.62 4.675 ;
      RECT 10.595 4.193 10.6 4.683 ;
      RECT 10.585 4.2 10.595 4.69 ;
      RECT 10.575 4.207 10.585 4.698 ;
      RECT 10.56 4.217 10.575 4.706 ;
      RECT 10.55 4.231 10.56 4.716 ;
      RECT 10.54 4.243 10.55 4.728 ;
      RECT 10.525 4.265 10.54 4.741 ;
      RECT 10.515 4.287 10.525 4.752 ;
      RECT 10.505 4.307 10.515 4.761 ;
      RECT 10.5 4.322 10.505 4.768 ;
      RECT 10.47 4.355 10.5 4.782 ;
      RECT 10.46 4.39 10.47 4.797 ;
      RECT 10.455 4.397 10.46 4.803 ;
      RECT 10.435 4.412 10.455 4.81 ;
      RECT 10.43 4.427 10.435 4.818 ;
      RECT 10.425 4.436 10.43 4.823 ;
      RECT 10.41 4.442 10.425 4.83 ;
      RECT 10.405 4.448 10.41 4.838 ;
      RECT 10.4 4.452 10.405 4.845 ;
      RECT 10.395 4.456 10.4 4.855 ;
      RECT 10.385 4.461 10.395 4.865 ;
      RECT 10.365 4.472 10.385 4.893 ;
      RECT 10.35 4.484 10.365 4.92 ;
      RECT 10.33 4.497 10.35 4.945 ;
      RECT 10.31 4.512 10.33 4.969 ;
      RECT 10.295 4.527 10.31 4.984 ;
      RECT 10.29 4.538 10.295 4.993 ;
      RECT 10.225 4.583 10.29 5.003 ;
      RECT 10.19 4.642 10.225 5.016 ;
      RECT 10.185 4.665 10.19 5.022 ;
      RECT 10.18 4.672 10.185 5.024 ;
      RECT 10.165 4.682 10.18 5.027 ;
      RECT 10.135 4.707 10.165 5.031 ;
      RECT 10.13 4.725 10.135 5.035 ;
      RECT 10.125 4.732 10.13 5.036 ;
      RECT 10.105 4.74 10.125 5.04 ;
      RECT 10.095 4.747 10.105 5.044 ;
      RECT 10.051 4.758 10.095 5.051 ;
      RECT 9.965 4.786 10.051 5.067 ;
      RECT 9.905 4.81 9.965 5.085 ;
      RECT 9.86 4.82 9.905 5.099 ;
      RECT 9.801 4.828 9.86 5.113 ;
      RECT 9.715 4.835 9.801 5.132 ;
      RECT 9.69 4.84 9.715 5.147 ;
      RECT 9.61 4.843 9.69 5.15 ;
      RECT 9.53 4.847 9.61 5.137 ;
      RECT 9.521 4.85 9.53 5.122 ;
      RECT 9.435 4.85 9.521 5.107 ;
      RECT 9.375 4.852 9.435 5.084 ;
      RECT 9.371 4.855 9.375 5.074 ;
      RECT 9.285 4.855 9.371 5.059 ;
      RECT 9.21 4.855 9.285 5.035 ;
      RECT 10.525 3.864 10.535 4.04 ;
      RECT 10.48 3.831 10.525 4.04 ;
      RECT 10.435 3.782 10.48 4.04 ;
      RECT 10.405 3.752 10.435 4.041 ;
      RECT 10.4 3.735 10.405 4.042 ;
      RECT 10.375 3.715 10.4 4.043 ;
      RECT 10.36 3.69 10.375 4.044 ;
      RECT 10.355 3.677 10.36 4.045 ;
      RECT 10.35 3.671 10.355 4.043 ;
      RECT 10.345 3.663 10.35 4.037 ;
      RECT 10.32 3.655 10.345 4.017 ;
      RECT 10.3 3.644 10.32 3.988 ;
      RECT 10.27 3.629 10.3 3.959 ;
      RECT 10.25 3.615 10.27 3.931 ;
      RECT 10.24 3.609 10.25 3.91 ;
      RECT 10.235 3.606 10.24 3.893 ;
      RECT 10.23 3.603 10.235 3.878 ;
      RECT 10.215 3.598 10.23 3.843 ;
      RECT 10.21 3.594 10.215 3.81 ;
      RECT 10.19 3.589 10.21 3.786 ;
      RECT 10.16 3.581 10.19 3.751 ;
      RECT 10.145 3.575 10.16 3.728 ;
      RECT 10.105 3.568 10.145 3.713 ;
      RECT 10.08 3.56 10.105 3.693 ;
      RECT 10.06 3.555 10.08 3.683 ;
      RECT 10.025 3.549 10.06 3.678 ;
      RECT 9.98 3.54 10.025 3.677 ;
      RECT 9.95 3.536 9.98 3.679 ;
      RECT 9.865 3.544 9.95 3.683 ;
      RECT 9.795 3.555 9.865 3.705 ;
      RECT 9.782 3.561 9.795 3.728 ;
      RECT 9.696 3.568 9.782 3.75 ;
      RECT 9.61 3.58 9.696 3.787 ;
      RECT 9.61 3.957 9.62 4.195 ;
      RECT 9.605 3.586 9.61 3.81 ;
      RECT 9.6 3.842 9.61 4.195 ;
      RECT 9.6 3.587 9.605 3.815 ;
      RECT 9.595 3.588 9.6 4.195 ;
      RECT 9.571 3.59 9.595 4.196 ;
      RECT 9.485 3.598 9.571 4.198 ;
      RECT 9.465 3.612 9.485 4.201 ;
      RECT 9.46 3.64 9.465 4.202 ;
      RECT 9.455 3.652 9.46 4.203 ;
      RECT 9.45 3.667 9.455 4.204 ;
      RECT 9.44 3.697 9.45 4.205 ;
      RECT 9.435 3.735 9.44 4.203 ;
      RECT 9.43 3.755 9.435 4.198 ;
      RECT 9.415 3.79 9.43 4.183 ;
      RECT 9.405 3.842 9.415 4.163 ;
      RECT 9.4 3.872 9.405 4.151 ;
      RECT 9.385 3.885 9.4 4.134 ;
      RECT 9.36 3.889 9.385 4.101 ;
      RECT 9.345 3.887 9.36 4.078 ;
      RECT 9.33 3.886 9.345 4.075 ;
      RECT 9.27 3.884 9.33 4.073 ;
      RECT 9.26 3.882 9.27 4.068 ;
      RECT 9.22 3.881 9.26 4.065 ;
      RECT 9.15 3.878 9.22 4.063 ;
      RECT 9.095 3.876 9.15 4.058 ;
      RECT 9.025 3.87 9.095 4.053 ;
      RECT 9.016 3.87 9.025 4.05 ;
      RECT 8.93 3.87 9.016 4.045 ;
      RECT 8.925 3.87 8.93 4.04 ;
      RECT 10.23 3.105 10.405 3.455 ;
      RECT 10.23 3.12 10.415 3.453 ;
      RECT 10.205 3.07 10.35 3.45 ;
      RECT 10.185 3.071 10.35 3.443 ;
      RECT 10.175 3.072 10.36 3.438 ;
      RECT 10.145 3.073 10.36 3.425 ;
      RECT 10.095 3.074 10.36 3.401 ;
      RECT 10.09 3.076 10.36 3.386 ;
      RECT 10.09 3.142 10.42 3.38 ;
      RECT 10.07 3.083 10.375 3.36 ;
      RECT 10.06 3.092 10.385 3.215 ;
      RECT 10.07 3.087 10.385 3.36 ;
      RECT 10.09 3.077 10.375 3.386 ;
      RECT 9.675 4.402 9.845 4.69 ;
      RECT 9.67 4.42 9.855 4.685 ;
      RECT 9.635 4.428 9.92 4.605 ;
      RECT 9.635 4.428 10.006 4.595 ;
      RECT 9.635 4.428 10.06 4.541 ;
      RECT 9.92 4.325 10.09 4.509 ;
      RECT 9.635 4.48 10.095 4.497 ;
      RECT 9.62 4.45 10.09 4.493 ;
      RECT 9.88 4.332 9.92 4.644 ;
      RECT 9.76 4.369 10.09 4.509 ;
      RECT 9.855 4.344 9.88 4.67 ;
      RECT 9.845 4.351 10.09 4.509 ;
      RECT 9.976 3.815 10.045 4.074 ;
      RECT 9.976 3.87 10.05 4.073 ;
      RECT 9.89 3.87 10.05 4.072 ;
      RECT 9.885 3.87 10.055 4.065 ;
      RECT 9.875 3.815 10.045 4.06 ;
      RECT 9.255 3.114 9.43 3.415 ;
      RECT 9.24 3.102 9.255 3.4 ;
      RECT 9.21 3.101 9.24 3.353 ;
      RECT 9.21 3.119 9.435 3.348 ;
      RECT 9.195 3.103 9.255 3.313 ;
      RECT 9.19 3.125 9.445 3.213 ;
      RECT 9.19 3.108 9.341 3.213 ;
      RECT 9.19 3.11 9.345 3.213 ;
      RECT 9.195 3.106 9.341 3.313 ;
      RECT 9.3 4.342 9.305 4.69 ;
      RECT 9.29 4.332 9.3 4.696 ;
      RECT 9.255 4.322 9.29 4.698 ;
      RECT 9.217 4.317 9.255 4.702 ;
      RECT 9.131 4.31 9.217 4.709 ;
      RECT 9.045 4.3 9.131 4.719 ;
      RECT 9 4.295 9.045 4.727 ;
      RECT 8.996 4.295 9 4.731 ;
      RECT 8.91 4.295 8.996 4.738 ;
      RECT 8.895 4.295 8.91 4.738 ;
      RECT 8.885 4.293 8.895 4.71 ;
      RECT 8.875 4.289 8.885 4.653 ;
      RECT 8.855 4.283 8.875 4.585 ;
      RECT 8.85 4.279 8.855 4.533 ;
      RECT 8.84 4.278 8.85 4.5 ;
      RECT 8.79 4.276 8.84 4.485 ;
      RECT 8.765 4.274 8.79 4.48 ;
      RECT 8.722 4.272 8.765 4.476 ;
      RECT 8.636 4.268 8.722 4.464 ;
      RECT 8.55 4.263 8.636 4.448 ;
      RECT 8.52 4.26 8.55 4.435 ;
      RECT 8.495 4.259 8.52 4.423 ;
      RECT 8.49 4.259 8.495 4.413 ;
      RECT 8.45 4.258 8.49 4.405 ;
      RECT 8.435 4.257 8.45 4.398 ;
      RECT 8.385 4.256 8.435 4.39 ;
      RECT 8.383 4.255 8.385 4.385 ;
      RECT 8.297 4.253 8.383 4.385 ;
      RECT 8.211 4.248 8.297 4.385 ;
      RECT 8.125 4.244 8.211 4.385 ;
      RECT 8.076 4.24 8.125 4.383 ;
      RECT 7.99 4.237 8.076 4.378 ;
      RECT 7.967 4.234 7.99 4.374 ;
      RECT 7.881 4.231 7.967 4.369 ;
      RECT 7.795 4.227 7.881 4.36 ;
      RECT 7.77 4.22 7.795 4.355 ;
      RECT 7.71 4.185 7.77 4.352 ;
      RECT 7.69 4.11 7.71 4.349 ;
      RECT 7.685 4.052 7.69 4.348 ;
      RECT 7.66 3.992 7.685 4.347 ;
      RECT 7.585 3.87 7.66 4.343 ;
      RECT 7.575 3.87 7.585 4.335 ;
      RECT 7.56 3.87 7.575 4.325 ;
      RECT 7.545 3.87 7.56 4.295 ;
      RECT 7.53 3.87 7.545 4.24 ;
      RECT 7.515 3.87 7.53 4.178 ;
      RECT 7.49 3.87 7.515 4.103 ;
      RECT 7.485 3.87 7.49 4.053 ;
      RECT 8.83 3.415 8.85 3.724 ;
      RECT 8.816 3.417 8.865 3.721 ;
      RECT 8.816 3.422 8.885 3.712 ;
      RECT 8.73 3.42 8.865 3.706 ;
      RECT 8.73 3.428 8.92 3.689 ;
      RECT 8.695 3.43 8.92 3.688 ;
      RECT 8.665 3.438 8.92 3.679 ;
      RECT 8.655 3.443 8.94 3.665 ;
      RECT 8.695 3.433 8.94 3.665 ;
      RECT 8.695 3.436 8.95 3.653 ;
      RECT 8.665 3.438 8.96 3.64 ;
      RECT 8.665 3.442 8.97 3.583 ;
      RECT 8.655 3.447 8.975 3.498 ;
      RECT 8.816 3.415 8.85 3.721 ;
      RECT 8.255 3.518 8.26 3.73 ;
      RECT 8.13 3.515 8.145 3.73 ;
      RECT 7.595 3.545 7.665 3.73 ;
      RECT 7.48 3.545 7.515 3.725 ;
      RECT 8.601 3.847 8.62 4.041 ;
      RECT 8.515 3.802 8.601 4.042 ;
      RECT 8.505 3.755 8.515 4.044 ;
      RECT 8.5 3.735 8.505 4.045 ;
      RECT 8.48 3.7 8.5 4.046 ;
      RECT 8.465 3.65 8.48 4.047 ;
      RECT 8.445 3.587 8.465 4.048 ;
      RECT 8.435 3.55 8.445 4.049 ;
      RECT 8.42 3.539 8.435 4.05 ;
      RECT 8.415 3.531 8.42 4.048 ;
      RECT 8.405 3.53 8.415 4.04 ;
      RECT 8.375 3.527 8.405 4.019 ;
      RECT 8.3 3.522 8.375 3.964 ;
      RECT 8.285 3.518 8.3 3.91 ;
      RECT 8.275 3.518 8.285 3.805 ;
      RECT 8.26 3.518 8.275 3.738 ;
      RECT 8.245 3.518 8.255 3.728 ;
      RECT 8.19 3.517 8.245 3.725 ;
      RECT 8.145 3.515 8.19 3.728 ;
      RECT 8.117 3.515 8.13 3.731 ;
      RECT 8.031 3.519 8.117 3.733 ;
      RECT 7.945 3.525 8.031 3.738 ;
      RECT 7.925 3.529 7.945 3.74 ;
      RECT 7.923 3.53 7.925 3.739 ;
      RECT 7.837 3.532 7.923 3.738 ;
      RECT 7.751 3.537 7.837 3.735 ;
      RECT 7.665 3.542 7.751 3.732 ;
      RECT 7.515 3.545 7.595 3.728 ;
      RECT 8.175 7.305 8.345 10.595 ;
      RECT 8.175 9.605 8.58 9.935 ;
      RECT 8.175 8.765 8.58 9.095 ;
      RECT 8.291 4.52 8.34 4.854 ;
      RECT 8.291 4.52 8.345 4.853 ;
      RECT 8.205 4.52 8.345 4.852 ;
      RECT 7.98 4.628 8.35 4.85 ;
      RECT 8.205 4.52 8.375 4.843 ;
      RECT 8.175 4.532 8.38 4.834 ;
      RECT 8.16 4.55 8.385 4.831 ;
      RECT 7.975 4.634 8.385 4.758 ;
      RECT 7.97 4.641 8.385 4.718 ;
      RECT 7.985 4.607 8.385 4.831 ;
      RECT 8.146 4.553 8.35 4.85 ;
      RECT 8.06 4.573 8.385 4.831 ;
      RECT 8.16 4.547 8.38 4.834 ;
      RECT 7.93 3.871 8.12 4.065 ;
      RECT 7.925 3.873 8.12 4.064 ;
      RECT 7.92 3.877 8.135 4.061 ;
      RECT 7.935 3.87 8.135 4.061 ;
      RECT 7.92 3.98 8.14 4.056 ;
      RECT 7.215 4.48 7.306 4.778 ;
      RECT 7.21 4.482 7.385 4.773 ;
      RECT 7.215 4.48 7.385 4.773 ;
      RECT 7.21 4.486 7.405 4.771 ;
      RECT 7.21 4.541 7.445 4.77 ;
      RECT 7.21 4.576 7.46 4.764 ;
      RECT 7.21 4.61 7.47 4.754 ;
      RECT 7.2 4.49 7.405 4.605 ;
      RECT 7.2 4.51 7.42 4.605 ;
      RECT 7.2 4.493 7.41 4.605 ;
      RECT 7.425 3.261 7.43 3.323 ;
      RECT 7.42 3.183 7.425 3.346 ;
      RECT 7.415 3.14 7.42 3.357 ;
      RECT 7.41 3.13 7.415 3.369 ;
      RECT 7.405 3.13 7.41 3.378 ;
      RECT 7.38 3.13 7.405 3.41 ;
      RECT 7.375 3.13 7.38 3.443 ;
      RECT 7.36 3.13 7.375 3.468 ;
      RECT 7.35 3.13 7.36 3.495 ;
      RECT 7.345 3.13 7.35 3.508 ;
      RECT 7.34 3.13 7.345 3.523 ;
      RECT 7.33 3.13 7.34 3.538 ;
      RECT 7.325 3.13 7.33 3.558 ;
      RECT 7.3 3.13 7.325 3.593 ;
      RECT 7.255 3.13 7.3 3.638 ;
      RECT 7.245 3.13 7.255 3.651 ;
      RECT 7.16 3.215 7.245 3.658 ;
      RECT 7.125 3.337 7.16 3.667 ;
      RECT 7.12 3.377 7.125 3.671 ;
      RECT 7.1 3.4 7.12 3.673 ;
      RECT 7.095 3.43 7.1 3.676 ;
      RECT 7.085 3.442 7.095 3.677 ;
      RECT 7.04 3.465 7.085 3.682 ;
      RECT 7 3.495 7.04 3.69 ;
      RECT 6.965 3.507 7 3.696 ;
      RECT 6.96 3.512 6.965 3.7 ;
      RECT 6.89 3.522 6.96 3.707 ;
      RECT 6.85 3.532 6.89 3.717 ;
      RECT 6.83 3.537 6.85 3.723 ;
      RECT 6.82 3.541 6.83 3.728 ;
      RECT 6.815 3.544 6.82 3.731 ;
      RECT 6.805 3.545 6.815 3.732 ;
      RECT 6.78 3.547 6.805 3.736 ;
      RECT 6.77 3.552 6.78 3.739 ;
      RECT 6.725 3.56 6.77 3.74 ;
      RECT 6.6 3.565 6.725 3.74 ;
      RECT 7.155 3.862 7.175 4.044 ;
      RECT 7.106 3.847 7.155 4.043 ;
      RECT 7.02 3.862 7.175 4.041 ;
      RECT 7.005 3.862 7.175 4.04 ;
      RECT 6.97 3.84 7.14 4.025 ;
      RECT 7.04 4.86 7.055 5.069 ;
      RECT 7.04 4.868 7.06 5.068 ;
      RECT 6.985 4.868 7.06 5.067 ;
      RECT 6.965 4.872 7.065 5.065 ;
      RECT 6.945 4.822 6.985 5.064 ;
      RECT 6.89 4.88 7.07 5.062 ;
      RECT 6.855 4.837 6.985 5.06 ;
      RECT 6.851 4.84 7.04 5.059 ;
      RECT 6.765 4.848 7.04 5.057 ;
      RECT 6.765 4.892 7.075 5.05 ;
      RECT 6.755 4.985 7.075 5.048 ;
      RECT 6.765 4.904 7.08 5.033 ;
      RECT 6.765 4.925 7.095 5.003 ;
      RECT 6.765 4.952 7.1 4.973 ;
      RECT 6.89 4.83 6.985 5.062 ;
      RECT 6.52 3.875 6.525 4.413 ;
      RECT 6.325 4.205 6.33 4.4 ;
      RECT 4.625 3.87 4.64 4.25 ;
      RECT 6.69 3.87 6.695 4.04 ;
      RECT 6.685 3.87 6.69 4.05 ;
      RECT 6.68 3.87 6.685 4.063 ;
      RECT 6.655 3.87 6.68 4.105 ;
      RECT 6.63 3.87 6.655 4.178 ;
      RECT 6.615 3.87 6.63 4.23 ;
      RECT 6.61 3.87 6.615 4.26 ;
      RECT 6.585 3.87 6.61 4.3 ;
      RECT 6.57 3.87 6.585 4.355 ;
      RECT 6.565 3.87 6.57 4.388 ;
      RECT 6.54 3.87 6.565 4.408 ;
      RECT 6.525 3.87 6.54 4.414 ;
      RECT 6.455 3.905 6.52 4.41 ;
      RECT 6.405 3.96 6.455 4.405 ;
      RECT 6.395 3.992 6.405 4.403 ;
      RECT 6.39 4.017 6.395 4.403 ;
      RECT 6.37 4.09 6.39 4.403 ;
      RECT 6.36 4.17 6.37 4.402 ;
      RECT 6.345 4.2 6.36 4.402 ;
      RECT 6.33 4.205 6.345 4.401 ;
      RECT 6.27 4.207 6.325 4.398 ;
      RECT 6.24 4.212 6.27 4.394 ;
      RECT 6.238 4.215 6.24 4.393 ;
      RECT 6.152 4.217 6.238 4.39 ;
      RECT 6.066 4.223 6.152 4.384 ;
      RECT 5.98 4.228 6.066 4.378 ;
      RECT 5.907 4.233 5.98 4.379 ;
      RECT 5.821 4.239 5.907 4.387 ;
      RECT 5.735 4.245 5.821 4.396 ;
      RECT 5.715 4.249 5.735 4.401 ;
      RECT 5.668 4.251 5.715 4.404 ;
      RECT 5.582 4.256 5.668 4.41 ;
      RECT 5.496 4.261 5.582 4.419 ;
      RECT 5.41 4.267 5.496 4.427 ;
      RECT 5.325 4.265 5.41 4.436 ;
      RECT 5.321 4.26 5.325 4.44 ;
      RECT 5.235 4.255 5.321 4.432 ;
      RECT 5.171 4.246 5.235 4.42 ;
      RECT 5.085 4.237 5.171 4.407 ;
      RECT 5.061 4.23 5.085 4.398 ;
      RECT 4.975 4.224 5.061 4.385 ;
      RECT 4.935 4.217 4.975 4.371 ;
      RECT 4.93 4.207 4.935 4.367 ;
      RECT 4.92 4.195 4.93 4.366 ;
      RECT 4.9 4.165 4.92 4.363 ;
      RECT 4.845 4.085 4.9 4.357 ;
      RECT 4.825 4.004 4.845 4.352 ;
      RECT 4.805 3.962 4.825 4.348 ;
      RECT 4.78 3.915 4.805 4.342 ;
      RECT 4.775 3.89 4.78 4.339 ;
      RECT 4.74 3.87 4.775 4.334 ;
      RECT 4.731 3.87 4.74 4.327 ;
      RECT 4.645 3.87 4.731 4.297 ;
      RECT 4.64 3.87 4.645 4.26 ;
      RECT 4.605 3.87 4.625 4.182 ;
      RECT 4.6 3.912 4.605 4.147 ;
      RECT 4.595 3.987 4.6 4.103 ;
      RECT 6.045 3.792 6.22 4.04 ;
      RECT 6.045 3.792 6.225 4.038 ;
      RECT 6.04 3.824 6.225 3.998 ;
      RECT 6.07 3.765 6.24 3.985 ;
      RECT 6.035 3.842 6.24 3.918 ;
      RECT 5.345 3.305 5.515 3.48 ;
      RECT 5.345 3.305 5.687 3.472 ;
      RECT 5.345 3.305 5.77 3.466 ;
      RECT 5.345 3.305 5.805 3.462 ;
      RECT 5.345 3.305 5.825 3.461 ;
      RECT 5.345 3.305 5.911 3.457 ;
      RECT 5.805 3.13 5.975 3.452 ;
      RECT 5.38 3.237 6.005 3.45 ;
      RECT 5.37 3.292 6.01 3.448 ;
      RECT 5.345 3.328 6.02 3.443 ;
      RECT 5.345 3.355 6.025 3.373 ;
      RECT 5.41 3.18 5.985 3.45 ;
      RECT 5.601 3.165 5.985 3.45 ;
      RECT 5.435 3.168 5.985 3.45 ;
      RECT 5.515 3.166 5.601 3.477 ;
      RECT 5.601 3.163 5.98 3.45 ;
      RECT 5.785 3.14 5.98 3.45 ;
      RECT 5.687 3.161 5.98 3.45 ;
      RECT 5.77 3.155 5.785 3.463 ;
      RECT 5.92 4.52 5.925 4.72 ;
      RECT 5.385 4.585 5.43 4.72 ;
      RECT 5.955 4.52 5.975 4.693 ;
      RECT 5.925 4.52 5.955 4.708 ;
      RECT 5.86 4.52 5.92 4.745 ;
      RECT 5.845 4.52 5.86 4.775 ;
      RECT 5.83 4.52 5.845 4.788 ;
      RECT 5.81 4.52 5.83 4.803 ;
      RECT 5.805 4.52 5.81 4.812 ;
      RECT 5.795 4.524 5.805 4.817 ;
      RECT 5.78 4.534 5.795 4.828 ;
      RECT 5.755 4.55 5.78 4.838 ;
      RECT 5.745 4.564 5.755 4.84 ;
      RECT 5.725 4.576 5.745 4.837 ;
      RECT 5.695 4.597 5.725 4.831 ;
      RECT 5.685 4.609 5.695 4.826 ;
      RECT 5.675 4.607 5.685 4.823 ;
      RECT 5.66 4.606 5.675 4.818 ;
      RECT 5.655 4.605 5.66 4.813 ;
      RECT 5.62 4.603 5.655 4.803 ;
      RECT 5.6 4.6 5.62 4.785 ;
      RECT 5.59 4.598 5.6 4.78 ;
      RECT 5.58 4.597 5.59 4.775 ;
      RECT 5.545 4.595 5.58 4.763 ;
      RECT 5.49 4.591 5.545 4.743 ;
      RECT 5.48 4.589 5.49 4.728 ;
      RECT 5.475 4.589 5.48 4.723 ;
      RECT 5.43 4.587 5.475 4.72 ;
      RECT 5.335 4.585 5.385 4.724 ;
      RECT 5.325 4.586 5.335 4.729 ;
      RECT 5.265 4.593 5.325 4.743 ;
      RECT 5.24 4.601 5.265 4.763 ;
      RECT 5.23 4.605 5.24 4.775 ;
      RECT 5.225 4.606 5.23 4.78 ;
      RECT 5.21 4.608 5.225 4.783 ;
      RECT 5.195 4.61 5.21 4.788 ;
      RECT 5.19 4.61 5.195 4.791 ;
      RECT 5.145 4.615 5.19 4.802 ;
      RECT 5.14 4.619 5.145 4.814 ;
      RECT 5.115 4.615 5.14 4.818 ;
      RECT 5.105 4.611 5.115 4.822 ;
      RECT 5.095 4.61 5.105 4.826 ;
      RECT 5.08 4.6 5.095 4.832 ;
      RECT 5.075 4.588 5.08 4.836 ;
      RECT 5.07 4.585 5.075 4.837 ;
      RECT 5.065 4.582 5.07 4.839 ;
      RECT 5.05 4.57 5.065 4.838 ;
      RECT 5.035 4.552 5.05 4.835 ;
      RECT 5.015 4.531 5.035 4.828 ;
      RECT 4.95 4.52 5.015 4.8 ;
      RECT 4.946 4.52 4.95 4.779 ;
      RECT 4.86 4.52 4.946 4.749 ;
      RECT 4.845 4.52 4.86 4.705 ;
      RECT 5.42 3.62 5.425 3.855 ;
      RECT 4.55 3.536 4.555 3.74 ;
      RECT 5.13 3.565 5.135 3.72 ;
      RECT 5.05 3.545 5.055 3.72 ;
      RECT 5.72 3.687 5.735 4.04 ;
      RECT 5.646 3.672 5.72 4.04 ;
      RECT 5.56 3.655 5.646 4.04 ;
      RECT 5.55 3.645 5.56 4.038 ;
      RECT 5.545 3.643 5.55 4.033 ;
      RECT 5.53 3.641 5.545 4.019 ;
      RECT 5.46 3.633 5.53 3.959 ;
      RECT 5.44 3.624 5.46 3.893 ;
      RECT 5.435 3.621 5.44 3.873 ;
      RECT 5.425 3.62 5.435 3.863 ;
      RECT 5.415 3.62 5.42 3.847 ;
      RECT 5.405 3.619 5.415 3.837 ;
      RECT 5.395 3.617 5.405 3.825 ;
      RECT 5.38 3.614 5.395 3.805 ;
      RECT 5.37 3.612 5.38 3.79 ;
      RECT 5.35 3.609 5.37 3.778 ;
      RECT 5.345 3.607 5.35 3.768 ;
      RECT 5.32 3.605 5.345 3.755 ;
      RECT 5.29 3.6 5.32 3.74 ;
      RECT 5.21 3.591 5.29 3.731 ;
      RECT 5.165 3.58 5.21 3.724 ;
      RECT 5.145 3.571 5.165 3.721 ;
      RECT 5.135 3.566 5.145 3.72 ;
      RECT 5.09 3.56 5.13 3.72 ;
      RECT 5.075 3.552 5.09 3.72 ;
      RECT 5.055 3.547 5.075 3.72 ;
      RECT 5.035 3.544 5.05 3.72 ;
      RECT 4.952 3.543 5.035 3.719 ;
      RECT 4.866 3.542 4.952 3.715 ;
      RECT 4.78 3.54 4.866 3.712 ;
      RECT 4.727 3.539 4.78 3.714 ;
      RECT 4.641 3.538 4.727 3.723 ;
      RECT 4.555 3.537 4.641 3.735 ;
      RECT 4.535 3.536 4.55 3.743 ;
      RECT 4.455 3.535 4.535 3.755 ;
      RECT 4.43 3.535 4.455 3.768 ;
      RECT 4.405 3.535 4.43 3.783 ;
      RECT 4.4 3.535 4.405 3.805 ;
      RECT 4.395 3.535 4.4 3.823 ;
      RECT 4.39 3.535 4.395 3.84 ;
      RECT 4.385 3.535 4.39 3.853 ;
      RECT 4.38 3.535 4.385 3.863 ;
      RECT 4.34 3.535 4.38 3.948 ;
      RECT 4.325 3.535 4.34 4.033 ;
      RECT 4.315 3.536 4.325 4.045 ;
      RECT 4.28 3.541 4.315 4.05 ;
      RECT 4.24 3.55 4.28 4.05 ;
      RECT 4.225 3.56 4.24 4.05 ;
      RECT 4.22 3.57 4.225 4.05 ;
      RECT 4.2 3.597 4.22 4.05 ;
      RECT 4.15 3.68 4.2 4.05 ;
      RECT 4.145 3.742 4.15 4.05 ;
      RECT 4.135 3.755 4.145 4.05 ;
      RECT 4.125 3.777 4.135 4.05 ;
      RECT 4.115 3.802 4.125 4.045 ;
      RECT 4.11 3.84 4.115 4.038 ;
      RECT 4.1 3.95 4.11 4.033 ;
      RECT 5.495 4.871 5.51 5.13 ;
      RECT 5.495 4.886 5.515 5.129 ;
      RECT 5.411 4.886 5.515 5.127 ;
      RECT 5.411 4.9 5.52 5.126 ;
      RECT 5.325 4.942 5.525 5.123 ;
      RECT 5.32 4.885 5.51 5.118 ;
      RECT 5.32 4.956 5.53 5.115 ;
      RECT 5.315 4.987 5.53 5.113 ;
      RECT 5.32 4.984 5.545 5.103 ;
      RECT 5.315 5.03 5.56 5.088 ;
      RECT 5.315 5.058 5.565 5.073 ;
      RECT 5.325 4.86 5.495 5.123 ;
      RECT 5.085 3.87 5.255 4.04 ;
      RECT 5.05 3.87 5.255 4.035 ;
      RECT 5.04 3.87 5.255 4.028 ;
      RECT 5.035 3.855 5.205 4.025 ;
      RECT 3.865 4.392 4.13 4.835 ;
      RECT 3.86 4.363 4.075 4.833 ;
      RECT 3.855 4.517 4.135 4.828 ;
      RECT 3.86 4.412 4.135 4.828 ;
      RECT 3.86 4.423 4.145 4.815 ;
      RECT 3.86 4.37 4.105 4.833 ;
      RECT 3.865 4.357 4.075 4.835 ;
      RECT 3.865 4.355 4.025 4.835 ;
      RECT 3.966 4.347 4.025 4.835 ;
      RECT 3.88 4.348 4.025 4.835 ;
      RECT 3.966 4.346 4.015 4.835 ;
      RECT 3.77 3.161 3.945 3.46 ;
      RECT 3.82 3.123 3.945 3.46 ;
      RECT 3.805 3.125 4.031 3.452 ;
      RECT 3.805 3.128 4.07 3.439 ;
      RECT 3.805 3.129 4.08 3.425 ;
      RECT 3.76 3.18 4.08 3.415 ;
      RECT 3.805 3.13 4.085 3.41 ;
      RECT 3.76 3.34 4.09 3.4 ;
      RECT 3.745 3.2 4.085 3.34 ;
      RECT 3.74 3.216 4.085 3.28 ;
      RECT 3.785 3.14 4.085 3.41 ;
      RECT 3.82 3.121 3.906 3.46 ;
      RECT 1.2 10.145 1.37 10.595 ;
      RECT 1.255 8.365 1.425 10.315 ;
      RECT 1.2 7.305 1.37 8.535 ;
      RECT 0.68 7.305 0.85 10.595 ;
      RECT 0.68 9.605 1.085 9.935 ;
      RECT 0.68 8.765 1.085 9.095 ;
      RECT 78.58 7.31 78.75 8.78 ;
      RECT 78.58 10.09 78.75 10.6 ;
      RECT 77.59 1.865 77.76 2.375 ;
      RECT 77.59 3.685 77.76 5.155 ;
      RECT 77.59 7.31 77.76 8.78 ;
      RECT 77.59 10.09 77.76 10.6 ;
      RECT 76.23 1.87 76.4 5.16 ;
      RECT 76.23 7.305 76.4 10.595 ;
      RECT 75.8 1.87 75.97 2.38 ;
      RECT 75.8 2.95 75.97 5.16 ;
      RECT 75.8 7.305 75.97 9.515 ;
      RECT 75.8 10.085 75.97 10.595 ;
      RECT 70.595 7.305 70.765 10.595 ;
      RECT 70.165 7.305 70.335 9.515 ;
      RECT 70.165 10.085 70.335 10.595 ;
      RECT 63.32 7.31 63.49 8.78 ;
      RECT 63.32 10.09 63.49 10.6 ;
      RECT 62.33 1.865 62.5 2.375 ;
      RECT 62.33 3.685 62.5 5.155 ;
      RECT 62.33 7.31 62.5 8.78 ;
      RECT 62.33 10.09 62.5 10.6 ;
      RECT 60.97 1.87 61.14 5.16 ;
      RECT 60.97 7.305 61.14 10.595 ;
      RECT 60.54 1.87 60.71 2.38 ;
      RECT 60.54 2.95 60.71 5.16 ;
      RECT 60.54 7.305 60.71 9.515 ;
      RECT 60.54 10.085 60.71 10.595 ;
      RECT 55.335 7.305 55.505 10.595 ;
      RECT 54.905 7.305 55.075 9.515 ;
      RECT 54.905 10.085 55.075 10.595 ;
      RECT 48.06 7.31 48.23 8.78 ;
      RECT 48.06 10.09 48.23 10.6 ;
      RECT 47.07 1.865 47.24 2.375 ;
      RECT 47.07 3.685 47.24 5.155 ;
      RECT 47.07 7.31 47.24 8.78 ;
      RECT 47.07 10.09 47.24 10.6 ;
      RECT 45.71 1.87 45.88 5.16 ;
      RECT 45.71 7.305 45.88 10.595 ;
      RECT 45.28 1.87 45.45 2.38 ;
      RECT 45.28 2.95 45.45 5.16 ;
      RECT 45.28 7.305 45.45 9.515 ;
      RECT 45.28 10.085 45.45 10.595 ;
      RECT 40.075 7.305 40.245 10.595 ;
      RECT 39.645 7.305 39.815 9.515 ;
      RECT 39.645 10.085 39.815 10.595 ;
      RECT 32.8 7.31 32.97 8.78 ;
      RECT 32.8 10.09 32.97 10.6 ;
      RECT 31.81 1.865 31.98 2.375 ;
      RECT 31.81 3.685 31.98 5.155 ;
      RECT 31.81 7.31 31.98 8.78 ;
      RECT 31.81 10.09 31.98 10.6 ;
      RECT 30.45 1.87 30.62 5.16 ;
      RECT 30.45 7.305 30.62 10.595 ;
      RECT 30.02 1.87 30.19 2.38 ;
      RECT 30.02 2.95 30.19 5.16 ;
      RECT 30.02 7.305 30.19 9.515 ;
      RECT 30.02 10.085 30.19 10.595 ;
      RECT 24.815 7.305 24.985 10.595 ;
      RECT 24.385 7.305 24.555 9.515 ;
      RECT 24.385 10.085 24.555 10.595 ;
      RECT 17.54 7.31 17.71 8.78 ;
      RECT 17.54 10.09 17.71 10.6 ;
      RECT 16.55 1.865 16.72 2.375 ;
      RECT 16.55 3.685 16.72 5.155 ;
      RECT 16.55 7.31 16.72 8.78 ;
      RECT 16.55 10.09 16.72 10.6 ;
      RECT 15.19 1.87 15.36 5.16 ;
      RECT 15.19 7.305 15.36 10.595 ;
      RECT 14.76 1.87 14.93 2.38 ;
      RECT 14.76 2.95 14.93 5.16 ;
      RECT 14.76 7.305 14.93 9.515 ;
      RECT 14.76 10.085 14.93 10.595 ;
      RECT 9.555 7.305 9.725 10.595 ;
      RECT 9.125 7.305 9.295 9.515 ;
      RECT 9.125 10.085 9.295 10.595 ;
      RECT 1.63 7.305 1.8 9.515 ;
      RECT 1.63 10.085 1.8 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r2 ;
  SIZE 79.105 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 17.515 1.865 17.685 2.375 ;
        RECT 17.515 3.685 17.685 5.155 ;
      LAYER met1 ;
        RECT 17.455 3.655 17.745 3.885 ;
        RECT 17.455 2.175 17.745 2.405 ;
        RECT 17.515 2.175 17.685 3.885 ;
      LAYER mcon ;
        RECT 17.515 3.685 17.685 3.855 ;
        RECT 17.515 2.205 17.685 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 32.775 1.865 32.945 2.375 ;
        RECT 32.775 3.685 32.945 5.155 ;
      LAYER met1 ;
        RECT 32.715 3.655 33.005 3.885 ;
        RECT 32.715 2.175 33.005 2.405 ;
        RECT 32.775 2.175 32.945 3.885 ;
      LAYER mcon ;
        RECT 32.775 3.685 32.945 3.855 ;
        RECT 32.775 2.205 32.945 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 48.035 1.865 48.205 2.375 ;
        RECT 48.035 3.685 48.205 5.155 ;
      LAYER met1 ;
        RECT 47.975 3.655 48.265 3.885 ;
        RECT 47.975 2.175 48.265 2.405 ;
        RECT 48.035 2.175 48.205 3.885 ;
      LAYER mcon ;
        RECT 48.035 3.685 48.205 3.855 ;
        RECT 48.035 2.205 48.205 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 63.295 1.865 63.465 2.375 ;
        RECT 63.295 3.685 63.465 5.155 ;
      LAYER met1 ;
        RECT 63.235 3.655 63.525 3.885 ;
        RECT 63.235 2.175 63.525 2.405 ;
        RECT 63.295 2.175 63.465 3.885 ;
      LAYER mcon ;
        RECT 63.295 3.685 63.465 3.855 ;
        RECT 63.295 2.205 63.465 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4706 ;
    PORT
      LAYER li1 ;
        RECT 78.555 1.865 78.725 2.375 ;
        RECT 78.555 3.685 78.725 5.155 ;
      LAYER met1 ;
        RECT 78.495 3.655 78.785 3.885 ;
        RECT 78.495 2.175 78.785 2.405 ;
        RECT 78.555 2.175 78.725 3.885 ;
      LAYER mcon ;
        RECT 78.555 3.685 78.725 3.855 ;
        RECT 78.555 2.205 78.725 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 13.285 4 13.625 4.35 ;
        RECT 13.28 8.15 13.62 8.5 ;
        RECT 13.36 4 13.535 8.5 ;
      LAYER li1 ;
        RECT 13.365 2.955 13.535 4.23 ;
        RECT 13.365 8.235 13.535 9.51 ;
        RECT 7.73 8.235 7.9 9.51 ;
      LAYER met1 ;
        RECT 13.285 4.06 13.765 4.23 ;
        RECT 13.285 4 13.625 4.35 ;
        RECT 7.67 8.235 13.765 8.405 ;
        RECT 13.28 8.15 13.62 8.5 ;
        RECT 7.67 8.205 7.96 8.435 ;
      LAYER via1 ;
        RECT 13.38 8.25 13.53 8.4 ;
        RECT 13.385 4.1 13.535 4.25 ;
      LAYER mcon ;
        RECT 7.73 8.235 7.9 8.405 ;
        RECT 13.365 8.235 13.535 8.405 ;
        RECT 13.365 4.06 13.535 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 28.545 4 28.885 4.35 ;
        RECT 28.54 8.15 28.88 8.5 ;
        RECT 28.62 4 28.795 8.5 ;
      LAYER li1 ;
        RECT 28.625 2.955 28.795 4.23 ;
        RECT 28.625 8.235 28.795 9.51 ;
        RECT 22.99 8.235 23.16 9.51 ;
      LAYER met1 ;
        RECT 28.545 4.06 29.025 4.23 ;
        RECT 28.545 4 28.885 4.35 ;
        RECT 22.93 8.235 29.025 8.405 ;
        RECT 28.54 8.15 28.88 8.5 ;
        RECT 22.93 8.205 23.22 8.435 ;
      LAYER via1 ;
        RECT 28.64 8.25 28.79 8.4 ;
        RECT 28.645 4.1 28.795 4.25 ;
      LAYER mcon ;
        RECT 22.99 8.235 23.16 8.405 ;
        RECT 28.625 8.235 28.795 8.405 ;
        RECT 28.625 4.06 28.795 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 43.805 4 44.145 4.35 ;
        RECT 43.8 8.15 44.14 8.5 ;
        RECT 43.88 4 44.055 8.5 ;
      LAYER li1 ;
        RECT 43.885 2.955 44.055 4.23 ;
        RECT 43.885 8.235 44.055 9.51 ;
        RECT 38.25 8.235 38.42 9.51 ;
      LAYER met1 ;
        RECT 43.805 4.06 44.285 4.23 ;
        RECT 43.805 4 44.145 4.35 ;
        RECT 38.19 8.235 44.285 8.405 ;
        RECT 43.8 8.15 44.14 8.5 ;
        RECT 38.19 8.205 38.48 8.435 ;
      LAYER via1 ;
        RECT 43.9 8.25 44.05 8.4 ;
        RECT 43.905 4.1 44.055 4.25 ;
      LAYER mcon ;
        RECT 38.25 8.235 38.42 8.405 ;
        RECT 43.885 8.235 44.055 8.405 ;
        RECT 43.885 4.06 44.055 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 59.065 4 59.405 4.35 ;
        RECT 59.06 8.15 59.4 8.5 ;
        RECT 59.14 4 59.315 8.5 ;
      LAYER li1 ;
        RECT 59.145 2.955 59.315 4.23 ;
        RECT 59.145 8.235 59.315 9.51 ;
        RECT 53.51 8.235 53.68 9.51 ;
      LAYER met1 ;
        RECT 59.065 4.06 59.545 4.23 ;
        RECT 59.065 4 59.405 4.35 ;
        RECT 53.45 8.235 59.545 8.405 ;
        RECT 59.06 8.15 59.4 8.5 ;
        RECT 53.45 8.205 53.74 8.435 ;
      LAYER via1 ;
        RECT 59.16 8.25 59.31 8.4 ;
        RECT 59.165 4.1 59.315 4.25 ;
      LAYER mcon ;
        RECT 53.51 8.235 53.68 8.405 ;
        RECT 59.145 8.235 59.315 8.405 ;
        RECT 59.145 4.06 59.315 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 74.325 4 74.665 4.35 ;
        RECT 74.32 8.15 74.66 8.5 ;
        RECT 74.4 4 74.575 8.5 ;
      LAYER li1 ;
        RECT 74.405 2.955 74.575 4.23 ;
        RECT 74.405 8.235 74.575 9.51 ;
        RECT 68.77 8.235 68.94 9.51 ;
      LAYER met1 ;
        RECT 74.325 4.06 74.805 4.23 ;
        RECT 74.325 4 74.665 4.35 ;
        RECT 68.71 8.235 74.805 8.405 ;
        RECT 74.32 8.15 74.66 8.5 ;
        RECT 68.71 8.205 69 8.435 ;
      LAYER via1 ;
        RECT 74.42 8.25 74.57 8.4 ;
        RECT 74.425 4.1 74.575 4.25 ;
      LAYER mcon ;
        RECT 68.77 8.235 68.94 8.405 ;
        RECT 74.405 8.235 74.575 8.405 ;
        RECT 74.405 4.06 74.575 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.235 8.235 0.405 9.51 ;
      LAYER met1 ;
        RECT 0.175 8.235 0.635 8.405 ;
        RECT 0.175 8.205 0.465 8.435 ;
      LAYER mcon ;
        RECT 0.235 8.235 0.405 8.405 ;
    END
  END start
  OBS
    LAYER met3 ;
      RECT 73.71 2.245 74.04 4.35 ;
      RECT 73.71 4.03 74.055 4.32 ;
      RECT 67.7 2.245 68.03 3.88 ;
      RECT 67.7 2.245 74.04 2.575 ;
      RECT 70.04 9.345 70.41 9.715 ;
      RECT 70.075 5.565 70.375 9.715 ;
      RECT 65.885 6.525 70.375 6.86 ;
      RECT 69.025 5.565 70.375 6.86 ;
      RECT 65.885 5.435 66.19 6.86 ;
      RECT 69.065 3.15 69.365 6.86 ;
      RECT 65.885 3.73 66.185 6.86 ;
      RECT 69.02 4.055 69.365 4.785 ;
      RECT 65.78 3.31 66.11 4.04 ;
      RECT 68.66 3.15 69.39 3.48 ;
      RECT 58.45 2.245 58.78 4.35 ;
      RECT 58.45 4.03 58.795 4.32 ;
      RECT 52.44 2.245 52.77 3.88 ;
      RECT 52.44 2.245 58.78 2.575 ;
      RECT 54.78 9.345 55.15 9.715 ;
      RECT 54.815 5.565 55.115 9.715 ;
      RECT 50.625 6.525 55.115 6.86 ;
      RECT 53.765 5.565 55.115 6.86 ;
      RECT 50.625 5.435 50.93 6.86 ;
      RECT 53.805 3.15 54.105 6.86 ;
      RECT 50.625 3.73 50.925 6.86 ;
      RECT 53.76 4.055 54.105 4.785 ;
      RECT 50.52 3.31 50.85 4.04 ;
      RECT 53.4 3.15 54.13 3.48 ;
      RECT 43.19 2.245 43.52 4.35 ;
      RECT 43.19 4.03 43.535 4.32 ;
      RECT 37.18 2.245 37.51 3.88 ;
      RECT 37.18 2.245 43.52 2.575 ;
      RECT 39.52 9.345 39.89 9.715 ;
      RECT 39.555 5.565 39.855 9.715 ;
      RECT 35.365 6.525 39.855 6.86 ;
      RECT 38.505 5.565 39.855 6.86 ;
      RECT 35.365 5.435 35.67 6.86 ;
      RECT 38.545 3.15 38.845 6.86 ;
      RECT 35.365 3.73 35.665 6.86 ;
      RECT 38.5 4.055 38.845 4.785 ;
      RECT 35.26 3.31 35.59 4.04 ;
      RECT 38.14 3.15 38.87 3.48 ;
      RECT 27.93 2.245 28.26 4.35 ;
      RECT 27.93 4.03 28.275 4.32 ;
      RECT 21.92 2.245 22.25 3.88 ;
      RECT 21.92 2.245 28.26 2.575 ;
      RECT 24.26 9.345 24.63 9.715 ;
      RECT 24.295 5.565 24.595 9.715 ;
      RECT 20.105 6.525 24.595 6.86 ;
      RECT 23.245 5.565 24.595 6.86 ;
      RECT 20.105 5.435 20.41 6.86 ;
      RECT 23.285 3.15 23.585 6.86 ;
      RECT 20.105 3.73 20.405 6.86 ;
      RECT 23.24 4.055 23.585 4.785 ;
      RECT 20 3.31 20.33 4.04 ;
      RECT 22.88 3.15 23.61 3.48 ;
      RECT 12.67 2.245 13 4.35 ;
      RECT 12.67 4.03 13.015 4.32 ;
      RECT 6.66 2.245 6.99 3.88 ;
      RECT 6.66 2.245 13 2.575 ;
      RECT 9 9.345 9.37 9.715 ;
      RECT 9.035 5.565 9.335 9.715 ;
      RECT 4.845 6.525 9.335 6.86 ;
      RECT 7.985 5.565 9.335 6.86 ;
      RECT 4.845 5.435 5.15 6.86 ;
      RECT 8.025 3.15 8.325 6.86 ;
      RECT 4.845 3.73 5.145 6.86 ;
      RECT 7.98 4.055 8.325 4.785 ;
      RECT 4.74 3.31 5.07 4.04 ;
      RECT 7.62 3.15 8.35 3.48 ;
      RECT 72.14 3.31 72.47 4.04 ;
      RECT 70.94 4.175 71.27 4.905 ;
      RECT 70.1 3.15 70.83 3.48 ;
      RECT 66.5 3.31 66.83 4.04 ;
      RECT 56.88 3.31 57.21 4.04 ;
      RECT 55.68 4.175 56.01 4.905 ;
      RECT 54.84 3.15 55.57 3.48 ;
      RECT 51.24 3.31 51.57 4.04 ;
      RECT 41.62 3.31 41.95 4.04 ;
      RECT 40.42 4.175 40.75 4.905 ;
      RECT 39.58 3.15 40.31 3.48 ;
      RECT 35.98 3.31 36.31 4.04 ;
      RECT 26.36 3.31 26.69 4.04 ;
      RECT 25.16 4.175 25.49 4.905 ;
      RECT 24.32 3.15 25.05 3.48 ;
      RECT 20.72 3.31 21.05 4.04 ;
      RECT 11.1 3.31 11.43 4.04 ;
      RECT 9.9 4.175 10.23 4.905 ;
      RECT 9.06 3.15 9.79 3.48 ;
      RECT 5.46 3.31 5.79 4.04 ;
    LAYER via2 ;
      RECT 73.81 4.075 74.01 4.275 ;
      RECT 72.205 3.775 72.405 3.975 ;
      RECT 71.005 4.335 71.205 4.535 ;
      RECT 70.165 3.215 70.365 3.415 ;
      RECT 70.125 9.43 70.325 9.63 ;
      RECT 69.085 4.12 69.285 4.32 ;
      RECT 68.725 3.215 68.925 3.415 ;
      RECT 67.765 3.215 67.965 3.415 ;
      RECT 66.565 3.775 66.765 3.975 ;
      RECT 65.845 3.775 66.045 3.975 ;
      RECT 58.55 4.075 58.75 4.275 ;
      RECT 56.945 3.775 57.145 3.975 ;
      RECT 55.745 4.335 55.945 4.535 ;
      RECT 54.905 3.215 55.105 3.415 ;
      RECT 54.865 9.43 55.065 9.63 ;
      RECT 53.825 4.12 54.025 4.32 ;
      RECT 53.465 3.215 53.665 3.415 ;
      RECT 52.505 3.215 52.705 3.415 ;
      RECT 51.305 3.775 51.505 3.975 ;
      RECT 50.585 3.775 50.785 3.975 ;
      RECT 43.29 4.075 43.49 4.275 ;
      RECT 41.685 3.775 41.885 3.975 ;
      RECT 40.485 4.335 40.685 4.535 ;
      RECT 39.645 3.215 39.845 3.415 ;
      RECT 39.605 9.43 39.805 9.63 ;
      RECT 38.565 4.12 38.765 4.32 ;
      RECT 38.205 3.215 38.405 3.415 ;
      RECT 37.245 3.215 37.445 3.415 ;
      RECT 36.045 3.775 36.245 3.975 ;
      RECT 35.325 3.775 35.525 3.975 ;
      RECT 28.03 4.075 28.23 4.275 ;
      RECT 26.425 3.775 26.625 3.975 ;
      RECT 25.225 4.335 25.425 4.535 ;
      RECT 24.385 3.215 24.585 3.415 ;
      RECT 24.345 9.43 24.545 9.63 ;
      RECT 23.305 4.12 23.505 4.32 ;
      RECT 22.945 3.215 23.145 3.415 ;
      RECT 21.985 3.215 22.185 3.415 ;
      RECT 20.785 3.775 20.985 3.975 ;
      RECT 20.065 3.775 20.265 3.975 ;
      RECT 12.77 4.075 12.97 4.275 ;
      RECT 11.165 3.775 11.365 3.975 ;
      RECT 9.965 4.335 10.165 4.535 ;
      RECT 9.125 3.215 9.325 3.415 ;
      RECT 9.085 9.43 9.285 9.63 ;
      RECT 8.045 4.12 8.245 4.32 ;
      RECT 7.685 3.215 7.885 3.415 ;
      RECT 6.725 3.215 6.925 3.415 ;
      RECT 5.525 3.775 5.725 3.975 ;
      RECT 4.805 3.775 5.005 3.975 ;
    LAYER met2 ;
      RECT 1.23 10.69 78.73 10.86 ;
      RECT 78.56 9.565 78.73 10.86 ;
      RECT 1.23 8.545 1.4 10.86 ;
      RECT 78.53 9.565 78.88 9.915 ;
      RECT 1.17 8.545 1.46 8.895 ;
      RECT 75.37 8.51 75.69 8.835 ;
      RECT 75.4 7.985 75.57 8.835 ;
      RECT 75.4 7.985 75.575 8.335 ;
      RECT 75.4 7.985 76.375 8.16 ;
      RECT 76.2 3.26 76.375 8.16 ;
      RECT 76.145 3.26 76.495 3.61 ;
      RECT 76.17 8.945 76.495 9.27 ;
      RECT 75.055 9.035 76.495 9.205 ;
      RECT 75.055 3.69 75.215 9.205 ;
      RECT 75.37 3.66 75.69 3.98 ;
      RECT 75.055 3.69 75.69 3.86 ;
      RECT 73.72 4 74.105 4.35 ;
      RECT 73.71 4.065 74.105 4.265 ;
      RECT 73.855 3.995 74.025 4.35 ;
      RECT 72.165 3.735 72.445 4.015 ;
      RECT 72.16 3.735 72.445 3.968 ;
      RECT 72.14 3.735 72.445 3.945 ;
      RECT 72.13 3.735 72.445 3.925 ;
      RECT 72.12 3.735 72.445 3.91 ;
      RECT 72.095 3.735 72.445 3.883 ;
      RECT 72.085 3.735 72.445 3.858 ;
      RECT 72.04 3.59 72.32 3.85 ;
      RECT 72.04 3.685 72.42 3.85 ;
      RECT 72.04 3.63 72.365 3.85 ;
      RECT 72.04 3.622 72.36 3.85 ;
      RECT 72.04 3.612 72.355 3.85 ;
      RECT 72.04 3.6 72.35 3.85 ;
      RECT 70.965 4.295 71.245 4.575 ;
      RECT 70.965 4.295 71.28 4.555 ;
      RECT 63.245 8.945 63.595 9.295 ;
      RECT 70.71 8.9 71.06 9.25 ;
      RECT 63.245 8.975 71.06 9.175 ;
      RECT 71 3.715 71.05 3.975 ;
      RECT 70.79 3.715 70.795 3.975 ;
      RECT 69.985 3.27 70.015 3.53 ;
      RECT 69.755 3.27 69.83 3.53 ;
      RECT 70.975 3.665 71 3.975 ;
      RECT 70.97 3.622 70.975 3.975 ;
      RECT 70.965 3.605 70.97 3.975 ;
      RECT 70.96 3.592 70.965 3.975 ;
      RECT 70.885 3.475 70.96 3.975 ;
      RECT 70.84 3.292 70.885 3.975 ;
      RECT 70.835 3.22 70.84 3.975 ;
      RECT 70.82 3.195 70.835 3.975 ;
      RECT 70.795 3.157 70.82 3.975 ;
      RECT 70.785 3.137 70.795 3.697 ;
      RECT 70.77 3.129 70.785 3.652 ;
      RECT 70.765 3.121 70.77 3.623 ;
      RECT 70.76 3.118 70.765 3.603 ;
      RECT 70.755 3.115 70.76 3.583 ;
      RECT 70.75 3.112 70.755 3.563 ;
      RECT 70.72 3.101 70.75 3.5 ;
      RECT 70.7 3.086 70.72 3.415 ;
      RECT 70.695 3.078 70.7 3.378 ;
      RECT 70.685 3.072 70.695 3.345 ;
      RECT 70.67 3.064 70.685 3.305 ;
      RECT 70.665 3.057 70.67 3.265 ;
      RECT 70.66 3.054 70.665 3.243 ;
      RECT 70.655 3.051 70.66 3.23 ;
      RECT 70.65 3.05 70.655 3.22 ;
      RECT 70.635 3.044 70.65 3.21 ;
      RECT 70.61 3.031 70.635 3.195 ;
      RECT 70.56 3.006 70.61 3.166 ;
      RECT 70.545 2.985 70.56 3.141 ;
      RECT 70.535 2.978 70.545 3.13 ;
      RECT 70.48 2.959 70.535 3.103 ;
      RECT 70.455 2.937 70.48 3.076 ;
      RECT 70.45 2.93 70.455 3.071 ;
      RECT 70.435 2.93 70.45 3.069 ;
      RECT 70.41 2.922 70.435 3.065 ;
      RECT 70.395 2.92 70.41 3.061 ;
      RECT 70.365 2.92 70.395 3.058 ;
      RECT 70.355 2.92 70.365 3.053 ;
      RECT 70.31 2.92 70.355 3.051 ;
      RECT 70.281 2.92 70.31 3.052 ;
      RECT 70.195 2.92 70.281 3.054 ;
      RECT 70.181 2.921 70.195 3.056 ;
      RECT 70.095 2.922 70.181 3.058 ;
      RECT 70.08 2.923 70.095 3.068 ;
      RECT 70.075 2.924 70.08 3.077 ;
      RECT 70.055 2.927 70.075 3.087 ;
      RECT 70.04 2.935 70.055 3.102 ;
      RECT 70.02 2.953 70.04 3.117 ;
      RECT 70.01 2.965 70.02 3.14 ;
      RECT 70 2.974 70.01 3.17 ;
      RECT 69.985 2.986 70 3.215 ;
      RECT 69.93 3.019 69.985 3.53 ;
      RECT 69.925 3.047 69.93 3.53 ;
      RECT 69.905 3.062 69.925 3.53 ;
      RECT 69.87 3.122 69.905 3.53 ;
      RECT 69.868 3.172 69.87 3.53 ;
      RECT 69.865 3.18 69.868 3.53 ;
      RECT 69.855 3.195 69.865 3.53 ;
      RECT 69.85 3.207 69.855 3.53 ;
      RECT 69.84 3.232 69.85 3.53 ;
      RECT 69.83 3.26 69.84 3.53 ;
      RECT 67.735 4.765 67.785 5.025 ;
      RECT 70.645 4.315 70.705 4.575 ;
      RECT 70.63 4.315 70.645 4.585 ;
      RECT 70.611 4.315 70.63 4.618 ;
      RECT 70.525 4.315 70.611 4.743 ;
      RECT 70.445 4.315 70.525 4.925 ;
      RECT 70.44 4.552 70.445 5.01 ;
      RECT 70.415 4.622 70.44 5.038 ;
      RECT 70.41 4.692 70.415 5.065 ;
      RECT 70.39 4.764 70.41 5.087 ;
      RECT 70.385 4.831 70.39 5.11 ;
      RECT 70.375 4.86 70.385 5.125 ;
      RECT 70.365 4.882 70.375 5.142 ;
      RECT 70.36 4.892 70.365 5.153 ;
      RECT 70.355 4.9 70.36 5.161 ;
      RECT 70.345 4.908 70.355 5.173 ;
      RECT 70.34 4.92 70.345 5.183 ;
      RECT 70.335 4.928 70.34 5.188 ;
      RECT 70.315 4.946 70.335 5.198 ;
      RECT 70.31 4.963 70.315 5.205 ;
      RECT 70.305 4.971 70.31 5.206 ;
      RECT 70.3 4.982 70.305 5.208 ;
      RECT 70.26 5.02 70.3 5.218 ;
      RECT 70.255 5.055 70.26 5.229 ;
      RECT 70.25 5.06 70.255 5.232 ;
      RECT 70.225 5.07 70.25 5.239 ;
      RECT 70.215 5.084 70.225 5.248 ;
      RECT 70.195 5.096 70.215 5.251 ;
      RECT 70.145 5.115 70.195 5.255 ;
      RECT 70.1 5.13 70.145 5.26 ;
      RECT 70.035 5.133 70.1 5.266 ;
      RECT 70.02 5.131 70.035 5.273 ;
      RECT 69.99 5.13 70.02 5.273 ;
      RECT 69.951 5.129 69.99 5.269 ;
      RECT 69.865 5.126 69.951 5.265 ;
      RECT 69.848 5.124 69.865 5.262 ;
      RECT 69.762 5.122 69.848 5.259 ;
      RECT 69.676 5.119 69.762 5.253 ;
      RECT 69.59 5.115 69.676 5.248 ;
      RECT 69.512 5.112 69.59 5.244 ;
      RECT 69.426 5.109 69.512 5.242 ;
      RECT 69.34 5.106 69.426 5.239 ;
      RECT 69.282 5.104 69.34 5.236 ;
      RECT 69.196 5.101 69.282 5.234 ;
      RECT 69.11 5.097 69.196 5.232 ;
      RECT 69.024 5.094 69.11 5.229 ;
      RECT 68.938 5.09 69.024 5.227 ;
      RECT 68.852 5.086 68.938 5.224 ;
      RECT 68.766 5.083 68.852 5.222 ;
      RECT 68.68 5.079 68.766 5.219 ;
      RECT 68.594 5.076 68.68 5.217 ;
      RECT 68.508 5.072 68.594 5.214 ;
      RECT 68.422 5.069 68.508 5.212 ;
      RECT 68.336 5.065 68.422 5.209 ;
      RECT 68.25 5.062 68.336 5.207 ;
      RECT 68.24 5.06 68.25 5.203 ;
      RECT 68.235 5.06 68.24 5.201 ;
      RECT 68.195 5.055 68.235 5.195 ;
      RECT 68.181 5.046 68.195 5.188 ;
      RECT 68.095 5.016 68.181 5.173 ;
      RECT 68.075 4.982 68.095 5.158 ;
      RECT 68.005 4.951 68.075 5.145 ;
      RECT 68 4.926 68.005 5.134 ;
      RECT 67.995 4.92 68 5.132 ;
      RECT 67.926 4.765 67.995 5.12 ;
      RECT 67.84 4.765 67.926 5.094 ;
      RECT 67.815 4.765 67.84 5.073 ;
      RECT 67.81 4.765 67.815 5.063 ;
      RECT 67.805 4.765 67.81 5.055 ;
      RECT 67.785 4.765 67.805 5.038 ;
      RECT 70.205 3.335 70.465 3.595 ;
      RECT 70.19 3.335 70.465 3.498 ;
      RECT 70.16 3.335 70.465 3.473 ;
      RECT 70.125 3.175 70.405 3.455 ;
      RECT 70.095 4.665 70.155 4.925 ;
      RECT 69.12 3.355 69.175 3.615 ;
      RECT 70.055 4.622 70.095 4.925 ;
      RECT 70.026 4.543 70.055 4.925 ;
      RECT 69.94 4.415 70.026 4.925 ;
      RECT 69.92 4.295 69.94 4.925 ;
      RECT 69.895 4.246 69.92 4.925 ;
      RECT 69.89 4.211 69.895 4.775 ;
      RECT 69.86 4.171 69.89 4.713 ;
      RECT 69.835 4.108 69.86 4.628 ;
      RECT 69.825 4.07 69.835 4.565 ;
      RECT 69.81 4.045 69.825 4.526 ;
      RECT 69.767 4.003 69.81 4.432 ;
      RECT 69.765 3.976 69.767 4.359 ;
      RECT 69.76 3.971 69.765 4.35 ;
      RECT 69.755 3.964 69.76 4.325 ;
      RECT 69.75 3.958 69.755 4.31 ;
      RECT 69.745 3.952 69.75 4.298 ;
      RECT 69.735 3.943 69.745 4.28 ;
      RECT 69.73 3.934 69.735 4.258 ;
      RECT 69.705 3.915 69.73 4.208 ;
      RECT 69.7 3.896 69.705 4.158 ;
      RECT 69.685 3.882 69.7 4.118 ;
      RECT 69.68 3.868 69.685 4.085 ;
      RECT 69.675 3.861 69.68 4.078 ;
      RECT 69.66 3.848 69.675 4.07 ;
      RECT 69.615 3.81 69.66 4.043 ;
      RECT 69.585 3.763 69.615 4.008 ;
      RECT 69.565 3.732 69.585 3.985 ;
      RECT 69.485 3.665 69.565 3.938 ;
      RECT 69.455 3.595 69.485 3.885 ;
      RECT 69.45 3.572 69.455 3.868 ;
      RECT 69.42 3.55 69.45 3.853 ;
      RECT 69.39 3.509 69.42 3.825 ;
      RECT 69.385 3.484 69.39 3.81 ;
      RECT 69.38 3.478 69.385 3.803 ;
      RECT 69.37 3.355 69.38 3.795 ;
      RECT 69.36 3.355 69.37 3.788 ;
      RECT 69.355 3.355 69.36 3.78 ;
      RECT 69.335 3.355 69.355 3.768 ;
      RECT 69.285 3.355 69.335 3.738 ;
      RECT 69.23 3.355 69.285 3.688 ;
      RECT 69.2 3.355 69.23 3.648 ;
      RECT 69.175 3.355 69.2 3.625 ;
      RECT 69.045 4.08 69.325 4.36 ;
      RECT 69.01 3.995 69.27 4.255 ;
      RECT 69.01 4.077 69.28 4.255 ;
      RECT 67.21 3.45 67.215 3.935 ;
      RECT 67.1 3.635 67.105 3.935 ;
      RECT 67.01 3.675 67.075 3.935 ;
      RECT 68.685 3.175 68.775 3.805 ;
      RECT 68.65 3.225 68.655 3.805 ;
      RECT 68.595 3.25 68.605 3.805 ;
      RECT 68.55 3.25 68.56 3.805 ;
      RECT 68.92 3.175 68.965 3.455 ;
      RECT 67.77 2.905 67.97 3.045 ;
      RECT 68.886 3.175 68.92 3.467 ;
      RECT 68.8 3.175 68.886 3.507 ;
      RECT 68.785 3.175 68.8 3.548 ;
      RECT 68.78 3.175 68.785 3.568 ;
      RECT 68.775 3.175 68.78 3.588 ;
      RECT 68.655 3.217 68.685 3.805 ;
      RECT 68.605 3.237 68.65 3.805 ;
      RECT 68.59 3.252 68.595 3.805 ;
      RECT 68.56 3.252 68.59 3.805 ;
      RECT 68.515 3.237 68.55 3.805 ;
      RECT 68.51 3.225 68.515 3.585 ;
      RECT 68.505 3.222 68.51 3.565 ;
      RECT 68.49 3.212 68.505 3.518 ;
      RECT 68.485 3.205 68.49 3.481 ;
      RECT 68.48 3.202 68.485 3.464 ;
      RECT 68.465 3.192 68.48 3.42 ;
      RECT 68.46 3.183 68.465 3.38 ;
      RECT 68.455 3.179 68.46 3.365 ;
      RECT 68.445 3.173 68.455 3.348 ;
      RECT 68.405 3.154 68.445 3.323 ;
      RECT 68.4 3.136 68.405 3.303 ;
      RECT 68.39 3.13 68.4 3.298 ;
      RECT 68.36 3.114 68.39 3.285 ;
      RECT 68.345 3.096 68.36 3.268 ;
      RECT 68.33 3.084 68.345 3.255 ;
      RECT 68.325 3.076 68.33 3.248 ;
      RECT 68.295 3.062 68.325 3.235 ;
      RECT 68.29 3.047 68.295 3.223 ;
      RECT 68.28 3.041 68.29 3.215 ;
      RECT 68.26 3.029 68.28 3.203 ;
      RECT 68.25 3.017 68.26 3.19 ;
      RECT 68.22 3.001 68.25 3.175 ;
      RECT 68.2 2.981 68.22 3.158 ;
      RECT 68.195 2.971 68.2 3.148 ;
      RECT 68.17 2.959 68.195 3.135 ;
      RECT 68.165 2.947 68.17 3.123 ;
      RECT 68.16 2.942 68.165 3.119 ;
      RECT 68.145 2.935 68.16 3.111 ;
      RECT 68.135 2.922 68.145 3.101 ;
      RECT 68.13 2.92 68.135 3.095 ;
      RECT 68.105 2.913 68.13 3.084 ;
      RECT 68.1 2.906 68.105 3.073 ;
      RECT 68.075 2.905 68.1 3.06 ;
      RECT 68.056 2.905 68.075 3.05 ;
      RECT 67.97 2.905 68.056 3.047 ;
      RECT 67.74 2.905 67.77 3.05 ;
      RECT 67.7 2.912 67.74 3.063 ;
      RECT 67.675 2.922 67.7 3.076 ;
      RECT 67.66 2.931 67.675 3.086 ;
      RECT 67.63 2.936 67.66 3.105 ;
      RECT 67.625 2.942 67.63 3.123 ;
      RECT 67.605 2.952 67.625 3.138 ;
      RECT 67.595 2.965 67.605 3.158 ;
      RECT 67.58 2.977 67.595 3.175 ;
      RECT 67.575 2.987 67.58 3.185 ;
      RECT 67.57 2.992 67.575 3.19 ;
      RECT 67.56 3 67.57 3.203 ;
      RECT 67.51 3.032 67.56 3.24 ;
      RECT 67.495 3.067 67.51 3.281 ;
      RECT 67.49 3.077 67.495 3.296 ;
      RECT 67.485 3.082 67.49 3.303 ;
      RECT 67.46 3.098 67.485 3.323 ;
      RECT 67.445 3.119 67.46 3.348 ;
      RECT 67.42 3.14 67.445 3.373 ;
      RECT 67.41 3.159 67.42 3.396 ;
      RECT 67.385 3.177 67.41 3.419 ;
      RECT 67.37 3.197 67.385 3.443 ;
      RECT 67.365 3.207 67.37 3.455 ;
      RECT 67.35 3.219 67.365 3.475 ;
      RECT 67.34 3.234 67.35 3.515 ;
      RECT 67.335 3.242 67.34 3.543 ;
      RECT 67.325 3.252 67.335 3.563 ;
      RECT 67.32 3.265 67.325 3.588 ;
      RECT 67.315 3.278 67.32 3.608 ;
      RECT 67.31 3.284 67.315 3.63 ;
      RECT 67.3 3.293 67.31 3.65 ;
      RECT 67.295 3.313 67.3 3.673 ;
      RECT 67.29 3.319 67.295 3.693 ;
      RECT 67.285 3.326 67.29 3.715 ;
      RECT 67.28 3.337 67.285 3.728 ;
      RECT 67.27 3.347 67.28 3.753 ;
      RECT 67.25 3.372 67.27 3.935 ;
      RECT 67.22 3.412 67.25 3.935 ;
      RECT 67.215 3.442 67.22 3.935 ;
      RECT 67.19 3.47 67.21 3.935 ;
      RECT 67.16 3.515 67.19 3.935 ;
      RECT 67.155 3.542 67.16 3.935 ;
      RECT 67.135 3.56 67.155 3.935 ;
      RECT 67.125 3.585 67.135 3.935 ;
      RECT 67.12 3.597 67.125 3.935 ;
      RECT 67.105 3.62 67.12 3.935 ;
      RECT 67.085 3.647 67.1 3.935 ;
      RECT 67.075 3.67 67.085 3.935 ;
      RECT 68.865 4.555 68.945 4.815 ;
      RECT 68.1 3.775 68.17 4.035 ;
      RECT 68.831 4.522 68.865 4.815 ;
      RECT 68.745 4.425 68.831 4.815 ;
      RECT 68.725 4.337 68.745 4.815 ;
      RECT 68.715 4.307 68.725 4.815 ;
      RECT 68.705 4.287 68.715 4.815 ;
      RECT 68.685 4.274 68.705 4.815 ;
      RECT 68.67 4.264 68.685 4.643 ;
      RECT 68.665 4.257 68.67 4.598 ;
      RECT 68.655 4.251 68.665 4.588 ;
      RECT 68.645 4.243 68.655 4.57 ;
      RECT 68.64 4.237 68.645 4.558 ;
      RECT 68.63 4.232 68.64 4.545 ;
      RECT 68.61 4.222 68.63 4.518 ;
      RECT 68.57 4.201 68.61 4.47 ;
      RECT 68.555 4.182 68.57 4.428 ;
      RECT 68.53 4.168 68.555 4.398 ;
      RECT 68.52 4.156 68.53 4.365 ;
      RECT 68.515 4.151 68.52 4.355 ;
      RECT 68.485 4.137 68.515 4.335 ;
      RECT 68.475 4.121 68.485 4.308 ;
      RECT 68.47 4.116 68.475 4.298 ;
      RECT 68.445 4.107 68.47 4.278 ;
      RECT 68.435 4.095 68.445 4.258 ;
      RECT 68.365 4.063 68.435 4.233 ;
      RECT 68.36 4.032 68.365 4.21 ;
      RECT 68.311 3.775 68.36 4.193 ;
      RECT 68.225 3.775 68.311 4.152 ;
      RECT 68.17 3.775 68.225 4.08 ;
      RECT 68.26 4.56 68.42 4.82 ;
      RECT 67.785 3.175 67.835 3.86 ;
      RECT 67.575 3.6 67.61 3.86 ;
      RECT 67.89 3.175 67.895 3.635 ;
      RECT 67.98 3.175 68.005 3.455 ;
      RECT 68.255 4.557 68.26 4.82 ;
      RECT 68.22 4.545 68.255 4.82 ;
      RECT 68.16 4.518 68.22 4.82 ;
      RECT 68.155 4.501 68.16 4.674 ;
      RECT 68.15 4.498 68.155 4.661 ;
      RECT 68.13 4.491 68.15 4.648 ;
      RECT 68.095 4.474 68.13 4.63 ;
      RECT 68.055 4.453 68.095 4.61 ;
      RECT 68.05 4.441 68.055 4.598 ;
      RECT 68.01 4.427 68.05 4.584 ;
      RECT 67.99 4.41 68.01 4.566 ;
      RECT 67.98 4.402 67.99 4.558 ;
      RECT 67.965 3.175 67.98 3.473 ;
      RECT 67.95 4.392 67.98 4.545 ;
      RECT 67.935 3.175 67.965 3.518 ;
      RECT 67.94 4.382 67.95 4.532 ;
      RECT 67.91 4.367 67.94 4.519 ;
      RECT 67.895 3.175 67.935 3.585 ;
      RECT 67.895 4.335 67.91 4.505 ;
      RECT 67.89 4.307 67.895 4.499 ;
      RECT 67.885 3.175 67.89 3.64 ;
      RECT 67.875 4.277 67.89 4.493 ;
      RECT 67.88 3.175 67.885 3.653 ;
      RECT 67.87 3.175 67.88 3.673 ;
      RECT 67.835 4.19 67.875 4.478 ;
      RECT 67.835 3.175 67.87 3.713 ;
      RECT 67.83 4.122 67.835 4.466 ;
      RECT 67.815 4.077 67.83 4.461 ;
      RECT 67.81 4.015 67.815 4.456 ;
      RECT 67.785 3.922 67.81 4.449 ;
      RECT 67.78 3.175 67.785 4.441 ;
      RECT 67.765 3.175 67.78 4.428 ;
      RECT 67.745 3.175 67.765 4.385 ;
      RECT 67.735 3.175 67.745 4.335 ;
      RECT 67.73 3.175 67.735 4.308 ;
      RECT 67.725 3.175 67.73 4.286 ;
      RECT 67.72 3.401 67.725 4.269 ;
      RECT 67.715 3.423 67.72 4.247 ;
      RECT 67.71 3.465 67.715 4.23 ;
      RECT 67.68 3.515 67.71 4.174 ;
      RECT 67.675 3.542 67.68 4.116 ;
      RECT 67.66 3.56 67.675 4.08 ;
      RECT 67.655 3.578 67.66 4.044 ;
      RECT 67.649 3.585 67.655 4.025 ;
      RECT 67.645 3.592 67.649 4.008 ;
      RECT 67.64 3.597 67.645 3.977 ;
      RECT 67.63 3.6 67.64 3.952 ;
      RECT 67.62 3.6 67.63 3.918 ;
      RECT 67.615 3.6 67.62 3.895 ;
      RECT 67.61 3.6 67.615 3.875 ;
      RECT 66.525 3.735 66.805 4.015 ;
      RECT 66.525 3.735 66.825 3.91 ;
      RECT 66.615 3.625 66.875 3.885 ;
      RECT 66.58 3.72 66.875 3.885 ;
      RECT 66.705 2.24 66.87 3.885 ;
      RECT 66.605 2.24 66.975 2.61 ;
      RECT 66.23 4.765 66.49 5.025 ;
      RECT 66.25 4.692 66.43 5.025 ;
      RECT 66.25 4.435 66.425 5.025 ;
      RECT 66.25 4.227 66.415 5.025 ;
      RECT 66.255 4.145 66.415 5.025 ;
      RECT 66.255 3.91 66.405 5.025 ;
      RECT 66.255 3.757 66.4 5.025 ;
      RECT 66.26 3.742 66.4 5.025 ;
      RECT 66.31 3.457 66.4 5.025 ;
      RECT 66.265 3.692 66.4 5.025 ;
      RECT 66.295 3.51 66.4 5.025 ;
      RECT 66.28 3.622 66.4 5.025 ;
      RECT 66.285 3.58 66.4 5.025 ;
      RECT 66.28 3.622 66.415 3.685 ;
      RECT 66.315 3.21 66.42 3.63 ;
      RECT 66.315 3.21 66.435 3.613 ;
      RECT 66.315 3.21 66.47 3.575 ;
      RECT 66.31 3.457 66.52 3.508 ;
      RECT 66.315 3.21 66.575 3.47 ;
      RECT 65.575 3.915 65.835 4.175 ;
      RECT 65.575 3.915 65.845 4.133 ;
      RECT 65.575 3.915 65.931 4.104 ;
      RECT 65.575 3.915 66 4.056 ;
      RECT 65.575 3.915 66.035 4.025 ;
      RECT 65.805 3.735 66.085 4.015 ;
      RECT 65.64 3.9 66.085 4.015 ;
      RECT 65.73 3.777 65.835 4.175 ;
      RECT 65.66 3.84 66.085 4.015 ;
      RECT 60.11 8.51 60.43 8.835 ;
      RECT 60.14 7.985 60.31 8.835 ;
      RECT 60.14 7.985 60.315 8.335 ;
      RECT 60.14 7.985 61.115 8.16 ;
      RECT 60.94 3.26 61.115 8.16 ;
      RECT 60.885 3.26 61.235 3.61 ;
      RECT 60.91 8.945 61.235 9.27 ;
      RECT 59.795 9.035 61.235 9.205 ;
      RECT 59.795 3.69 59.955 9.205 ;
      RECT 60.11 3.66 60.43 3.98 ;
      RECT 59.795 3.69 60.43 3.86 ;
      RECT 58.46 4 58.845 4.35 ;
      RECT 58.45 4.065 58.845 4.265 ;
      RECT 58.595 3.995 58.765 4.35 ;
      RECT 56.905 3.735 57.185 4.015 ;
      RECT 56.9 3.735 57.185 3.968 ;
      RECT 56.88 3.735 57.185 3.945 ;
      RECT 56.87 3.735 57.185 3.925 ;
      RECT 56.86 3.735 57.185 3.91 ;
      RECT 56.835 3.735 57.185 3.883 ;
      RECT 56.825 3.735 57.185 3.858 ;
      RECT 56.78 3.59 57.06 3.85 ;
      RECT 56.78 3.685 57.16 3.85 ;
      RECT 56.78 3.63 57.105 3.85 ;
      RECT 56.78 3.622 57.1 3.85 ;
      RECT 56.78 3.612 57.095 3.85 ;
      RECT 56.78 3.6 57.09 3.85 ;
      RECT 55.705 4.295 55.985 4.575 ;
      RECT 55.705 4.295 56.02 4.555 ;
      RECT 47.985 8.945 48.335 9.295 ;
      RECT 55.45 8.9 55.8 9.25 ;
      RECT 47.985 8.975 55.8 9.175 ;
      RECT 55.74 3.715 55.79 3.975 ;
      RECT 55.53 3.715 55.535 3.975 ;
      RECT 54.725 3.27 54.755 3.53 ;
      RECT 54.495 3.27 54.57 3.53 ;
      RECT 55.715 3.665 55.74 3.975 ;
      RECT 55.71 3.622 55.715 3.975 ;
      RECT 55.705 3.605 55.71 3.975 ;
      RECT 55.7 3.592 55.705 3.975 ;
      RECT 55.625 3.475 55.7 3.975 ;
      RECT 55.58 3.292 55.625 3.975 ;
      RECT 55.575 3.22 55.58 3.975 ;
      RECT 55.56 3.195 55.575 3.975 ;
      RECT 55.535 3.157 55.56 3.975 ;
      RECT 55.525 3.137 55.535 3.697 ;
      RECT 55.51 3.129 55.525 3.652 ;
      RECT 55.505 3.121 55.51 3.623 ;
      RECT 55.5 3.118 55.505 3.603 ;
      RECT 55.495 3.115 55.5 3.583 ;
      RECT 55.49 3.112 55.495 3.563 ;
      RECT 55.46 3.101 55.49 3.5 ;
      RECT 55.44 3.086 55.46 3.415 ;
      RECT 55.435 3.078 55.44 3.378 ;
      RECT 55.425 3.072 55.435 3.345 ;
      RECT 55.41 3.064 55.425 3.305 ;
      RECT 55.405 3.057 55.41 3.265 ;
      RECT 55.4 3.054 55.405 3.243 ;
      RECT 55.395 3.051 55.4 3.23 ;
      RECT 55.39 3.05 55.395 3.22 ;
      RECT 55.375 3.044 55.39 3.21 ;
      RECT 55.35 3.031 55.375 3.195 ;
      RECT 55.3 3.006 55.35 3.166 ;
      RECT 55.285 2.985 55.3 3.141 ;
      RECT 55.275 2.978 55.285 3.13 ;
      RECT 55.22 2.959 55.275 3.103 ;
      RECT 55.195 2.937 55.22 3.076 ;
      RECT 55.19 2.93 55.195 3.071 ;
      RECT 55.175 2.93 55.19 3.069 ;
      RECT 55.15 2.922 55.175 3.065 ;
      RECT 55.135 2.92 55.15 3.061 ;
      RECT 55.105 2.92 55.135 3.058 ;
      RECT 55.095 2.92 55.105 3.053 ;
      RECT 55.05 2.92 55.095 3.051 ;
      RECT 55.021 2.92 55.05 3.052 ;
      RECT 54.935 2.92 55.021 3.054 ;
      RECT 54.921 2.921 54.935 3.056 ;
      RECT 54.835 2.922 54.921 3.058 ;
      RECT 54.82 2.923 54.835 3.068 ;
      RECT 54.815 2.924 54.82 3.077 ;
      RECT 54.795 2.927 54.815 3.087 ;
      RECT 54.78 2.935 54.795 3.102 ;
      RECT 54.76 2.953 54.78 3.117 ;
      RECT 54.75 2.965 54.76 3.14 ;
      RECT 54.74 2.974 54.75 3.17 ;
      RECT 54.725 2.986 54.74 3.215 ;
      RECT 54.67 3.019 54.725 3.53 ;
      RECT 54.665 3.047 54.67 3.53 ;
      RECT 54.645 3.062 54.665 3.53 ;
      RECT 54.61 3.122 54.645 3.53 ;
      RECT 54.608 3.172 54.61 3.53 ;
      RECT 54.605 3.18 54.608 3.53 ;
      RECT 54.595 3.195 54.605 3.53 ;
      RECT 54.59 3.207 54.595 3.53 ;
      RECT 54.58 3.232 54.59 3.53 ;
      RECT 54.57 3.26 54.58 3.53 ;
      RECT 52.475 4.765 52.525 5.025 ;
      RECT 55.385 4.315 55.445 4.575 ;
      RECT 55.37 4.315 55.385 4.585 ;
      RECT 55.351 4.315 55.37 4.618 ;
      RECT 55.265 4.315 55.351 4.743 ;
      RECT 55.185 4.315 55.265 4.925 ;
      RECT 55.18 4.552 55.185 5.01 ;
      RECT 55.155 4.622 55.18 5.038 ;
      RECT 55.15 4.692 55.155 5.065 ;
      RECT 55.13 4.764 55.15 5.087 ;
      RECT 55.125 4.831 55.13 5.11 ;
      RECT 55.115 4.86 55.125 5.125 ;
      RECT 55.105 4.882 55.115 5.142 ;
      RECT 55.1 4.892 55.105 5.153 ;
      RECT 55.095 4.9 55.1 5.161 ;
      RECT 55.085 4.908 55.095 5.173 ;
      RECT 55.08 4.92 55.085 5.183 ;
      RECT 55.075 4.928 55.08 5.188 ;
      RECT 55.055 4.946 55.075 5.198 ;
      RECT 55.05 4.963 55.055 5.205 ;
      RECT 55.045 4.971 55.05 5.206 ;
      RECT 55.04 4.982 55.045 5.208 ;
      RECT 55 5.02 55.04 5.218 ;
      RECT 54.995 5.055 55 5.229 ;
      RECT 54.99 5.06 54.995 5.232 ;
      RECT 54.965 5.07 54.99 5.239 ;
      RECT 54.955 5.084 54.965 5.248 ;
      RECT 54.935 5.096 54.955 5.251 ;
      RECT 54.885 5.115 54.935 5.255 ;
      RECT 54.84 5.13 54.885 5.26 ;
      RECT 54.775 5.133 54.84 5.266 ;
      RECT 54.76 5.131 54.775 5.273 ;
      RECT 54.73 5.13 54.76 5.273 ;
      RECT 54.691 5.129 54.73 5.269 ;
      RECT 54.605 5.126 54.691 5.265 ;
      RECT 54.588 5.124 54.605 5.262 ;
      RECT 54.502 5.122 54.588 5.259 ;
      RECT 54.416 5.119 54.502 5.253 ;
      RECT 54.33 5.115 54.416 5.248 ;
      RECT 54.252 5.112 54.33 5.244 ;
      RECT 54.166 5.109 54.252 5.242 ;
      RECT 54.08 5.106 54.166 5.239 ;
      RECT 54.022 5.104 54.08 5.236 ;
      RECT 53.936 5.101 54.022 5.234 ;
      RECT 53.85 5.097 53.936 5.232 ;
      RECT 53.764 5.094 53.85 5.229 ;
      RECT 53.678 5.09 53.764 5.227 ;
      RECT 53.592 5.086 53.678 5.224 ;
      RECT 53.506 5.083 53.592 5.222 ;
      RECT 53.42 5.079 53.506 5.219 ;
      RECT 53.334 5.076 53.42 5.217 ;
      RECT 53.248 5.072 53.334 5.214 ;
      RECT 53.162 5.069 53.248 5.212 ;
      RECT 53.076 5.065 53.162 5.209 ;
      RECT 52.99 5.062 53.076 5.207 ;
      RECT 52.98 5.06 52.99 5.203 ;
      RECT 52.975 5.06 52.98 5.201 ;
      RECT 52.935 5.055 52.975 5.195 ;
      RECT 52.921 5.046 52.935 5.188 ;
      RECT 52.835 5.016 52.921 5.173 ;
      RECT 52.815 4.982 52.835 5.158 ;
      RECT 52.745 4.951 52.815 5.145 ;
      RECT 52.74 4.926 52.745 5.134 ;
      RECT 52.735 4.92 52.74 5.132 ;
      RECT 52.666 4.765 52.735 5.12 ;
      RECT 52.58 4.765 52.666 5.094 ;
      RECT 52.555 4.765 52.58 5.073 ;
      RECT 52.55 4.765 52.555 5.063 ;
      RECT 52.545 4.765 52.55 5.055 ;
      RECT 52.525 4.765 52.545 5.038 ;
      RECT 54.945 3.335 55.205 3.595 ;
      RECT 54.93 3.335 55.205 3.498 ;
      RECT 54.9 3.335 55.205 3.473 ;
      RECT 54.865 3.175 55.145 3.455 ;
      RECT 54.835 4.665 54.895 4.925 ;
      RECT 53.86 3.355 53.915 3.615 ;
      RECT 54.795 4.622 54.835 4.925 ;
      RECT 54.766 4.543 54.795 4.925 ;
      RECT 54.68 4.415 54.766 4.925 ;
      RECT 54.66 4.295 54.68 4.925 ;
      RECT 54.635 4.246 54.66 4.925 ;
      RECT 54.63 4.211 54.635 4.775 ;
      RECT 54.6 4.171 54.63 4.713 ;
      RECT 54.575 4.108 54.6 4.628 ;
      RECT 54.565 4.07 54.575 4.565 ;
      RECT 54.55 4.045 54.565 4.526 ;
      RECT 54.507 4.003 54.55 4.432 ;
      RECT 54.505 3.976 54.507 4.359 ;
      RECT 54.5 3.971 54.505 4.35 ;
      RECT 54.495 3.964 54.5 4.325 ;
      RECT 54.49 3.958 54.495 4.31 ;
      RECT 54.485 3.952 54.49 4.298 ;
      RECT 54.475 3.943 54.485 4.28 ;
      RECT 54.47 3.934 54.475 4.258 ;
      RECT 54.445 3.915 54.47 4.208 ;
      RECT 54.44 3.896 54.445 4.158 ;
      RECT 54.425 3.882 54.44 4.118 ;
      RECT 54.42 3.868 54.425 4.085 ;
      RECT 54.415 3.861 54.42 4.078 ;
      RECT 54.4 3.848 54.415 4.07 ;
      RECT 54.355 3.81 54.4 4.043 ;
      RECT 54.325 3.763 54.355 4.008 ;
      RECT 54.305 3.732 54.325 3.985 ;
      RECT 54.225 3.665 54.305 3.938 ;
      RECT 54.195 3.595 54.225 3.885 ;
      RECT 54.19 3.572 54.195 3.868 ;
      RECT 54.16 3.55 54.19 3.853 ;
      RECT 54.13 3.509 54.16 3.825 ;
      RECT 54.125 3.484 54.13 3.81 ;
      RECT 54.12 3.478 54.125 3.803 ;
      RECT 54.11 3.355 54.12 3.795 ;
      RECT 54.1 3.355 54.11 3.788 ;
      RECT 54.095 3.355 54.1 3.78 ;
      RECT 54.075 3.355 54.095 3.768 ;
      RECT 54.025 3.355 54.075 3.738 ;
      RECT 53.97 3.355 54.025 3.688 ;
      RECT 53.94 3.355 53.97 3.648 ;
      RECT 53.915 3.355 53.94 3.625 ;
      RECT 53.785 4.08 54.065 4.36 ;
      RECT 53.75 3.995 54.01 4.255 ;
      RECT 53.75 4.077 54.02 4.255 ;
      RECT 51.95 3.45 51.955 3.935 ;
      RECT 51.84 3.635 51.845 3.935 ;
      RECT 51.75 3.675 51.815 3.935 ;
      RECT 53.425 3.175 53.515 3.805 ;
      RECT 53.39 3.225 53.395 3.805 ;
      RECT 53.335 3.25 53.345 3.805 ;
      RECT 53.29 3.25 53.3 3.805 ;
      RECT 53.66 3.175 53.705 3.455 ;
      RECT 52.51 2.905 52.71 3.045 ;
      RECT 53.626 3.175 53.66 3.467 ;
      RECT 53.54 3.175 53.626 3.507 ;
      RECT 53.525 3.175 53.54 3.548 ;
      RECT 53.52 3.175 53.525 3.568 ;
      RECT 53.515 3.175 53.52 3.588 ;
      RECT 53.395 3.217 53.425 3.805 ;
      RECT 53.345 3.237 53.39 3.805 ;
      RECT 53.33 3.252 53.335 3.805 ;
      RECT 53.3 3.252 53.33 3.805 ;
      RECT 53.255 3.237 53.29 3.805 ;
      RECT 53.25 3.225 53.255 3.585 ;
      RECT 53.245 3.222 53.25 3.565 ;
      RECT 53.23 3.212 53.245 3.518 ;
      RECT 53.225 3.205 53.23 3.481 ;
      RECT 53.22 3.202 53.225 3.464 ;
      RECT 53.205 3.192 53.22 3.42 ;
      RECT 53.2 3.183 53.205 3.38 ;
      RECT 53.195 3.179 53.2 3.365 ;
      RECT 53.185 3.173 53.195 3.348 ;
      RECT 53.145 3.154 53.185 3.323 ;
      RECT 53.14 3.136 53.145 3.303 ;
      RECT 53.13 3.13 53.14 3.298 ;
      RECT 53.1 3.114 53.13 3.285 ;
      RECT 53.085 3.096 53.1 3.268 ;
      RECT 53.07 3.084 53.085 3.255 ;
      RECT 53.065 3.076 53.07 3.248 ;
      RECT 53.035 3.062 53.065 3.235 ;
      RECT 53.03 3.047 53.035 3.223 ;
      RECT 53.02 3.041 53.03 3.215 ;
      RECT 53 3.029 53.02 3.203 ;
      RECT 52.99 3.017 53 3.19 ;
      RECT 52.96 3.001 52.99 3.175 ;
      RECT 52.94 2.981 52.96 3.158 ;
      RECT 52.935 2.971 52.94 3.148 ;
      RECT 52.91 2.959 52.935 3.135 ;
      RECT 52.905 2.947 52.91 3.123 ;
      RECT 52.9 2.942 52.905 3.119 ;
      RECT 52.885 2.935 52.9 3.111 ;
      RECT 52.875 2.922 52.885 3.101 ;
      RECT 52.87 2.92 52.875 3.095 ;
      RECT 52.845 2.913 52.87 3.084 ;
      RECT 52.84 2.906 52.845 3.073 ;
      RECT 52.815 2.905 52.84 3.06 ;
      RECT 52.796 2.905 52.815 3.05 ;
      RECT 52.71 2.905 52.796 3.047 ;
      RECT 52.48 2.905 52.51 3.05 ;
      RECT 52.44 2.912 52.48 3.063 ;
      RECT 52.415 2.922 52.44 3.076 ;
      RECT 52.4 2.931 52.415 3.086 ;
      RECT 52.37 2.936 52.4 3.105 ;
      RECT 52.365 2.942 52.37 3.123 ;
      RECT 52.345 2.952 52.365 3.138 ;
      RECT 52.335 2.965 52.345 3.158 ;
      RECT 52.32 2.977 52.335 3.175 ;
      RECT 52.315 2.987 52.32 3.185 ;
      RECT 52.31 2.992 52.315 3.19 ;
      RECT 52.3 3 52.31 3.203 ;
      RECT 52.25 3.032 52.3 3.24 ;
      RECT 52.235 3.067 52.25 3.281 ;
      RECT 52.23 3.077 52.235 3.296 ;
      RECT 52.225 3.082 52.23 3.303 ;
      RECT 52.2 3.098 52.225 3.323 ;
      RECT 52.185 3.119 52.2 3.348 ;
      RECT 52.16 3.14 52.185 3.373 ;
      RECT 52.15 3.159 52.16 3.396 ;
      RECT 52.125 3.177 52.15 3.419 ;
      RECT 52.11 3.197 52.125 3.443 ;
      RECT 52.105 3.207 52.11 3.455 ;
      RECT 52.09 3.219 52.105 3.475 ;
      RECT 52.08 3.234 52.09 3.515 ;
      RECT 52.075 3.242 52.08 3.543 ;
      RECT 52.065 3.252 52.075 3.563 ;
      RECT 52.06 3.265 52.065 3.588 ;
      RECT 52.055 3.278 52.06 3.608 ;
      RECT 52.05 3.284 52.055 3.63 ;
      RECT 52.04 3.293 52.05 3.65 ;
      RECT 52.035 3.313 52.04 3.673 ;
      RECT 52.03 3.319 52.035 3.693 ;
      RECT 52.025 3.326 52.03 3.715 ;
      RECT 52.02 3.337 52.025 3.728 ;
      RECT 52.01 3.347 52.02 3.753 ;
      RECT 51.99 3.372 52.01 3.935 ;
      RECT 51.96 3.412 51.99 3.935 ;
      RECT 51.955 3.442 51.96 3.935 ;
      RECT 51.93 3.47 51.95 3.935 ;
      RECT 51.9 3.515 51.93 3.935 ;
      RECT 51.895 3.542 51.9 3.935 ;
      RECT 51.875 3.56 51.895 3.935 ;
      RECT 51.865 3.585 51.875 3.935 ;
      RECT 51.86 3.597 51.865 3.935 ;
      RECT 51.845 3.62 51.86 3.935 ;
      RECT 51.825 3.647 51.84 3.935 ;
      RECT 51.815 3.67 51.825 3.935 ;
      RECT 53.605 4.555 53.685 4.815 ;
      RECT 52.84 3.775 52.91 4.035 ;
      RECT 53.571 4.522 53.605 4.815 ;
      RECT 53.485 4.425 53.571 4.815 ;
      RECT 53.465 4.337 53.485 4.815 ;
      RECT 53.455 4.307 53.465 4.815 ;
      RECT 53.445 4.287 53.455 4.815 ;
      RECT 53.425 4.274 53.445 4.815 ;
      RECT 53.41 4.264 53.425 4.643 ;
      RECT 53.405 4.257 53.41 4.598 ;
      RECT 53.395 4.251 53.405 4.588 ;
      RECT 53.385 4.243 53.395 4.57 ;
      RECT 53.38 4.237 53.385 4.558 ;
      RECT 53.37 4.232 53.38 4.545 ;
      RECT 53.35 4.222 53.37 4.518 ;
      RECT 53.31 4.201 53.35 4.47 ;
      RECT 53.295 4.182 53.31 4.428 ;
      RECT 53.27 4.168 53.295 4.398 ;
      RECT 53.26 4.156 53.27 4.365 ;
      RECT 53.255 4.151 53.26 4.355 ;
      RECT 53.225 4.137 53.255 4.335 ;
      RECT 53.215 4.121 53.225 4.308 ;
      RECT 53.21 4.116 53.215 4.298 ;
      RECT 53.185 4.107 53.21 4.278 ;
      RECT 53.175 4.095 53.185 4.258 ;
      RECT 53.105 4.063 53.175 4.233 ;
      RECT 53.1 4.032 53.105 4.21 ;
      RECT 53.051 3.775 53.1 4.193 ;
      RECT 52.965 3.775 53.051 4.152 ;
      RECT 52.91 3.775 52.965 4.08 ;
      RECT 53 4.56 53.16 4.82 ;
      RECT 52.525 3.175 52.575 3.86 ;
      RECT 52.315 3.6 52.35 3.86 ;
      RECT 52.63 3.175 52.635 3.635 ;
      RECT 52.72 3.175 52.745 3.455 ;
      RECT 52.995 4.557 53 4.82 ;
      RECT 52.96 4.545 52.995 4.82 ;
      RECT 52.9 4.518 52.96 4.82 ;
      RECT 52.895 4.501 52.9 4.674 ;
      RECT 52.89 4.498 52.895 4.661 ;
      RECT 52.87 4.491 52.89 4.648 ;
      RECT 52.835 4.474 52.87 4.63 ;
      RECT 52.795 4.453 52.835 4.61 ;
      RECT 52.79 4.441 52.795 4.598 ;
      RECT 52.75 4.427 52.79 4.584 ;
      RECT 52.73 4.41 52.75 4.566 ;
      RECT 52.72 4.402 52.73 4.558 ;
      RECT 52.705 3.175 52.72 3.473 ;
      RECT 52.69 4.392 52.72 4.545 ;
      RECT 52.675 3.175 52.705 3.518 ;
      RECT 52.68 4.382 52.69 4.532 ;
      RECT 52.65 4.367 52.68 4.519 ;
      RECT 52.635 3.175 52.675 3.585 ;
      RECT 52.635 4.335 52.65 4.505 ;
      RECT 52.63 4.307 52.635 4.499 ;
      RECT 52.625 3.175 52.63 3.64 ;
      RECT 52.615 4.277 52.63 4.493 ;
      RECT 52.62 3.175 52.625 3.653 ;
      RECT 52.61 3.175 52.62 3.673 ;
      RECT 52.575 4.19 52.615 4.478 ;
      RECT 52.575 3.175 52.61 3.713 ;
      RECT 52.57 4.122 52.575 4.466 ;
      RECT 52.555 4.077 52.57 4.461 ;
      RECT 52.55 4.015 52.555 4.456 ;
      RECT 52.525 3.922 52.55 4.449 ;
      RECT 52.52 3.175 52.525 4.441 ;
      RECT 52.505 3.175 52.52 4.428 ;
      RECT 52.485 3.175 52.505 4.385 ;
      RECT 52.475 3.175 52.485 4.335 ;
      RECT 52.47 3.175 52.475 4.308 ;
      RECT 52.465 3.175 52.47 4.286 ;
      RECT 52.46 3.401 52.465 4.269 ;
      RECT 52.455 3.423 52.46 4.247 ;
      RECT 52.45 3.465 52.455 4.23 ;
      RECT 52.42 3.515 52.45 4.174 ;
      RECT 52.415 3.542 52.42 4.116 ;
      RECT 52.4 3.56 52.415 4.08 ;
      RECT 52.395 3.578 52.4 4.044 ;
      RECT 52.389 3.585 52.395 4.025 ;
      RECT 52.385 3.592 52.389 4.008 ;
      RECT 52.38 3.597 52.385 3.977 ;
      RECT 52.37 3.6 52.38 3.952 ;
      RECT 52.36 3.6 52.37 3.918 ;
      RECT 52.355 3.6 52.36 3.895 ;
      RECT 52.35 3.6 52.355 3.875 ;
      RECT 51.265 3.735 51.545 4.015 ;
      RECT 51.265 3.735 51.565 3.91 ;
      RECT 51.355 3.625 51.615 3.885 ;
      RECT 51.32 3.72 51.615 3.885 ;
      RECT 51.445 2.24 51.61 3.885 ;
      RECT 51.345 2.24 51.715 2.61 ;
      RECT 50.97 4.765 51.23 5.025 ;
      RECT 50.99 4.692 51.17 5.025 ;
      RECT 50.99 4.435 51.165 5.025 ;
      RECT 50.99 4.227 51.155 5.025 ;
      RECT 50.995 4.145 51.155 5.025 ;
      RECT 50.995 3.91 51.145 5.025 ;
      RECT 50.995 3.757 51.14 5.025 ;
      RECT 51 3.742 51.14 5.025 ;
      RECT 51.05 3.457 51.14 5.025 ;
      RECT 51.005 3.692 51.14 5.025 ;
      RECT 51.035 3.51 51.14 5.025 ;
      RECT 51.02 3.622 51.14 5.025 ;
      RECT 51.025 3.58 51.14 5.025 ;
      RECT 51.02 3.622 51.155 3.685 ;
      RECT 51.055 3.21 51.16 3.63 ;
      RECT 51.055 3.21 51.175 3.613 ;
      RECT 51.055 3.21 51.21 3.575 ;
      RECT 51.05 3.457 51.26 3.508 ;
      RECT 51.055 3.21 51.315 3.47 ;
      RECT 50.315 3.915 50.575 4.175 ;
      RECT 50.315 3.915 50.585 4.133 ;
      RECT 50.315 3.915 50.671 4.104 ;
      RECT 50.315 3.915 50.74 4.056 ;
      RECT 50.315 3.915 50.775 4.025 ;
      RECT 50.545 3.735 50.825 4.015 ;
      RECT 50.38 3.9 50.825 4.015 ;
      RECT 50.47 3.777 50.575 4.175 ;
      RECT 50.4 3.84 50.825 4.015 ;
      RECT 44.85 8.51 45.17 8.835 ;
      RECT 44.88 7.985 45.05 8.835 ;
      RECT 44.88 7.985 45.055 8.335 ;
      RECT 44.88 7.985 45.855 8.16 ;
      RECT 45.68 3.26 45.855 8.16 ;
      RECT 45.625 3.26 45.975 3.61 ;
      RECT 45.65 8.945 45.975 9.27 ;
      RECT 44.535 9.035 45.975 9.205 ;
      RECT 44.535 3.69 44.695 9.205 ;
      RECT 44.85 3.66 45.17 3.98 ;
      RECT 44.535 3.69 45.17 3.86 ;
      RECT 43.2 4 43.585 4.35 ;
      RECT 43.19 4.065 43.585 4.265 ;
      RECT 43.335 3.995 43.505 4.35 ;
      RECT 41.645 3.735 41.925 4.015 ;
      RECT 41.64 3.735 41.925 3.968 ;
      RECT 41.62 3.735 41.925 3.945 ;
      RECT 41.61 3.735 41.925 3.925 ;
      RECT 41.6 3.735 41.925 3.91 ;
      RECT 41.575 3.735 41.925 3.883 ;
      RECT 41.565 3.735 41.925 3.858 ;
      RECT 41.52 3.59 41.8 3.85 ;
      RECT 41.52 3.685 41.9 3.85 ;
      RECT 41.52 3.63 41.845 3.85 ;
      RECT 41.52 3.622 41.84 3.85 ;
      RECT 41.52 3.612 41.835 3.85 ;
      RECT 41.52 3.6 41.83 3.85 ;
      RECT 40.445 4.295 40.725 4.575 ;
      RECT 40.445 4.295 40.76 4.555 ;
      RECT 32.77 8.95 33.12 9.3 ;
      RECT 40.19 8.905 40.54 9.255 ;
      RECT 32.77 8.98 40.54 9.18 ;
      RECT 40.48 3.715 40.53 3.975 ;
      RECT 40.27 3.715 40.275 3.975 ;
      RECT 39.465 3.27 39.495 3.53 ;
      RECT 39.235 3.27 39.31 3.53 ;
      RECT 40.455 3.665 40.48 3.975 ;
      RECT 40.45 3.622 40.455 3.975 ;
      RECT 40.445 3.605 40.45 3.975 ;
      RECT 40.44 3.592 40.445 3.975 ;
      RECT 40.365 3.475 40.44 3.975 ;
      RECT 40.32 3.292 40.365 3.975 ;
      RECT 40.315 3.22 40.32 3.975 ;
      RECT 40.3 3.195 40.315 3.975 ;
      RECT 40.275 3.157 40.3 3.975 ;
      RECT 40.265 3.137 40.275 3.697 ;
      RECT 40.25 3.129 40.265 3.652 ;
      RECT 40.245 3.121 40.25 3.623 ;
      RECT 40.24 3.118 40.245 3.603 ;
      RECT 40.235 3.115 40.24 3.583 ;
      RECT 40.23 3.112 40.235 3.563 ;
      RECT 40.2 3.101 40.23 3.5 ;
      RECT 40.18 3.086 40.2 3.415 ;
      RECT 40.175 3.078 40.18 3.378 ;
      RECT 40.165 3.072 40.175 3.345 ;
      RECT 40.15 3.064 40.165 3.305 ;
      RECT 40.145 3.057 40.15 3.265 ;
      RECT 40.14 3.054 40.145 3.243 ;
      RECT 40.135 3.051 40.14 3.23 ;
      RECT 40.13 3.05 40.135 3.22 ;
      RECT 40.115 3.044 40.13 3.21 ;
      RECT 40.09 3.031 40.115 3.195 ;
      RECT 40.04 3.006 40.09 3.166 ;
      RECT 40.025 2.985 40.04 3.141 ;
      RECT 40.015 2.978 40.025 3.13 ;
      RECT 39.96 2.959 40.015 3.103 ;
      RECT 39.935 2.937 39.96 3.076 ;
      RECT 39.93 2.93 39.935 3.071 ;
      RECT 39.915 2.93 39.93 3.069 ;
      RECT 39.89 2.922 39.915 3.065 ;
      RECT 39.875 2.92 39.89 3.061 ;
      RECT 39.845 2.92 39.875 3.058 ;
      RECT 39.835 2.92 39.845 3.053 ;
      RECT 39.79 2.92 39.835 3.051 ;
      RECT 39.761 2.92 39.79 3.052 ;
      RECT 39.675 2.92 39.761 3.054 ;
      RECT 39.661 2.921 39.675 3.056 ;
      RECT 39.575 2.922 39.661 3.058 ;
      RECT 39.56 2.923 39.575 3.068 ;
      RECT 39.555 2.924 39.56 3.077 ;
      RECT 39.535 2.927 39.555 3.087 ;
      RECT 39.52 2.935 39.535 3.102 ;
      RECT 39.5 2.953 39.52 3.117 ;
      RECT 39.49 2.965 39.5 3.14 ;
      RECT 39.48 2.974 39.49 3.17 ;
      RECT 39.465 2.986 39.48 3.215 ;
      RECT 39.41 3.019 39.465 3.53 ;
      RECT 39.405 3.047 39.41 3.53 ;
      RECT 39.385 3.062 39.405 3.53 ;
      RECT 39.35 3.122 39.385 3.53 ;
      RECT 39.348 3.172 39.35 3.53 ;
      RECT 39.345 3.18 39.348 3.53 ;
      RECT 39.335 3.195 39.345 3.53 ;
      RECT 39.33 3.207 39.335 3.53 ;
      RECT 39.32 3.232 39.33 3.53 ;
      RECT 39.31 3.26 39.32 3.53 ;
      RECT 37.215 4.765 37.265 5.025 ;
      RECT 40.125 4.315 40.185 4.575 ;
      RECT 40.11 4.315 40.125 4.585 ;
      RECT 40.091 4.315 40.11 4.618 ;
      RECT 40.005 4.315 40.091 4.743 ;
      RECT 39.925 4.315 40.005 4.925 ;
      RECT 39.92 4.552 39.925 5.01 ;
      RECT 39.895 4.622 39.92 5.038 ;
      RECT 39.89 4.692 39.895 5.065 ;
      RECT 39.87 4.764 39.89 5.087 ;
      RECT 39.865 4.831 39.87 5.11 ;
      RECT 39.855 4.86 39.865 5.125 ;
      RECT 39.845 4.882 39.855 5.142 ;
      RECT 39.84 4.892 39.845 5.153 ;
      RECT 39.835 4.9 39.84 5.161 ;
      RECT 39.825 4.908 39.835 5.173 ;
      RECT 39.82 4.92 39.825 5.183 ;
      RECT 39.815 4.928 39.82 5.188 ;
      RECT 39.795 4.946 39.815 5.198 ;
      RECT 39.79 4.963 39.795 5.205 ;
      RECT 39.785 4.971 39.79 5.206 ;
      RECT 39.78 4.982 39.785 5.208 ;
      RECT 39.74 5.02 39.78 5.218 ;
      RECT 39.735 5.055 39.74 5.229 ;
      RECT 39.73 5.06 39.735 5.232 ;
      RECT 39.705 5.07 39.73 5.239 ;
      RECT 39.695 5.084 39.705 5.248 ;
      RECT 39.675 5.096 39.695 5.251 ;
      RECT 39.625 5.115 39.675 5.255 ;
      RECT 39.58 5.13 39.625 5.26 ;
      RECT 39.515 5.133 39.58 5.266 ;
      RECT 39.5 5.131 39.515 5.273 ;
      RECT 39.47 5.13 39.5 5.273 ;
      RECT 39.431 5.129 39.47 5.269 ;
      RECT 39.345 5.126 39.431 5.265 ;
      RECT 39.328 5.124 39.345 5.262 ;
      RECT 39.242 5.122 39.328 5.259 ;
      RECT 39.156 5.119 39.242 5.253 ;
      RECT 39.07 5.115 39.156 5.248 ;
      RECT 38.992 5.112 39.07 5.244 ;
      RECT 38.906 5.109 38.992 5.242 ;
      RECT 38.82 5.106 38.906 5.239 ;
      RECT 38.762 5.104 38.82 5.236 ;
      RECT 38.676 5.101 38.762 5.234 ;
      RECT 38.59 5.097 38.676 5.232 ;
      RECT 38.504 5.094 38.59 5.229 ;
      RECT 38.418 5.09 38.504 5.227 ;
      RECT 38.332 5.086 38.418 5.224 ;
      RECT 38.246 5.083 38.332 5.222 ;
      RECT 38.16 5.079 38.246 5.219 ;
      RECT 38.074 5.076 38.16 5.217 ;
      RECT 37.988 5.072 38.074 5.214 ;
      RECT 37.902 5.069 37.988 5.212 ;
      RECT 37.816 5.065 37.902 5.209 ;
      RECT 37.73 5.062 37.816 5.207 ;
      RECT 37.72 5.06 37.73 5.203 ;
      RECT 37.715 5.06 37.72 5.201 ;
      RECT 37.675 5.055 37.715 5.195 ;
      RECT 37.661 5.046 37.675 5.188 ;
      RECT 37.575 5.016 37.661 5.173 ;
      RECT 37.555 4.982 37.575 5.158 ;
      RECT 37.485 4.951 37.555 5.145 ;
      RECT 37.48 4.926 37.485 5.134 ;
      RECT 37.475 4.92 37.48 5.132 ;
      RECT 37.406 4.765 37.475 5.12 ;
      RECT 37.32 4.765 37.406 5.094 ;
      RECT 37.295 4.765 37.32 5.073 ;
      RECT 37.29 4.765 37.295 5.063 ;
      RECT 37.285 4.765 37.29 5.055 ;
      RECT 37.265 4.765 37.285 5.038 ;
      RECT 39.685 3.335 39.945 3.595 ;
      RECT 39.67 3.335 39.945 3.498 ;
      RECT 39.64 3.335 39.945 3.473 ;
      RECT 39.605 3.175 39.885 3.455 ;
      RECT 39.575 4.665 39.635 4.925 ;
      RECT 38.6 3.355 38.655 3.615 ;
      RECT 39.535 4.622 39.575 4.925 ;
      RECT 39.506 4.543 39.535 4.925 ;
      RECT 39.42 4.415 39.506 4.925 ;
      RECT 39.4 4.295 39.42 4.925 ;
      RECT 39.375 4.246 39.4 4.925 ;
      RECT 39.37 4.211 39.375 4.775 ;
      RECT 39.34 4.171 39.37 4.713 ;
      RECT 39.315 4.108 39.34 4.628 ;
      RECT 39.305 4.07 39.315 4.565 ;
      RECT 39.29 4.045 39.305 4.526 ;
      RECT 39.247 4.003 39.29 4.432 ;
      RECT 39.245 3.976 39.247 4.359 ;
      RECT 39.24 3.971 39.245 4.35 ;
      RECT 39.235 3.964 39.24 4.325 ;
      RECT 39.23 3.958 39.235 4.31 ;
      RECT 39.225 3.952 39.23 4.298 ;
      RECT 39.215 3.943 39.225 4.28 ;
      RECT 39.21 3.934 39.215 4.258 ;
      RECT 39.185 3.915 39.21 4.208 ;
      RECT 39.18 3.896 39.185 4.158 ;
      RECT 39.165 3.882 39.18 4.118 ;
      RECT 39.16 3.868 39.165 4.085 ;
      RECT 39.155 3.861 39.16 4.078 ;
      RECT 39.14 3.848 39.155 4.07 ;
      RECT 39.095 3.81 39.14 4.043 ;
      RECT 39.065 3.763 39.095 4.008 ;
      RECT 39.045 3.732 39.065 3.985 ;
      RECT 38.965 3.665 39.045 3.938 ;
      RECT 38.935 3.595 38.965 3.885 ;
      RECT 38.93 3.572 38.935 3.868 ;
      RECT 38.9 3.55 38.93 3.853 ;
      RECT 38.87 3.509 38.9 3.825 ;
      RECT 38.865 3.484 38.87 3.81 ;
      RECT 38.86 3.478 38.865 3.803 ;
      RECT 38.85 3.355 38.86 3.795 ;
      RECT 38.84 3.355 38.85 3.788 ;
      RECT 38.835 3.355 38.84 3.78 ;
      RECT 38.815 3.355 38.835 3.768 ;
      RECT 38.765 3.355 38.815 3.738 ;
      RECT 38.71 3.355 38.765 3.688 ;
      RECT 38.68 3.355 38.71 3.648 ;
      RECT 38.655 3.355 38.68 3.625 ;
      RECT 38.525 4.08 38.805 4.36 ;
      RECT 38.49 3.995 38.75 4.255 ;
      RECT 38.49 4.077 38.76 4.255 ;
      RECT 36.69 3.45 36.695 3.935 ;
      RECT 36.58 3.635 36.585 3.935 ;
      RECT 36.49 3.675 36.555 3.935 ;
      RECT 38.165 3.175 38.255 3.805 ;
      RECT 38.13 3.225 38.135 3.805 ;
      RECT 38.075 3.25 38.085 3.805 ;
      RECT 38.03 3.25 38.04 3.805 ;
      RECT 38.4 3.175 38.445 3.455 ;
      RECT 37.25 2.905 37.45 3.045 ;
      RECT 38.366 3.175 38.4 3.467 ;
      RECT 38.28 3.175 38.366 3.507 ;
      RECT 38.265 3.175 38.28 3.548 ;
      RECT 38.26 3.175 38.265 3.568 ;
      RECT 38.255 3.175 38.26 3.588 ;
      RECT 38.135 3.217 38.165 3.805 ;
      RECT 38.085 3.237 38.13 3.805 ;
      RECT 38.07 3.252 38.075 3.805 ;
      RECT 38.04 3.252 38.07 3.805 ;
      RECT 37.995 3.237 38.03 3.805 ;
      RECT 37.99 3.225 37.995 3.585 ;
      RECT 37.985 3.222 37.99 3.565 ;
      RECT 37.97 3.212 37.985 3.518 ;
      RECT 37.965 3.205 37.97 3.481 ;
      RECT 37.96 3.202 37.965 3.464 ;
      RECT 37.945 3.192 37.96 3.42 ;
      RECT 37.94 3.183 37.945 3.38 ;
      RECT 37.935 3.179 37.94 3.365 ;
      RECT 37.925 3.173 37.935 3.348 ;
      RECT 37.885 3.154 37.925 3.323 ;
      RECT 37.88 3.136 37.885 3.303 ;
      RECT 37.87 3.13 37.88 3.298 ;
      RECT 37.84 3.114 37.87 3.285 ;
      RECT 37.825 3.096 37.84 3.268 ;
      RECT 37.81 3.084 37.825 3.255 ;
      RECT 37.805 3.076 37.81 3.248 ;
      RECT 37.775 3.062 37.805 3.235 ;
      RECT 37.77 3.047 37.775 3.223 ;
      RECT 37.76 3.041 37.77 3.215 ;
      RECT 37.74 3.029 37.76 3.203 ;
      RECT 37.73 3.017 37.74 3.19 ;
      RECT 37.7 3.001 37.73 3.175 ;
      RECT 37.68 2.981 37.7 3.158 ;
      RECT 37.675 2.971 37.68 3.148 ;
      RECT 37.65 2.959 37.675 3.135 ;
      RECT 37.645 2.947 37.65 3.123 ;
      RECT 37.64 2.942 37.645 3.119 ;
      RECT 37.625 2.935 37.64 3.111 ;
      RECT 37.615 2.922 37.625 3.101 ;
      RECT 37.61 2.92 37.615 3.095 ;
      RECT 37.585 2.913 37.61 3.084 ;
      RECT 37.58 2.906 37.585 3.073 ;
      RECT 37.555 2.905 37.58 3.06 ;
      RECT 37.536 2.905 37.555 3.05 ;
      RECT 37.45 2.905 37.536 3.047 ;
      RECT 37.22 2.905 37.25 3.05 ;
      RECT 37.18 2.912 37.22 3.063 ;
      RECT 37.155 2.922 37.18 3.076 ;
      RECT 37.14 2.931 37.155 3.086 ;
      RECT 37.11 2.936 37.14 3.105 ;
      RECT 37.105 2.942 37.11 3.123 ;
      RECT 37.085 2.952 37.105 3.138 ;
      RECT 37.075 2.965 37.085 3.158 ;
      RECT 37.06 2.977 37.075 3.175 ;
      RECT 37.055 2.987 37.06 3.185 ;
      RECT 37.05 2.992 37.055 3.19 ;
      RECT 37.04 3 37.05 3.203 ;
      RECT 36.99 3.032 37.04 3.24 ;
      RECT 36.975 3.067 36.99 3.281 ;
      RECT 36.97 3.077 36.975 3.296 ;
      RECT 36.965 3.082 36.97 3.303 ;
      RECT 36.94 3.098 36.965 3.323 ;
      RECT 36.925 3.119 36.94 3.348 ;
      RECT 36.9 3.14 36.925 3.373 ;
      RECT 36.89 3.159 36.9 3.396 ;
      RECT 36.865 3.177 36.89 3.419 ;
      RECT 36.85 3.197 36.865 3.443 ;
      RECT 36.845 3.207 36.85 3.455 ;
      RECT 36.83 3.219 36.845 3.475 ;
      RECT 36.82 3.234 36.83 3.515 ;
      RECT 36.815 3.242 36.82 3.543 ;
      RECT 36.805 3.252 36.815 3.563 ;
      RECT 36.8 3.265 36.805 3.588 ;
      RECT 36.795 3.278 36.8 3.608 ;
      RECT 36.79 3.284 36.795 3.63 ;
      RECT 36.78 3.293 36.79 3.65 ;
      RECT 36.775 3.313 36.78 3.673 ;
      RECT 36.77 3.319 36.775 3.693 ;
      RECT 36.765 3.326 36.77 3.715 ;
      RECT 36.76 3.337 36.765 3.728 ;
      RECT 36.75 3.347 36.76 3.753 ;
      RECT 36.73 3.372 36.75 3.935 ;
      RECT 36.7 3.412 36.73 3.935 ;
      RECT 36.695 3.442 36.7 3.935 ;
      RECT 36.67 3.47 36.69 3.935 ;
      RECT 36.64 3.515 36.67 3.935 ;
      RECT 36.635 3.542 36.64 3.935 ;
      RECT 36.615 3.56 36.635 3.935 ;
      RECT 36.605 3.585 36.615 3.935 ;
      RECT 36.6 3.597 36.605 3.935 ;
      RECT 36.585 3.62 36.6 3.935 ;
      RECT 36.565 3.647 36.58 3.935 ;
      RECT 36.555 3.67 36.565 3.935 ;
      RECT 38.345 4.555 38.425 4.815 ;
      RECT 37.58 3.775 37.65 4.035 ;
      RECT 38.311 4.522 38.345 4.815 ;
      RECT 38.225 4.425 38.311 4.815 ;
      RECT 38.205 4.337 38.225 4.815 ;
      RECT 38.195 4.307 38.205 4.815 ;
      RECT 38.185 4.287 38.195 4.815 ;
      RECT 38.165 4.274 38.185 4.815 ;
      RECT 38.15 4.264 38.165 4.643 ;
      RECT 38.145 4.257 38.15 4.598 ;
      RECT 38.135 4.251 38.145 4.588 ;
      RECT 38.125 4.243 38.135 4.57 ;
      RECT 38.12 4.237 38.125 4.558 ;
      RECT 38.11 4.232 38.12 4.545 ;
      RECT 38.09 4.222 38.11 4.518 ;
      RECT 38.05 4.201 38.09 4.47 ;
      RECT 38.035 4.182 38.05 4.428 ;
      RECT 38.01 4.168 38.035 4.398 ;
      RECT 38 4.156 38.01 4.365 ;
      RECT 37.995 4.151 38 4.355 ;
      RECT 37.965 4.137 37.995 4.335 ;
      RECT 37.955 4.121 37.965 4.308 ;
      RECT 37.95 4.116 37.955 4.298 ;
      RECT 37.925 4.107 37.95 4.278 ;
      RECT 37.915 4.095 37.925 4.258 ;
      RECT 37.845 4.063 37.915 4.233 ;
      RECT 37.84 4.032 37.845 4.21 ;
      RECT 37.791 3.775 37.84 4.193 ;
      RECT 37.705 3.775 37.791 4.152 ;
      RECT 37.65 3.775 37.705 4.08 ;
      RECT 37.74 4.56 37.9 4.82 ;
      RECT 37.265 3.175 37.315 3.86 ;
      RECT 37.055 3.6 37.09 3.86 ;
      RECT 37.37 3.175 37.375 3.635 ;
      RECT 37.46 3.175 37.485 3.455 ;
      RECT 37.735 4.557 37.74 4.82 ;
      RECT 37.7 4.545 37.735 4.82 ;
      RECT 37.64 4.518 37.7 4.82 ;
      RECT 37.635 4.501 37.64 4.674 ;
      RECT 37.63 4.498 37.635 4.661 ;
      RECT 37.61 4.491 37.63 4.648 ;
      RECT 37.575 4.474 37.61 4.63 ;
      RECT 37.535 4.453 37.575 4.61 ;
      RECT 37.53 4.441 37.535 4.598 ;
      RECT 37.49 4.427 37.53 4.584 ;
      RECT 37.47 4.41 37.49 4.566 ;
      RECT 37.46 4.402 37.47 4.558 ;
      RECT 37.445 3.175 37.46 3.473 ;
      RECT 37.43 4.392 37.46 4.545 ;
      RECT 37.415 3.175 37.445 3.518 ;
      RECT 37.42 4.382 37.43 4.532 ;
      RECT 37.39 4.367 37.42 4.519 ;
      RECT 37.375 3.175 37.415 3.585 ;
      RECT 37.375 4.335 37.39 4.505 ;
      RECT 37.37 4.307 37.375 4.499 ;
      RECT 37.365 3.175 37.37 3.64 ;
      RECT 37.355 4.277 37.37 4.493 ;
      RECT 37.36 3.175 37.365 3.653 ;
      RECT 37.35 3.175 37.36 3.673 ;
      RECT 37.315 4.19 37.355 4.478 ;
      RECT 37.315 3.175 37.35 3.713 ;
      RECT 37.31 4.122 37.315 4.466 ;
      RECT 37.295 4.077 37.31 4.461 ;
      RECT 37.29 4.015 37.295 4.456 ;
      RECT 37.265 3.922 37.29 4.449 ;
      RECT 37.26 3.175 37.265 4.441 ;
      RECT 37.245 3.175 37.26 4.428 ;
      RECT 37.225 3.175 37.245 4.385 ;
      RECT 37.215 3.175 37.225 4.335 ;
      RECT 37.21 3.175 37.215 4.308 ;
      RECT 37.205 3.175 37.21 4.286 ;
      RECT 37.2 3.401 37.205 4.269 ;
      RECT 37.195 3.423 37.2 4.247 ;
      RECT 37.19 3.465 37.195 4.23 ;
      RECT 37.16 3.515 37.19 4.174 ;
      RECT 37.155 3.542 37.16 4.116 ;
      RECT 37.14 3.56 37.155 4.08 ;
      RECT 37.135 3.578 37.14 4.044 ;
      RECT 37.129 3.585 37.135 4.025 ;
      RECT 37.125 3.592 37.129 4.008 ;
      RECT 37.12 3.597 37.125 3.977 ;
      RECT 37.11 3.6 37.12 3.952 ;
      RECT 37.1 3.6 37.11 3.918 ;
      RECT 37.095 3.6 37.1 3.895 ;
      RECT 37.09 3.6 37.095 3.875 ;
      RECT 36.005 3.735 36.285 4.015 ;
      RECT 36.005 3.735 36.305 3.91 ;
      RECT 36.095 3.625 36.355 3.885 ;
      RECT 36.06 3.72 36.355 3.885 ;
      RECT 36.185 2.24 36.35 3.885 ;
      RECT 36.085 2.24 36.455 2.61 ;
      RECT 35.71 4.765 35.97 5.025 ;
      RECT 35.73 4.692 35.91 5.025 ;
      RECT 35.73 4.435 35.905 5.025 ;
      RECT 35.73 4.227 35.895 5.025 ;
      RECT 35.735 4.145 35.895 5.025 ;
      RECT 35.735 3.91 35.885 5.025 ;
      RECT 35.735 3.757 35.88 5.025 ;
      RECT 35.74 3.742 35.88 5.025 ;
      RECT 35.79 3.457 35.88 5.025 ;
      RECT 35.745 3.692 35.88 5.025 ;
      RECT 35.775 3.51 35.88 5.025 ;
      RECT 35.76 3.622 35.88 5.025 ;
      RECT 35.765 3.58 35.88 5.025 ;
      RECT 35.76 3.622 35.895 3.685 ;
      RECT 35.795 3.21 35.9 3.63 ;
      RECT 35.795 3.21 35.915 3.613 ;
      RECT 35.795 3.21 35.95 3.575 ;
      RECT 35.79 3.457 36 3.508 ;
      RECT 35.795 3.21 36.055 3.47 ;
      RECT 35.055 3.915 35.315 4.175 ;
      RECT 35.055 3.915 35.325 4.133 ;
      RECT 35.055 3.915 35.411 4.104 ;
      RECT 35.055 3.915 35.48 4.056 ;
      RECT 35.055 3.915 35.515 4.025 ;
      RECT 35.285 3.735 35.565 4.015 ;
      RECT 35.12 3.9 35.565 4.015 ;
      RECT 35.21 3.777 35.315 4.175 ;
      RECT 35.14 3.84 35.565 4.015 ;
      RECT 29.59 8.51 29.91 8.835 ;
      RECT 29.62 7.985 29.79 8.835 ;
      RECT 29.62 7.985 29.795 8.335 ;
      RECT 29.62 7.985 30.595 8.16 ;
      RECT 30.42 3.26 30.595 8.16 ;
      RECT 30.365 3.26 30.715 3.61 ;
      RECT 30.39 8.945 30.715 9.27 ;
      RECT 29.275 9.035 30.715 9.205 ;
      RECT 29.275 3.69 29.435 9.205 ;
      RECT 29.59 3.66 29.91 3.98 ;
      RECT 29.275 3.69 29.91 3.86 ;
      RECT 27.94 4 28.325 4.35 ;
      RECT 27.93 4.065 28.325 4.265 ;
      RECT 28.075 3.995 28.245 4.35 ;
      RECT 26.385 3.735 26.665 4.015 ;
      RECT 26.38 3.735 26.665 3.968 ;
      RECT 26.36 3.735 26.665 3.945 ;
      RECT 26.35 3.735 26.665 3.925 ;
      RECT 26.34 3.735 26.665 3.91 ;
      RECT 26.315 3.735 26.665 3.883 ;
      RECT 26.305 3.735 26.665 3.858 ;
      RECT 26.26 3.59 26.54 3.85 ;
      RECT 26.26 3.685 26.64 3.85 ;
      RECT 26.26 3.63 26.585 3.85 ;
      RECT 26.26 3.622 26.58 3.85 ;
      RECT 26.26 3.612 26.575 3.85 ;
      RECT 26.26 3.6 26.57 3.85 ;
      RECT 25.185 4.295 25.465 4.575 ;
      RECT 25.185 4.295 25.5 4.555 ;
      RECT 17.51 8.945 17.86 9.295 ;
      RECT 24.93 8.9 25.28 9.25 ;
      RECT 17.51 8.975 25.28 9.175 ;
      RECT 25.22 3.715 25.27 3.975 ;
      RECT 25.01 3.715 25.015 3.975 ;
      RECT 24.205 3.27 24.235 3.53 ;
      RECT 23.975 3.27 24.05 3.53 ;
      RECT 25.195 3.665 25.22 3.975 ;
      RECT 25.19 3.622 25.195 3.975 ;
      RECT 25.185 3.605 25.19 3.975 ;
      RECT 25.18 3.592 25.185 3.975 ;
      RECT 25.105 3.475 25.18 3.975 ;
      RECT 25.06 3.292 25.105 3.975 ;
      RECT 25.055 3.22 25.06 3.975 ;
      RECT 25.04 3.195 25.055 3.975 ;
      RECT 25.015 3.157 25.04 3.975 ;
      RECT 25.005 3.137 25.015 3.697 ;
      RECT 24.99 3.129 25.005 3.652 ;
      RECT 24.985 3.121 24.99 3.623 ;
      RECT 24.98 3.118 24.985 3.603 ;
      RECT 24.975 3.115 24.98 3.583 ;
      RECT 24.97 3.112 24.975 3.563 ;
      RECT 24.94 3.101 24.97 3.5 ;
      RECT 24.92 3.086 24.94 3.415 ;
      RECT 24.915 3.078 24.92 3.378 ;
      RECT 24.905 3.072 24.915 3.345 ;
      RECT 24.89 3.064 24.905 3.305 ;
      RECT 24.885 3.057 24.89 3.265 ;
      RECT 24.88 3.054 24.885 3.243 ;
      RECT 24.875 3.051 24.88 3.23 ;
      RECT 24.87 3.05 24.875 3.22 ;
      RECT 24.855 3.044 24.87 3.21 ;
      RECT 24.83 3.031 24.855 3.195 ;
      RECT 24.78 3.006 24.83 3.166 ;
      RECT 24.765 2.985 24.78 3.141 ;
      RECT 24.755 2.978 24.765 3.13 ;
      RECT 24.7 2.959 24.755 3.103 ;
      RECT 24.675 2.937 24.7 3.076 ;
      RECT 24.67 2.93 24.675 3.071 ;
      RECT 24.655 2.93 24.67 3.069 ;
      RECT 24.63 2.922 24.655 3.065 ;
      RECT 24.615 2.92 24.63 3.061 ;
      RECT 24.585 2.92 24.615 3.058 ;
      RECT 24.575 2.92 24.585 3.053 ;
      RECT 24.53 2.92 24.575 3.051 ;
      RECT 24.501 2.92 24.53 3.052 ;
      RECT 24.415 2.92 24.501 3.054 ;
      RECT 24.401 2.921 24.415 3.056 ;
      RECT 24.315 2.922 24.401 3.058 ;
      RECT 24.3 2.923 24.315 3.068 ;
      RECT 24.295 2.924 24.3 3.077 ;
      RECT 24.275 2.927 24.295 3.087 ;
      RECT 24.26 2.935 24.275 3.102 ;
      RECT 24.24 2.953 24.26 3.117 ;
      RECT 24.23 2.965 24.24 3.14 ;
      RECT 24.22 2.974 24.23 3.17 ;
      RECT 24.205 2.986 24.22 3.215 ;
      RECT 24.15 3.019 24.205 3.53 ;
      RECT 24.145 3.047 24.15 3.53 ;
      RECT 24.125 3.062 24.145 3.53 ;
      RECT 24.09 3.122 24.125 3.53 ;
      RECT 24.088 3.172 24.09 3.53 ;
      RECT 24.085 3.18 24.088 3.53 ;
      RECT 24.075 3.195 24.085 3.53 ;
      RECT 24.07 3.207 24.075 3.53 ;
      RECT 24.06 3.232 24.07 3.53 ;
      RECT 24.05 3.26 24.06 3.53 ;
      RECT 21.955 4.765 22.005 5.025 ;
      RECT 24.865 4.315 24.925 4.575 ;
      RECT 24.85 4.315 24.865 4.585 ;
      RECT 24.831 4.315 24.85 4.618 ;
      RECT 24.745 4.315 24.831 4.743 ;
      RECT 24.665 4.315 24.745 4.925 ;
      RECT 24.66 4.552 24.665 5.01 ;
      RECT 24.635 4.622 24.66 5.038 ;
      RECT 24.63 4.692 24.635 5.065 ;
      RECT 24.61 4.764 24.63 5.087 ;
      RECT 24.605 4.831 24.61 5.11 ;
      RECT 24.595 4.86 24.605 5.125 ;
      RECT 24.585 4.882 24.595 5.142 ;
      RECT 24.58 4.892 24.585 5.153 ;
      RECT 24.575 4.9 24.58 5.161 ;
      RECT 24.565 4.908 24.575 5.173 ;
      RECT 24.56 4.92 24.565 5.183 ;
      RECT 24.555 4.928 24.56 5.188 ;
      RECT 24.535 4.946 24.555 5.198 ;
      RECT 24.53 4.963 24.535 5.205 ;
      RECT 24.525 4.971 24.53 5.206 ;
      RECT 24.52 4.982 24.525 5.208 ;
      RECT 24.48 5.02 24.52 5.218 ;
      RECT 24.475 5.055 24.48 5.229 ;
      RECT 24.47 5.06 24.475 5.232 ;
      RECT 24.445 5.07 24.47 5.239 ;
      RECT 24.435 5.084 24.445 5.248 ;
      RECT 24.415 5.096 24.435 5.251 ;
      RECT 24.365 5.115 24.415 5.255 ;
      RECT 24.32 5.13 24.365 5.26 ;
      RECT 24.255 5.133 24.32 5.266 ;
      RECT 24.24 5.131 24.255 5.273 ;
      RECT 24.21 5.13 24.24 5.273 ;
      RECT 24.171 5.129 24.21 5.269 ;
      RECT 24.085 5.126 24.171 5.265 ;
      RECT 24.068 5.124 24.085 5.262 ;
      RECT 23.982 5.122 24.068 5.259 ;
      RECT 23.896 5.119 23.982 5.253 ;
      RECT 23.81 5.115 23.896 5.248 ;
      RECT 23.732 5.112 23.81 5.244 ;
      RECT 23.646 5.109 23.732 5.242 ;
      RECT 23.56 5.106 23.646 5.239 ;
      RECT 23.502 5.104 23.56 5.236 ;
      RECT 23.416 5.101 23.502 5.234 ;
      RECT 23.33 5.097 23.416 5.232 ;
      RECT 23.244 5.094 23.33 5.229 ;
      RECT 23.158 5.09 23.244 5.227 ;
      RECT 23.072 5.086 23.158 5.224 ;
      RECT 22.986 5.083 23.072 5.222 ;
      RECT 22.9 5.079 22.986 5.219 ;
      RECT 22.814 5.076 22.9 5.217 ;
      RECT 22.728 5.072 22.814 5.214 ;
      RECT 22.642 5.069 22.728 5.212 ;
      RECT 22.556 5.065 22.642 5.209 ;
      RECT 22.47 5.062 22.556 5.207 ;
      RECT 22.46 5.06 22.47 5.203 ;
      RECT 22.455 5.06 22.46 5.201 ;
      RECT 22.415 5.055 22.455 5.195 ;
      RECT 22.401 5.046 22.415 5.188 ;
      RECT 22.315 5.016 22.401 5.173 ;
      RECT 22.295 4.982 22.315 5.158 ;
      RECT 22.225 4.951 22.295 5.145 ;
      RECT 22.22 4.926 22.225 5.134 ;
      RECT 22.215 4.92 22.22 5.132 ;
      RECT 22.146 4.765 22.215 5.12 ;
      RECT 22.06 4.765 22.146 5.094 ;
      RECT 22.035 4.765 22.06 5.073 ;
      RECT 22.03 4.765 22.035 5.063 ;
      RECT 22.025 4.765 22.03 5.055 ;
      RECT 22.005 4.765 22.025 5.038 ;
      RECT 24.425 3.335 24.685 3.595 ;
      RECT 24.41 3.335 24.685 3.498 ;
      RECT 24.38 3.335 24.685 3.473 ;
      RECT 24.345 3.175 24.625 3.455 ;
      RECT 24.315 4.665 24.375 4.925 ;
      RECT 23.34 3.355 23.395 3.615 ;
      RECT 24.275 4.622 24.315 4.925 ;
      RECT 24.246 4.543 24.275 4.925 ;
      RECT 24.16 4.415 24.246 4.925 ;
      RECT 24.14 4.295 24.16 4.925 ;
      RECT 24.115 4.246 24.14 4.925 ;
      RECT 24.11 4.211 24.115 4.775 ;
      RECT 24.08 4.171 24.11 4.713 ;
      RECT 24.055 4.108 24.08 4.628 ;
      RECT 24.045 4.07 24.055 4.565 ;
      RECT 24.03 4.045 24.045 4.526 ;
      RECT 23.987 4.003 24.03 4.432 ;
      RECT 23.985 3.976 23.987 4.359 ;
      RECT 23.98 3.971 23.985 4.35 ;
      RECT 23.975 3.964 23.98 4.325 ;
      RECT 23.97 3.958 23.975 4.31 ;
      RECT 23.965 3.952 23.97 4.298 ;
      RECT 23.955 3.943 23.965 4.28 ;
      RECT 23.95 3.934 23.955 4.258 ;
      RECT 23.925 3.915 23.95 4.208 ;
      RECT 23.92 3.896 23.925 4.158 ;
      RECT 23.905 3.882 23.92 4.118 ;
      RECT 23.9 3.868 23.905 4.085 ;
      RECT 23.895 3.861 23.9 4.078 ;
      RECT 23.88 3.848 23.895 4.07 ;
      RECT 23.835 3.81 23.88 4.043 ;
      RECT 23.805 3.763 23.835 4.008 ;
      RECT 23.785 3.732 23.805 3.985 ;
      RECT 23.705 3.665 23.785 3.938 ;
      RECT 23.675 3.595 23.705 3.885 ;
      RECT 23.67 3.572 23.675 3.868 ;
      RECT 23.64 3.55 23.67 3.853 ;
      RECT 23.61 3.509 23.64 3.825 ;
      RECT 23.605 3.484 23.61 3.81 ;
      RECT 23.6 3.478 23.605 3.803 ;
      RECT 23.59 3.355 23.6 3.795 ;
      RECT 23.58 3.355 23.59 3.788 ;
      RECT 23.575 3.355 23.58 3.78 ;
      RECT 23.555 3.355 23.575 3.768 ;
      RECT 23.505 3.355 23.555 3.738 ;
      RECT 23.45 3.355 23.505 3.688 ;
      RECT 23.42 3.355 23.45 3.648 ;
      RECT 23.395 3.355 23.42 3.625 ;
      RECT 23.265 4.08 23.545 4.36 ;
      RECT 23.23 3.995 23.49 4.255 ;
      RECT 23.23 4.077 23.5 4.255 ;
      RECT 21.43 3.45 21.435 3.935 ;
      RECT 21.32 3.635 21.325 3.935 ;
      RECT 21.23 3.675 21.295 3.935 ;
      RECT 22.905 3.175 22.995 3.805 ;
      RECT 22.87 3.225 22.875 3.805 ;
      RECT 22.815 3.25 22.825 3.805 ;
      RECT 22.77 3.25 22.78 3.805 ;
      RECT 23.14 3.175 23.185 3.455 ;
      RECT 21.99 2.905 22.19 3.045 ;
      RECT 23.106 3.175 23.14 3.467 ;
      RECT 23.02 3.175 23.106 3.507 ;
      RECT 23.005 3.175 23.02 3.548 ;
      RECT 23 3.175 23.005 3.568 ;
      RECT 22.995 3.175 23 3.588 ;
      RECT 22.875 3.217 22.905 3.805 ;
      RECT 22.825 3.237 22.87 3.805 ;
      RECT 22.81 3.252 22.815 3.805 ;
      RECT 22.78 3.252 22.81 3.805 ;
      RECT 22.735 3.237 22.77 3.805 ;
      RECT 22.73 3.225 22.735 3.585 ;
      RECT 22.725 3.222 22.73 3.565 ;
      RECT 22.71 3.212 22.725 3.518 ;
      RECT 22.705 3.205 22.71 3.481 ;
      RECT 22.7 3.202 22.705 3.464 ;
      RECT 22.685 3.192 22.7 3.42 ;
      RECT 22.68 3.183 22.685 3.38 ;
      RECT 22.675 3.179 22.68 3.365 ;
      RECT 22.665 3.173 22.675 3.348 ;
      RECT 22.625 3.154 22.665 3.323 ;
      RECT 22.62 3.136 22.625 3.303 ;
      RECT 22.61 3.13 22.62 3.298 ;
      RECT 22.58 3.114 22.61 3.285 ;
      RECT 22.565 3.096 22.58 3.268 ;
      RECT 22.55 3.084 22.565 3.255 ;
      RECT 22.545 3.076 22.55 3.248 ;
      RECT 22.515 3.062 22.545 3.235 ;
      RECT 22.51 3.047 22.515 3.223 ;
      RECT 22.5 3.041 22.51 3.215 ;
      RECT 22.48 3.029 22.5 3.203 ;
      RECT 22.47 3.017 22.48 3.19 ;
      RECT 22.44 3.001 22.47 3.175 ;
      RECT 22.42 2.981 22.44 3.158 ;
      RECT 22.415 2.971 22.42 3.148 ;
      RECT 22.39 2.959 22.415 3.135 ;
      RECT 22.385 2.947 22.39 3.123 ;
      RECT 22.38 2.942 22.385 3.119 ;
      RECT 22.365 2.935 22.38 3.111 ;
      RECT 22.355 2.922 22.365 3.101 ;
      RECT 22.35 2.92 22.355 3.095 ;
      RECT 22.325 2.913 22.35 3.084 ;
      RECT 22.32 2.906 22.325 3.073 ;
      RECT 22.295 2.905 22.32 3.06 ;
      RECT 22.276 2.905 22.295 3.05 ;
      RECT 22.19 2.905 22.276 3.047 ;
      RECT 21.96 2.905 21.99 3.05 ;
      RECT 21.92 2.912 21.96 3.063 ;
      RECT 21.895 2.922 21.92 3.076 ;
      RECT 21.88 2.931 21.895 3.086 ;
      RECT 21.85 2.936 21.88 3.105 ;
      RECT 21.845 2.942 21.85 3.123 ;
      RECT 21.825 2.952 21.845 3.138 ;
      RECT 21.815 2.965 21.825 3.158 ;
      RECT 21.8 2.977 21.815 3.175 ;
      RECT 21.795 2.987 21.8 3.185 ;
      RECT 21.79 2.992 21.795 3.19 ;
      RECT 21.78 3 21.79 3.203 ;
      RECT 21.73 3.032 21.78 3.24 ;
      RECT 21.715 3.067 21.73 3.281 ;
      RECT 21.71 3.077 21.715 3.296 ;
      RECT 21.705 3.082 21.71 3.303 ;
      RECT 21.68 3.098 21.705 3.323 ;
      RECT 21.665 3.119 21.68 3.348 ;
      RECT 21.64 3.14 21.665 3.373 ;
      RECT 21.63 3.159 21.64 3.396 ;
      RECT 21.605 3.177 21.63 3.419 ;
      RECT 21.59 3.197 21.605 3.443 ;
      RECT 21.585 3.207 21.59 3.455 ;
      RECT 21.57 3.219 21.585 3.475 ;
      RECT 21.56 3.234 21.57 3.515 ;
      RECT 21.555 3.242 21.56 3.543 ;
      RECT 21.545 3.252 21.555 3.563 ;
      RECT 21.54 3.265 21.545 3.588 ;
      RECT 21.535 3.278 21.54 3.608 ;
      RECT 21.53 3.284 21.535 3.63 ;
      RECT 21.52 3.293 21.53 3.65 ;
      RECT 21.515 3.313 21.52 3.673 ;
      RECT 21.51 3.319 21.515 3.693 ;
      RECT 21.505 3.326 21.51 3.715 ;
      RECT 21.5 3.337 21.505 3.728 ;
      RECT 21.49 3.347 21.5 3.753 ;
      RECT 21.47 3.372 21.49 3.935 ;
      RECT 21.44 3.412 21.47 3.935 ;
      RECT 21.435 3.442 21.44 3.935 ;
      RECT 21.41 3.47 21.43 3.935 ;
      RECT 21.38 3.515 21.41 3.935 ;
      RECT 21.375 3.542 21.38 3.935 ;
      RECT 21.355 3.56 21.375 3.935 ;
      RECT 21.345 3.585 21.355 3.935 ;
      RECT 21.34 3.597 21.345 3.935 ;
      RECT 21.325 3.62 21.34 3.935 ;
      RECT 21.305 3.647 21.32 3.935 ;
      RECT 21.295 3.67 21.305 3.935 ;
      RECT 23.085 4.555 23.165 4.815 ;
      RECT 22.32 3.775 22.39 4.035 ;
      RECT 23.051 4.522 23.085 4.815 ;
      RECT 22.965 4.425 23.051 4.815 ;
      RECT 22.945 4.337 22.965 4.815 ;
      RECT 22.935 4.307 22.945 4.815 ;
      RECT 22.925 4.287 22.935 4.815 ;
      RECT 22.905 4.274 22.925 4.815 ;
      RECT 22.89 4.264 22.905 4.643 ;
      RECT 22.885 4.257 22.89 4.598 ;
      RECT 22.875 4.251 22.885 4.588 ;
      RECT 22.865 4.243 22.875 4.57 ;
      RECT 22.86 4.237 22.865 4.558 ;
      RECT 22.85 4.232 22.86 4.545 ;
      RECT 22.83 4.222 22.85 4.518 ;
      RECT 22.79 4.201 22.83 4.47 ;
      RECT 22.775 4.182 22.79 4.428 ;
      RECT 22.75 4.168 22.775 4.398 ;
      RECT 22.74 4.156 22.75 4.365 ;
      RECT 22.735 4.151 22.74 4.355 ;
      RECT 22.705 4.137 22.735 4.335 ;
      RECT 22.695 4.121 22.705 4.308 ;
      RECT 22.69 4.116 22.695 4.298 ;
      RECT 22.665 4.107 22.69 4.278 ;
      RECT 22.655 4.095 22.665 4.258 ;
      RECT 22.585 4.063 22.655 4.233 ;
      RECT 22.58 4.032 22.585 4.21 ;
      RECT 22.531 3.775 22.58 4.193 ;
      RECT 22.445 3.775 22.531 4.152 ;
      RECT 22.39 3.775 22.445 4.08 ;
      RECT 22.48 4.56 22.64 4.82 ;
      RECT 22.005 3.175 22.055 3.86 ;
      RECT 21.795 3.6 21.83 3.86 ;
      RECT 22.11 3.175 22.115 3.635 ;
      RECT 22.2 3.175 22.225 3.455 ;
      RECT 22.475 4.557 22.48 4.82 ;
      RECT 22.44 4.545 22.475 4.82 ;
      RECT 22.38 4.518 22.44 4.82 ;
      RECT 22.375 4.501 22.38 4.674 ;
      RECT 22.37 4.498 22.375 4.661 ;
      RECT 22.35 4.491 22.37 4.648 ;
      RECT 22.315 4.474 22.35 4.63 ;
      RECT 22.275 4.453 22.315 4.61 ;
      RECT 22.27 4.441 22.275 4.598 ;
      RECT 22.23 4.427 22.27 4.584 ;
      RECT 22.21 4.41 22.23 4.566 ;
      RECT 22.2 4.402 22.21 4.558 ;
      RECT 22.185 3.175 22.2 3.473 ;
      RECT 22.17 4.392 22.2 4.545 ;
      RECT 22.155 3.175 22.185 3.518 ;
      RECT 22.16 4.382 22.17 4.532 ;
      RECT 22.13 4.367 22.16 4.519 ;
      RECT 22.115 3.175 22.155 3.585 ;
      RECT 22.115 4.335 22.13 4.505 ;
      RECT 22.11 4.307 22.115 4.499 ;
      RECT 22.105 3.175 22.11 3.64 ;
      RECT 22.095 4.277 22.11 4.493 ;
      RECT 22.1 3.175 22.105 3.653 ;
      RECT 22.09 3.175 22.1 3.673 ;
      RECT 22.055 4.19 22.095 4.478 ;
      RECT 22.055 3.175 22.09 3.713 ;
      RECT 22.05 4.122 22.055 4.466 ;
      RECT 22.035 4.077 22.05 4.461 ;
      RECT 22.03 4.015 22.035 4.456 ;
      RECT 22.005 3.922 22.03 4.449 ;
      RECT 22 3.175 22.005 4.441 ;
      RECT 21.985 3.175 22 4.428 ;
      RECT 21.965 3.175 21.985 4.385 ;
      RECT 21.955 3.175 21.965 4.335 ;
      RECT 21.95 3.175 21.955 4.308 ;
      RECT 21.945 3.175 21.95 4.286 ;
      RECT 21.94 3.401 21.945 4.269 ;
      RECT 21.935 3.423 21.94 4.247 ;
      RECT 21.93 3.465 21.935 4.23 ;
      RECT 21.9 3.515 21.93 4.174 ;
      RECT 21.895 3.542 21.9 4.116 ;
      RECT 21.88 3.56 21.895 4.08 ;
      RECT 21.875 3.578 21.88 4.044 ;
      RECT 21.869 3.585 21.875 4.025 ;
      RECT 21.865 3.592 21.869 4.008 ;
      RECT 21.86 3.597 21.865 3.977 ;
      RECT 21.85 3.6 21.86 3.952 ;
      RECT 21.84 3.6 21.85 3.918 ;
      RECT 21.835 3.6 21.84 3.895 ;
      RECT 21.83 3.6 21.835 3.875 ;
      RECT 20.745 3.735 21.025 4.015 ;
      RECT 20.745 3.735 21.045 3.91 ;
      RECT 20.835 3.625 21.095 3.885 ;
      RECT 20.8 3.72 21.095 3.885 ;
      RECT 20.925 2.24 21.09 3.885 ;
      RECT 20.825 2.24 21.195 2.61 ;
      RECT 20.45 4.765 20.71 5.025 ;
      RECT 20.47 4.692 20.65 5.025 ;
      RECT 20.47 4.435 20.645 5.025 ;
      RECT 20.47 4.227 20.635 5.025 ;
      RECT 20.475 4.145 20.635 5.025 ;
      RECT 20.475 3.91 20.625 5.025 ;
      RECT 20.475 3.757 20.62 5.025 ;
      RECT 20.48 3.742 20.62 5.025 ;
      RECT 20.53 3.457 20.62 5.025 ;
      RECT 20.485 3.692 20.62 5.025 ;
      RECT 20.515 3.51 20.62 5.025 ;
      RECT 20.5 3.622 20.62 5.025 ;
      RECT 20.505 3.58 20.62 5.025 ;
      RECT 20.5 3.622 20.635 3.685 ;
      RECT 20.535 3.21 20.64 3.63 ;
      RECT 20.535 3.21 20.655 3.613 ;
      RECT 20.535 3.21 20.69 3.575 ;
      RECT 20.53 3.457 20.74 3.508 ;
      RECT 20.535 3.21 20.795 3.47 ;
      RECT 19.795 3.915 20.055 4.175 ;
      RECT 19.795 3.915 20.065 4.133 ;
      RECT 19.795 3.915 20.151 4.104 ;
      RECT 19.795 3.915 20.22 4.056 ;
      RECT 19.795 3.915 20.255 4.025 ;
      RECT 20.025 3.735 20.305 4.015 ;
      RECT 19.86 3.9 20.305 4.015 ;
      RECT 19.95 3.777 20.055 4.175 ;
      RECT 19.88 3.84 20.305 4.015 ;
      RECT 14.33 8.51 14.65 8.835 ;
      RECT 14.36 7.985 14.53 8.835 ;
      RECT 14.36 7.985 14.535 8.335 ;
      RECT 14.36 7.985 15.335 8.16 ;
      RECT 15.16 3.26 15.335 8.16 ;
      RECT 15.105 3.26 15.455 3.61 ;
      RECT 15.13 8.945 15.455 9.27 ;
      RECT 14.015 9.035 15.455 9.205 ;
      RECT 14.015 3.69 14.175 9.205 ;
      RECT 14.33 3.66 14.65 3.98 ;
      RECT 14.015 3.69 14.65 3.86 ;
      RECT 12.68 4 13.065 4.35 ;
      RECT 12.67 4.065 13.065 4.265 ;
      RECT 12.815 3.995 12.985 4.35 ;
      RECT 11.125 3.735 11.405 4.015 ;
      RECT 11.12 3.735 11.405 3.968 ;
      RECT 11.1 3.735 11.405 3.945 ;
      RECT 11.09 3.735 11.405 3.925 ;
      RECT 11.08 3.735 11.405 3.91 ;
      RECT 11.055 3.735 11.405 3.883 ;
      RECT 11.045 3.735 11.405 3.858 ;
      RECT 11 3.59 11.28 3.85 ;
      RECT 11 3.685 11.38 3.85 ;
      RECT 11 3.63 11.325 3.85 ;
      RECT 11 3.622 11.32 3.85 ;
      RECT 11 3.612 11.315 3.85 ;
      RECT 11 3.6 11.31 3.85 ;
      RECT 9.925 4.295 10.205 4.575 ;
      RECT 9.925 4.295 10.24 4.555 ;
      RECT 1.545 9.285 1.835 9.635 ;
      RECT 1.545 9.36 2.91 9.53 ;
      RECT 2.74 8.975 2.91 9.53 ;
      RECT 9.67 8.895 10.02 9.245 ;
      RECT 2.74 8.975 10.02 9.145 ;
      RECT 9.96 3.715 10.01 3.975 ;
      RECT 9.75 3.715 9.755 3.975 ;
      RECT 8.945 3.27 8.975 3.53 ;
      RECT 8.715 3.27 8.79 3.53 ;
      RECT 9.935 3.665 9.96 3.975 ;
      RECT 9.93 3.622 9.935 3.975 ;
      RECT 9.925 3.605 9.93 3.975 ;
      RECT 9.92 3.592 9.925 3.975 ;
      RECT 9.845 3.475 9.92 3.975 ;
      RECT 9.8 3.292 9.845 3.975 ;
      RECT 9.795 3.22 9.8 3.975 ;
      RECT 9.78 3.195 9.795 3.975 ;
      RECT 9.755 3.157 9.78 3.975 ;
      RECT 9.745 3.137 9.755 3.697 ;
      RECT 9.73 3.129 9.745 3.652 ;
      RECT 9.725 3.121 9.73 3.623 ;
      RECT 9.72 3.118 9.725 3.603 ;
      RECT 9.715 3.115 9.72 3.583 ;
      RECT 9.71 3.112 9.715 3.563 ;
      RECT 9.68 3.101 9.71 3.5 ;
      RECT 9.66 3.086 9.68 3.415 ;
      RECT 9.655 3.078 9.66 3.378 ;
      RECT 9.645 3.072 9.655 3.345 ;
      RECT 9.63 3.064 9.645 3.305 ;
      RECT 9.625 3.057 9.63 3.265 ;
      RECT 9.62 3.054 9.625 3.243 ;
      RECT 9.615 3.051 9.62 3.23 ;
      RECT 9.61 3.05 9.615 3.22 ;
      RECT 9.595 3.044 9.61 3.21 ;
      RECT 9.57 3.031 9.595 3.195 ;
      RECT 9.52 3.006 9.57 3.166 ;
      RECT 9.505 2.985 9.52 3.141 ;
      RECT 9.495 2.978 9.505 3.13 ;
      RECT 9.44 2.959 9.495 3.103 ;
      RECT 9.415 2.937 9.44 3.076 ;
      RECT 9.41 2.93 9.415 3.071 ;
      RECT 9.395 2.93 9.41 3.069 ;
      RECT 9.37 2.922 9.395 3.065 ;
      RECT 9.355 2.92 9.37 3.061 ;
      RECT 9.325 2.92 9.355 3.058 ;
      RECT 9.315 2.92 9.325 3.053 ;
      RECT 9.27 2.92 9.315 3.051 ;
      RECT 9.241 2.92 9.27 3.052 ;
      RECT 9.155 2.92 9.241 3.054 ;
      RECT 9.141 2.921 9.155 3.056 ;
      RECT 9.055 2.922 9.141 3.058 ;
      RECT 9.04 2.923 9.055 3.068 ;
      RECT 9.035 2.924 9.04 3.077 ;
      RECT 9.015 2.927 9.035 3.087 ;
      RECT 9 2.935 9.015 3.102 ;
      RECT 8.98 2.953 9 3.117 ;
      RECT 8.97 2.965 8.98 3.14 ;
      RECT 8.96 2.974 8.97 3.17 ;
      RECT 8.945 2.986 8.96 3.215 ;
      RECT 8.89 3.019 8.945 3.53 ;
      RECT 8.885 3.047 8.89 3.53 ;
      RECT 8.865 3.062 8.885 3.53 ;
      RECT 8.83 3.122 8.865 3.53 ;
      RECT 8.828 3.172 8.83 3.53 ;
      RECT 8.825 3.18 8.828 3.53 ;
      RECT 8.815 3.195 8.825 3.53 ;
      RECT 8.81 3.207 8.815 3.53 ;
      RECT 8.8 3.232 8.81 3.53 ;
      RECT 8.79 3.26 8.8 3.53 ;
      RECT 6.695 4.765 6.745 5.025 ;
      RECT 9.605 4.315 9.665 4.575 ;
      RECT 9.59 4.315 9.605 4.585 ;
      RECT 9.571 4.315 9.59 4.618 ;
      RECT 9.485 4.315 9.571 4.743 ;
      RECT 9.405 4.315 9.485 4.925 ;
      RECT 9.4 4.552 9.405 5.01 ;
      RECT 9.375 4.622 9.4 5.038 ;
      RECT 9.37 4.692 9.375 5.065 ;
      RECT 9.35 4.764 9.37 5.087 ;
      RECT 9.345 4.831 9.35 5.11 ;
      RECT 9.335 4.86 9.345 5.125 ;
      RECT 9.325 4.882 9.335 5.142 ;
      RECT 9.32 4.892 9.325 5.153 ;
      RECT 9.315 4.9 9.32 5.161 ;
      RECT 9.305 4.908 9.315 5.173 ;
      RECT 9.3 4.92 9.305 5.183 ;
      RECT 9.295 4.928 9.3 5.188 ;
      RECT 9.275 4.946 9.295 5.198 ;
      RECT 9.27 4.963 9.275 5.205 ;
      RECT 9.265 4.971 9.27 5.206 ;
      RECT 9.26 4.982 9.265 5.208 ;
      RECT 9.22 5.02 9.26 5.218 ;
      RECT 9.215 5.055 9.22 5.229 ;
      RECT 9.21 5.06 9.215 5.232 ;
      RECT 9.185 5.07 9.21 5.239 ;
      RECT 9.175 5.084 9.185 5.248 ;
      RECT 9.155 5.096 9.175 5.251 ;
      RECT 9.105 5.115 9.155 5.255 ;
      RECT 9.06 5.13 9.105 5.26 ;
      RECT 8.995 5.133 9.06 5.266 ;
      RECT 8.98 5.131 8.995 5.273 ;
      RECT 8.95 5.13 8.98 5.273 ;
      RECT 8.911 5.129 8.95 5.269 ;
      RECT 8.825 5.126 8.911 5.265 ;
      RECT 8.808 5.124 8.825 5.262 ;
      RECT 8.722 5.122 8.808 5.259 ;
      RECT 8.636 5.119 8.722 5.253 ;
      RECT 8.55 5.115 8.636 5.248 ;
      RECT 8.472 5.112 8.55 5.244 ;
      RECT 8.386 5.109 8.472 5.242 ;
      RECT 8.3 5.106 8.386 5.239 ;
      RECT 8.242 5.104 8.3 5.236 ;
      RECT 8.156 5.101 8.242 5.234 ;
      RECT 8.07 5.097 8.156 5.232 ;
      RECT 7.984 5.094 8.07 5.229 ;
      RECT 7.898 5.09 7.984 5.227 ;
      RECT 7.812 5.086 7.898 5.224 ;
      RECT 7.726 5.083 7.812 5.222 ;
      RECT 7.64 5.079 7.726 5.219 ;
      RECT 7.554 5.076 7.64 5.217 ;
      RECT 7.468 5.072 7.554 5.214 ;
      RECT 7.382 5.069 7.468 5.212 ;
      RECT 7.296 5.065 7.382 5.209 ;
      RECT 7.21 5.062 7.296 5.207 ;
      RECT 7.2 5.06 7.21 5.203 ;
      RECT 7.195 5.06 7.2 5.201 ;
      RECT 7.155 5.055 7.195 5.195 ;
      RECT 7.141 5.046 7.155 5.188 ;
      RECT 7.055 5.016 7.141 5.173 ;
      RECT 7.035 4.982 7.055 5.158 ;
      RECT 6.965 4.951 7.035 5.145 ;
      RECT 6.96 4.926 6.965 5.134 ;
      RECT 6.955 4.92 6.96 5.132 ;
      RECT 6.886 4.765 6.955 5.12 ;
      RECT 6.8 4.765 6.886 5.094 ;
      RECT 6.775 4.765 6.8 5.073 ;
      RECT 6.77 4.765 6.775 5.063 ;
      RECT 6.765 4.765 6.77 5.055 ;
      RECT 6.745 4.765 6.765 5.038 ;
      RECT 9.165 3.335 9.425 3.595 ;
      RECT 9.15 3.335 9.425 3.498 ;
      RECT 9.12 3.335 9.425 3.473 ;
      RECT 9.085 3.175 9.365 3.455 ;
      RECT 9.055 4.665 9.115 4.925 ;
      RECT 8.08 3.355 8.135 3.615 ;
      RECT 9.015 4.622 9.055 4.925 ;
      RECT 8.986 4.543 9.015 4.925 ;
      RECT 8.9 4.415 8.986 4.925 ;
      RECT 8.88 4.295 8.9 4.925 ;
      RECT 8.855 4.246 8.88 4.925 ;
      RECT 8.85 4.211 8.855 4.775 ;
      RECT 8.82 4.171 8.85 4.713 ;
      RECT 8.795 4.108 8.82 4.628 ;
      RECT 8.785 4.07 8.795 4.565 ;
      RECT 8.77 4.045 8.785 4.526 ;
      RECT 8.727 4.003 8.77 4.432 ;
      RECT 8.725 3.976 8.727 4.359 ;
      RECT 8.72 3.971 8.725 4.35 ;
      RECT 8.715 3.964 8.72 4.325 ;
      RECT 8.71 3.958 8.715 4.31 ;
      RECT 8.705 3.952 8.71 4.298 ;
      RECT 8.695 3.943 8.705 4.28 ;
      RECT 8.69 3.934 8.695 4.258 ;
      RECT 8.665 3.915 8.69 4.208 ;
      RECT 8.66 3.896 8.665 4.158 ;
      RECT 8.645 3.882 8.66 4.118 ;
      RECT 8.64 3.868 8.645 4.085 ;
      RECT 8.635 3.861 8.64 4.078 ;
      RECT 8.62 3.848 8.635 4.07 ;
      RECT 8.575 3.81 8.62 4.043 ;
      RECT 8.545 3.763 8.575 4.008 ;
      RECT 8.525 3.732 8.545 3.985 ;
      RECT 8.445 3.665 8.525 3.938 ;
      RECT 8.415 3.595 8.445 3.885 ;
      RECT 8.41 3.572 8.415 3.868 ;
      RECT 8.38 3.55 8.41 3.853 ;
      RECT 8.35 3.509 8.38 3.825 ;
      RECT 8.345 3.484 8.35 3.81 ;
      RECT 8.34 3.478 8.345 3.803 ;
      RECT 8.33 3.355 8.34 3.795 ;
      RECT 8.32 3.355 8.33 3.788 ;
      RECT 8.315 3.355 8.32 3.78 ;
      RECT 8.295 3.355 8.315 3.768 ;
      RECT 8.245 3.355 8.295 3.738 ;
      RECT 8.19 3.355 8.245 3.688 ;
      RECT 8.16 3.355 8.19 3.648 ;
      RECT 8.135 3.355 8.16 3.625 ;
      RECT 8.005 4.08 8.285 4.36 ;
      RECT 7.97 3.995 8.23 4.255 ;
      RECT 7.97 4.077 8.24 4.255 ;
      RECT 6.17 3.45 6.175 3.935 ;
      RECT 6.06 3.635 6.065 3.935 ;
      RECT 5.97 3.675 6.035 3.935 ;
      RECT 7.645 3.175 7.735 3.805 ;
      RECT 7.61 3.225 7.615 3.805 ;
      RECT 7.555 3.25 7.565 3.805 ;
      RECT 7.51 3.25 7.52 3.805 ;
      RECT 7.88 3.175 7.925 3.455 ;
      RECT 6.73 2.905 6.93 3.045 ;
      RECT 7.846 3.175 7.88 3.467 ;
      RECT 7.76 3.175 7.846 3.507 ;
      RECT 7.745 3.175 7.76 3.548 ;
      RECT 7.74 3.175 7.745 3.568 ;
      RECT 7.735 3.175 7.74 3.588 ;
      RECT 7.615 3.217 7.645 3.805 ;
      RECT 7.565 3.237 7.61 3.805 ;
      RECT 7.55 3.252 7.555 3.805 ;
      RECT 7.52 3.252 7.55 3.805 ;
      RECT 7.475 3.237 7.51 3.805 ;
      RECT 7.47 3.225 7.475 3.585 ;
      RECT 7.465 3.222 7.47 3.565 ;
      RECT 7.45 3.212 7.465 3.518 ;
      RECT 7.445 3.205 7.45 3.481 ;
      RECT 7.44 3.202 7.445 3.464 ;
      RECT 7.425 3.192 7.44 3.42 ;
      RECT 7.42 3.183 7.425 3.38 ;
      RECT 7.415 3.179 7.42 3.365 ;
      RECT 7.405 3.173 7.415 3.348 ;
      RECT 7.365 3.154 7.405 3.323 ;
      RECT 7.36 3.136 7.365 3.303 ;
      RECT 7.35 3.13 7.36 3.298 ;
      RECT 7.32 3.114 7.35 3.285 ;
      RECT 7.305 3.096 7.32 3.268 ;
      RECT 7.29 3.084 7.305 3.255 ;
      RECT 7.285 3.076 7.29 3.248 ;
      RECT 7.255 3.062 7.285 3.235 ;
      RECT 7.25 3.047 7.255 3.223 ;
      RECT 7.24 3.041 7.25 3.215 ;
      RECT 7.22 3.029 7.24 3.203 ;
      RECT 7.21 3.017 7.22 3.19 ;
      RECT 7.18 3.001 7.21 3.175 ;
      RECT 7.16 2.981 7.18 3.158 ;
      RECT 7.155 2.971 7.16 3.148 ;
      RECT 7.13 2.959 7.155 3.135 ;
      RECT 7.125 2.947 7.13 3.123 ;
      RECT 7.12 2.942 7.125 3.119 ;
      RECT 7.105 2.935 7.12 3.111 ;
      RECT 7.095 2.922 7.105 3.101 ;
      RECT 7.09 2.92 7.095 3.095 ;
      RECT 7.065 2.913 7.09 3.084 ;
      RECT 7.06 2.906 7.065 3.073 ;
      RECT 7.035 2.905 7.06 3.06 ;
      RECT 7.016 2.905 7.035 3.05 ;
      RECT 6.93 2.905 7.016 3.047 ;
      RECT 6.7 2.905 6.73 3.05 ;
      RECT 6.66 2.912 6.7 3.063 ;
      RECT 6.635 2.922 6.66 3.076 ;
      RECT 6.62 2.931 6.635 3.086 ;
      RECT 6.59 2.936 6.62 3.105 ;
      RECT 6.585 2.942 6.59 3.123 ;
      RECT 6.565 2.952 6.585 3.138 ;
      RECT 6.555 2.965 6.565 3.158 ;
      RECT 6.54 2.977 6.555 3.175 ;
      RECT 6.535 2.987 6.54 3.185 ;
      RECT 6.53 2.992 6.535 3.19 ;
      RECT 6.52 3 6.53 3.203 ;
      RECT 6.47 3.032 6.52 3.24 ;
      RECT 6.455 3.067 6.47 3.281 ;
      RECT 6.45 3.077 6.455 3.296 ;
      RECT 6.445 3.082 6.45 3.303 ;
      RECT 6.42 3.098 6.445 3.323 ;
      RECT 6.405 3.119 6.42 3.348 ;
      RECT 6.38 3.14 6.405 3.373 ;
      RECT 6.37 3.159 6.38 3.396 ;
      RECT 6.345 3.177 6.37 3.419 ;
      RECT 6.33 3.197 6.345 3.443 ;
      RECT 6.325 3.207 6.33 3.455 ;
      RECT 6.31 3.219 6.325 3.475 ;
      RECT 6.3 3.234 6.31 3.515 ;
      RECT 6.295 3.242 6.3 3.543 ;
      RECT 6.285 3.252 6.295 3.563 ;
      RECT 6.28 3.265 6.285 3.588 ;
      RECT 6.275 3.278 6.28 3.608 ;
      RECT 6.27 3.284 6.275 3.63 ;
      RECT 6.26 3.293 6.27 3.65 ;
      RECT 6.255 3.313 6.26 3.673 ;
      RECT 6.25 3.319 6.255 3.693 ;
      RECT 6.245 3.326 6.25 3.715 ;
      RECT 6.24 3.337 6.245 3.728 ;
      RECT 6.23 3.347 6.24 3.753 ;
      RECT 6.21 3.372 6.23 3.935 ;
      RECT 6.18 3.412 6.21 3.935 ;
      RECT 6.175 3.442 6.18 3.935 ;
      RECT 6.15 3.47 6.17 3.935 ;
      RECT 6.12 3.515 6.15 3.935 ;
      RECT 6.115 3.542 6.12 3.935 ;
      RECT 6.095 3.56 6.115 3.935 ;
      RECT 6.085 3.585 6.095 3.935 ;
      RECT 6.08 3.597 6.085 3.935 ;
      RECT 6.065 3.62 6.08 3.935 ;
      RECT 6.045 3.647 6.06 3.935 ;
      RECT 6.035 3.67 6.045 3.935 ;
      RECT 7.825 4.555 7.905 4.815 ;
      RECT 7.06 3.775 7.13 4.035 ;
      RECT 7.791 4.522 7.825 4.815 ;
      RECT 7.705 4.425 7.791 4.815 ;
      RECT 7.685 4.337 7.705 4.815 ;
      RECT 7.675 4.307 7.685 4.815 ;
      RECT 7.665 4.287 7.675 4.815 ;
      RECT 7.645 4.274 7.665 4.815 ;
      RECT 7.63 4.264 7.645 4.643 ;
      RECT 7.625 4.257 7.63 4.598 ;
      RECT 7.615 4.251 7.625 4.588 ;
      RECT 7.605 4.243 7.615 4.57 ;
      RECT 7.6 4.237 7.605 4.558 ;
      RECT 7.59 4.232 7.6 4.545 ;
      RECT 7.57 4.222 7.59 4.518 ;
      RECT 7.53 4.201 7.57 4.47 ;
      RECT 7.515 4.182 7.53 4.428 ;
      RECT 7.49 4.168 7.515 4.398 ;
      RECT 7.48 4.156 7.49 4.365 ;
      RECT 7.475 4.151 7.48 4.355 ;
      RECT 7.445 4.137 7.475 4.335 ;
      RECT 7.435 4.121 7.445 4.308 ;
      RECT 7.43 4.116 7.435 4.298 ;
      RECT 7.405 4.107 7.43 4.278 ;
      RECT 7.395 4.095 7.405 4.258 ;
      RECT 7.325 4.063 7.395 4.233 ;
      RECT 7.32 4.032 7.325 4.21 ;
      RECT 7.271 3.775 7.32 4.193 ;
      RECT 7.185 3.775 7.271 4.152 ;
      RECT 7.13 3.775 7.185 4.08 ;
      RECT 7.22 4.56 7.38 4.82 ;
      RECT 6.745 3.175 6.795 3.86 ;
      RECT 6.535 3.6 6.57 3.86 ;
      RECT 6.85 3.175 6.855 3.635 ;
      RECT 6.94 3.175 6.965 3.455 ;
      RECT 7.215 4.557 7.22 4.82 ;
      RECT 7.18 4.545 7.215 4.82 ;
      RECT 7.12 4.518 7.18 4.82 ;
      RECT 7.115 4.501 7.12 4.674 ;
      RECT 7.11 4.498 7.115 4.661 ;
      RECT 7.09 4.491 7.11 4.648 ;
      RECT 7.055 4.474 7.09 4.63 ;
      RECT 7.015 4.453 7.055 4.61 ;
      RECT 7.01 4.441 7.015 4.598 ;
      RECT 6.97 4.427 7.01 4.584 ;
      RECT 6.95 4.41 6.97 4.566 ;
      RECT 6.94 4.402 6.95 4.558 ;
      RECT 6.925 3.175 6.94 3.473 ;
      RECT 6.91 4.392 6.94 4.545 ;
      RECT 6.895 3.175 6.925 3.518 ;
      RECT 6.9 4.382 6.91 4.532 ;
      RECT 6.87 4.367 6.9 4.519 ;
      RECT 6.855 3.175 6.895 3.585 ;
      RECT 6.855 4.335 6.87 4.505 ;
      RECT 6.85 4.307 6.855 4.499 ;
      RECT 6.845 3.175 6.85 3.64 ;
      RECT 6.835 4.277 6.85 4.493 ;
      RECT 6.84 3.175 6.845 3.653 ;
      RECT 6.83 3.175 6.84 3.673 ;
      RECT 6.795 4.19 6.835 4.478 ;
      RECT 6.795 3.175 6.83 3.713 ;
      RECT 6.79 4.122 6.795 4.466 ;
      RECT 6.775 4.077 6.79 4.461 ;
      RECT 6.77 4.015 6.775 4.456 ;
      RECT 6.745 3.922 6.77 4.449 ;
      RECT 6.74 3.175 6.745 4.441 ;
      RECT 6.725 3.175 6.74 4.428 ;
      RECT 6.705 3.175 6.725 4.385 ;
      RECT 6.695 3.175 6.705 4.335 ;
      RECT 6.69 3.175 6.695 4.308 ;
      RECT 6.685 3.175 6.69 4.286 ;
      RECT 6.68 3.401 6.685 4.269 ;
      RECT 6.675 3.423 6.68 4.247 ;
      RECT 6.67 3.465 6.675 4.23 ;
      RECT 6.64 3.515 6.67 4.174 ;
      RECT 6.635 3.542 6.64 4.116 ;
      RECT 6.62 3.56 6.635 4.08 ;
      RECT 6.615 3.578 6.62 4.044 ;
      RECT 6.609 3.585 6.615 4.025 ;
      RECT 6.605 3.592 6.609 4.008 ;
      RECT 6.6 3.597 6.605 3.977 ;
      RECT 6.59 3.6 6.6 3.952 ;
      RECT 6.58 3.6 6.59 3.918 ;
      RECT 6.575 3.6 6.58 3.895 ;
      RECT 6.57 3.6 6.575 3.875 ;
      RECT 5.485 3.735 5.765 4.015 ;
      RECT 5.485 3.735 5.785 3.91 ;
      RECT 5.575 3.625 5.835 3.885 ;
      RECT 5.54 3.72 5.835 3.885 ;
      RECT 5.665 2.24 5.83 3.885 ;
      RECT 5.565 2.24 5.935 2.61 ;
      RECT 5.19 4.765 5.45 5.025 ;
      RECT 5.21 4.692 5.39 5.025 ;
      RECT 5.21 4.435 5.385 5.025 ;
      RECT 5.21 4.227 5.375 5.025 ;
      RECT 5.215 4.145 5.375 5.025 ;
      RECT 5.215 3.91 5.365 5.025 ;
      RECT 5.215 3.757 5.36 5.025 ;
      RECT 5.22 3.742 5.36 5.025 ;
      RECT 5.27 3.457 5.36 5.025 ;
      RECT 5.225 3.692 5.36 5.025 ;
      RECT 5.255 3.51 5.36 5.025 ;
      RECT 5.24 3.622 5.36 5.025 ;
      RECT 5.245 3.58 5.36 5.025 ;
      RECT 5.24 3.622 5.375 3.685 ;
      RECT 5.275 3.21 5.38 3.63 ;
      RECT 5.275 3.21 5.395 3.613 ;
      RECT 5.275 3.21 5.43 3.575 ;
      RECT 5.27 3.457 5.48 3.508 ;
      RECT 5.275 3.21 5.535 3.47 ;
      RECT 4.535 3.915 4.795 4.175 ;
      RECT 4.535 3.915 4.805 4.133 ;
      RECT 4.535 3.915 4.891 4.104 ;
      RECT 4.535 3.915 4.96 4.056 ;
      RECT 4.535 3.915 4.995 4.025 ;
      RECT 4.765 3.735 5.045 4.015 ;
      RECT 4.6 3.9 5.045 4.015 ;
      RECT 4.69 3.777 4.795 4.175 ;
      RECT 4.62 3.84 5.045 4.015 ;
      RECT 70.04 9.345 70.41 9.715 ;
      RECT 54.78 9.345 55.15 9.715 ;
      RECT 39.52 9.345 39.89 9.715 ;
      RECT 24.26 9.345 24.63 9.715 ;
      RECT 9 9.345 9.37 9.715 ;
    LAYER via1 ;
      RECT 78.63 9.665 78.78 9.815 ;
      RECT 76.26 9.03 76.41 9.18 ;
      RECT 76.245 3.36 76.395 3.51 ;
      RECT 75.455 3.745 75.605 3.895 ;
      RECT 75.455 8.615 75.605 8.765 ;
      RECT 73.865 4.1 74.015 4.25 ;
      RECT 72.095 3.645 72.245 3.795 ;
      RECT 71.075 4.35 71.225 4.5 ;
      RECT 70.845 3.77 70.995 3.92 ;
      RECT 70.81 9 70.96 9.15 ;
      RECT 70.5 4.37 70.65 4.52 ;
      RECT 70.26 3.39 70.41 3.54 ;
      RECT 70.15 9.455 70.3 9.605 ;
      RECT 69.95 4.72 70.1 4.87 ;
      RECT 69.81 3.325 69.96 3.475 ;
      RECT 69.175 3.41 69.325 3.56 ;
      RECT 69.065 4.05 69.215 4.2 ;
      RECT 68.74 4.61 68.89 4.76 ;
      RECT 68.57 3.6 68.72 3.75 ;
      RECT 68.215 4.615 68.365 4.765 ;
      RECT 68.155 3.83 68.305 3.98 ;
      RECT 67.79 4.82 67.94 4.97 ;
      RECT 67.63 3.655 67.78 3.805 ;
      RECT 67.065 3.73 67.215 3.88 ;
      RECT 66.715 2.35 66.865 2.5 ;
      RECT 66.67 3.68 66.82 3.83 ;
      RECT 66.37 3.265 66.52 3.415 ;
      RECT 66.285 4.82 66.435 4.97 ;
      RECT 65.63 3.97 65.78 4.12 ;
      RECT 63.345 9.045 63.495 9.195 ;
      RECT 61 9.03 61.15 9.18 ;
      RECT 60.985 3.36 61.135 3.51 ;
      RECT 60.195 3.745 60.345 3.895 ;
      RECT 60.195 8.615 60.345 8.765 ;
      RECT 58.605 4.1 58.755 4.25 ;
      RECT 56.835 3.645 56.985 3.795 ;
      RECT 55.815 4.35 55.965 4.5 ;
      RECT 55.585 3.77 55.735 3.92 ;
      RECT 55.55 9 55.7 9.15 ;
      RECT 55.24 4.37 55.39 4.52 ;
      RECT 55 3.39 55.15 3.54 ;
      RECT 54.89 9.455 55.04 9.605 ;
      RECT 54.69 4.72 54.84 4.87 ;
      RECT 54.55 3.325 54.7 3.475 ;
      RECT 53.915 3.41 54.065 3.56 ;
      RECT 53.805 4.05 53.955 4.2 ;
      RECT 53.48 4.61 53.63 4.76 ;
      RECT 53.31 3.6 53.46 3.75 ;
      RECT 52.955 4.615 53.105 4.765 ;
      RECT 52.895 3.83 53.045 3.98 ;
      RECT 52.53 4.82 52.68 4.97 ;
      RECT 52.37 3.655 52.52 3.805 ;
      RECT 51.805 3.73 51.955 3.88 ;
      RECT 51.455 2.35 51.605 2.5 ;
      RECT 51.41 3.68 51.56 3.83 ;
      RECT 51.11 3.265 51.26 3.415 ;
      RECT 51.025 4.82 51.175 4.97 ;
      RECT 50.37 3.97 50.52 4.12 ;
      RECT 48.085 9.045 48.235 9.195 ;
      RECT 45.74 9.03 45.89 9.18 ;
      RECT 45.725 3.36 45.875 3.51 ;
      RECT 44.935 3.745 45.085 3.895 ;
      RECT 44.935 8.615 45.085 8.765 ;
      RECT 43.345 4.1 43.495 4.25 ;
      RECT 41.575 3.645 41.725 3.795 ;
      RECT 40.555 4.35 40.705 4.5 ;
      RECT 40.325 3.77 40.475 3.92 ;
      RECT 40.29 9.005 40.44 9.155 ;
      RECT 39.98 4.37 40.13 4.52 ;
      RECT 39.74 3.39 39.89 3.54 ;
      RECT 39.63 9.455 39.78 9.605 ;
      RECT 39.43 4.72 39.58 4.87 ;
      RECT 39.29 3.325 39.44 3.475 ;
      RECT 38.655 3.41 38.805 3.56 ;
      RECT 38.545 4.05 38.695 4.2 ;
      RECT 38.22 4.61 38.37 4.76 ;
      RECT 38.05 3.6 38.2 3.75 ;
      RECT 37.695 4.615 37.845 4.765 ;
      RECT 37.635 3.83 37.785 3.98 ;
      RECT 37.27 4.82 37.42 4.97 ;
      RECT 37.11 3.655 37.26 3.805 ;
      RECT 36.545 3.73 36.695 3.88 ;
      RECT 36.195 2.35 36.345 2.5 ;
      RECT 36.15 3.68 36.3 3.83 ;
      RECT 35.85 3.265 36 3.415 ;
      RECT 35.765 4.82 35.915 4.97 ;
      RECT 35.11 3.97 35.26 4.12 ;
      RECT 32.87 9.05 33.02 9.2 ;
      RECT 30.48 9.03 30.63 9.18 ;
      RECT 30.465 3.36 30.615 3.51 ;
      RECT 29.675 3.745 29.825 3.895 ;
      RECT 29.675 8.615 29.825 8.765 ;
      RECT 28.085 4.1 28.235 4.25 ;
      RECT 26.315 3.645 26.465 3.795 ;
      RECT 25.295 4.35 25.445 4.5 ;
      RECT 25.065 3.77 25.215 3.92 ;
      RECT 25.03 9 25.18 9.15 ;
      RECT 24.72 4.37 24.87 4.52 ;
      RECT 24.48 3.39 24.63 3.54 ;
      RECT 24.37 9.455 24.52 9.605 ;
      RECT 24.17 4.72 24.32 4.87 ;
      RECT 24.03 3.325 24.18 3.475 ;
      RECT 23.395 3.41 23.545 3.56 ;
      RECT 23.285 4.05 23.435 4.2 ;
      RECT 22.96 4.61 23.11 4.76 ;
      RECT 22.79 3.6 22.94 3.75 ;
      RECT 22.435 4.615 22.585 4.765 ;
      RECT 22.375 3.83 22.525 3.98 ;
      RECT 22.01 4.82 22.16 4.97 ;
      RECT 21.85 3.655 22 3.805 ;
      RECT 21.285 3.73 21.435 3.88 ;
      RECT 20.935 2.35 21.085 2.5 ;
      RECT 20.89 3.68 21.04 3.83 ;
      RECT 20.59 3.265 20.74 3.415 ;
      RECT 20.505 4.82 20.655 4.97 ;
      RECT 19.85 3.97 20 4.12 ;
      RECT 17.61 9.045 17.76 9.195 ;
      RECT 15.22 9.03 15.37 9.18 ;
      RECT 15.205 3.36 15.355 3.51 ;
      RECT 14.415 3.745 14.565 3.895 ;
      RECT 14.415 8.615 14.565 8.765 ;
      RECT 12.825 4.1 12.975 4.25 ;
      RECT 11.055 3.645 11.205 3.795 ;
      RECT 10.035 4.35 10.185 4.5 ;
      RECT 9.805 3.77 9.955 3.92 ;
      RECT 9.77 8.995 9.92 9.145 ;
      RECT 9.46 4.37 9.61 4.52 ;
      RECT 9.22 3.39 9.37 3.54 ;
      RECT 9.11 9.455 9.26 9.605 ;
      RECT 8.91 4.72 9.06 4.87 ;
      RECT 8.77 3.325 8.92 3.475 ;
      RECT 8.135 3.41 8.285 3.56 ;
      RECT 8.025 4.05 8.175 4.2 ;
      RECT 7.7 4.61 7.85 4.76 ;
      RECT 7.53 3.6 7.68 3.75 ;
      RECT 7.175 4.615 7.325 4.765 ;
      RECT 7.115 3.83 7.265 3.98 ;
      RECT 6.75 4.82 6.9 4.97 ;
      RECT 6.59 3.655 6.74 3.805 ;
      RECT 6.025 3.73 6.175 3.88 ;
      RECT 5.675 2.35 5.825 2.5 ;
      RECT 5.63 3.68 5.78 3.83 ;
      RECT 5.33 3.265 5.48 3.415 ;
      RECT 5.245 4.82 5.395 4.97 ;
      RECT 4.59 3.97 4.74 4.12 ;
      RECT 1.615 9.385 1.765 9.535 ;
      RECT 1.24 8.645 1.39 8.795 ;
    LAYER met1 ;
      RECT 76.965 5.425 78.945 7.04 ;
      RECT 61.705 5.425 63.685 7.04 ;
      RECT 46.445 5.425 48.425 7.04 ;
      RECT 31.185 5.425 33.165 7.04 ;
      RECT 15.925 5.425 17.905 7.04 ;
      RECT 74.22 5.43 78.945 7.035 ;
      RECT 72.26 5.275 73.14 7.035 ;
      RECT 71.405 5.275 71.625 7.035 ;
      RECT 68.585 5.275 71.335 7.035 ;
      RECT 58.96 5.43 63.685 7.035 ;
      RECT 57 5.275 57.88 7.035 ;
      RECT 56.145 5.275 56.365 7.035 ;
      RECT 53.325 5.275 56.075 7.035 ;
      RECT 43.7 5.43 48.425 7.035 ;
      RECT 41.74 5.275 42.62 7.035 ;
      RECT 40.885 5.275 41.105 7.035 ;
      RECT 38.065 5.275 40.815 7.035 ;
      RECT 28.44 5.43 33.165 7.035 ;
      RECT 26.48 5.275 27.36 7.035 ;
      RECT 25.625 5.275 25.845 7.035 ;
      RECT 22.805 5.275 25.555 7.035 ;
      RECT 13.18 5.43 17.905 7.035 ;
      RECT 11.22 5.275 12.1 7.035 ;
      RECT 10.365 5.275 10.585 7.035 ;
      RECT 7.545 5.275 10.295 7.035 ;
      RECT 0 5.435 3.695 7.035 ;
      RECT 2.805 5.43 79.105 7.03 ;
      RECT 64.59 5.275 73.33 7.03 ;
      RECT 49.33 5.275 58.07 7.03 ;
      RECT 34.07 5.275 42.81 7.03 ;
      RECT 18.81 5.275 27.55 7.03 ;
      RECT 3.55 5.275 12.29 7.03 ;
      RECT 64.59 0 73.33 3.035 ;
      RECT 49.33 0 58.07 3.035 ;
      RECT 34.07 0 42.81 3.035 ;
      RECT 18.81 0 27.55 3.035 ;
      RECT 3.55 0 12.29 3.035 ;
      RECT 0.005 0 79.1 1.6 ;
      RECT 0.005 10.865 79.1 12.465 ;
      RECT 69.535 8.605 69.705 12.465 ;
      RECT 54.275 8.605 54.445 12.465 ;
      RECT 39.015 8.605 39.185 12.465 ;
      RECT 23.755 8.605 23.925 12.465 ;
      RECT 8.495 8.605 8.665 12.465 ;
      RECT 69.705 8.575 69.995 8.805 ;
      RECT 54.445 8.575 54.735 8.805 ;
      RECT 39.185 8.575 39.475 8.805 ;
      RECT 23.925 8.575 24.215 8.805 ;
      RECT 8.665 8.575 8.955 8.805 ;
      RECT 78.495 10.06 78.785 10.29 ;
      RECT 78.555 8.58 78.725 10.29 ;
      RECT 78.53 9.565 78.88 9.915 ;
      RECT 78.495 8.58 78.785 8.81 ;
      RECT 78.09 3.69 78.195 4.26 ;
      RECT 78.09 4.025 78.415 4.255 ;
      RECT 78.09 4.055 78.585 4.225 ;
      RECT 78.09 3.69 78.28 4.255 ;
      RECT 77.505 3.655 77.795 3.885 ;
      RECT 77.505 3.69 78.28 3.86 ;
      RECT 77.565 2.175 77.735 3.885 ;
      RECT 77.505 2.175 77.795 2.405 ;
      RECT 77.505 10.06 77.795 10.29 ;
      RECT 77.565 8.58 77.735 10.29 ;
      RECT 77.505 8.58 77.795 8.81 ;
      RECT 77.505 8.615 78.355 8.775 ;
      RECT 78.19 8.21 78.355 8.775 ;
      RECT 77.505 8.61 77.9 8.775 ;
      RECT 78.125 8.21 78.415 8.44 ;
      RECT 78.125 8.24 78.585 8.41 ;
      RECT 77.135 4.025 77.425 4.255 ;
      RECT 77.135 4.055 77.595 4.225 ;
      RECT 77.2 2.95 77.365 4.255 ;
      RECT 75.715 2.92 76.005 3.15 ;
      RECT 75.715 2.95 77.365 3.12 ;
      RECT 75.775 2.18 75.945 3.15 ;
      RECT 75.715 2.18 76.005 2.41 ;
      RECT 75.715 10.055 76.005 10.285 ;
      RECT 75.775 9.315 75.945 10.285 ;
      RECT 75.775 9.41 77.365 9.58 ;
      RECT 77.195 8.21 77.365 9.58 ;
      RECT 75.715 9.315 76.005 9.545 ;
      RECT 77.135 8.21 77.425 8.44 ;
      RECT 77.135 8.24 77.595 8.41 ;
      RECT 73.765 4 74.105 4.35 ;
      RECT 73.855 3.32 74.025 4.35 ;
      RECT 76.145 3.26 76.495 3.61 ;
      RECT 73.855 3.32 76.495 3.49 ;
      RECT 76.17 8.945 76.495 9.27 ;
      RECT 70.71 8.9 71.06 9.25 ;
      RECT 76.145 8.945 76.495 9.175 ;
      RECT 70.51 8.945 71.06 9.175 ;
      RECT 70.34 8.975 76.495 9.145 ;
      RECT 75.37 3.66 75.69 3.98 ;
      RECT 75.34 3.66 75.69 3.89 ;
      RECT 75.17 3.69 75.69 3.86 ;
      RECT 75.37 8.545 75.69 8.835 ;
      RECT 75.34 8.575 75.69 8.805 ;
      RECT 75.17 8.605 75.69 8.775 ;
      RECT 71.06 4.28 71.21 4.555 ;
      RECT 71.6 3.36 71.605 3.58 ;
      RECT 72.75 3.56 72.765 3.758 ;
      RECT 72.715 3.552 72.75 3.765 ;
      RECT 72.685 3.545 72.715 3.765 ;
      RECT 72.63 3.51 72.685 3.765 ;
      RECT 72.565 3.447 72.63 3.765 ;
      RECT 72.56 3.412 72.565 3.763 ;
      RECT 72.555 3.407 72.56 3.755 ;
      RECT 72.55 3.402 72.555 3.741 ;
      RECT 72.545 3.399 72.55 3.734 ;
      RECT 72.5 3.389 72.545 3.685 ;
      RECT 72.48 3.376 72.5 3.62 ;
      RECT 72.475 3.371 72.48 3.593 ;
      RECT 72.47 3.37 72.475 3.586 ;
      RECT 72.465 3.369 72.47 3.579 ;
      RECT 72.38 3.354 72.465 3.525 ;
      RECT 72.35 3.335 72.38 3.475 ;
      RECT 72.27 3.318 72.35 3.46 ;
      RECT 72.235 3.305 72.27 3.445 ;
      RECT 72.227 3.305 72.235 3.44 ;
      RECT 72.141 3.306 72.227 3.44 ;
      RECT 72.055 3.308 72.141 3.44 ;
      RECT 72.03 3.309 72.055 3.444 ;
      RECT 71.955 3.315 72.03 3.459 ;
      RECT 71.872 3.327 71.955 3.483 ;
      RECT 71.786 3.34 71.872 3.509 ;
      RECT 71.7 3.353 71.786 3.535 ;
      RECT 71.665 3.362 71.7 3.554 ;
      RECT 71.615 3.362 71.665 3.567 ;
      RECT 71.605 3.36 71.615 3.578 ;
      RECT 71.59 3.357 71.6 3.58 ;
      RECT 71.575 3.349 71.59 3.588 ;
      RECT 71.56 3.341 71.575 3.608 ;
      RECT 71.555 3.336 71.56 3.665 ;
      RECT 71.54 3.331 71.555 3.738 ;
      RECT 71.535 3.326 71.54 3.78 ;
      RECT 71.53 3.324 71.535 3.808 ;
      RECT 71.525 3.322 71.53 3.83 ;
      RECT 71.515 3.318 71.525 3.873 ;
      RECT 71.51 3.315 71.515 3.898 ;
      RECT 71.505 3.313 71.51 3.918 ;
      RECT 71.5 3.311 71.505 3.942 ;
      RECT 71.495 3.307 71.5 3.965 ;
      RECT 71.49 3.303 71.495 3.988 ;
      RECT 71.455 3.293 71.49 4.095 ;
      RECT 71.45 3.283 71.455 4.193 ;
      RECT 71.445 3.281 71.45 4.22 ;
      RECT 71.44 3.28 71.445 4.24 ;
      RECT 71.435 3.272 71.44 4.26 ;
      RECT 71.43 3.267 71.435 4.295 ;
      RECT 71.425 3.265 71.43 4.313 ;
      RECT 71.42 3.265 71.425 4.338 ;
      RECT 71.415 3.265 71.42 4.36 ;
      RECT 71.38 3.265 71.415 4.403 ;
      RECT 71.355 3.265 71.38 4.432 ;
      RECT 71.345 3.265 71.355 3.618 ;
      RECT 71.348 3.675 71.355 4.442 ;
      RECT 71.345 3.732 71.348 4.445 ;
      RECT 71.34 3.265 71.345 3.59 ;
      RECT 71.34 3.782 71.345 4.448 ;
      RECT 71.33 3.265 71.34 3.58 ;
      RECT 71.335 3.835 71.34 4.451 ;
      RECT 71.33 3.92 71.335 4.455 ;
      RECT 71.32 3.265 71.33 3.568 ;
      RECT 71.325 3.967 71.33 4.459 ;
      RECT 71.32 4.042 71.325 4.463 ;
      RECT 71.285 3.265 71.32 3.543 ;
      RECT 71.31 4.125 71.32 4.468 ;
      RECT 71.3 4.192 71.31 4.475 ;
      RECT 71.295 4.22 71.3 4.48 ;
      RECT 71.285 4.233 71.295 4.486 ;
      RECT 71.24 3.265 71.285 3.5 ;
      RECT 71.28 4.238 71.285 4.493 ;
      RECT 71.24 4.255 71.28 4.555 ;
      RECT 71.235 3.267 71.24 3.473 ;
      RECT 71.21 4.275 71.24 4.555 ;
      RECT 71.23 3.272 71.235 3.445 ;
      RECT 71.02 4.284 71.06 4.555 ;
      RECT 70.995 4.292 71.02 4.525 ;
      RECT 70.95 4.3 70.995 4.525 ;
      RECT 70.935 4.305 70.95 4.52 ;
      RECT 70.925 4.305 70.935 4.514 ;
      RECT 70.915 4.312 70.925 4.511 ;
      RECT 70.91 4.35 70.915 4.5 ;
      RECT 70.905 4.412 70.91 4.478 ;
      RECT 72.175 4.287 72.36 4.51 ;
      RECT 72.175 4.302 72.365 4.506 ;
      RECT 72.165 3.575 72.25 4.505 ;
      RECT 72.165 4.302 72.37 4.499 ;
      RECT 72.16 4.31 72.37 4.498 ;
      RECT 72.365 4.03 72.685 4.35 ;
      RECT 72.16 4.202 72.33 4.293 ;
      RECT 72.155 4.202 72.33 4.275 ;
      RECT 72.145 4.01 72.28 4.25 ;
      RECT 72.14 4.01 72.28 4.195 ;
      RECT 72.1 3.59 72.27 4.095 ;
      RECT 72.085 3.59 72.27 3.965 ;
      RECT 72.08 3.59 72.27 3.918 ;
      RECT 72.075 3.59 72.27 3.898 ;
      RECT 72.07 3.59 72.27 3.873 ;
      RECT 72.04 3.59 72.3 3.85 ;
      RECT 72.05 3.587 72.26 3.85 ;
      RECT 72.175 3.582 72.26 4.51 ;
      RECT 72.06 3.575 72.25 3.85 ;
      RECT 72.055 3.58 72.25 3.85 ;
      RECT 70.885 3.792 71.07 4.005 ;
      RECT 70.885 3.8 71.08 3.998 ;
      RECT 70.865 3.8 71.08 3.995 ;
      RECT 70.86 3.8 71.08 3.98 ;
      RECT 70.79 3.715 71.05 3.975 ;
      RECT 70.79 3.86 71.085 3.888 ;
      RECT 70.445 4.315 70.705 4.575 ;
      RECT 70.47 4.26 70.665 4.575 ;
      RECT 70.465 4.009 70.645 4.303 ;
      RECT 70.465 4.015 70.655 4.303 ;
      RECT 70.445 4.017 70.655 4.248 ;
      RECT 70.44 4.027 70.655 4.115 ;
      RECT 70.47 4.007 70.645 4.575 ;
      RECT 70.556 4.005 70.645 4.575 ;
      RECT 70.415 3.225 70.45 3.595 ;
      RECT 70.205 3.335 70.21 3.595 ;
      RECT 70.45 3.232 70.465 3.595 ;
      RECT 70.34 3.225 70.415 3.673 ;
      RECT 70.33 3.225 70.34 3.758 ;
      RECT 70.305 3.225 70.33 3.793 ;
      RECT 70.265 3.225 70.305 3.861 ;
      RECT 70.255 3.232 70.265 3.913 ;
      RECT 70.225 3.335 70.255 3.954 ;
      RECT 70.22 3.335 70.225 3.993 ;
      RECT 70.21 3.335 70.22 4.013 ;
      RECT 70.205 3.63 70.21 4.05 ;
      RECT 70.2 3.647 70.205 4.07 ;
      RECT 70.185 3.71 70.2 4.11 ;
      RECT 70.18 3.753 70.185 4.145 ;
      RECT 70.175 3.761 70.18 4.158 ;
      RECT 70.165 3.775 70.175 4.18 ;
      RECT 70.14 3.81 70.165 4.245 ;
      RECT 70.13 3.845 70.14 4.308 ;
      RECT 70.11 3.875 70.13 4.369 ;
      RECT 70.095 3.911 70.11 4.436 ;
      RECT 70.085 3.939 70.095 4.475 ;
      RECT 70.075 3.961 70.085 4.495 ;
      RECT 70.07 3.971 70.075 4.506 ;
      RECT 70.065 3.98 70.07 4.509 ;
      RECT 70.055 3.998 70.065 4.513 ;
      RECT 70.045 4.016 70.055 4.514 ;
      RECT 70.02 4.055 70.045 4.511 ;
      RECT 70 4.097 70.02 4.508 ;
      RECT 69.985 4.135 70 4.507 ;
      RECT 69.95 4.17 69.985 4.504 ;
      RECT 69.945 4.192 69.95 4.502 ;
      RECT 69.88 4.232 69.945 4.499 ;
      RECT 69.875 4.272 69.88 4.495 ;
      RECT 69.86 4.282 69.875 4.486 ;
      RECT 69.85 4.402 69.86 4.471 ;
      RECT 70.33 4.815 70.34 5.075 ;
      RECT 70.33 4.818 70.35 5.074 ;
      RECT 70.32 4.808 70.33 5.073 ;
      RECT 70.31 4.823 70.39 5.069 ;
      RECT 70.295 4.802 70.31 5.067 ;
      RECT 70.27 4.827 70.395 5.063 ;
      RECT 70.255 4.787 70.27 5.058 ;
      RECT 70.255 4.829 70.405 5.057 ;
      RECT 70.255 4.837 70.42 5.05 ;
      RECT 70.195 4.774 70.255 5.04 ;
      RECT 70.185 4.761 70.195 5.022 ;
      RECT 70.16 4.751 70.185 5.012 ;
      RECT 70.155 4.741 70.16 5.004 ;
      RECT 70.09 4.837 70.42 4.986 ;
      RECT 70.005 4.837 70.42 4.948 ;
      RECT 69.895 4.665 70.155 4.925 ;
      RECT 70.27 4.795 70.295 5.063 ;
      RECT 70.31 4.805 70.32 5.069 ;
      RECT 69.895 4.813 70.335 4.925 ;
      RECT 70.08 10.055 70.37 10.285 ;
      RECT 70.14 9.315 70.31 10.285 ;
      RECT 70.04 9.345 70.41 9.715 ;
      RECT 70.08 9.315 70.37 9.715 ;
      RECT 69.11 4.57 69.14 4.87 ;
      RECT 68.885 4.555 68.89 4.83 ;
      RECT 68.685 4.555 68.84 4.815 ;
      RECT 69.985 3.27 70.015 3.53 ;
      RECT 69.975 3.27 69.985 3.638 ;
      RECT 69.955 3.27 69.975 3.648 ;
      RECT 69.94 3.27 69.955 3.66 ;
      RECT 69.885 3.27 69.94 3.71 ;
      RECT 69.87 3.27 69.885 3.758 ;
      RECT 69.84 3.27 69.87 3.793 ;
      RECT 69.785 3.27 69.84 3.855 ;
      RECT 69.765 3.27 69.785 3.923 ;
      RECT 69.76 3.27 69.765 3.953 ;
      RECT 69.755 3.27 69.76 3.965 ;
      RECT 69.75 3.387 69.755 3.983 ;
      RECT 69.73 3.405 69.75 4.008 ;
      RECT 69.71 3.432 69.73 4.058 ;
      RECT 69.705 3.452 69.71 4.089 ;
      RECT 69.7 3.46 69.705 4.106 ;
      RECT 69.685 3.486 69.7 4.135 ;
      RECT 69.67 3.528 69.685 4.17 ;
      RECT 69.665 3.557 69.67 4.193 ;
      RECT 69.66 3.572 69.665 4.206 ;
      RECT 69.655 3.595 69.66 4.217 ;
      RECT 69.645 3.615 69.655 4.235 ;
      RECT 69.635 3.645 69.645 4.258 ;
      RECT 69.63 3.667 69.635 4.278 ;
      RECT 69.625 3.682 69.63 4.293 ;
      RECT 69.61 3.712 69.625 4.32 ;
      RECT 69.605 3.742 69.61 4.346 ;
      RECT 69.6 3.76 69.605 4.358 ;
      RECT 69.59 3.79 69.6 4.377 ;
      RECT 69.58 3.815 69.59 4.402 ;
      RECT 69.575 3.835 69.58 4.421 ;
      RECT 69.57 3.852 69.575 4.434 ;
      RECT 69.56 3.878 69.57 4.453 ;
      RECT 69.55 3.916 69.56 4.48 ;
      RECT 69.545 3.942 69.55 4.5 ;
      RECT 69.54 3.952 69.545 4.51 ;
      RECT 69.535 3.965 69.54 4.525 ;
      RECT 69.53 3.98 69.535 4.535 ;
      RECT 69.525 4.002 69.53 4.55 ;
      RECT 69.52 4.02 69.525 4.561 ;
      RECT 69.515 4.03 69.52 4.572 ;
      RECT 69.51 4.038 69.515 4.584 ;
      RECT 69.505 4.046 69.51 4.595 ;
      RECT 69.5 4.072 69.505 4.608 ;
      RECT 69.49 4.1 69.5 4.621 ;
      RECT 69.485 4.13 69.49 4.63 ;
      RECT 69.48 4.145 69.485 4.637 ;
      RECT 69.465 4.17 69.48 4.644 ;
      RECT 69.46 4.192 69.465 4.65 ;
      RECT 69.455 4.217 69.46 4.653 ;
      RECT 69.446 4.245 69.455 4.657 ;
      RECT 69.44 4.262 69.446 4.662 ;
      RECT 69.435 4.28 69.44 4.666 ;
      RECT 69.43 4.292 69.435 4.669 ;
      RECT 69.425 4.313 69.43 4.673 ;
      RECT 69.42 4.331 69.425 4.676 ;
      RECT 69.415 4.345 69.42 4.679 ;
      RECT 69.41 4.362 69.415 4.682 ;
      RECT 69.405 4.375 69.41 4.685 ;
      RECT 69.38 4.412 69.405 4.693 ;
      RECT 69.375 4.457 69.38 4.702 ;
      RECT 69.37 4.485 69.375 4.705 ;
      RECT 69.36 4.505 69.37 4.709 ;
      RECT 69.355 4.525 69.36 4.714 ;
      RECT 69.35 4.54 69.355 4.717 ;
      RECT 69.33 4.55 69.35 4.724 ;
      RECT 69.265 4.557 69.33 4.75 ;
      RECT 69.23 4.56 69.265 4.778 ;
      RECT 69.215 4.563 69.23 4.793 ;
      RECT 69.205 4.564 69.215 4.808 ;
      RECT 69.195 4.565 69.205 4.825 ;
      RECT 69.19 4.565 69.195 4.84 ;
      RECT 69.185 4.565 69.19 4.848 ;
      RECT 69.17 4.566 69.185 4.863 ;
      RECT 69.14 4.568 69.17 4.87 ;
      RECT 69.03 4.575 69.11 4.87 ;
      RECT 68.985 4.58 69.03 4.87 ;
      RECT 68.975 4.581 68.985 4.86 ;
      RECT 68.965 4.582 68.975 4.853 ;
      RECT 68.945 4.584 68.965 4.848 ;
      RECT 68.935 4.555 68.945 4.843 ;
      RECT 68.89 4.555 68.935 4.835 ;
      RECT 68.86 4.555 68.885 4.825 ;
      RECT 68.84 4.555 68.86 4.818 ;
      RECT 69.12 3.355 69.38 3.615 ;
      RECT 69 3.37 69.01 3.535 ;
      RECT 68.985 3.37 68.99 3.53 ;
      RECT 66.35 3.21 66.535 3.5 ;
      RECT 68.165 3.335 68.18 3.49 ;
      RECT 66.315 3.21 66.34 3.47 ;
      RECT 68.73 3.26 68.735 3.402 ;
      RECT 68.645 3.255 68.67 3.395 ;
      RECT 69.045 3.372 69.12 3.565 ;
      RECT 69.03 3.37 69.045 3.548 ;
      RECT 69.01 3.37 69.03 3.54 ;
      RECT 68.99 3.37 69 3.533 ;
      RECT 68.945 3.365 68.985 3.523 ;
      RECT 68.905 3.34 68.945 3.508 ;
      RECT 68.89 3.315 68.905 3.498 ;
      RECT 68.885 3.309 68.89 3.496 ;
      RECT 68.85 3.301 68.885 3.479 ;
      RECT 68.845 3.294 68.85 3.467 ;
      RECT 68.825 3.289 68.845 3.455 ;
      RECT 68.815 3.283 68.825 3.44 ;
      RECT 68.795 3.278 68.815 3.425 ;
      RECT 68.785 3.273 68.795 3.418 ;
      RECT 68.78 3.271 68.785 3.413 ;
      RECT 68.775 3.27 68.78 3.41 ;
      RECT 68.735 3.265 68.775 3.406 ;
      RECT 68.715 3.259 68.73 3.401 ;
      RECT 68.68 3.256 68.715 3.398 ;
      RECT 68.67 3.255 68.68 3.396 ;
      RECT 68.61 3.255 68.645 3.393 ;
      RECT 68.565 3.255 68.61 3.393 ;
      RECT 68.515 3.255 68.565 3.396 ;
      RECT 68.5 3.257 68.515 3.398 ;
      RECT 68.485 3.26 68.5 3.399 ;
      RECT 68.475 3.265 68.485 3.4 ;
      RECT 68.445 3.27 68.475 3.405 ;
      RECT 68.435 3.276 68.445 3.413 ;
      RECT 68.425 3.278 68.435 3.417 ;
      RECT 68.415 3.282 68.425 3.421 ;
      RECT 68.39 3.288 68.415 3.429 ;
      RECT 68.38 3.293 68.39 3.437 ;
      RECT 68.365 3.297 68.38 3.441 ;
      RECT 68.33 3.303 68.365 3.449 ;
      RECT 68.31 3.308 68.33 3.459 ;
      RECT 68.28 3.315 68.31 3.468 ;
      RECT 68.235 3.324 68.28 3.482 ;
      RECT 68.23 3.329 68.235 3.493 ;
      RECT 68.21 3.332 68.23 3.494 ;
      RECT 68.18 3.335 68.21 3.492 ;
      RECT 68.145 3.335 68.165 3.488 ;
      RECT 68.075 3.335 68.145 3.479 ;
      RECT 68.06 3.332 68.075 3.471 ;
      RECT 68.02 3.325 68.06 3.466 ;
      RECT 67.995 3.315 68.02 3.459 ;
      RECT 67.99 3.309 67.995 3.456 ;
      RECT 67.95 3.303 67.99 3.453 ;
      RECT 67.935 3.296 67.95 3.448 ;
      RECT 67.915 3.292 67.935 3.443 ;
      RECT 67.9 3.287 67.915 3.439 ;
      RECT 67.885 3.282 67.9 3.437 ;
      RECT 67.87 3.278 67.885 3.436 ;
      RECT 67.855 3.276 67.87 3.432 ;
      RECT 67.845 3.274 67.855 3.427 ;
      RECT 67.83 3.271 67.845 3.423 ;
      RECT 67.82 3.269 67.83 3.418 ;
      RECT 67.8 3.266 67.82 3.414 ;
      RECT 67.755 3.265 67.8 3.412 ;
      RECT 67.695 3.267 67.755 3.413 ;
      RECT 67.675 3.269 67.695 3.415 ;
      RECT 67.645 3.272 67.675 3.416 ;
      RECT 67.595 3.277 67.645 3.418 ;
      RECT 67.59 3.28 67.595 3.42 ;
      RECT 67.58 3.282 67.59 3.423 ;
      RECT 67.575 3.284 67.58 3.426 ;
      RECT 67.525 3.287 67.575 3.433 ;
      RECT 67.505 3.291 67.525 3.445 ;
      RECT 67.495 3.294 67.505 3.451 ;
      RECT 67.485 3.295 67.495 3.454 ;
      RECT 67.446 3.298 67.485 3.456 ;
      RECT 67.36 3.305 67.446 3.459 ;
      RECT 67.286 3.315 67.36 3.463 ;
      RECT 67.2 3.326 67.286 3.468 ;
      RECT 67.185 3.333 67.2 3.47 ;
      RECT 67.13 3.337 67.185 3.471 ;
      RECT 67.116 3.34 67.13 3.473 ;
      RECT 67.03 3.34 67.116 3.475 ;
      RECT 66.99 3.337 67.03 3.478 ;
      RECT 66.966 3.333 66.99 3.48 ;
      RECT 66.88 3.323 66.966 3.483 ;
      RECT 66.85 3.312 66.88 3.484 ;
      RECT 66.831 3.308 66.85 3.483 ;
      RECT 66.745 3.301 66.831 3.48 ;
      RECT 66.685 3.29 66.745 3.477 ;
      RECT 66.665 3.282 66.685 3.475 ;
      RECT 66.63 3.277 66.665 3.474 ;
      RECT 66.605 3.272 66.63 3.473 ;
      RECT 66.575 3.267 66.605 3.472 ;
      RECT 66.55 3.21 66.575 3.471 ;
      RECT 66.535 3.21 66.55 3.495 ;
      RECT 66.34 3.21 66.35 3.495 ;
      RECT 68.115 4.23 68.12 4.37 ;
      RECT 67.775 4.23 67.81 4.368 ;
      RECT 67.35 4.215 67.365 4.36 ;
      RECT 69.18 3.995 69.27 4.255 ;
      RECT 69.01 3.86 69.11 4.255 ;
      RECT 66.045 3.835 66.125 4.045 ;
      RECT 69.135 3.972 69.18 4.255 ;
      RECT 69.125 3.942 69.135 4.255 ;
      RECT 69.11 3.865 69.125 4.255 ;
      RECT 68.925 3.86 69.01 4.22 ;
      RECT 68.92 3.862 68.925 4.215 ;
      RECT 68.915 3.867 68.92 4.215 ;
      RECT 68.88 3.967 68.915 4.215 ;
      RECT 68.87 3.995 68.88 4.215 ;
      RECT 68.86 4.01 68.87 4.215 ;
      RECT 68.85 4.022 68.86 4.215 ;
      RECT 68.845 4.032 68.85 4.215 ;
      RECT 68.83 4.042 68.845 4.217 ;
      RECT 68.825 4.057 68.83 4.219 ;
      RECT 68.81 4.07 68.825 4.221 ;
      RECT 68.805 4.085 68.81 4.224 ;
      RECT 68.785 4.095 68.805 4.228 ;
      RECT 68.77 4.105 68.785 4.231 ;
      RECT 68.735 4.112 68.77 4.236 ;
      RECT 68.691 4.119 68.735 4.244 ;
      RECT 68.605 4.131 68.691 4.257 ;
      RECT 68.58 4.142 68.605 4.268 ;
      RECT 68.55 4.147 68.58 4.273 ;
      RECT 68.515 4.152 68.55 4.281 ;
      RECT 68.485 4.157 68.515 4.288 ;
      RECT 68.46 4.162 68.485 4.293 ;
      RECT 68.395 4.169 68.46 4.302 ;
      RECT 68.325 4.182 68.395 4.318 ;
      RECT 68.295 4.192 68.325 4.33 ;
      RECT 68.27 4.197 68.295 4.337 ;
      RECT 68.215 4.204 68.27 4.345 ;
      RECT 68.21 4.211 68.215 4.35 ;
      RECT 68.205 4.213 68.21 4.351 ;
      RECT 68.19 4.215 68.205 4.353 ;
      RECT 68.185 4.215 68.19 4.356 ;
      RECT 68.12 4.222 68.185 4.363 ;
      RECT 68.085 4.232 68.115 4.373 ;
      RECT 68.068 4.235 68.085 4.375 ;
      RECT 67.982 4.234 68.068 4.374 ;
      RECT 67.896 4.232 67.982 4.371 ;
      RECT 67.81 4.231 67.896 4.369 ;
      RECT 67.709 4.229 67.775 4.368 ;
      RECT 67.623 4.226 67.709 4.366 ;
      RECT 67.537 4.222 67.623 4.364 ;
      RECT 67.451 4.219 67.537 4.363 ;
      RECT 67.365 4.216 67.451 4.361 ;
      RECT 67.265 4.215 67.35 4.358 ;
      RECT 67.215 4.213 67.265 4.356 ;
      RECT 67.195 4.21 67.215 4.354 ;
      RECT 67.175 4.208 67.195 4.351 ;
      RECT 67.15 4.204 67.175 4.348 ;
      RECT 67.105 4.198 67.15 4.343 ;
      RECT 67.065 4.192 67.105 4.335 ;
      RECT 67.04 4.187 67.065 4.328 ;
      RECT 66.985 4.18 67.04 4.32 ;
      RECT 66.961 4.173 66.985 4.313 ;
      RECT 66.875 4.164 66.961 4.303 ;
      RECT 66.845 4.156 66.875 4.293 ;
      RECT 66.815 4.152 66.845 4.288 ;
      RECT 66.81 4.149 66.815 4.285 ;
      RECT 66.805 4.148 66.81 4.285 ;
      RECT 66.73 4.141 66.805 4.278 ;
      RECT 66.691 4.132 66.73 4.267 ;
      RECT 66.605 4.122 66.691 4.255 ;
      RECT 66.565 4.112 66.605 4.243 ;
      RECT 66.526 4.107 66.565 4.236 ;
      RECT 66.44 4.097 66.526 4.225 ;
      RECT 66.4 4.085 66.44 4.214 ;
      RECT 66.365 4.07 66.4 4.207 ;
      RECT 66.355 4.06 66.365 4.204 ;
      RECT 66.335 4.045 66.355 4.202 ;
      RECT 66.305 4.015 66.335 4.198 ;
      RECT 66.295 3.995 66.305 4.193 ;
      RECT 66.29 3.987 66.295 4.19 ;
      RECT 66.285 3.98 66.29 4.188 ;
      RECT 66.27 3.967 66.285 4.181 ;
      RECT 66.265 3.957 66.27 4.173 ;
      RECT 66.26 3.95 66.265 4.168 ;
      RECT 66.255 3.945 66.26 4.164 ;
      RECT 66.24 3.932 66.255 4.156 ;
      RECT 66.235 3.842 66.24 4.145 ;
      RECT 66.23 3.837 66.235 4.138 ;
      RECT 66.155 3.835 66.23 4.098 ;
      RECT 66.125 3.835 66.155 4.053 ;
      RECT 66.03 3.84 66.045 4.04 ;
      RECT 68.515 3.545 68.775 3.805 ;
      RECT 68.5 3.533 68.68 3.77 ;
      RECT 68.495 3.534 68.68 3.768 ;
      RECT 68.48 3.538 68.69 3.758 ;
      RECT 68.475 3.543 68.695 3.728 ;
      RECT 68.48 3.54 68.695 3.758 ;
      RECT 68.495 3.535 68.69 3.768 ;
      RECT 68.515 3.532 68.68 3.805 ;
      RECT 68.515 3.531 68.67 3.805 ;
      RECT 68.54 3.53 68.67 3.805 ;
      RECT 68.1 3.775 68.36 4.035 ;
      RECT 67.975 3.82 68.36 4.03 ;
      RECT 67.965 3.825 68.36 4.025 ;
      RECT 67.98 4.765 67.995 5.075 ;
      RECT 66.575 4.535 66.585 4.665 ;
      RECT 66.355 4.53 66.46 4.665 ;
      RECT 66.27 4.535 66.32 4.665 ;
      RECT 64.82 3.27 64.825 4.375 ;
      RECT 68.075 4.857 68.08 4.993 ;
      RECT 68.07 4.852 68.075 5.053 ;
      RECT 68.065 4.85 68.07 5.066 ;
      RECT 68.05 4.847 68.065 5.068 ;
      RECT 68.045 4.842 68.05 5.07 ;
      RECT 68.04 4.838 68.045 5.073 ;
      RECT 68.025 4.833 68.04 5.075 ;
      RECT 67.995 4.825 68.025 5.075 ;
      RECT 67.956 4.765 67.98 5.075 ;
      RECT 67.87 4.765 67.956 5.072 ;
      RECT 67.84 4.765 67.87 5.065 ;
      RECT 67.815 4.765 67.84 5.058 ;
      RECT 67.79 4.765 67.815 5.05 ;
      RECT 67.775 4.765 67.79 5.043 ;
      RECT 67.75 4.765 67.775 5.035 ;
      RECT 67.735 4.765 67.75 5.028 ;
      RECT 67.695 4.775 67.735 5.017 ;
      RECT 67.685 4.77 67.695 5.007 ;
      RECT 67.681 4.769 67.685 5.004 ;
      RECT 67.595 4.761 67.681 4.987 ;
      RECT 67.562 4.75 67.595 4.964 ;
      RECT 67.476 4.739 67.562 4.942 ;
      RECT 67.39 4.723 67.476 4.911 ;
      RECT 67.32 4.708 67.39 4.883 ;
      RECT 67.31 4.701 67.32 4.87 ;
      RECT 67.28 4.698 67.31 4.86 ;
      RECT 67.255 4.694 67.28 4.853 ;
      RECT 67.24 4.691 67.255 4.848 ;
      RECT 67.235 4.69 67.24 4.843 ;
      RECT 67.205 4.685 67.235 4.836 ;
      RECT 67.2 4.68 67.205 4.831 ;
      RECT 67.185 4.677 67.2 4.826 ;
      RECT 67.18 4.672 67.185 4.821 ;
      RECT 67.16 4.667 67.18 4.818 ;
      RECT 67.145 4.662 67.16 4.81 ;
      RECT 67.13 4.656 67.145 4.805 ;
      RECT 67.1 4.647 67.13 4.798 ;
      RECT 67.095 4.64 67.1 4.79 ;
      RECT 67.09 4.638 67.095 4.788 ;
      RECT 67.085 4.637 67.09 4.785 ;
      RECT 67.045 4.63 67.085 4.778 ;
      RECT 67.031 4.62 67.045 4.768 ;
      RECT 66.98 4.609 67.031 4.756 ;
      RECT 66.955 4.595 66.98 4.742 ;
      RECT 66.93 4.584 66.955 4.734 ;
      RECT 66.91 4.573 66.93 4.728 ;
      RECT 66.9 4.567 66.91 4.723 ;
      RECT 66.895 4.565 66.9 4.719 ;
      RECT 66.875 4.56 66.895 4.714 ;
      RECT 66.845 4.55 66.875 4.704 ;
      RECT 66.84 4.542 66.845 4.697 ;
      RECT 66.825 4.54 66.84 4.693 ;
      RECT 66.805 4.54 66.825 4.688 ;
      RECT 66.8 4.539 66.805 4.686 ;
      RECT 66.795 4.539 66.8 4.683 ;
      RECT 66.755 4.538 66.795 4.678 ;
      RECT 66.73 4.537 66.755 4.673 ;
      RECT 66.67 4.536 66.73 4.67 ;
      RECT 66.585 4.535 66.67 4.668 ;
      RECT 66.546 4.534 66.575 4.665 ;
      RECT 66.46 4.532 66.546 4.665 ;
      RECT 66.32 4.532 66.355 4.665 ;
      RECT 66.23 4.536 66.27 4.668 ;
      RECT 66.215 4.539 66.23 4.675 ;
      RECT 66.205 4.54 66.215 4.682 ;
      RECT 66.18 4.543 66.205 4.687 ;
      RECT 66.175 4.545 66.18 4.69 ;
      RECT 66.125 4.547 66.175 4.691 ;
      RECT 66.086 4.551 66.125 4.693 ;
      RECT 66 4.553 66.086 4.696 ;
      RECT 65.982 4.555 66 4.698 ;
      RECT 65.896 4.558 65.982 4.7 ;
      RECT 65.81 4.562 65.896 4.703 ;
      RECT 65.773 4.566 65.81 4.706 ;
      RECT 65.687 4.569 65.773 4.709 ;
      RECT 65.601 4.573 65.687 4.712 ;
      RECT 65.515 4.578 65.601 4.716 ;
      RECT 65.495 4.58 65.515 4.719 ;
      RECT 65.475 4.579 65.495 4.72 ;
      RECT 65.426 4.576 65.475 4.721 ;
      RECT 65.34 4.571 65.426 4.724 ;
      RECT 65.29 4.566 65.34 4.726 ;
      RECT 65.266 4.564 65.29 4.727 ;
      RECT 65.18 4.559 65.266 4.729 ;
      RECT 65.155 4.555 65.18 4.728 ;
      RECT 65.145 4.552 65.155 4.726 ;
      RECT 65.135 4.545 65.145 4.723 ;
      RECT 65.13 4.525 65.135 4.718 ;
      RECT 65.12 4.495 65.13 4.713 ;
      RECT 65.105 4.365 65.12 4.704 ;
      RECT 65.1 4.357 65.105 4.697 ;
      RECT 65.08 4.35 65.1 4.689 ;
      RECT 65.075 4.332 65.08 4.681 ;
      RECT 65.065 4.312 65.075 4.676 ;
      RECT 65.06 4.285 65.065 4.672 ;
      RECT 65.055 4.262 65.06 4.669 ;
      RECT 65.035 4.22 65.055 4.661 ;
      RECT 65 4.135 65.035 4.645 ;
      RECT 64.995 4.067 65 4.633 ;
      RECT 64.98 4.037 64.995 4.627 ;
      RECT 64.975 3.282 64.98 3.528 ;
      RECT 64.965 4.007 64.98 4.618 ;
      RECT 64.97 3.277 64.975 3.56 ;
      RECT 64.965 3.272 64.97 3.603 ;
      RECT 64.96 3.27 64.965 3.638 ;
      RECT 64.945 3.97 64.965 4.608 ;
      RECT 64.955 3.27 64.96 3.675 ;
      RECT 64.94 3.27 64.955 3.773 ;
      RECT 64.94 3.943 64.945 4.601 ;
      RECT 64.935 3.27 64.94 3.848 ;
      RECT 64.935 3.931 64.94 4.598 ;
      RECT 64.93 3.27 64.935 3.88 ;
      RECT 64.93 3.91 64.935 4.595 ;
      RECT 64.925 3.27 64.93 4.592 ;
      RECT 64.89 3.27 64.925 4.578 ;
      RECT 64.875 3.27 64.89 4.56 ;
      RECT 64.855 3.27 64.875 4.55 ;
      RECT 64.83 3.27 64.855 4.533 ;
      RECT 64.825 3.27 64.83 4.483 ;
      RECT 64.815 3.27 64.82 4.313 ;
      RECT 64.81 3.27 64.815 4.22 ;
      RECT 64.805 3.27 64.81 4.133 ;
      RECT 64.8 3.27 64.805 4.065 ;
      RECT 64.795 3.27 64.8 4.008 ;
      RECT 64.785 3.27 64.795 3.903 ;
      RECT 64.78 3.27 64.785 3.775 ;
      RECT 64.775 3.27 64.78 3.693 ;
      RECT 64.77 3.272 64.775 3.61 ;
      RECT 64.765 3.277 64.77 3.543 ;
      RECT 64.76 3.282 64.765 3.47 ;
      RECT 67.575 3.6 67.835 3.86 ;
      RECT 67.595 3.567 67.805 3.86 ;
      RECT 67.595 3.565 67.795 3.86 ;
      RECT 67.605 3.552 67.795 3.86 ;
      RECT 67.605 3.55 67.72 3.86 ;
      RECT 67.08 3.675 67.255 3.955 ;
      RECT 67.075 3.675 67.255 3.953 ;
      RECT 67.075 3.675 67.27 3.95 ;
      RECT 67.065 3.675 67.27 3.948 ;
      RECT 67.01 3.675 67.27 3.935 ;
      RECT 67.01 3.75 67.275 3.913 ;
      RECT 66.555 3.687 66.575 3.93 ;
      RECT 66.555 3.687 66.615 3.929 ;
      RECT 66.55 3.689 66.615 3.928 ;
      RECT 66.55 3.689 66.701 3.927 ;
      RECT 66.55 3.689 66.77 3.926 ;
      RECT 66.55 3.689 66.79 3.918 ;
      RECT 66.53 3.692 66.79 3.916 ;
      RECT 66.515 3.702 66.79 3.901 ;
      RECT 66.515 3.702 66.805 3.9 ;
      RECT 66.51 3.711 66.805 3.892 ;
      RECT 66.51 3.711 66.81 3.888 ;
      RECT 66.615 3.625 66.875 3.885 ;
      RECT 66.505 3.713 66.875 3.77 ;
      RECT 66.575 3.68 66.875 3.885 ;
      RECT 66.54 4.873 66.545 5.08 ;
      RECT 66.49 4.867 66.54 5.079 ;
      RECT 66.457 4.881 66.55 5.078 ;
      RECT 66.371 4.881 66.55 5.077 ;
      RECT 66.285 4.881 66.55 5.076 ;
      RECT 66.285 4.98 66.555 5.073 ;
      RECT 66.28 4.98 66.555 5.068 ;
      RECT 66.275 4.98 66.555 5.05 ;
      RECT 66.27 4.98 66.555 5.033 ;
      RECT 66.23 4.765 66.49 5.025 ;
      RECT 65.69 3.915 65.776 4.329 ;
      RECT 65.69 3.915 65.815 4.326 ;
      RECT 65.69 3.915 65.835 4.316 ;
      RECT 65.645 3.915 65.835 4.313 ;
      RECT 65.645 4.067 65.845 4.303 ;
      RECT 65.645 4.088 65.85 4.297 ;
      RECT 65.645 4.106 65.855 4.293 ;
      RECT 65.645 4.126 65.865 4.288 ;
      RECT 65.62 4.126 65.865 4.285 ;
      RECT 65.61 4.126 65.865 4.263 ;
      RECT 65.61 4.142 65.87 4.233 ;
      RECT 65.575 3.915 65.835 4.22 ;
      RECT 65.575 4.154 65.875 4.175 ;
      RECT 63.235 10.06 63.525 10.29 ;
      RECT 63.295 8.58 63.465 10.29 ;
      RECT 63.245 8.945 63.595 9.295 ;
      RECT 63.235 8.58 63.525 8.81 ;
      RECT 62.83 3.69 62.935 4.26 ;
      RECT 62.83 4.025 63.155 4.255 ;
      RECT 62.83 4.055 63.325 4.225 ;
      RECT 62.83 3.69 63.02 4.255 ;
      RECT 62.245 3.655 62.535 3.885 ;
      RECT 62.245 3.69 63.02 3.86 ;
      RECT 62.305 2.175 62.475 3.885 ;
      RECT 62.245 2.175 62.535 2.405 ;
      RECT 62.245 10.06 62.535 10.29 ;
      RECT 62.305 8.58 62.475 10.29 ;
      RECT 62.245 8.58 62.535 8.81 ;
      RECT 62.245 8.615 63.095 8.775 ;
      RECT 62.93 8.21 63.095 8.775 ;
      RECT 62.245 8.61 62.64 8.775 ;
      RECT 62.865 8.21 63.155 8.44 ;
      RECT 62.865 8.24 63.325 8.41 ;
      RECT 61.875 4.025 62.165 4.255 ;
      RECT 61.875 4.055 62.335 4.225 ;
      RECT 61.94 2.95 62.105 4.255 ;
      RECT 60.455 2.92 60.745 3.15 ;
      RECT 60.455 2.95 62.105 3.12 ;
      RECT 60.515 2.18 60.685 3.15 ;
      RECT 60.455 2.18 60.745 2.41 ;
      RECT 60.455 10.055 60.745 10.285 ;
      RECT 60.515 9.315 60.685 10.285 ;
      RECT 60.515 9.41 62.105 9.58 ;
      RECT 61.935 8.21 62.105 9.58 ;
      RECT 60.455 9.315 60.745 9.545 ;
      RECT 61.875 8.21 62.165 8.44 ;
      RECT 61.875 8.24 62.335 8.41 ;
      RECT 58.505 4 58.845 4.35 ;
      RECT 58.595 3.32 58.765 4.35 ;
      RECT 60.885 3.26 61.235 3.61 ;
      RECT 58.595 3.32 61.235 3.49 ;
      RECT 60.91 8.945 61.235 9.27 ;
      RECT 55.45 8.9 55.8 9.25 ;
      RECT 60.885 8.945 61.235 9.175 ;
      RECT 55.25 8.945 55.8 9.175 ;
      RECT 55.08 8.975 61.235 9.145 ;
      RECT 60.11 3.66 60.43 3.98 ;
      RECT 60.08 3.66 60.43 3.89 ;
      RECT 59.91 3.69 60.43 3.86 ;
      RECT 60.11 8.545 60.43 8.835 ;
      RECT 60.08 8.575 60.43 8.805 ;
      RECT 59.91 8.605 60.43 8.775 ;
      RECT 55.8 4.28 55.95 4.555 ;
      RECT 56.34 3.36 56.345 3.58 ;
      RECT 57.49 3.56 57.505 3.758 ;
      RECT 57.455 3.552 57.49 3.765 ;
      RECT 57.425 3.545 57.455 3.765 ;
      RECT 57.37 3.51 57.425 3.765 ;
      RECT 57.305 3.447 57.37 3.765 ;
      RECT 57.3 3.412 57.305 3.763 ;
      RECT 57.295 3.407 57.3 3.755 ;
      RECT 57.29 3.402 57.295 3.741 ;
      RECT 57.285 3.399 57.29 3.734 ;
      RECT 57.24 3.389 57.285 3.685 ;
      RECT 57.22 3.376 57.24 3.62 ;
      RECT 57.215 3.371 57.22 3.593 ;
      RECT 57.21 3.37 57.215 3.586 ;
      RECT 57.205 3.369 57.21 3.579 ;
      RECT 57.12 3.354 57.205 3.525 ;
      RECT 57.09 3.335 57.12 3.475 ;
      RECT 57.01 3.318 57.09 3.46 ;
      RECT 56.975 3.305 57.01 3.445 ;
      RECT 56.967 3.305 56.975 3.44 ;
      RECT 56.881 3.306 56.967 3.44 ;
      RECT 56.795 3.308 56.881 3.44 ;
      RECT 56.77 3.309 56.795 3.444 ;
      RECT 56.695 3.315 56.77 3.459 ;
      RECT 56.612 3.327 56.695 3.483 ;
      RECT 56.526 3.34 56.612 3.509 ;
      RECT 56.44 3.353 56.526 3.535 ;
      RECT 56.405 3.362 56.44 3.554 ;
      RECT 56.355 3.362 56.405 3.567 ;
      RECT 56.345 3.36 56.355 3.578 ;
      RECT 56.33 3.357 56.34 3.58 ;
      RECT 56.315 3.349 56.33 3.588 ;
      RECT 56.3 3.341 56.315 3.608 ;
      RECT 56.295 3.336 56.3 3.665 ;
      RECT 56.28 3.331 56.295 3.738 ;
      RECT 56.275 3.326 56.28 3.78 ;
      RECT 56.27 3.324 56.275 3.808 ;
      RECT 56.265 3.322 56.27 3.83 ;
      RECT 56.255 3.318 56.265 3.873 ;
      RECT 56.25 3.315 56.255 3.898 ;
      RECT 56.245 3.313 56.25 3.918 ;
      RECT 56.24 3.311 56.245 3.942 ;
      RECT 56.235 3.307 56.24 3.965 ;
      RECT 56.23 3.303 56.235 3.988 ;
      RECT 56.195 3.293 56.23 4.095 ;
      RECT 56.19 3.283 56.195 4.193 ;
      RECT 56.185 3.281 56.19 4.22 ;
      RECT 56.18 3.28 56.185 4.24 ;
      RECT 56.175 3.272 56.18 4.26 ;
      RECT 56.17 3.267 56.175 4.295 ;
      RECT 56.165 3.265 56.17 4.313 ;
      RECT 56.16 3.265 56.165 4.338 ;
      RECT 56.155 3.265 56.16 4.36 ;
      RECT 56.12 3.265 56.155 4.403 ;
      RECT 56.095 3.265 56.12 4.432 ;
      RECT 56.085 3.265 56.095 3.618 ;
      RECT 56.088 3.675 56.095 4.442 ;
      RECT 56.085 3.732 56.088 4.445 ;
      RECT 56.08 3.265 56.085 3.59 ;
      RECT 56.08 3.782 56.085 4.448 ;
      RECT 56.07 3.265 56.08 3.58 ;
      RECT 56.075 3.835 56.08 4.451 ;
      RECT 56.07 3.92 56.075 4.455 ;
      RECT 56.06 3.265 56.07 3.568 ;
      RECT 56.065 3.967 56.07 4.459 ;
      RECT 56.06 4.042 56.065 4.463 ;
      RECT 56.025 3.265 56.06 3.543 ;
      RECT 56.05 4.125 56.06 4.468 ;
      RECT 56.04 4.192 56.05 4.475 ;
      RECT 56.035 4.22 56.04 4.48 ;
      RECT 56.025 4.233 56.035 4.486 ;
      RECT 55.98 3.265 56.025 3.5 ;
      RECT 56.02 4.238 56.025 4.493 ;
      RECT 55.98 4.255 56.02 4.555 ;
      RECT 55.975 3.267 55.98 3.473 ;
      RECT 55.95 4.275 55.98 4.555 ;
      RECT 55.97 3.272 55.975 3.445 ;
      RECT 55.76 4.284 55.8 4.555 ;
      RECT 55.735 4.292 55.76 4.525 ;
      RECT 55.69 4.3 55.735 4.525 ;
      RECT 55.675 4.305 55.69 4.52 ;
      RECT 55.665 4.305 55.675 4.514 ;
      RECT 55.655 4.312 55.665 4.511 ;
      RECT 55.65 4.35 55.655 4.5 ;
      RECT 55.645 4.412 55.65 4.478 ;
      RECT 56.915 4.287 57.1 4.51 ;
      RECT 56.915 4.302 57.105 4.506 ;
      RECT 56.905 3.575 56.99 4.505 ;
      RECT 56.905 4.302 57.11 4.499 ;
      RECT 56.9 4.31 57.11 4.498 ;
      RECT 57.105 4.03 57.425 4.35 ;
      RECT 56.9 4.202 57.07 4.293 ;
      RECT 56.895 4.202 57.07 4.275 ;
      RECT 56.885 4.01 57.02 4.25 ;
      RECT 56.88 4.01 57.02 4.195 ;
      RECT 56.84 3.59 57.01 4.095 ;
      RECT 56.825 3.59 57.01 3.965 ;
      RECT 56.82 3.59 57.01 3.918 ;
      RECT 56.815 3.59 57.01 3.898 ;
      RECT 56.81 3.59 57.01 3.873 ;
      RECT 56.78 3.59 57.04 3.85 ;
      RECT 56.79 3.587 57 3.85 ;
      RECT 56.915 3.582 57 4.51 ;
      RECT 56.8 3.575 56.99 3.85 ;
      RECT 56.795 3.58 56.99 3.85 ;
      RECT 55.625 3.792 55.81 4.005 ;
      RECT 55.625 3.8 55.82 3.998 ;
      RECT 55.605 3.8 55.82 3.995 ;
      RECT 55.6 3.8 55.82 3.98 ;
      RECT 55.53 3.715 55.79 3.975 ;
      RECT 55.53 3.86 55.825 3.888 ;
      RECT 55.185 4.315 55.445 4.575 ;
      RECT 55.21 4.26 55.405 4.575 ;
      RECT 55.205 4.009 55.385 4.303 ;
      RECT 55.205 4.015 55.395 4.303 ;
      RECT 55.185 4.017 55.395 4.248 ;
      RECT 55.18 4.027 55.395 4.115 ;
      RECT 55.21 4.007 55.385 4.575 ;
      RECT 55.296 4.005 55.385 4.575 ;
      RECT 55.155 3.225 55.19 3.595 ;
      RECT 54.945 3.335 54.95 3.595 ;
      RECT 55.19 3.232 55.205 3.595 ;
      RECT 55.08 3.225 55.155 3.673 ;
      RECT 55.07 3.225 55.08 3.758 ;
      RECT 55.045 3.225 55.07 3.793 ;
      RECT 55.005 3.225 55.045 3.861 ;
      RECT 54.995 3.232 55.005 3.913 ;
      RECT 54.965 3.335 54.995 3.954 ;
      RECT 54.96 3.335 54.965 3.993 ;
      RECT 54.95 3.335 54.96 4.013 ;
      RECT 54.945 3.63 54.95 4.05 ;
      RECT 54.94 3.647 54.945 4.07 ;
      RECT 54.925 3.71 54.94 4.11 ;
      RECT 54.92 3.753 54.925 4.145 ;
      RECT 54.915 3.761 54.92 4.158 ;
      RECT 54.905 3.775 54.915 4.18 ;
      RECT 54.88 3.81 54.905 4.245 ;
      RECT 54.87 3.845 54.88 4.308 ;
      RECT 54.85 3.875 54.87 4.369 ;
      RECT 54.835 3.911 54.85 4.436 ;
      RECT 54.825 3.939 54.835 4.475 ;
      RECT 54.815 3.961 54.825 4.495 ;
      RECT 54.81 3.971 54.815 4.506 ;
      RECT 54.805 3.98 54.81 4.509 ;
      RECT 54.795 3.998 54.805 4.513 ;
      RECT 54.785 4.016 54.795 4.514 ;
      RECT 54.76 4.055 54.785 4.511 ;
      RECT 54.74 4.097 54.76 4.508 ;
      RECT 54.725 4.135 54.74 4.507 ;
      RECT 54.69 4.17 54.725 4.504 ;
      RECT 54.685 4.192 54.69 4.502 ;
      RECT 54.62 4.232 54.685 4.499 ;
      RECT 54.615 4.272 54.62 4.495 ;
      RECT 54.6 4.282 54.615 4.486 ;
      RECT 54.59 4.402 54.6 4.471 ;
      RECT 55.07 4.815 55.08 5.075 ;
      RECT 55.07 4.818 55.09 5.074 ;
      RECT 55.06 4.808 55.07 5.073 ;
      RECT 55.05 4.823 55.13 5.069 ;
      RECT 55.035 4.802 55.05 5.067 ;
      RECT 55.01 4.827 55.135 5.063 ;
      RECT 54.995 4.787 55.01 5.058 ;
      RECT 54.995 4.829 55.145 5.057 ;
      RECT 54.995 4.837 55.16 5.05 ;
      RECT 54.935 4.774 54.995 5.04 ;
      RECT 54.925 4.761 54.935 5.022 ;
      RECT 54.9 4.751 54.925 5.012 ;
      RECT 54.895 4.741 54.9 5.004 ;
      RECT 54.83 4.837 55.16 4.986 ;
      RECT 54.745 4.837 55.16 4.948 ;
      RECT 54.635 4.665 54.895 4.925 ;
      RECT 55.01 4.795 55.035 5.063 ;
      RECT 55.05 4.805 55.06 5.069 ;
      RECT 54.635 4.813 55.075 4.925 ;
      RECT 54.82 10.055 55.11 10.285 ;
      RECT 54.88 9.315 55.05 10.285 ;
      RECT 54.78 9.345 55.15 9.715 ;
      RECT 54.82 9.315 55.11 9.715 ;
      RECT 53.85 4.57 53.88 4.87 ;
      RECT 53.625 4.555 53.63 4.83 ;
      RECT 53.425 4.555 53.58 4.815 ;
      RECT 54.725 3.27 54.755 3.53 ;
      RECT 54.715 3.27 54.725 3.638 ;
      RECT 54.695 3.27 54.715 3.648 ;
      RECT 54.68 3.27 54.695 3.66 ;
      RECT 54.625 3.27 54.68 3.71 ;
      RECT 54.61 3.27 54.625 3.758 ;
      RECT 54.58 3.27 54.61 3.793 ;
      RECT 54.525 3.27 54.58 3.855 ;
      RECT 54.505 3.27 54.525 3.923 ;
      RECT 54.5 3.27 54.505 3.953 ;
      RECT 54.495 3.27 54.5 3.965 ;
      RECT 54.49 3.387 54.495 3.983 ;
      RECT 54.47 3.405 54.49 4.008 ;
      RECT 54.45 3.432 54.47 4.058 ;
      RECT 54.445 3.452 54.45 4.089 ;
      RECT 54.44 3.46 54.445 4.106 ;
      RECT 54.425 3.486 54.44 4.135 ;
      RECT 54.41 3.528 54.425 4.17 ;
      RECT 54.405 3.557 54.41 4.193 ;
      RECT 54.4 3.572 54.405 4.206 ;
      RECT 54.395 3.595 54.4 4.217 ;
      RECT 54.385 3.615 54.395 4.235 ;
      RECT 54.375 3.645 54.385 4.258 ;
      RECT 54.37 3.667 54.375 4.278 ;
      RECT 54.365 3.682 54.37 4.293 ;
      RECT 54.35 3.712 54.365 4.32 ;
      RECT 54.345 3.742 54.35 4.346 ;
      RECT 54.34 3.76 54.345 4.358 ;
      RECT 54.33 3.79 54.34 4.377 ;
      RECT 54.32 3.815 54.33 4.402 ;
      RECT 54.315 3.835 54.32 4.421 ;
      RECT 54.31 3.852 54.315 4.434 ;
      RECT 54.3 3.878 54.31 4.453 ;
      RECT 54.29 3.916 54.3 4.48 ;
      RECT 54.285 3.942 54.29 4.5 ;
      RECT 54.28 3.952 54.285 4.51 ;
      RECT 54.275 3.965 54.28 4.525 ;
      RECT 54.27 3.98 54.275 4.535 ;
      RECT 54.265 4.002 54.27 4.55 ;
      RECT 54.26 4.02 54.265 4.561 ;
      RECT 54.255 4.03 54.26 4.572 ;
      RECT 54.25 4.038 54.255 4.584 ;
      RECT 54.245 4.046 54.25 4.595 ;
      RECT 54.24 4.072 54.245 4.608 ;
      RECT 54.23 4.1 54.24 4.621 ;
      RECT 54.225 4.13 54.23 4.63 ;
      RECT 54.22 4.145 54.225 4.637 ;
      RECT 54.205 4.17 54.22 4.644 ;
      RECT 54.2 4.192 54.205 4.65 ;
      RECT 54.195 4.217 54.2 4.653 ;
      RECT 54.186 4.245 54.195 4.657 ;
      RECT 54.18 4.262 54.186 4.662 ;
      RECT 54.175 4.28 54.18 4.666 ;
      RECT 54.17 4.292 54.175 4.669 ;
      RECT 54.165 4.313 54.17 4.673 ;
      RECT 54.16 4.331 54.165 4.676 ;
      RECT 54.155 4.345 54.16 4.679 ;
      RECT 54.15 4.362 54.155 4.682 ;
      RECT 54.145 4.375 54.15 4.685 ;
      RECT 54.12 4.412 54.145 4.693 ;
      RECT 54.115 4.457 54.12 4.702 ;
      RECT 54.11 4.485 54.115 4.705 ;
      RECT 54.1 4.505 54.11 4.709 ;
      RECT 54.095 4.525 54.1 4.714 ;
      RECT 54.09 4.54 54.095 4.717 ;
      RECT 54.07 4.55 54.09 4.724 ;
      RECT 54.005 4.557 54.07 4.75 ;
      RECT 53.97 4.56 54.005 4.778 ;
      RECT 53.955 4.563 53.97 4.793 ;
      RECT 53.945 4.564 53.955 4.808 ;
      RECT 53.935 4.565 53.945 4.825 ;
      RECT 53.93 4.565 53.935 4.84 ;
      RECT 53.925 4.565 53.93 4.848 ;
      RECT 53.91 4.566 53.925 4.863 ;
      RECT 53.88 4.568 53.91 4.87 ;
      RECT 53.77 4.575 53.85 4.87 ;
      RECT 53.725 4.58 53.77 4.87 ;
      RECT 53.715 4.581 53.725 4.86 ;
      RECT 53.705 4.582 53.715 4.853 ;
      RECT 53.685 4.584 53.705 4.848 ;
      RECT 53.675 4.555 53.685 4.843 ;
      RECT 53.63 4.555 53.675 4.835 ;
      RECT 53.6 4.555 53.625 4.825 ;
      RECT 53.58 4.555 53.6 4.818 ;
      RECT 53.86 3.355 54.12 3.615 ;
      RECT 53.74 3.37 53.75 3.535 ;
      RECT 53.725 3.37 53.73 3.53 ;
      RECT 51.09 3.21 51.275 3.5 ;
      RECT 52.905 3.335 52.92 3.49 ;
      RECT 51.055 3.21 51.08 3.47 ;
      RECT 53.47 3.26 53.475 3.402 ;
      RECT 53.385 3.255 53.41 3.395 ;
      RECT 53.785 3.372 53.86 3.565 ;
      RECT 53.77 3.37 53.785 3.548 ;
      RECT 53.75 3.37 53.77 3.54 ;
      RECT 53.73 3.37 53.74 3.533 ;
      RECT 53.685 3.365 53.725 3.523 ;
      RECT 53.645 3.34 53.685 3.508 ;
      RECT 53.63 3.315 53.645 3.498 ;
      RECT 53.625 3.309 53.63 3.496 ;
      RECT 53.59 3.301 53.625 3.479 ;
      RECT 53.585 3.294 53.59 3.467 ;
      RECT 53.565 3.289 53.585 3.455 ;
      RECT 53.555 3.283 53.565 3.44 ;
      RECT 53.535 3.278 53.555 3.425 ;
      RECT 53.525 3.273 53.535 3.418 ;
      RECT 53.52 3.271 53.525 3.413 ;
      RECT 53.515 3.27 53.52 3.41 ;
      RECT 53.475 3.265 53.515 3.406 ;
      RECT 53.455 3.259 53.47 3.401 ;
      RECT 53.42 3.256 53.455 3.398 ;
      RECT 53.41 3.255 53.42 3.396 ;
      RECT 53.35 3.255 53.385 3.393 ;
      RECT 53.305 3.255 53.35 3.393 ;
      RECT 53.255 3.255 53.305 3.396 ;
      RECT 53.24 3.257 53.255 3.398 ;
      RECT 53.225 3.26 53.24 3.399 ;
      RECT 53.215 3.265 53.225 3.4 ;
      RECT 53.185 3.27 53.215 3.405 ;
      RECT 53.175 3.276 53.185 3.413 ;
      RECT 53.165 3.278 53.175 3.417 ;
      RECT 53.155 3.282 53.165 3.421 ;
      RECT 53.13 3.288 53.155 3.429 ;
      RECT 53.12 3.293 53.13 3.437 ;
      RECT 53.105 3.297 53.12 3.441 ;
      RECT 53.07 3.303 53.105 3.449 ;
      RECT 53.05 3.308 53.07 3.459 ;
      RECT 53.02 3.315 53.05 3.468 ;
      RECT 52.975 3.324 53.02 3.482 ;
      RECT 52.97 3.329 52.975 3.493 ;
      RECT 52.95 3.332 52.97 3.494 ;
      RECT 52.92 3.335 52.95 3.492 ;
      RECT 52.885 3.335 52.905 3.488 ;
      RECT 52.815 3.335 52.885 3.479 ;
      RECT 52.8 3.332 52.815 3.471 ;
      RECT 52.76 3.325 52.8 3.466 ;
      RECT 52.735 3.315 52.76 3.459 ;
      RECT 52.73 3.309 52.735 3.456 ;
      RECT 52.69 3.303 52.73 3.453 ;
      RECT 52.675 3.296 52.69 3.448 ;
      RECT 52.655 3.292 52.675 3.443 ;
      RECT 52.64 3.287 52.655 3.439 ;
      RECT 52.625 3.282 52.64 3.437 ;
      RECT 52.61 3.278 52.625 3.436 ;
      RECT 52.595 3.276 52.61 3.432 ;
      RECT 52.585 3.274 52.595 3.427 ;
      RECT 52.57 3.271 52.585 3.423 ;
      RECT 52.56 3.269 52.57 3.418 ;
      RECT 52.54 3.266 52.56 3.414 ;
      RECT 52.495 3.265 52.54 3.412 ;
      RECT 52.435 3.267 52.495 3.413 ;
      RECT 52.415 3.269 52.435 3.415 ;
      RECT 52.385 3.272 52.415 3.416 ;
      RECT 52.335 3.277 52.385 3.418 ;
      RECT 52.33 3.28 52.335 3.42 ;
      RECT 52.32 3.282 52.33 3.423 ;
      RECT 52.315 3.284 52.32 3.426 ;
      RECT 52.265 3.287 52.315 3.433 ;
      RECT 52.245 3.291 52.265 3.445 ;
      RECT 52.235 3.294 52.245 3.451 ;
      RECT 52.225 3.295 52.235 3.454 ;
      RECT 52.186 3.298 52.225 3.456 ;
      RECT 52.1 3.305 52.186 3.459 ;
      RECT 52.026 3.315 52.1 3.463 ;
      RECT 51.94 3.326 52.026 3.468 ;
      RECT 51.925 3.333 51.94 3.47 ;
      RECT 51.87 3.337 51.925 3.471 ;
      RECT 51.856 3.34 51.87 3.473 ;
      RECT 51.77 3.34 51.856 3.475 ;
      RECT 51.73 3.337 51.77 3.478 ;
      RECT 51.706 3.333 51.73 3.48 ;
      RECT 51.62 3.323 51.706 3.483 ;
      RECT 51.59 3.312 51.62 3.484 ;
      RECT 51.571 3.308 51.59 3.483 ;
      RECT 51.485 3.301 51.571 3.48 ;
      RECT 51.425 3.29 51.485 3.477 ;
      RECT 51.405 3.282 51.425 3.475 ;
      RECT 51.37 3.277 51.405 3.474 ;
      RECT 51.345 3.272 51.37 3.473 ;
      RECT 51.315 3.267 51.345 3.472 ;
      RECT 51.29 3.21 51.315 3.471 ;
      RECT 51.275 3.21 51.29 3.495 ;
      RECT 51.08 3.21 51.09 3.495 ;
      RECT 52.855 4.23 52.86 4.37 ;
      RECT 52.515 4.23 52.55 4.368 ;
      RECT 52.09 4.215 52.105 4.36 ;
      RECT 53.92 3.995 54.01 4.255 ;
      RECT 53.75 3.86 53.85 4.255 ;
      RECT 50.785 3.835 50.865 4.045 ;
      RECT 53.875 3.972 53.92 4.255 ;
      RECT 53.865 3.942 53.875 4.255 ;
      RECT 53.85 3.865 53.865 4.255 ;
      RECT 53.665 3.86 53.75 4.22 ;
      RECT 53.66 3.862 53.665 4.215 ;
      RECT 53.655 3.867 53.66 4.215 ;
      RECT 53.62 3.967 53.655 4.215 ;
      RECT 53.61 3.995 53.62 4.215 ;
      RECT 53.6 4.01 53.61 4.215 ;
      RECT 53.59 4.022 53.6 4.215 ;
      RECT 53.585 4.032 53.59 4.215 ;
      RECT 53.57 4.042 53.585 4.217 ;
      RECT 53.565 4.057 53.57 4.219 ;
      RECT 53.55 4.07 53.565 4.221 ;
      RECT 53.545 4.085 53.55 4.224 ;
      RECT 53.525 4.095 53.545 4.228 ;
      RECT 53.51 4.105 53.525 4.231 ;
      RECT 53.475 4.112 53.51 4.236 ;
      RECT 53.431 4.119 53.475 4.244 ;
      RECT 53.345 4.131 53.431 4.257 ;
      RECT 53.32 4.142 53.345 4.268 ;
      RECT 53.29 4.147 53.32 4.273 ;
      RECT 53.255 4.152 53.29 4.281 ;
      RECT 53.225 4.157 53.255 4.288 ;
      RECT 53.2 4.162 53.225 4.293 ;
      RECT 53.135 4.169 53.2 4.302 ;
      RECT 53.065 4.182 53.135 4.318 ;
      RECT 53.035 4.192 53.065 4.33 ;
      RECT 53.01 4.197 53.035 4.337 ;
      RECT 52.955 4.204 53.01 4.345 ;
      RECT 52.95 4.211 52.955 4.35 ;
      RECT 52.945 4.213 52.95 4.351 ;
      RECT 52.93 4.215 52.945 4.353 ;
      RECT 52.925 4.215 52.93 4.356 ;
      RECT 52.86 4.222 52.925 4.363 ;
      RECT 52.825 4.232 52.855 4.373 ;
      RECT 52.808 4.235 52.825 4.375 ;
      RECT 52.722 4.234 52.808 4.374 ;
      RECT 52.636 4.232 52.722 4.371 ;
      RECT 52.55 4.231 52.636 4.369 ;
      RECT 52.449 4.229 52.515 4.368 ;
      RECT 52.363 4.226 52.449 4.366 ;
      RECT 52.277 4.222 52.363 4.364 ;
      RECT 52.191 4.219 52.277 4.363 ;
      RECT 52.105 4.216 52.191 4.361 ;
      RECT 52.005 4.215 52.09 4.358 ;
      RECT 51.955 4.213 52.005 4.356 ;
      RECT 51.935 4.21 51.955 4.354 ;
      RECT 51.915 4.208 51.935 4.351 ;
      RECT 51.89 4.204 51.915 4.348 ;
      RECT 51.845 4.198 51.89 4.343 ;
      RECT 51.805 4.192 51.845 4.335 ;
      RECT 51.78 4.187 51.805 4.328 ;
      RECT 51.725 4.18 51.78 4.32 ;
      RECT 51.701 4.173 51.725 4.313 ;
      RECT 51.615 4.164 51.701 4.303 ;
      RECT 51.585 4.156 51.615 4.293 ;
      RECT 51.555 4.152 51.585 4.288 ;
      RECT 51.55 4.149 51.555 4.285 ;
      RECT 51.545 4.148 51.55 4.285 ;
      RECT 51.47 4.141 51.545 4.278 ;
      RECT 51.431 4.132 51.47 4.267 ;
      RECT 51.345 4.122 51.431 4.255 ;
      RECT 51.305 4.112 51.345 4.243 ;
      RECT 51.266 4.107 51.305 4.236 ;
      RECT 51.18 4.097 51.266 4.225 ;
      RECT 51.14 4.085 51.18 4.214 ;
      RECT 51.105 4.07 51.14 4.207 ;
      RECT 51.095 4.06 51.105 4.204 ;
      RECT 51.075 4.045 51.095 4.202 ;
      RECT 51.045 4.015 51.075 4.198 ;
      RECT 51.035 3.995 51.045 4.193 ;
      RECT 51.03 3.987 51.035 4.19 ;
      RECT 51.025 3.98 51.03 4.188 ;
      RECT 51.01 3.967 51.025 4.181 ;
      RECT 51.005 3.957 51.01 4.173 ;
      RECT 51 3.95 51.005 4.168 ;
      RECT 50.995 3.945 51 4.164 ;
      RECT 50.98 3.932 50.995 4.156 ;
      RECT 50.975 3.842 50.98 4.145 ;
      RECT 50.97 3.837 50.975 4.138 ;
      RECT 50.895 3.835 50.97 4.098 ;
      RECT 50.865 3.835 50.895 4.053 ;
      RECT 50.77 3.84 50.785 4.04 ;
      RECT 53.255 3.545 53.515 3.805 ;
      RECT 53.24 3.533 53.42 3.77 ;
      RECT 53.235 3.534 53.42 3.768 ;
      RECT 53.22 3.538 53.43 3.758 ;
      RECT 53.215 3.543 53.435 3.728 ;
      RECT 53.22 3.54 53.435 3.758 ;
      RECT 53.235 3.535 53.43 3.768 ;
      RECT 53.255 3.532 53.42 3.805 ;
      RECT 53.255 3.531 53.41 3.805 ;
      RECT 53.28 3.53 53.41 3.805 ;
      RECT 52.84 3.775 53.1 4.035 ;
      RECT 52.715 3.82 53.1 4.03 ;
      RECT 52.705 3.825 53.1 4.025 ;
      RECT 52.72 4.765 52.735 5.075 ;
      RECT 51.315 4.535 51.325 4.665 ;
      RECT 51.095 4.53 51.2 4.665 ;
      RECT 51.01 4.535 51.06 4.665 ;
      RECT 49.56 3.27 49.565 4.375 ;
      RECT 52.815 4.857 52.82 4.993 ;
      RECT 52.81 4.852 52.815 5.053 ;
      RECT 52.805 4.85 52.81 5.066 ;
      RECT 52.79 4.847 52.805 5.068 ;
      RECT 52.785 4.842 52.79 5.07 ;
      RECT 52.78 4.838 52.785 5.073 ;
      RECT 52.765 4.833 52.78 5.075 ;
      RECT 52.735 4.825 52.765 5.075 ;
      RECT 52.696 4.765 52.72 5.075 ;
      RECT 52.61 4.765 52.696 5.072 ;
      RECT 52.58 4.765 52.61 5.065 ;
      RECT 52.555 4.765 52.58 5.058 ;
      RECT 52.53 4.765 52.555 5.05 ;
      RECT 52.515 4.765 52.53 5.043 ;
      RECT 52.49 4.765 52.515 5.035 ;
      RECT 52.475 4.765 52.49 5.028 ;
      RECT 52.435 4.775 52.475 5.017 ;
      RECT 52.425 4.77 52.435 5.007 ;
      RECT 52.421 4.769 52.425 5.004 ;
      RECT 52.335 4.761 52.421 4.987 ;
      RECT 52.302 4.75 52.335 4.964 ;
      RECT 52.216 4.739 52.302 4.942 ;
      RECT 52.13 4.723 52.216 4.911 ;
      RECT 52.06 4.708 52.13 4.883 ;
      RECT 52.05 4.701 52.06 4.87 ;
      RECT 52.02 4.698 52.05 4.86 ;
      RECT 51.995 4.694 52.02 4.853 ;
      RECT 51.98 4.691 51.995 4.848 ;
      RECT 51.975 4.69 51.98 4.843 ;
      RECT 51.945 4.685 51.975 4.836 ;
      RECT 51.94 4.68 51.945 4.831 ;
      RECT 51.925 4.677 51.94 4.826 ;
      RECT 51.92 4.672 51.925 4.821 ;
      RECT 51.9 4.667 51.92 4.818 ;
      RECT 51.885 4.662 51.9 4.81 ;
      RECT 51.87 4.656 51.885 4.805 ;
      RECT 51.84 4.647 51.87 4.798 ;
      RECT 51.835 4.64 51.84 4.79 ;
      RECT 51.83 4.638 51.835 4.788 ;
      RECT 51.825 4.637 51.83 4.785 ;
      RECT 51.785 4.63 51.825 4.778 ;
      RECT 51.771 4.62 51.785 4.768 ;
      RECT 51.72 4.609 51.771 4.756 ;
      RECT 51.695 4.595 51.72 4.742 ;
      RECT 51.67 4.584 51.695 4.734 ;
      RECT 51.65 4.573 51.67 4.728 ;
      RECT 51.64 4.567 51.65 4.723 ;
      RECT 51.635 4.565 51.64 4.719 ;
      RECT 51.615 4.56 51.635 4.714 ;
      RECT 51.585 4.55 51.615 4.704 ;
      RECT 51.58 4.542 51.585 4.697 ;
      RECT 51.565 4.54 51.58 4.693 ;
      RECT 51.545 4.54 51.565 4.688 ;
      RECT 51.54 4.539 51.545 4.686 ;
      RECT 51.535 4.539 51.54 4.683 ;
      RECT 51.495 4.538 51.535 4.678 ;
      RECT 51.47 4.537 51.495 4.673 ;
      RECT 51.41 4.536 51.47 4.67 ;
      RECT 51.325 4.535 51.41 4.668 ;
      RECT 51.286 4.534 51.315 4.665 ;
      RECT 51.2 4.532 51.286 4.665 ;
      RECT 51.06 4.532 51.095 4.665 ;
      RECT 50.97 4.536 51.01 4.668 ;
      RECT 50.955 4.539 50.97 4.675 ;
      RECT 50.945 4.54 50.955 4.682 ;
      RECT 50.92 4.543 50.945 4.687 ;
      RECT 50.915 4.545 50.92 4.69 ;
      RECT 50.865 4.547 50.915 4.691 ;
      RECT 50.826 4.551 50.865 4.693 ;
      RECT 50.74 4.553 50.826 4.696 ;
      RECT 50.722 4.555 50.74 4.698 ;
      RECT 50.636 4.558 50.722 4.7 ;
      RECT 50.55 4.562 50.636 4.703 ;
      RECT 50.513 4.566 50.55 4.706 ;
      RECT 50.427 4.569 50.513 4.709 ;
      RECT 50.341 4.573 50.427 4.712 ;
      RECT 50.255 4.578 50.341 4.716 ;
      RECT 50.235 4.58 50.255 4.719 ;
      RECT 50.215 4.579 50.235 4.72 ;
      RECT 50.166 4.576 50.215 4.721 ;
      RECT 50.08 4.571 50.166 4.724 ;
      RECT 50.03 4.566 50.08 4.726 ;
      RECT 50.006 4.564 50.03 4.727 ;
      RECT 49.92 4.559 50.006 4.729 ;
      RECT 49.895 4.555 49.92 4.728 ;
      RECT 49.885 4.552 49.895 4.726 ;
      RECT 49.875 4.545 49.885 4.723 ;
      RECT 49.87 4.525 49.875 4.718 ;
      RECT 49.86 4.495 49.87 4.713 ;
      RECT 49.845 4.365 49.86 4.704 ;
      RECT 49.84 4.357 49.845 4.697 ;
      RECT 49.82 4.35 49.84 4.689 ;
      RECT 49.815 4.332 49.82 4.681 ;
      RECT 49.805 4.312 49.815 4.676 ;
      RECT 49.8 4.285 49.805 4.672 ;
      RECT 49.795 4.262 49.8 4.669 ;
      RECT 49.775 4.22 49.795 4.661 ;
      RECT 49.74 4.135 49.775 4.645 ;
      RECT 49.735 4.067 49.74 4.633 ;
      RECT 49.72 4.037 49.735 4.627 ;
      RECT 49.715 3.282 49.72 3.528 ;
      RECT 49.705 4.007 49.72 4.618 ;
      RECT 49.71 3.277 49.715 3.56 ;
      RECT 49.705 3.272 49.71 3.603 ;
      RECT 49.7 3.27 49.705 3.638 ;
      RECT 49.685 3.97 49.705 4.608 ;
      RECT 49.695 3.27 49.7 3.675 ;
      RECT 49.68 3.27 49.695 3.773 ;
      RECT 49.68 3.943 49.685 4.601 ;
      RECT 49.675 3.27 49.68 3.848 ;
      RECT 49.675 3.931 49.68 4.598 ;
      RECT 49.67 3.27 49.675 3.88 ;
      RECT 49.67 3.91 49.675 4.595 ;
      RECT 49.665 3.27 49.67 4.592 ;
      RECT 49.63 3.27 49.665 4.578 ;
      RECT 49.615 3.27 49.63 4.56 ;
      RECT 49.595 3.27 49.615 4.55 ;
      RECT 49.57 3.27 49.595 4.533 ;
      RECT 49.565 3.27 49.57 4.483 ;
      RECT 49.555 3.27 49.56 4.313 ;
      RECT 49.55 3.27 49.555 4.22 ;
      RECT 49.545 3.27 49.55 4.133 ;
      RECT 49.54 3.27 49.545 4.065 ;
      RECT 49.535 3.27 49.54 4.008 ;
      RECT 49.525 3.27 49.535 3.903 ;
      RECT 49.52 3.27 49.525 3.775 ;
      RECT 49.515 3.27 49.52 3.693 ;
      RECT 49.51 3.272 49.515 3.61 ;
      RECT 49.505 3.277 49.51 3.543 ;
      RECT 49.5 3.282 49.505 3.47 ;
      RECT 52.315 3.6 52.575 3.86 ;
      RECT 52.335 3.567 52.545 3.86 ;
      RECT 52.335 3.565 52.535 3.86 ;
      RECT 52.345 3.552 52.535 3.86 ;
      RECT 52.345 3.55 52.46 3.86 ;
      RECT 51.82 3.675 51.995 3.955 ;
      RECT 51.815 3.675 51.995 3.953 ;
      RECT 51.815 3.675 52.01 3.95 ;
      RECT 51.805 3.675 52.01 3.948 ;
      RECT 51.75 3.675 52.01 3.935 ;
      RECT 51.75 3.75 52.015 3.913 ;
      RECT 51.295 3.687 51.315 3.93 ;
      RECT 51.295 3.687 51.355 3.929 ;
      RECT 51.29 3.689 51.355 3.928 ;
      RECT 51.29 3.689 51.441 3.927 ;
      RECT 51.29 3.689 51.51 3.926 ;
      RECT 51.29 3.689 51.53 3.918 ;
      RECT 51.27 3.692 51.53 3.916 ;
      RECT 51.255 3.702 51.53 3.901 ;
      RECT 51.255 3.702 51.545 3.9 ;
      RECT 51.25 3.711 51.545 3.892 ;
      RECT 51.25 3.711 51.55 3.888 ;
      RECT 51.355 3.625 51.615 3.885 ;
      RECT 51.245 3.713 51.615 3.77 ;
      RECT 51.315 3.68 51.615 3.885 ;
      RECT 51.28 4.873 51.285 5.08 ;
      RECT 51.23 4.867 51.28 5.079 ;
      RECT 51.197 4.881 51.29 5.078 ;
      RECT 51.111 4.881 51.29 5.077 ;
      RECT 51.025 4.881 51.29 5.076 ;
      RECT 51.025 4.98 51.295 5.073 ;
      RECT 51.02 4.98 51.295 5.068 ;
      RECT 51.015 4.98 51.295 5.05 ;
      RECT 51.01 4.98 51.295 5.033 ;
      RECT 50.97 4.765 51.23 5.025 ;
      RECT 50.43 3.915 50.516 4.329 ;
      RECT 50.43 3.915 50.555 4.326 ;
      RECT 50.43 3.915 50.575 4.316 ;
      RECT 50.385 3.915 50.575 4.313 ;
      RECT 50.385 4.067 50.585 4.303 ;
      RECT 50.385 4.088 50.59 4.297 ;
      RECT 50.385 4.106 50.595 4.293 ;
      RECT 50.385 4.126 50.605 4.288 ;
      RECT 50.36 4.126 50.605 4.285 ;
      RECT 50.35 4.126 50.605 4.263 ;
      RECT 50.35 4.142 50.61 4.233 ;
      RECT 50.315 3.915 50.575 4.22 ;
      RECT 50.315 4.154 50.615 4.175 ;
      RECT 47.975 10.06 48.265 10.29 ;
      RECT 48.035 8.58 48.205 10.29 ;
      RECT 47.985 8.945 48.335 9.295 ;
      RECT 47.975 8.58 48.265 8.81 ;
      RECT 47.57 3.69 47.675 4.26 ;
      RECT 47.57 4.025 47.895 4.255 ;
      RECT 47.57 4.055 48.065 4.225 ;
      RECT 47.57 3.69 47.76 4.255 ;
      RECT 46.985 3.655 47.275 3.885 ;
      RECT 46.985 3.69 47.76 3.86 ;
      RECT 47.045 2.175 47.215 3.885 ;
      RECT 46.985 2.175 47.275 2.405 ;
      RECT 46.985 10.06 47.275 10.29 ;
      RECT 47.045 8.58 47.215 10.29 ;
      RECT 46.985 8.58 47.275 8.81 ;
      RECT 46.985 8.615 47.835 8.775 ;
      RECT 47.67 8.21 47.835 8.775 ;
      RECT 46.985 8.61 47.38 8.775 ;
      RECT 47.605 8.21 47.895 8.44 ;
      RECT 47.605 8.24 48.065 8.41 ;
      RECT 46.615 4.025 46.905 4.255 ;
      RECT 46.615 4.055 47.075 4.225 ;
      RECT 46.68 2.95 46.845 4.255 ;
      RECT 45.195 2.92 45.485 3.15 ;
      RECT 45.195 2.95 46.845 3.12 ;
      RECT 45.255 2.18 45.425 3.15 ;
      RECT 45.195 2.18 45.485 2.41 ;
      RECT 45.195 10.055 45.485 10.285 ;
      RECT 45.255 9.315 45.425 10.285 ;
      RECT 45.255 9.41 46.845 9.58 ;
      RECT 46.675 8.21 46.845 9.58 ;
      RECT 45.195 9.315 45.485 9.545 ;
      RECT 46.615 8.21 46.905 8.44 ;
      RECT 46.615 8.24 47.075 8.41 ;
      RECT 43.245 4 43.585 4.35 ;
      RECT 43.335 3.32 43.505 4.35 ;
      RECT 45.625 3.26 45.975 3.61 ;
      RECT 43.335 3.32 45.975 3.49 ;
      RECT 45.65 8.945 45.975 9.27 ;
      RECT 40.19 8.905 40.54 9.255 ;
      RECT 45.625 8.945 45.975 9.175 ;
      RECT 39.99 8.945 40.54 9.175 ;
      RECT 39.82 8.975 45.975 9.145 ;
      RECT 44.85 3.66 45.17 3.98 ;
      RECT 44.82 3.66 45.17 3.89 ;
      RECT 44.65 3.69 45.17 3.86 ;
      RECT 44.85 8.545 45.17 8.835 ;
      RECT 44.82 8.575 45.17 8.805 ;
      RECT 44.65 8.605 45.17 8.775 ;
      RECT 40.54 4.28 40.69 4.555 ;
      RECT 41.08 3.36 41.085 3.58 ;
      RECT 42.23 3.56 42.245 3.758 ;
      RECT 42.195 3.552 42.23 3.765 ;
      RECT 42.165 3.545 42.195 3.765 ;
      RECT 42.11 3.51 42.165 3.765 ;
      RECT 42.045 3.447 42.11 3.765 ;
      RECT 42.04 3.412 42.045 3.763 ;
      RECT 42.035 3.407 42.04 3.755 ;
      RECT 42.03 3.402 42.035 3.741 ;
      RECT 42.025 3.399 42.03 3.734 ;
      RECT 41.98 3.389 42.025 3.685 ;
      RECT 41.96 3.376 41.98 3.62 ;
      RECT 41.955 3.371 41.96 3.593 ;
      RECT 41.95 3.37 41.955 3.586 ;
      RECT 41.945 3.369 41.95 3.579 ;
      RECT 41.86 3.354 41.945 3.525 ;
      RECT 41.83 3.335 41.86 3.475 ;
      RECT 41.75 3.318 41.83 3.46 ;
      RECT 41.715 3.305 41.75 3.445 ;
      RECT 41.707 3.305 41.715 3.44 ;
      RECT 41.621 3.306 41.707 3.44 ;
      RECT 41.535 3.308 41.621 3.44 ;
      RECT 41.51 3.309 41.535 3.444 ;
      RECT 41.435 3.315 41.51 3.459 ;
      RECT 41.352 3.327 41.435 3.483 ;
      RECT 41.266 3.34 41.352 3.509 ;
      RECT 41.18 3.353 41.266 3.535 ;
      RECT 41.145 3.362 41.18 3.554 ;
      RECT 41.095 3.362 41.145 3.567 ;
      RECT 41.085 3.36 41.095 3.578 ;
      RECT 41.07 3.357 41.08 3.58 ;
      RECT 41.055 3.349 41.07 3.588 ;
      RECT 41.04 3.341 41.055 3.608 ;
      RECT 41.035 3.336 41.04 3.665 ;
      RECT 41.02 3.331 41.035 3.738 ;
      RECT 41.015 3.326 41.02 3.78 ;
      RECT 41.01 3.324 41.015 3.808 ;
      RECT 41.005 3.322 41.01 3.83 ;
      RECT 40.995 3.318 41.005 3.873 ;
      RECT 40.99 3.315 40.995 3.898 ;
      RECT 40.985 3.313 40.99 3.918 ;
      RECT 40.98 3.311 40.985 3.942 ;
      RECT 40.975 3.307 40.98 3.965 ;
      RECT 40.97 3.303 40.975 3.988 ;
      RECT 40.935 3.293 40.97 4.095 ;
      RECT 40.93 3.283 40.935 4.193 ;
      RECT 40.925 3.281 40.93 4.22 ;
      RECT 40.92 3.28 40.925 4.24 ;
      RECT 40.915 3.272 40.92 4.26 ;
      RECT 40.91 3.267 40.915 4.295 ;
      RECT 40.905 3.265 40.91 4.313 ;
      RECT 40.9 3.265 40.905 4.338 ;
      RECT 40.895 3.265 40.9 4.36 ;
      RECT 40.86 3.265 40.895 4.403 ;
      RECT 40.835 3.265 40.86 4.432 ;
      RECT 40.825 3.265 40.835 3.618 ;
      RECT 40.828 3.675 40.835 4.442 ;
      RECT 40.825 3.732 40.828 4.445 ;
      RECT 40.82 3.265 40.825 3.59 ;
      RECT 40.82 3.782 40.825 4.448 ;
      RECT 40.81 3.265 40.82 3.58 ;
      RECT 40.815 3.835 40.82 4.451 ;
      RECT 40.81 3.92 40.815 4.455 ;
      RECT 40.8 3.265 40.81 3.568 ;
      RECT 40.805 3.967 40.81 4.459 ;
      RECT 40.8 4.042 40.805 4.463 ;
      RECT 40.765 3.265 40.8 3.543 ;
      RECT 40.79 4.125 40.8 4.468 ;
      RECT 40.78 4.192 40.79 4.475 ;
      RECT 40.775 4.22 40.78 4.48 ;
      RECT 40.765 4.233 40.775 4.486 ;
      RECT 40.72 3.265 40.765 3.5 ;
      RECT 40.76 4.238 40.765 4.493 ;
      RECT 40.72 4.255 40.76 4.555 ;
      RECT 40.715 3.267 40.72 3.473 ;
      RECT 40.69 4.275 40.72 4.555 ;
      RECT 40.71 3.272 40.715 3.445 ;
      RECT 40.5 4.284 40.54 4.555 ;
      RECT 40.475 4.292 40.5 4.525 ;
      RECT 40.43 4.3 40.475 4.525 ;
      RECT 40.415 4.305 40.43 4.52 ;
      RECT 40.405 4.305 40.415 4.514 ;
      RECT 40.395 4.312 40.405 4.511 ;
      RECT 40.39 4.35 40.395 4.5 ;
      RECT 40.385 4.412 40.39 4.478 ;
      RECT 41.655 4.287 41.84 4.51 ;
      RECT 41.655 4.302 41.845 4.506 ;
      RECT 41.645 3.575 41.73 4.505 ;
      RECT 41.645 4.302 41.85 4.499 ;
      RECT 41.64 4.31 41.85 4.498 ;
      RECT 41.845 4.03 42.165 4.35 ;
      RECT 41.64 4.202 41.81 4.293 ;
      RECT 41.635 4.202 41.81 4.275 ;
      RECT 41.625 4.01 41.76 4.25 ;
      RECT 41.62 4.01 41.76 4.195 ;
      RECT 41.58 3.59 41.75 4.095 ;
      RECT 41.565 3.59 41.75 3.965 ;
      RECT 41.56 3.59 41.75 3.918 ;
      RECT 41.555 3.59 41.75 3.898 ;
      RECT 41.55 3.59 41.75 3.873 ;
      RECT 41.52 3.59 41.78 3.85 ;
      RECT 41.53 3.587 41.74 3.85 ;
      RECT 41.655 3.582 41.74 4.51 ;
      RECT 41.54 3.575 41.73 3.85 ;
      RECT 41.535 3.58 41.73 3.85 ;
      RECT 40.365 3.792 40.55 4.005 ;
      RECT 40.365 3.8 40.56 3.998 ;
      RECT 40.345 3.8 40.56 3.995 ;
      RECT 40.34 3.8 40.56 3.98 ;
      RECT 40.27 3.715 40.53 3.975 ;
      RECT 40.27 3.86 40.565 3.888 ;
      RECT 39.925 4.315 40.185 4.575 ;
      RECT 39.95 4.26 40.145 4.575 ;
      RECT 39.945 4.009 40.125 4.303 ;
      RECT 39.945 4.015 40.135 4.303 ;
      RECT 39.925 4.017 40.135 4.248 ;
      RECT 39.92 4.027 40.135 4.115 ;
      RECT 39.95 4.007 40.125 4.575 ;
      RECT 40.036 4.005 40.125 4.575 ;
      RECT 39.895 3.225 39.93 3.595 ;
      RECT 39.685 3.335 39.69 3.595 ;
      RECT 39.93 3.232 39.945 3.595 ;
      RECT 39.82 3.225 39.895 3.673 ;
      RECT 39.81 3.225 39.82 3.758 ;
      RECT 39.785 3.225 39.81 3.793 ;
      RECT 39.745 3.225 39.785 3.861 ;
      RECT 39.735 3.232 39.745 3.913 ;
      RECT 39.705 3.335 39.735 3.954 ;
      RECT 39.7 3.335 39.705 3.993 ;
      RECT 39.69 3.335 39.7 4.013 ;
      RECT 39.685 3.63 39.69 4.05 ;
      RECT 39.68 3.647 39.685 4.07 ;
      RECT 39.665 3.71 39.68 4.11 ;
      RECT 39.66 3.753 39.665 4.145 ;
      RECT 39.655 3.761 39.66 4.158 ;
      RECT 39.645 3.775 39.655 4.18 ;
      RECT 39.62 3.81 39.645 4.245 ;
      RECT 39.61 3.845 39.62 4.308 ;
      RECT 39.59 3.875 39.61 4.369 ;
      RECT 39.575 3.911 39.59 4.436 ;
      RECT 39.565 3.939 39.575 4.475 ;
      RECT 39.555 3.961 39.565 4.495 ;
      RECT 39.55 3.971 39.555 4.506 ;
      RECT 39.545 3.98 39.55 4.509 ;
      RECT 39.535 3.998 39.545 4.513 ;
      RECT 39.525 4.016 39.535 4.514 ;
      RECT 39.5 4.055 39.525 4.511 ;
      RECT 39.48 4.097 39.5 4.508 ;
      RECT 39.465 4.135 39.48 4.507 ;
      RECT 39.43 4.17 39.465 4.504 ;
      RECT 39.425 4.192 39.43 4.502 ;
      RECT 39.36 4.232 39.425 4.499 ;
      RECT 39.355 4.272 39.36 4.495 ;
      RECT 39.34 4.282 39.355 4.486 ;
      RECT 39.33 4.402 39.34 4.471 ;
      RECT 39.81 4.815 39.82 5.075 ;
      RECT 39.81 4.818 39.83 5.074 ;
      RECT 39.8 4.808 39.81 5.073 ;
      RECT 39.79 4.823 39.87 5.069 ;
      RECT 39.775 4.802 39.79 5.067 ;
      RECT 39.75 4.827 39.875 5.063 ;
      RECT 39.735 4.787 39.75 5.058 ;
      RECT 39.735 4.829 39.885 5.057 ;
      RECT 39.735 4.837 39.9 5.05 ;
      RECT 39.675 4.774 39.735 5.04 ;
      RECT 39.665 4.761 39.675 5.022 ;
      RECT 39.64 4.751 39.665 5.012 ;
      RECT 39.635 4.741 39.64 5.004 ;
      RECT 39.57 4.837 39.9 4.986 ;
      RECT 39.485 4.837 39.9 4.948 ;
      RECT 39.375 4.665 39.635 4.925 ;
      RECT 39.75 4.795 39.775 5.063 ;
      RECT 39.79 4.805 39.8 5.069 ;
      RECT 39.375 4.813 39.815 4.925 ;
      RECT 39.56 10.055 39.85 10.285 ;
      RECT 39.62 9.315 39.79 10.285 ;
      RECT 39.52 9.345 39.89 9.715 ;
      RECT 39.56 9.315 39.85 9.715 ;
      RECT 38.59 4.57 38.62 4.87 ;
      RECT 38.365 4.555 38.37 4.83 ;
      RECT 38.165 4.555 38.32 4.815 ;
      RECT 39.465 3.27 39.495 3.53 ;
      RECT 39.455 3.27 39.465 3.638 ;
      RECT 39.435 3.27 39.455 3.648 ;
      RECT 39.42 3.27 39.435 3.66 ;
      RECT 39.365 3.27 39.42 3.71 ;
      RECT 39.35 3.27 39.365 3.758 ;
      RECT 39.32 3.27 39.35 3.793 ;
      RECT 39.265 3.27 39.32 3.855 ;
      RECT 39.245 3.27 39.265 3.923 ;
      RECT 39.24 3.27 39.245 3.953 ;
      RECT 39.235 3.27 39.24 3.965 ;
      RECT 39.23 3.387 39.235 3.983 ;
      RECT 39.21 3.405 39.23 4.008 ;
      RECT 39.19 3.432 39.21 4.058 ;
      RECT 39.185 3.452 39.19 4.089 ;
      RECT 39.18 3.46 39.185 4.106 ;
      RECT 39.165 3.486 39.18 4.135 ;
      RECT 39.15 3.528 39.165 4.17 ;
      RECT 39.145 3.557 39.15 4.193 ;
      RECT 39.14 3.572 39.145 4.206 ;
      RECT 39.135 3.595 39.14 4.217 ;
      RECT 39.125 3.615 39.135 4.235 ;
      RECT 39.115 3.645 39.125 4.258 ;
      RECT 39.11 3.667 39.115 4.278 ;
      RECT 39.105 3.682 39.11 4.293 ;
      RECT 39.09 3.712 39.105 4.32 ;
      RECT 39.085 3.742 39.09 4.346 ;
      RECT 39.08 3.76 39.085 4.358 ;
      RECT 39.07 3.79 39.08 4.377 ;
      RECT 39.06 3.815 39.07 4.402 ;
      RECT 39.055 3.835 39.06 4.421 ;
      RECT 39.05 3.852 39.055 4.434 ;
      RECT 39.04 3.878 39.05 4.453 ;
      RECT 39.03 3.916 39.04 4.48 ;
      RECT 39.025 3.942 39.03 4.5 ;
      RECT 39.02 3.952 39.025 4.51 ;
      RECT 39.015 3.965 39.02 4.525 ;
      RECT 39.01 3.98 39.015 4.535 ;
      RECT 39.005 4.002 39.01 4.55 ;
      RECT 39 4.02 39.005 4.561 ;
      RECT 38.995 4.03 39 4.572 ;
      RECT 38.99 4.038 38.995 4.584 ;
      RECT 38.985 4.046 38.99 4.595 ;
      RECT 38.98 4.072 38.985 4.608 ;
      RECT 38.97 4.1 38.98 4.621 ;
      RECT 38.965 4.13 38.97 4.63 ;
      RECT 38.96 4.145 38.965 4.637 ;
      RECT 38.945 4.17 38.96 4.644 ;
      RECT 38.94 4.192 38.945 4.65 ;
      RECT 38.935 4.217 38.94 4.653 ;
      RECT 38.926 4.245 38.935 4.657 ;
      RECT 38.92 4.262 38.926 4.662 ;
      RECT 38.915 4.28 38.92 4.666 ;
      RECT 38.91 4.292 38.915 4.669 ;
      RECT 38.905 4.313 38.91 4.673 ;
      RECT 38.9 4.331 38.905 4.676 ;
      RECT 38.895 4.345 38.9 4.679 ;
      RECT 38.89 4.362 38.895 4.682 ;
      RECT 38.885 4.375 38.89 4.685 ;
      RECT 38.86 4.412 38.885 4.693 ;
      RECT 38.855 4.457 38.86 4.702 ;
      RECT 38.85 4.485 38.855 4.705 ;
      RECT 38.84 4.505 38.85 4.709 ;
      RECT 38.835 4.525 38.84 4.714 ;
      RECT 38.83 4.54 38.835 4.717 ;
      RECT 38.81 4.55 38.83 4.724 ;
      RECT 38.745 4.557 38.81 4.75 ;
      RECT 38.71 4.56 38.745 4.778 ;
      RECT 38.695 4.563 38.71 4.793 ;
      RECT 38.685 4.564 38.695 4.808 ;
      RECT 38.675 4.565 38.685 4.825 ;
      RECT 38.67 4.565 38.675 4.84 ;
      RECT 38.665 4.565 38.67 4.848 ;
      RECT 38.65 4.566 38.665 4.863 ;
      RECT 38.62 4.568 38.65 4.87 ;
      RECT 38.51 4.575 38.59 4.87 ;
      RECT 38.465 4.58 38.51 4.87 ;
      RECT 38.455 4.581 38.465 4.86 ;
      RECT 38.445 4.582 38.455 4.853 ;
      RECT 38.425 4.584 38.445 4.848 ;
      RECT 38.415 4.555 38.425 4.843 ;
      RECT 38.37 4.555 38.415 4.835 ;
      RECT 38.34 4.555 38.365 4.825 ;
      RECT 38.32 4.555 38.34 4.818 ;
      RECT 38.6 3.355 38.86 3.615 ;
      RECT 38.48 3.37 38.49 3.535 ;
      RECT 38.465 3.37 38.47 3.53 ;
      RECT 35.83 3.21 36.015 3.5 ;
      RECT 37.645 3.335 37.66 3.49 ;
      RECT 35.795 3.21 35.82 3.47 ;
      RECT 38.21 3.26 38.215 3.402 ;
      RECT 38.125 3.255 38.15 3.395 ;
      RECT 38.525 3.372 38.6 3.565 ;
      RECT 38.51 3.37 38.525 3.548 ;
      RECT 38.49 3.37 38.51 3.54 ;
      RECT 38.47 3.37 38.48 3.533 ;
      RECT 38.425 3.365 38.465 3.523 ;
      RECT 38.385 3.34 38.425 3.508 ;
      RECT 38.37 3.315 38.385 3.498 ;
      RECT 38.365 3.309 38.37 3.496 ;
      RECT 38.33 3.301 38.365 3.479 ;
      RECT 38.325 3.294 38.33 3.467 ;
      RECT 38.305 3.289 38.325 3.455 ;
      RECT 38.295 3.283 38.305 3.44 ;
      RECT 38.275 3.278 38.295 3.425 ;
      RECT 38.265 3.273 38.275 3.418 ;
      RECT 38.26 3.271 38.265 3.413 ;
      RECT 38.255 3.27 38.26 3.41 ;
      RECT 38.215 3.265 38.255 3.406 ;
      RECT 38.195 3.259 38.21 3.401 ;
      RECT 38.16 3.256 38.195 3.398 ;
      RECT 38.15 3.255 38.16 3.396 ;
      RECT 38.09 3.255 38.125 3.393 ;
      RECT 38.045 3.255 38.09 3.393 ;
      RECT 37.995 3.255 38.045 3.396 ;
      RECT 37.98 3.257 37.995 3.398 ;
      RECT 37.965 3.26 37.98 3.399 ;
      RECT 37.955 3.265 37.965 3.4 ;
      RECT 37.925 3.27 37.955 3.405 ;
      RECT 37.915 3.276 37.925 3.413 ;
      RECT 37.905 3.278 37.915 3.417 ;
      RECT 37.895 3.282 37.905 3.421 ;
      RECT 37.87 3.288 37.895 3.429 ;
      RECT 37.86 3.293 37.87 3.437 ;
      RECT 37.845 3.297 37.86 3.441 ;
      RECT 37.81 3.303 37.845 3.449 ;
      RECT 37.79 3.308 37.81 3.459 ;
      RECT 37.76 3.315 37.79 3.468 ;
      RECT 37.715 3.324 37.76 3.482 ;
      RECT 37.71 3.329 37.715 3.493 ;
      RECT 37.69 3.332 37.71 3.494 ;
      RECT 37.66 3.335 37.69 3.492 ;
      RECT 37.625 3.335 37.645 3.488 ;
      RECT 37.555 3.335 37.625 3.479 ;
      RECT 37.54 3.332 37.555 3.471 ;
      RECT 37.5 3.325 37.54 3.466 ;
      RECT 37.475 3.315 37.5 3.459 ;
      RECT 37.47 3.309 37.475 3.456 ;
      RECT 37.43 3.303 37.47 3.453 ;
      RECT 37.415 3.296 37.43 3.448 ;
      RECT 37.395 3.292 37.415 3.443 ;
      RECT 37.38 3.287 37.395 3.439 ;
      RECT 37.365 3.282 37.38 3.437 ;
      RECT 37.35 3.278 37.365 3.436 ;
      RECT 37.335 3.276 37.35 3.432 ;
      RECT 37.325 3.274 37.335 3.427 ;
      RECT 37.31 3.271 37.325 3.423 ;
      RECT 37.3 3.269 37.31 3.418 ;
      RECT 37.28 3.266 37.3 3.414 ;
      RECT 37.235 3.265 37.28 3.412 ;
      RECT 37.175 3.267 37.235 3.413 ;
      RECT 37.155 3.269 37.175 3.415 ;
      RECT 37.125 3.272 37.155 3.416 ;
      RECT 37.075 3.277 37.125 3.418 ;
      RECT 37.07 3.28 37.075 3.42 ;
      RECT 37.06 3.282 37.07 3.423 ;
      RECT 37.055 3.284 37.06 3.426 ;
      RECT 37.005 3.287 37.055 3.433 ;
      RECT 36.985 3.291 37.005 3.445 ;
      RECT 36.975 3.294 36.985 3.451 ;
      RECT 36.965 3.295 36.975 3.454 ;
      RECT 36.926 3.298 36.965 3.456 ;
      RECT 36.84 3.305 36.926 3.459 ;
      RECT 36.766 3.315 36.84 3.463 ;
      RECT 36.68 3.326 36.766 3.468 ;
      RECT 36.665 3.333 36.68 3.47 ;
      RECT 36.61 3.337 36.665 3.471 ;
      RECT 36.596 3.34 36.61 3.473 ;
      RECT 36.51 3.34 36.596 3.475 ;
      RECT 36.47 3.337 36.51 3.478 ;
      RECT 36.446 3.333 36.47 3.48 ;
      RECT 36.36 3.323 36.446 3.483 ;
      RECT 36.33 3.312 36.36 3.484 ;
      RECT 36.311 3.308 36.33 3.483 ;
      RECT 36.225 3.301 36.311 3.48 ;
      RECT 36.165 3.29 36.225 3.477 ;
      RECT 36.145 3.282 36.165 3.475 ;
      RECT 36.11 3.277 36.145 3.474 ;
      RECT 36.085 3.272 36.11 3.473 ;
      RECT 36.055 3.267 36.085 3.472 ;
      RECT 36.03 3.21 36.055 3.471 ;
      RECT 36.015 3.21 36.03 3.495 ;
      RECT 35.82 3.21 35.83 3.495 ;
      RECT 37.595 4.23 37.6 4.37 ;
      RECT 37.255 4.23 37.29 4.368 ;
      RECT 36.83 4.215 36.845 4.36 ;
      RECT 38.66 3.995 38.75 4.255 ;
      RECT 38.49 3.86 38.59 4.255 ;
      RECT 35.525 3.835 35.605 4.045 ;
      RECT 38.615 3.972 38.66 4.255 ;
      RECT 38.605 3.942 38.615 4.255 ;
      RECT 38.59 3.865 38.605 4.255 ;
      RECT 38.405 3.86 38.49 4.22 ;
      RECT 38.4 3.862 38.405 4.215 ;
      RECT 38.395 3.867 38.4 4.215 ;
      RECT 38.36 3.967 38.395 4.215 ;
      RECT 38.35 3.995 38.36 4.215 ;
      RECT 38.34 4.01 38.35 4.215 ;
      RECT 38.33 4.022 38.34 4.215 ;
      RECT 38.325 4.032 38.33 4.215 ;
      RECT 38.31 4.042 38.325 4.217 ;
      RECT 38.305 4.057 38.31 4.219 ;
      RECT 38.29 4.07 38.305 4.221 ;
      RECT 38.285 4.085 38.29 4.224 ;
      RECT 38.265 4.095 38.285 4.228 ;
      RECT 38.25 4.105 38.265 4.231 ;
      RECT 38.215 4.112 38.25 4.236 ;
      RECT 38.171 4.119 38.215 4.244 ;
      RECT 38.085 4.131 38.171 4.257 ;
      RECT 38.06 4.142 38.085 4.268 ;
      RECT 38.03 4.147 38.06 4.273 ;
      RECT 37.995 4.152 38.03 4.281 ;
      RECT 37.965 4.157 37.995 4.288 ;
      RECT 37.94 4.162 37.965 4.293 ;
      RECT 37.875 4.169 37.94 4.302 ;
      RECT 37.805 4.182 37.875 4.318 ;
      RECT 37.775 4.192 37.805 4.33 ;
      RECT 37.75 4.197 37.775 4.337 ;
      RECT 37.695 4.204 37.75 4.345 ;
      RECT 37.69 4.211 37.695 4.35 ;
      RECT 37.685 4.213 37.69 4.351 ;
      RECT 37.67 4.215 37.685 4.353 ;
      RECT 37.665 4.215 37.67 4.356 ;
      RECT 37.6 4.222 37.665 4.363 ;
      RECT 37.565 4.232 37.595 4.373 ;
      RECT 37.548 4.235 37.565 4.375 ;
      RECT 37.462 4.234 37.548 4.374 ;
      RECT 37.376 4.232 37.462 4.371 ;
      RECT 37.29 4.231 37.376 4.369 ;
      RECT 37.189 4.229 37.255 4.368 ;
      RECT 37.103 4.226 37.189 4.366 ;
      RECT 37.017 4.222 37.103 4.364 ;
      RECT 36.931 4.219 37.017 4.363 ;
      RECT 36.845 4.216 36.931 4.361 ;
      RECT 36.745 4.215 36.83 4.358 ;
      RECT 36.695 4.213 36.745 4.356 ;
      RECT 36.675 4.21 36.695 4.354 ;
      RECT 36.655 4.208 36.675 4.351 ;
      RECT 36.63 4.204 36.655 4.348 ;
      RECT 36.585 4.198 36.63 4.343 ;
      RECT 36.545 4.192 36.585 4.335 ;
      RECT 36.52 4.187 36.545 4.328 ;
      RECT 36.465 4.18 36.52 4.32 ;
      RECT 36.441 4.173 36.465 4.313 ;
      RECT 36.355 4.164 36.441 4.303 ;
      RECT 36.325 4.156 36.355 4.293 ;
      RECT 36.295 4.152 36.325 4.288 ;
      RECT 36.29 4.149 36.295 4.285 ;
      RECT 36.285 4.148 36.29 4.285 ;
      RECT 36.21 4.141 36.285 4.278 ;
      RECT 36.171 4.132 36.21 4.267 ;
      RECT 36.085 4.122 36.171 4.255 ;
      RECT 36.045 4.112 36.085 4.243 ;
      RECT 36.006 4.107 36.045 4.236 ;
      RECT 35.92 4.097 36.006 4.225 ;
      RECT 35.88 4.085 35.92 4.214 ;
      RECT 35.845 4.07 35.88 4.207 ;
      RECT 35.835 4.06 35.845 4.204 ;
      RECT 35.815 4.045 35.835 4.202 ;
      RECT 35.785 4.015 35.815 4.198 ;
      RECT 35.775 3.995 35.785 4.193 ;
      RECT 35.77 3.987 35.775 4.19 ;
      RECT 35.765 3.98 35.77 4.188 ;
      RECT 35.75 3.967 35.765 4.181 ;
      RECT 35.745 3.957 35.75 4.173 ;
      RECT 35.74 3.95 35.745 4.168 ;
      RECT 35.735 3.945 35.74 4.164 ;
      RECT 35.72 3.932 35.735 4.156 ;
      RECT 35.715 3.842 35.72 4.145 ;
      RECT 35.71 3.837 35.715 4.138 ;
      RECT 35.635 3.835 35.71 4.098 ;
      RECT 35.605 3.835 35.635 4.053 ;
      RECT 35.51 3.84 35.525 4.04 ;
      RECT 37.995 3.545 38.255 3.805 ;
      RECT 37.98 3.533 38.16 3.77 ;
      RECT 37.975 3.534 38.16 3.768 ;
      RECT 37.96 3.538 38.17 3.758 ;
      RECT 37.955 3.543 38.175 3.728 ;
      RECT 37.96 3.54 38.175 3.758 ;
      RECT 37.975 3.535 38.17 3.768 ;
      RECT 37.995 3.532 38.16 3.805 ;
      RECT 37.995 3.531 38.15 3.805 ;
      RECT 38.02 3.53 38.15 3.805 ;
      RECT 37.58 3.775 37.84 4.035 ;
      RECT 37.455 3.82 37.84 4.03 ;
      RECT 37.445 3.825 37.84 4.025 ;
      RECT 37.46 4.765 37.475 5.075 ;
      RECT 36.055 4.535 36.065 4.665 ;
      RECT 35.835 4.53 35.94 4.665 ;
      RECT 35.75 4.535 35.8 4.665 ;
      RECT 34.3 3.27 34.305 4.375 ;
      RECT 37.555 4.857 37.56 4.993 ;
      RECT 37.55 4.852 37.555 5.053 ;
      RECT 37.545 4.85 37.55 5.066 ;
      RECT 37.53 4.847 37.545 5.068 ;
      RECT 37.525 4.842 37.53 5.07 ;
      RECT 37.52 4.838 37.525 5.073 ;
      RECT 37.505 4.833 37.52 5.075 ;
      RECT 37.475 4.825 37.505 5.075 ;
      RECT 37.436 4.765 37.46 5.075 ;
      RECT 37.35 4.765 37.436 5.072 ;
      RECT 37.32 4.765 37.35 5.065 ;
      RECT 37.295 4.765 37.32 5.058 ;
      RECT 37.27 4.765 37.295 5.05 ;
      RECT 37.255 4.765 37.27 5.043 ;
      RECT 37.23 4.765 37.255 5.035 ;
      RECT 37.215 4.765 37.23 5.028 ;
      RECT 37.175 4.775 37.215 5.017 ;
      RECT 37.165 4.77 37.175 5.007 ;
      RECT 37.161 4.769 37.165 5.004 ;
      RECT 37.075 4.761 37.161 4.987 ;
      RECT 37.042 4.75 37.075 4.964 ;
      RECT 36.956 4.739 37.042 4.942 ;
      RECT 36.87 4.723 36.956 4.911 ;
      RECT 36.8 4.708 36.87 4.883 ;
      RECT 36.79 4.701 36.8 4.87 ;
      RECT 36.76 4.698 36.79 4.86 ;
      RECT 36.735 4.694 36.76 4.853 ;
      RECT 36.72 4.691 36.735 4.848 ;
      RECT 36.715 4.69 36.72 4.843 ;
      RECT 36.685 4.685 36.715 4.836 ;
      RECT 36.68 4.68 36.685 4.831 ;
      RECT 36.665 4.677 36.68 4.826 ;
      RECT 36.66 4.672 36.665 4.821 ;
      RECT 36.64 4.667 36.66 4.818 ;
      RECT 36.625 4.662 36.64 4.81 ;
      RECT 36.61 4.656 36.625 4.805 ;
      RECT 36.58 4.647 36.61 4.798 ;
      RECT 36.575 4.64 36.58 4.79 ;
      RECT 36.57 4.638 36.575 4.788 ;
      RECT 36.565 4.637 36.57 4.785 ;
      RECT 36.525 4.63 36.565 4.778 ;
      RECT 36.511 4.62 36.525 4.768 ;
      RECT 36.46 4.609 36.511 4.756 ;
      RECT 36.435 4.595 36.46 4.742 ;
      RECT 36.41 4.584 36.435 4.734 ;
      RECT 36.39 4.573 36.41 4.728 ;
      RECT 36.38 4.567 36.39 4.723 ;
      RECT 36.375 4.565 36.38 4.719 ;
      RECT 36.355 4.56 36.375 4.714 ;
      RECT 36.325 4.55 36.355 4.704 ;
      RECT 36.32 4.542 36.325 4.697 ;
      RECT 36.305 4.54 36.32 4.693 ;
      RECT 36.285 4.54 36.305 4.688 ;
      RECT 36.28 4.539 36.285 4.686 ;
      RECT 36.275 4.539 36.28 4.683 ;
      RECT 36.235 4.538 36.275 4.678 ;
      RECT 36.21 4.537 36.235 4.673 ;
      RECT 36.15 4.536 36.21 4.67 ;
      RECT 36.065 4.535 36.15 4.668 ;
      RECT 36.026 4.534 36.055 4.665 ;
      RECT 35.94 4.532 36.026 4.665 ;
      RECT 35.8 4.532 35.835 4.665 ;
      RECT 35.71 4.536 35.75 4.668 ;
      RECT 35.695 4.539 35.71 4.675 ;
      RECT 35.685 4.54 35.695 4.682 ;
      RECT 35.66 4.543 35.685 4.687 ;
      RECT 35.655 4.545 35.66 4.69 ;
      RECT 35.605 4.547 35.655 4.691 ;
      RECT 35.566 4.551 35.605 4.693 ;
      RECT 35.48 4.553 35.566 4.696 ;
      RECT 35.462 4.555 35.48 4.698 ;
      RECT 35.376 4.558 35.462 4.7 ;
      RECT 35.29 4.562 35.376 4.703 ;
      RECT 35.253 4.566 35.29 4.706 ;
      RECT 35.167 4.569 35.253 4.709 ;
      RECT 35.081 4.573 35.167 4.712 ;
      RECT 34.995 4.578 35.081 4.716 ;
      RECT 34.975 4.58 34.995 4.719 ;
      RECT 34.955 4.579 34.975 4.72 ;
      RECT 34.906 4.576 34.955 4.721 ;
      RECT 34.82 4.571 34.906 4.724 ;
      RECT 34.77 4.566 34.82 4.726 ;
      RECT 34.746 4.564 34.77 4.727 ;
      RECT 34.66 4.559 34.746 4.729 ;
      RECT 34.635 4.555 34.66 4.728 ;
      RECT 34.625 4.552 34.635 4.726 ;
      RECT 34.615 4.545 34.625 4.723 ;
      RECT 34.61 4.525 34.615 4.718 ;
      RECT 34.6 4.495 34.61 4.713 ;
      RECT 34.585 4.365 34.6 4.704 ;
      RECT 34.58 4.357 34.585 4.697 ;
      RECT 34.56 4.35 34.58 4.689 ;
      RECT 34.555 4.332 34.56 4.681 ;
      RECT 34.545 4.312 34.555 4.676 ;
      RECT 34.54 4.285 34.545 4.672 ;
      RECT 34.535 4.262 34.54 4.669 ;
      RECT 34.515 4.22 34.535 4.661 ;
      RECT 34.48 4.135 34.515 4.645 ;
      RECT 34.475 4.067 34.48 4.633 ;
      RECT 34.46 4.037 34.475 4.627 ;
      RECT 34.455 3.282 34.46 3.528 ;
      RECT 34.445 4.007 34.46 4.618 ;
      RECT 34.45 3.277 34.455 3.56 ;
      RECT 34.445 3.272 34.45 3.603 ;
      RECT 34.44 3.27 34.445 3.638 ;
      RECT 34.425 3.97 34.445 4.608 ;
      RECT 34.435 3.27 34.44 3.675 ;
      RECT 34.42 3.27 34.435 3.773 ;
      RECT 34.42 3.943 34.425 4.601 ;
      RECT 34.415 3.27 34.42 3.848 ;
      RECT 34.415 3.931 34.42 4.598 ;
      RECT 34.41 3.27 34.415 3.88 ;
      RECT 34.41 3.91 34.415 4.595 ;
      RECT 34.405 3.27 34.41 4.592 ;
      RECT 34.37 3.27 34.405 4.578 ;
      RECT 34.355 3.27 34.37 4.56 ;
      RECT 34.335 3.27 34.355 4.55 ;
      RECT 34.31 3.27 34.335 4.533 ;
      RECT 34.305 3.27 34.31 4.483 ;
      RECT 34.295 3.27 34.3 4.313 ;
      RECT 34.29 3.27 34.295 4.22 ;
      RECT 34.285 3.27 34.29 4.133 ;
      RECT 34.28 3.27 34.285 4.065 ;
      RECT 34.275 3.27 34.28 4.008 ;
      RECT 34.265 3.27 34.275 3.903 ;
      RECT 34.26 3.27 34.265 3.775 ;
      RECT 34.255 3.27 34.26 3.693 ;
      RECT 34.25 3.272 34.255 3.61 ;
      RECT 34.245 3.277 34.25 3.543 ;
      RECT 34.24 3.282 34.245 3.47 ;
      RECT 37.055 3.6 37.315 3.86 ;
      RECT 37.075 3.567 37.285 3.86 ;
      RECT 37.075 3.565 37.275 3.86 ;
      RECT 37.085 3.552 37.275 3.86 ;
      RECT 37.085 3.55 37.2 3.86 ;
      RECT 36.56 3.675 36.735 3.955 ;
      RECT 36.555 3.675 36.735 3.953 ;
      RECT 36.555 3.675 36.75 3.95 ;
      RECT 36.545 3.675 36.75 3.948 ;
      RECT 36.49 3.675 36.75 3.935 ;
      RECT 36.49 3.75 36.755 3.913 ;
      RECT 36.035 3.687 36.055 3.93 ;
      RECT 36.035 3.687 36.095 3.929 ;
      RECT 36.03 3.689 36.095 3.928 ;
      RECT 36.03 3.689 36.181 3.927 ;
      RECT 36.03 3.689 36.25 3.926 ;
      RECT 36.03 3.689 36.27 3.918 ;
      RECT 36.01 3.692 36.27 3.916 ;
      RECT 35.995 3.702 36.27 3.901 ;
      RECT 35.995 3.702 36.285 3.9 ;
      RECT 35.99 3.711 36.285 3.892 ;
      RECT 35.99 3.711 36.29 3.888 ;
      RECT 36.095 3.625 36.355 3.885 ;
      RECT 35.985 3.713 36.355 3.77 ;
      RECT 36.055 3.68 36.355 3.885 ;
      RECT 36.02 4.873 36.025 5.08 ;
      RECT 35.97 4.867 36.02 5.079 ;
      RECT 35.937 4.881 36.03 5.078 ;
      RECT 35.851 4.881 36.03 5.077 ;
      RECT 35.765 4.881 36.03 5.076 ;
      RECT 35.765 4.98 36.035 5.073 ;
      RECT 35.76 4.98 36.035 5.068 ;
      RECT 35.755 4.98 36.035 5.05 ;
      RECT 35.75 4.98 36.035 5.033 ;
      RECT 35.71 4.765 35.97 5.025 ;
      RECT 35.17 3.915 35.256 4.329 ;
      RECT 35.17 3.915 35.295 4.326 ;
      RECT 35.17 3.915 35.315 4.316 ;
      RECT 35.125 3.915 35.315 4.313 ;
      RECT 35.125 4.067 35.325 4.303 ;
      RECT 35.125 4.088 35.33 4.297 ;
      RECT 35.125 4.106 35.335 4.293 ;
      RECT 35.125 4.126 35.345 4.288 ;
      RECT 35.1 4.126 35.345 4.285 ;
      RECT 35.09 4.126 35.345 4.263 ;
      RECT 35.09 4.142 35.35 4.233 ;
      RECT 35.055 3.915 35.315 4.22 ;
      RECT 35.055 4.154 35.355 4.175 ;
      RECT 32.715 10.06 33.005 10.29 ;
      RECT 32.775 8.58 32.945 10.29 ;
      RECT 32.765 8.95 33.12 9.305 ;
      RECT 32.715 8.58 33.005 8.81 ;
      RECT 32.31 3.69 32.415 4.26 ;
      RECT 32.31 4.025 32.635 4.255 ;
      RECT 32.31 4.055 32.805 4.225 ;
      RECT 32.31 3.69 32.5 4.255 ;
      RECT 31.725 3.655 32.015 3.885 ;
      RECT 31.725 3.69 32.5 3.86 ;
      RECT 31.785 2.175 31.955 3.885 ;
      RECT 31.725 2.175 32.015 2.405 ;
      RECT 31.725 10.06 32.015 10.29 ;
      RECT 31.785 8.58 31.955 10.29 ;
      RECT 31.725 8.58 32.015 8.81 ;
      RECT 31.725 8.615 32.575 8.775 ;
      RECT 32.41 8.21 32.575 8.775 ;
      RECT 31.725 8.61 32.12 8.775 ;
      RECT 32.345 8.21 32.635 8.44 ;
      RECT 32.345 8.24 32.805 8.41 ;
      RECT 31.355 4.025 31.645 4.255 ;
      RECT 31.355 4.055 31.815 4.225 ;
      RECT 31.42 2.95 31.585 4.255 ;
      RECT 29.935 2.92 30.225 3.15 ;
      RECT 29.935 2.95 31.585 3.12 ;
      RECT 29.995 2.18 30.165 3.15 ;
      RECT 29.935 2.18 30.225 2.41 ;
      RECT 29.935 10.055 30.225 10.285 ;
      RECT 29.995 9.315 30.165 10.285 ;
      RECT 29.995 9.41 31.585 9.58 ;
      RECT 31.415 8.21 31.585 9.58 ;
      RECT 29.935 9.315 30.225 9.545 ;
      RECT 31.355 8.21 31.645 8.44 ;
      RECT 31.355 8.24 31.815 8.41 ;
      RECT 27.985 4 28.325 4.35 ;
      RECT 28.075 3.32 28.245 4.35 ;
      RECT 30.365 3.26 30.715 3.61 ;
      RECT 28.075 3.32 30.715 3.49 ;
      RECT 30.39 8.945 30.715 9.27 ;
      RECT 24.93 8.9 25.28 9.25 ;
      RECT 30.365 8.945 30.715 9.175 ;
      RECT 24.73 8.945 25.28 9.175 ;
      RECT 24.56 8.975 30.715 9.145 ;
      RECT 29.59 3.66 29.91 3.98 ;
      RECT 29.56 3.66 29.91 3.89 ;
      RECT 29.39 3.69 29.91 3.86 ;
      RECT 29.59 8.545 29.91 8.835 ;
      RECT 29.56 8.575 29.91 8.805 ;
      RECT 29.39 8.605 29.91 8.775 ;
      RECT 25.28 4.28 25.43 4.555 ;
      RECT 25.82 3.36 25.825 3.58 ;
      RECT 26.97 3.56 26.985 3.758 ;
      RECT 26.935 3.552 26.97 3.765 ;
      RECT 26.905 3.545 26.935 3.765 ;
      RECT 26.85 3.51 26.905 3.765 ;
      RECT 26.785 3.447 26.85 3.765 ;
      RECT 26.78 3.412 26.785 3.763 ;
      RECT 26.775 3.407 26.78 3.755 ;
      RECT 26.77 3.402 26.775 3.741 ;
      RECT 26.765 3.399 26.77 3.734 ;
      RECT 26.72 3.389 26.765 3.685 ;
      RECT 26.7 3.376 26.72 3.62 ;
      RECT 26.695 3.371 26.7 3.593 ;
      RECT 26.69 3.37 26.695 3.586 ;
      RECT 26.685 3.369 26.69 3.579 ;
      RECT 26.6 3.354 26.685 3.525 ;
      RECT 26.57 3.335 26.6 3.475 ;
      RECT 26.49 3.318 26.57 3.46 ;
      RECT 26.455 3.305 26.49 3.445 ;
      RECT 26.447 3.305 26.455 3.44 ;
      RECT 26.361 3.306 26.447 3.44 ;
      RECT 26.275 3.308 26.361 3.44 ;
      RECT 26.25 3.309 26.275 3.444 ;
      RECT 26.175 3.315 26.25 3.459 ;
      RECT 26.092 3.327 26.175 3.483 ;
      RECT 26.006 3.34 26.092 3.509 ;
      RECT 25.92 3.353 26.006 3.535 ;
      RECT 25.885 3.362 25.92 3.554 ;
      RECT 25.835 3.362 25.885 3.567 ;
      RECT 25.825 3.36 25.835 3.578 ;
      RECT 25.81 3.357 25.82 3.58 ;
      RECT 25.795 3.349 25.81 3.588 ;
      RECT 25.78 3.341 25.795 3.608 ;
      RECT 25.775 3.336 25.78 3.665 ;
      RECT 25.76 3.331 25.775 3.738 ;
      RECT 25.755 3.326 25.76 3.78 ;
      RECT 25.75 3.324 25.755 3.808 ;
      RECT 25.745 3.322 25.75 3.83 ;
      RECT 25.735 3.318 25.745 3.873 ;
      RECT 25.73 3.315 25.735 3.898 ;
      RECT 25.725 3.313 25.73 3.918 ;
      RECT 25.72 3.311 25.725 3.942 ;
      RECT 25.715 3.307 25.72 3.965 ;
      RECT 25.71 3.303 25.715 3.988 ;
      RECT 25.675 3.293 25.71 4.095 ;
      RECT 25.67 3.283 25.675 4.193 ;
      RECT 25.665 3.281 25.67 4.22 ;
      RECT 25.66 3.28 25.665 4.24 ;
      RECT 25.655 3.272 25.66 4.26 ;
      RECT 25.65 3.267 25.655 4.295 ;
      RECT 25.645 3.265 25.65 4.313 ;
      RECT 25.64 3.265 25.645 4.338 ;
      RECT 25.635 3.265 25.64 4.36 ;
      RECT 25.6 3.265 25.635 4.403 ;
      RECT 25.575 3.265 25.6 4.432 ;
      RECT 25.565 3.265 25.575 3.618 ;
      RECT 25.568 3.675 25.575 4.442 ;
      RECT 25.565 3.732 25.568 4.445 ;
      RECT 25.56 3.265 25.565 3.59 ;
      RECT 25.56 3.782 25.565 4.448 ;
      RECT 25.55 3.265 25.56 3.58 ;
      RECT 25.555 3.835 25.56 4.451 ;
      RECT 25.55 3.92 25.555 4.455 ;
      RECT 25.54 3.265 25.55 3.568 ;
      RECT 25.545 3.967 25.55 4.459 ;
      RECT 25.54 4.042 25.545 4.463 ;
      RECT 25.505 3.265 25.54 3.543 ;
      RECT 25.53 4.125 25.54 4.468 ;
      RECT 25.52 4.192 25.53 4.475 ;
      RECT 25.515 4.22 25.52 4.48 ;
      RECT 25.505 4.233 25.515 4.486 ;
      RECT 25.46 3.265 25.505 3.5 ;
      RECT 25.5 4.238 25.505 4.493 ;
      RECT 25.46 4.255 25.5 4.555 ;
      RECT 25.455 3.267 25.46 3.473 ;
      RECT 25.43 4.275 25.46 4.555 ;
      RECT 25.45 3.272 25.455 3.445 ;
      RECT 25.24 4.284 25.28 4.555 ;
      RECT 25.215 4.292 25.24 4.525 ;
      RECT 25.17 4.3 25.215 4.525 ;
      RECT 25.155 4.305 25.17 4.52 ;
      RECT 25.145 4.305 25.155 4.514 ;
      RECT 25.135 4.312 25.145 4.511 ;
      RECT 25.13 4.35 25.135 4.5 ;
      RECT 25.125 4.412 25.13 4.478 ;
      RECT 26.395 4.287 26.58 4.51 ;
      RECT 26.395 4.302 26.585 4.506 ;
      RECT 26.385 3.575 26.47 4.505 ;
      RECT 26.385 4.302 26.59 4.499 ;
      RECT 26.38 4.31 26.59 4.498 ;
      RECT 26.585 4.03 26.905 4.35 ;
      RECT 26.38 4.202 26.55 4.293 ;
      RECT 26.375 4.202 26.55 4.275 ;
      RECT 26.365 4.01 26.5 4.25 ;
      RECT 26.36 4.01 26.5 4.195 ;
      RECT 26.32 3.59 26.49 4.095 ;
      RECT 26.305 3.59 26.49 3.965 ;
      RECT 26.3 3.59 26.49 3.918 ;
      RECT 26.295 3.59 26.49 3.898 ;
      RECT 26.29 3.59 26.49 3.873 ;
      RECT 26.26 3.59 26.52 3.85 ;
      RECT 26.27 3.587 26.48 3.85 ;
      RECT 26.395 3.582 26.48 4.51 ;
      RECT 26.28 3.575 26.47 3.85 ;
      RECT 26.275 3.58 26.47 3.85 ;
      RECT 25.105 3.792 25.29 4.005 ;
      RECT 25.105 3.8 25.3 3.998 ;
      RECT 25.085 3.8 25.3 3.995 ;
      RECT 25.08 3.8 25.3 3.98 ;
      RECT 25.01 3.715 25.27 3.975 ;
      RECT 25.01 3.86 25.305 3.888 ;
      RECT 24.665 4.315 24.925 4.575 ;
      RECT 24.69 4.26 24.885 4.575 ;
      RECT 24.685 4.009 24.865 4.303 ;
      RECT 24.685 4.015 24.875 4.303 ;
      RECT 24.665 4.017 24.875 4.248 ;
      RECT 24.66 4.027 24.875 4.115 ;
      RECT 24.69 4.007 24.865 4.575 ;
      RECT 24.776 4.005 24.865 4.575 ;
      RECT 24.635 3.225 24.67 3.595 ;
      RECT 24.425 3.335 24.43 3.595 ;
      RECT 24.67 3.232 24.685 3.595 ;
      RECT 24.56 3.225 24.635 3.673 ;
      RECT 24.55 3.225 24.56 3.758 ;
      RECT 24.525 3.225 24.55 3.793 ;
      RECT 24.485 3.225 24.525 3.861 ;
      RECT 24.475 3.232 24.485 3.913 ;
      RECT 24.445 3.335 24.475 3.954 ;
      RECT 24.44 3.335 24.445 3.993 ;
      RECT 24.43 3.335 24.44 4.013 ;
      RECT 24.425 3.63 24.43 4.05 ;
      RECT 24.42 3.647 24.425 4.07 ;
      RECT 24.405 3.71 24.42 4.11 ;
      RECT 24.4 3.753 24.405 4.145 ;
      RECT 24.395 3.761 24.4 4.158 ;
      RECT 24.385 3.775 24.395 4.18 ;
      RECT 24.36 3.81 24.385 4.245 ;
      RECT 24.35 3.845 24.36 4.308 ;
      RECT 24.33 3.875 24.35 4.369 ;
      RECT 24.315 3.911 24.33 4.436 ;
      RECT 24.305 3.939 24.315 4.475 ;
      RECT 24.295 3.961 24.305 4.495 ;
      RECT 24.29 3.971 24.295 4.506 ;
      RECT 24.285 3.98 24.29 4.509 ;
      RECT 24.275 3.998 24.285 4.513 ;
      RECT 24.265 4.016 24.275 4.514 ;
      RECT 24.24 4.055 24.265 4.511 ;
      RECT 24.22 4.097 24.24 4.508 ;
      RECT 24.205 4.135 24.22 4.507 ;
      RECT 24.17 4.17 24.205 4.504 ;
      RECT 24.165 4.192 24.17 4.502 ;
      RECT 24.1 4.232 24.165 4.499 ;
      RECT 24.095 4.272 24.1 4.495 ;
      RECT 24.08 4.282 24.095 4.486 ;
      RECT 24.07 4.402 24.08 4.471 ;
      RECT 24.55 4.815 24.56 5.075 ;
      RECT 24.55 4.818 24.57 5.074 ;
      RECT 24.54 4.808 24.55 5.073 ;
      RECT 24.53 4.823 24.61 5.069 ;
      RECT 24.515 4.802 24.53 5.067 ;
      RECT 24.49 4.827 24.615 5.063 ;
      RECT 24.475 4.787 24.49 5.058 ;
      RECT 24.475 4.829 24.625 5.057 ;
      RECT 24.475 4.837 24.64 5.05 ;
      RECT 24.415 4.774 24.475 5.04 ;
      RECT 24.405 4.761 24.415 5.022 ;
      RECT 24.38 4.751 24.405 5.012 ;
      RECT 24.375 4.741 24.38 5.004 ;
      RECT 24.31 4.837 24.64 4.986 ;
      RECT 24.225 4.837 24.64 4.948 ;
      RECT 24.115 4.665 24.375 4.925 ;
      RECT 24.49 4.795 24.515 5.063 ;
      RECT 24.53 4.805 24.54 5.069 ;
      RECT 24.115 4.813 24.555 4.925 ;
      RECT 24.3 10.055 24.59 10.285 ;
      RECT 24.36 9.315 24.53 10.285 ;
      RECT 24.26 9.345 24.63 9.715 ;
      RECT 24.3 9.315 24.59 9.715 ;
      RECT 23.33 4.57 23.36 4.87 ;
      RECT 23.105 4.555 23.11 4.83 ;
      RECT 22.905 4.555 23.06 4.815 ;
      RECT 24.205 3.27 24.235 3.53 ;
      RECT 24.195 3.27 24.205 3.638 ;
      RECT 24.175 3.27 24.195 3.648 ;
      RECT 24.16 3.27 24.175 3.66 ;
      RECT 24.105 3.27 24.16 3.71 ;
      RECT 24.09 3.27 24.105 3.758 ;
      RECT 24.06 3.27 24.09 3.793 ;
      RECT 24.005 3.27 24.06 3.855 ;
      RECT 23.985 3.27 24.005 3.923 ;
      RECT 23.98 3.27 23.985 3.953 ;
      RECT 23.975 3.27 23.98 3.965 ;
      RECT 23.97 3.387 23.975 3.983 ;
      RECT 23.95 3.405 23.97 4.008 ;
      RECT 23.93 3.432 23.95 4.058 ;
      RECT 23.925 3.452 23.93 4.089 ;
      RECT 23.92 3.46 23.925 4.106 ;
      RECT 23.905 3.486 23.92 4.135 ;
      RECT 23.89 3.528 23.905 4.17 ;
      RECT 23.885 3.557 23.89 4.193 ;
      RECT 23.88 3.572 23.885 4.206 ;
      RECT 23.875 3.595 23.88 4.217 ;
      RECT 23.865 3.615 23.875 4.235 ;
      RECT 23.855 3.645 23.865 4.258 ;
      RECT 23.85 3.667 23.855 4.278 ;
      RECT 23.845 3.682 23.85 4.293 ;
      RECT 23.83 3.712 23.845 4.32 ;
      RECT 23.825 3.742 23.83 4.346 ;
      RECT 23.82 3.76 23.825 4.358 ;
      RECT 23.81 3.79 23.82 4.377 ;
      RECT 23.8 3.815 23.81 4.402 ;
      RECT 23.795 3.835 23.8 4.421 ;
      RECT 23.79 3.852 23.795 4.434 ;
      RECT 23.78 3.878 23.79 4.453 ;
      RECT 23.77 3.916 23.78 4.48 ;
      RECT 23.765 3.942 23.77 4.5 ;
      RECT 23.76 3.952 23.765 4.51 ;
      RECT 23.755 3.965 23.76 4.525 ;
      RECT 23.75 3.98 23.755 4.535 ;
      RECT 23.745 4.002 23.75 4.55 ;
      RECT 23.74 4.02 23.745 4.561 ;
      RECT 23.735 4.03 23.74 4.572 ;
      RECT 23.73 4.038 23.735 4.584 ;
      RECT 23.725 4.046 23.73 4.595 ;
      RECT 23.72 4.072 23.725 4.608 ;
      RECT 23.71 4.1 23.72 4.621 ;
      RECT 23.705 4.13 23.71 4.63 ;
      RECT 23.7 4.145 23.705 4.637 ;
      RECT 23.685 4.17 23.7 4.644 ;
      RECT 23.68 4.192 23.685 4.65 ;
      RECT 23.675 4.217 23.68 4.653 ;
      RECT 23.666 4.245 23.675 4.657 ;
      RECT 23.66 4.262 23.666 4.662 ;
      RECT 23.655 4.28 23.66 4.666 ;
      RECT 23.65 4.292 23.655 4.669 ;
      RECT 23.645 4.313 23.65 4.673 ;
      RECT 23.64 4.331 23.645 4.676 ;
      RECT 23.635 4.345 23.64 4.679 ;
      RECT 23.63 4.362 23.635 4.682 ;
      RECT 23.625 4.375 23.63 4.685 ;
      RECT 23.6 4.412 23.625 4.693 ;
      RECT 23.595 4.457 23.6 4.702 ;
      RECT 23.59 4.485 23.595 4.705 ;
      RECT 23.58 4.505 23.59 4.709 ;
      RECT 23.575 4.525 23.58 4.714 ;
      RECT 23.57 4.54 23.575 4.717 ;
      RECT 23.55 4.55 23.57 4.724 ;
      RECT 23.485 4.557 23.55 4.75 ;
      RECT 23.45 4.56 23.485 4.778 ;
      RECT 23.435 4.563 23.45 4.793 ;
      RECT 23.425 4.564 23.435 4.808 ;
      RECT 23.415 4.565 23.425 4.825 ;
      RECT 23.41 4.565 23.415 4.84 ;
      RECT 23.405 4.565 23.41 4.848 ;
      RECT 23.39 4.566 23.405 4.863 ;
      RECT 23.36 4.568 23.39 4.87 ;
      RECT 23.25 4.575 23.33 4.87 ;
      RECT 23.205 4.58 23.25 4.87 ;
      RECT 23.195 4.581 23.205 4.86 ;
      RECT 23.185 4.582 23.195 4.853 ;
      RECT 23.165 4.584 23.185 4.848 ;
      RECT 23.155 4.555 23.165 4.843 ;
      RECT 23.11 4.555 23.155 4.835 ;
      RECT 23.08 4.555 23.105 4.825 ;
      RECT 23.06 4.555 23.08 4.818 ;
      RECT 23.34 3.355 23.6 3.615 ;
      RECT 23.22 3.37 23.23 3.535 ;
      RECT 23.205 3.37 23.21 3.53 ;
      RECT 20.57 3.21 20.755 3.5 ;
      RECT 22.385 3.335 22.4 3.49 ;
      RECT 20.535 3.21 20.56 3.47 ;
      RECT 22.95 3.26 22.955 3.402 ;
      RECT 22.865 3.255 22.89 3.395 ;
      RECT 23.265 3.372 23.34 3.565 ;
      RECT 23.25 3.37 23.265 3.548 ;
      RECT 23.23 3.37 23.25 3.54 ;
      RECT 23.21 3.37 23.22 3.533 ;
      RECT 23.165 3.365 23.205 3.523 ;
      RECT 23.125 3.34 23.165 3.508 ;
      RECT 23.11 3.315 23.125 3.498 ;
      RECT 23.105 3.309 23.11 3.496 ;
      RECT 23.07 3.301 23.105 3.479 ;
      RECT 23.065 3.294 23.07 3.467 ;
      RECT 23.045 3.289 23.065 3.455 ;
      RECT 23.035 3.283 23.045 3.44 ;
      RECT 23.015 3.278 23.035 3.425 ;
      RECT 23.005 3.273 23.015 3.418 ;
      RECT 23 3.271 23.005 3.413 ;
      RECT 22.995 3.27 23 3.41 ;
      RECT 22.955 3.265 22.995 3.406 ;
      RECT 22.935 3.259 22.95 3.401 ;
      RECT 22.9 3.256 22.935 3.398 ;
      RECT 22.89 3.255 22.9 3.396 ;
      RECT 22.83 3.255 22.865 3.393 ;
      RECT 22.785 3.255 22.83 3.393 ;
      RECT 22.735 3.255 22.785 3.396 ;
      RECT 22.72 3.257 22.735 3.398 ;
      RECT 22.705 3.26 22.72 3.399 ;
      RECT 22.695 3.265 22.705 3.4 ;
      RECT 22.665 3.27 22.695 3.405 ;
      RECT 22.655 3.276 22.665 3.413 ;
      RECT 22.645 3.278 22.655 3.417 ;
      RECT 22.635 3.282 22.645 3.421 ;
      RECT 22.61 3.288 22.635 3.429 ;
      RECT 22.6 3.293 22.61 3.437 ;
      RECT 22.585 3.297 22.6 3.441 ;
      RECT 22.55 3.303 22.585 3.449 ;
      RECT 22.53 3.308 22.55 3.459 ;
      RECT 22.5 3.315 22.53 3.468 ;
      RECT 22.455 3.324 22.5 3.482 ;
      RECT 22.45 3.329 22.455 3.493 ;
      RECT 22.43 3.332 22.45 3.494 ;
      RECT 22.4 3.335 22.43 3.492 ;
      RECT 22.365 3.335 22.385 3.488 ;
      RECT 22.295 3.335 22.365 3.479 ;
      RECT 22.28 3.332 22.295 3.471 ;
      RECT 22.24 3.325 22.28 3.466 ;
      RECT 22.215 3.315 22.24 3.459 ;
      RECT 22.21 3.309 22.215 3.456 ;
      RECT 22.17 3.303 22.21 3.453 ;
      RECT 22.155 3.296 22.17 3.448 ;
      RECT 22.135 3.292 22.155 3.443 ;
      RECT 22.12 3.287 22.135 3.439 ;
      RECT 22.105 3.282 22.12 3.437 ;
      RECT 22.09 3.278 22.105 3.436 ;
      RECT 22.075 3.276 22.09 3.432 ;
      RECT 22.065 3.274 22.075 3.427 ;
      RECT 22.05 3.271 22.065 3.423 ;
      RECT 22.04 3.269 22.05 3.418 ;
      RECT 22.02 3.266 22.04 3.414 ;
      RECT 21.975 3.265 22.02 3.412 ;
      RECT 21.915 3.267 21.975 3.413 ;
      RECT 21.895 3.269 21.915 3.415 ;
      RECT 21.865 3.272 21.895 3.416 ;
      RECT 21.815 3.277 21.865 3.418 ;
      RECT 21.81 3.28 21.815 3.42 ;
      RECT 21.8 3.282 21.81 3.423 ;
      RECT 21.795 3.284 21.8 3.426 ;
      RECT 21.745 3.287 21.795 3.433 ;
      RECT 21.725 3.291 21.745 3.445 ;
      RECT 21.715 3.294 21.725 3.451 ;
      RECT 21.705 3.295 21.715 3.454 ;
      RECT 21.666 3.298 21.705 3.456 ;
      RECT 21.58 3.305 21.666 3.459 ;
      RECT 21.506 3.315 21.58 3.463 ;
      RECT 21.42 3.326 21.506 3.468 ;
      RECT 21.405 3.333 21.42 3.47 ;
      RECT 21.35 3.337 21.405 3.471 ;
      RECT 21.336 3.34 21.35 3.473 ;
      RECT 21.25 3.34 21.336 3.475 ;
      RECT 21.21 3.337 21.25 3.478 ;
      RECT 21.186 3.333 21.21 3.48 ;
      RECT 21.1 3.323 21.186 3.483 ;
      RECT 21.07 3.312 21.1 3.484 ;
      RECT 21.051 3.308 21.07 3.483 ;
      RECT 20.965 3.301 21.051 3.48 ;
      RECT 20.905 3.29 20.965 3.477 ;
      RECT 20.885 3.282 20.905 3.475 ;
      RECT 20.85 3.277 20.885 3.474 ;
      RECT 20.825 3.272 20.85 3.473 ;
      RECT 20.795 3.267 20.825 3.472 ;
      RECT 20.77 3.21 20.795 3.471 ;
      RECT 20.755 3.21 20.77 3.495 ;
      RECT 20.56 3.21 20.57 3.495 ;
      RECT 22.335 4.23 22.34 4.37 ;
      RECT 21.995 4.23 22.03 4.368 ;
      RECT 21.57 4.215 21.585 4.36 ;
      RECT 23.4 3.995 23.49 4.255 ;
      RECT 23.23 3.86 23.33 4.255 ;
      RECT 20.265 3.835 20.345 4.045 ;
      RECT 23.355 3.972 23.4 4.255 ;
      RECT 23.345 3.942 23.355 4.255 ;
      RECT 23.33 3.865 23.345 4.255 ;
      RECT 23.145 3.86 23.23 4.22 ;
      RECT 23.14 3.862 23.145 4.215 ;
      RECT 23.135 3.867 23.14 4.215 ;
      RECT 23.1 3.967 23.135 4.215 ;
      RECT 23.09 3.995 23.1 4.215 ;
      RECT 23.08 4.01 23.09 4.215 ;
      RECT 23.07 4.022 23.08 4.215 ;
      RECT 23.065 4.032 23.07 4.215 ;
      RECT 23.05 4.042 23.065 4.217 ;
      RECT 23.045 4.057 23.05 4.219 ;
      RECT 23.03 4.07 23.045 4.221 ;
      RECT 23.025 4.085 23.03 4.224 ;
      RECT 23.005 4.095 23.025 4.228 ;
      RECT 22.99 4.105 23.005 4.231 ;
      RECT 22.955 4.112 22.99 4.236 ;
      RECT 22.911 4.119 22.955 4.244 ;
      RECT 22.825 4.131 22.911 4.257 ;
      RECT 22.8 4.142 22.825 4.268 ;
      RECT 22.77 4.147 22.8 4.273 ;
      RECT 22.735 4.152 22.77 4.281 ;
      RECT 22.705 4.157 22.735 4.288 ;
      RECT 22.68 4.162 22.705 4.293 ;
      RECT 22.615 4.169 22.68 4.302 ;
      RECT 22.545 4.182 22.615 4.318 ;
      RECT 22.515 4.192 22.545 4.33 ;
      RECT 22.49 4.197 22.515 4.337 ;
      RECT 22.435 4.204 22.49 4.345 ;
      RECT 22.43 4.211 22.435 4.35 ;
      RECT 22.425 4.213 22.43 4.351 ;
      RECT 22.41 4.215 22.425 4.353 ;
      RECT 22.405 4.215 22.41 4.356 ;
      RECT 22.34 4.222 22.405 4.363 ;
      RECT 22.305 4.232 22.335 4.373 ;
      RECT 22.288 4.235 22.305 4.375 ;
      RECT 22.202 4.234 22.288 4.374 ;
      RECT 22.116 4.232 22.202 4.371 ;
      RECT 22.03 4.231 22.116 4.369 ;
      RECT 21.929 4.229 21.995 4.368 ;
      RECT 21.843 4.226 21.929 4.366 ;
      RECT 21.757 4.222 21.843 4.364 ;
      RECT 21.671 4.219 21.757 4.363 ;
      RECT 21.585 4.216 21.671 4.361 ;
      RECT 21.485 4.215 21.57 4.358 ;
      RECT 21.435 4.213 21.485 4.356 ;
      RECT 21.415 4.21 21.435 4.354 ;
      RECT 21.395 4.208 21.415 4.351 ;
      RECT 21.37 4.204 21.395 4.348 ;
      RECT 21.325 4.198 21.37 4.343 ;
      RECT 21.285 4.192 21.325 4.335 ;
      RECT 21.26 4.187 21.285 4.328 ;
      RECT 21.205 4.18 21.26 4.32 ;
      RECT 21.181 4.173 21.205 4.313 ;
      RECT 21.095 4.164 21.181 4.303 ;
      RECT 21.065 4.156 21.095 4.293 ;
      RECT 21.035 4.152 21.065 4.288 ;
      RECT 21.03 4.149 21.035 4.285 ;
      RECT 21.025 4.148 21.03 4.285 ;
      RECT 20.95 4.141 21.025 4.278 ;
      RECT 20.911 4.132 20.95 4.267 ;
      RECT 20.825 4.122 20.911 4.255 ;
      RECT 20.785 4.112 20.825 4.243 ;
      RECT 20.746 4.107 20.785 4.236 ;
      RECT 20.66 4.097 20.746 4.225 ;
      RECT 20.62 4.085 20.66 4.214 ;
      RECT 20.585 4.07 20.62 4.207 ;
      RECT 20.575 4.06 20.585 4.204 ;
      RECT 20.555 4.045 20.575 4.202 ;
      RECT 20.525 4.015 20.555 4.198 ;
      RECT 20.515 3.995 20.525 4.193 ;
      RECT 20.51 3.987 20.515 4.19 ;
      RECT 20.505 3.98 20.51 4.188 ;
      RECT 20.49 3.967 20.505 4.181 ;
      RECT 20.485 3.957 20.49 4.173 ;
      RECT 20.48 3.95 20.485 4.168 ;
      RECT 20.475 3.945 20.48 4.164 ;
      RECT 20.46 3.932 20.475 4.156 ;
      RECT 20.455 3.842 20.46 4.145 ;
      RECT 20.45 3.837 20.455 4.138 ;
      RECT 20.375 3.835 20.45 4.098 ;
      RECT 20.345 3.835 20.375 4.053 ;
      RECT 20.25 3.84 20.265 4.04 ;
      RECT 22.735 3.545 22.995 3.805 ;
      RECT 22.72 3.533 22.9 3.77 ;
      RECT 22.715 3.534 22.9 3.768 ;
      RECT 22.7 3.538 22.91 3.758 ;
      RECT 22.695 3.543 22.915 3.728 ;
      RECT 22.7 3.54 22.915 3.758 ;
      RECT 22.715 3.535 22.91 3.768 ;
      RECT 22.735 3.532 22.9 3.805 ;
      RECT 22.735 3.531 22.89 3.805 ;
      RECT 22.76 3.53 22.89 3.805 ;
      RECT 22.32 3.775 22.58 4.035 ;
      RECT 22.195 3.82 22.58 4.03 ;
      RECT 22.185 3.825 22.58 4.025 ;
      RECT 22.2 4.765 22.215 5.075 ;
      RECT 20.795 4.535 20.805 4.665 ;
      RECT 20.575 4.53 20.68 4.665 ;
      RECT 20.49 4.535 20.54 4.665 ;
      RECT 19.04 3.27 19.045 4.375 ;
      RECT 22.295 4.857 22.3 4.993 ;
      RECT 22.29 4.852 22.295 5.053 ;
      RECT 22.285 4.85 22.29 5.066 ;
      RECT 22.27 4.847 22.285 5.068 ;
      RECT 22.265 4.842 22.27 5.07 ;
      RECT 22.26 4.838 22.265 5.073 ;
      RECT 22.245 4.833 22.26 5.075 ;
      RECT 22.215 4.825 22.245 5.075 ;
      RECT 22.176 4.765 22.2 5.075 ;
      RECT 22.09 4.765 22.176 5.072 ;
      RECT 22.06 4.765 22.09 5.065 ;
      RECT 22.035 4.765 22.06 5.058 ;
      RECT 22.01 4.765 22.035 5.05 ;
      RECT 21.995 4.765 22.01 5.043 ;
      RECT 21.97 4.765 21.995 5.035 ;
      RECT 21.955 4.765 21.97 5.028 ;
      RECT 21.915 4.775 21.955 5.017 ;
      RECT 21.905 4.77 21.915 5.007 ;
      RECT 21.901 4.769 21.905 5.004 ;
      RECT 21.815 4.761 21.901 4.987 ;
      RECT 21.782 4.75 21.815 4.964 ;
      RECT 21.696 4.739 21.782 4.942 ;
      RECT 21.61 4.723 21.696 4.911 ;
      RECT 21.54 4.708 21.61 4.883 ;
      RECT 21.53 4.701 21.54 4.87 ;
      RECT 21.5 4.698 21.53 4.86 ;
      RECT 21.475 4.694 21.5 4.853 ;
      RECT 21.46 4.691 21.475 4.848 ;
      RECT 21.455 4.69 21.46 4.843 ;
      RECT 21.425 4.685 21.455 4.836 ;
      RECT 21.42 4.68 21.425 4.831 ;
      RECT 21.405 4.677 21.42 4.826 ;
      RECT 21.4 4.672 21.405 4.821 ;
      RECT 21.38 4.667 21.4 4.818 ;
      RECT 21.365 4.662 21.38 4.81 ;
      RECT 21.35 4.656 21.365 4.805 ;
      RECT 21.32 4.647 21.35 4.798 ;
      RECT 21.315 4.64 21.32 4.79 ;
      RECT 21.31 4.638 21.315 4.788 ;
      RECT 21.305 4.637 21.31 4.785 ;
      RECT 21.265 4.63 21.305 4.778 ;
      RECT 21.251 4.62 21.265 4.768 ;
      RECT 21.2 4.609 21.251 4.756 ;
      RECT 21.175 4.595 21.2 4.742 ;
      RECT 21.15 4.584 21.175 4.734 ;
      RECT 21.13 4.573 21.15 4.728 ;
      RECT 21.12 4.567 21.13 4.723 ;
      RECT 21.115 4.565 21.12 4.719 ;
      RECT 21.095 4.56 21.115 4.714 ;
      RECT 21.065 4.55 21.095 4.704 ;
      RECT 21.06 4.542 21.065 4.697 ;
      RECT 21.045 4.54 21.06 4.693 ;
      RECT 21.025 4.54 21.045 4.688 ;
      RECT 21.02 4.539 21.025 4.686 ;
      RECT 21.015 4.539 21.02 4.683 ;
      RECT 20.975 4.538 21.015 4.678 ;
      RECT 20.95 4.537 20.975 4.673 ;
      RECT 20.89 4.536 20.95 4.67 ;
      RECT 20.805 4.535 20.89 4.668 ;
      RECT 20.766 4.534 20.795 4.665 ;
      RECT 20.68 4.532 20.766 4.665 ;
      RECT 20.54 4.532 20.575 4.665 ;
      RECT 20.45 4.536 20.49 4.668 ;
      RECT 20.435 4.539 20.45 4.675 ;
      RECT 20.425 4.54 20.435 4.682 ;
      RECT 20.4 4.543 20.425 4.687 ;
      RECT 20.395 4.545 20.4 4.69 ;
      RECT 20.345 4.547 20.395 4.691 ;
      RECT 20.306 4.551 20.345 4.693 ;
      RECT 20.22 4.553 20.306 4.696 ;
      RECT 20.202 4.555 20.22 4.698 ;
      RECT 20.116 4.558 20.202 4.7 ;
      RECT 20.03 4.562 20.116 4.703 ;
      RECT 19.993 4.566 20.03 4.706 ;
      RECT 19.907 4.569 19.993 4.709 ;
      RECT 19.821 4.573 19.907 4.712 ;
      RECT 19.735 4.578 19.821 4.716 ;
      RECT 19.715 4.58 19.735 4.719 ;
      RECT 19.695 4.579 19.715 4.72 ;
      RECT 19.646 4.576 19.695 4.721 ;
      RECT 19.56 4.571 19.646 4.724 ;
      RECT 19.51 4.566 19.56 4.726 ;
      RECT 19.486 4.564 19.51 4.727 ;
      RECT 19.4 4.559 19.486 4.729 ;
      RECT 19.375 4.555 19.4 4.728 ;
      RECT 19.365 4.552 19.375 4.726 ;
      RECT 19.355 4.545 19.365 4.723 ;
      RECT 19.35 4.525 19.355 4.718 ;
      RECT 19.34 4.495 19.35 4.713 ;
      RECT 19.325 4.365 19.34 4.704 ;
      RECT 19.32 4.357 19.325 4.697 ;
      RECT 19.3 4.35 19.32 4.689 ;
      RECT 19.295 4.332 19.3 4.681 ;
      RECT 19.285 4.312 19.295 4.676 ;
      RECT 19.28 4.285 19.285 4.672 ;
      RECT 19.275 4.262 19.28 4.669 ;
      RECT 19.255 4.22 19.275 4.661 ;
      RECT 19.22 4.135 19.255 4.645 ;
      RECT 19.215 4.067 19.22 4.633 ;
      RECT 19.2 4.037 19.215 4.627 ;
      RECT 19.195 3.282 19.2 3.528 ;
      RECT 19.185 4.007 19.2 4.618 ;
      RECT 19.19 3.277 19.195 3.56 ;
      RECT 19.185 3.272 19.19 3.603 ;
      RECT 19.18 3.27 19.185 3.638 ;
      RECT 19.165 3.97 19.185 4.608 ;
      RECT 19.175 3.27 19.18 3.675 ;
      RECT 19.16 3.27 19.175 3.773 ;
      RECT 19.16 3.943 19.165 4.601 ;
      RECT 19.155 3.27 19.16 3.848 ;
      RECT 19.155 3.931 19.16 4.598 ;
      RECT 19.15 3.27 19.155 3.88 ;
      RECT 19.15 3.91 19.155 4.595 ;
      RECT 19.145 3.27 19.15 4.592 ;
      RECT 19.11 3.27 19.145 4.578 ;
      RECT 19.095 3.27 19.11 4.56 ;
      RECT 19.075 3.27 19.095 4.55 ;
      RECT 19.05 3.27 19.075 4.533 ;
      RECT 19.045 3.27 19.05 4.483 ;
      RECT 19.035 3.27 19.04 4.313 ;
      RECT 19.03 3.27 19.035 4.22 ;
      RECT 19.025 3.27 19.03 4.133 ;
      RECT 19.02 3.27 19.025 4.065 ;
      RECT 19.015 3.27 19.02 4.008 ;
      RECT 19.005 3.27 19.015 3.903 ;
      RECT 19 3.27 19.005 3.775 ;
      RECT 18.995 3.27 19 3.693 ;
      RECT 18.99 3.272 18.995 3.61 ;
      RECT 18.985 3.277 18.99 3.543 ;
      RECT 18.98 3.282 18.985 3.47 ;
      RECT 21.795 3.6 22.055 3.86 ;
      RECT 21.815 3.567 22.025 3.86 ;
      RECT 21.815 3.565 22.015 3.86 ;
      RECT 21.825 3.552 22.015 3.86 ;
      RECT 21.825 3.55 21.94 3.86 ;
      RECT 21.3 3.675 21.475 3.955 ;
      RECT 21.295 3.675 21.475 3.953 ;
      RECT 21.295 3.675 21.49 3.95 ;
      RECT 21.285 3.675 21.49 3.948 ;
      RECT 21.23 3.675 21.49 3.935 ;
      RECT 21.23 3.75 21.495 3.913 ;
      RECT 20.775 3.687 20.795 3.93 ;
      RECT 20.775 3.687 20.835 3.929 ;
      RECT 20.77 3.689 20.835 3.928 ;
      RECT 20.77 3.689 20.921 3.927 ;
      RECT 20.77 3.689 20.99 3.926 ;
      RECT 20.77 3.689 21.01 3.918 ;
      RECT 20.75 3.692 21.01 3.916 ;
      RECT 20.735 3.702 21.01 3.901 ;
      RECT 20.735 3.702 21.025 3.9 ;
      RECT 20.73 3.711 21.025 3.892 ;
      RECT 20.73 3.711 21.03 3.888 ;
      RECT 20.835 3.625 21.095 3.885 ;
      RECT 20.725 3.713 21.095 3.77 ;
      RECT 20.795 3.68 21.095 3.885 ;
      RECT 20.76 4.873 20.765 5.08 ;
      RECT 20.71 4.867 20.76 5.079 ;
      RECT 20.677 4.881 20.77 5.078 ;
      RECT 20.591 4.881 20.77 5.077 ;
      RECT 20.505 4.881 20.77 5.076 ;
      RECT 20.505 4.98 20.775 5.073 ;
      RECT 20.5 4.98 20.775 5.068 ;
      RECT 20.495 4.98 20.775 5.05 ;
      RECT 20.49 4.98 20.775 5.033 ;
      RECT 20.45 4.765 20.71 5.025 ;
      RECT 19.91 3.915 19.996 4.329 ;
      RECT 19.91 3.915 20.035 4.326 ;
      RECT 19.91 3.915 20.055 4.316 ;
      RECT 19.865 3.915 20.055 4.313 ;
      RECT 19.865 4.067 20.065 4.303 ;
      RECT 19.865 4.088 20.07 4.297 ;
      RECT 19.865 4.106 20.075 4.293 ;
      RECT 19.865 4.126 20.085 4.288 ;
      RECT 19.84 4.126 20.085 4.285 ;
      RECT 19.83 4.126 20.085 4.263 ;
      RECT 19.83 4.142 20.09 4.233 ;
      RECT 19.795 3.915 20.055 4.22 ;
      RECT 19.795 4.154 20.095 4.175 ;
      RECT 17.455 10.06 17.745 10.29 ;
      RECT 17.515 8.58 17.685 10.29 ;
      RECT 17.51 8.945 17.86 9.295 ;
      RECT 17.455 8.58 17.745 8.81 ;
      RECT 17.05 3.69 17.155 4.26 ;
      RECT 17.05 4.025 17.375 4.255 ;
      RECT 17.05 4.055 17.545 4.225 ;
      RECT 17.05 3.69 17.24 4.255 ;
      RECT 16.465 3.655 16.755 3.885 ;
      RECT 16.465 3.69 17.24 3.86 ;
      RECT 16.525 2.175 16.695 3.885 ;
      RECT 16.465 2.175 16.755 2.405 ;
      RECT 16.465 10.06 16.755 10.29 ;
      RECT 16.525 8.58 16.695 10.29 ;
      RECT 16.465 8.58 16.755 8.81 ;
      RECT 16.465 8.615 17.315 8.775 ;
      RECT 17.15 8.21 17.315 8.775 ;
      RECT 16.465 8.61 16.86 8.775 ;
      RECT 17.085 8.21 17.375 8.44 ;
      RECT 17.085 8.24 17.545 8.41 ;
      RECT 16.095 4.025 16.385 4.255 ;
      RECT 16.095 4.055 16.555 4.225 ;
      RECT 16.16 2.95 16.325 4.255 ;
      RECT 14.675 2.92 14.965 3.15 ;
      RECT 14.675 2.95 16.325 3.12 ;
      RECT 14.735 2.18 14.905 3.15 ;
      RECT 14.675 2.18 14.965 2.41 ;
      RECT 14.675 10.055 14.965 10.285 ;
      RECT 14.735 9.315 14.905 10.285 ;
      RECT 14.735 9.41 16.325 9.58 ;
      RECT 16.155 8.21 16.325 9.58 ;
      RECT 14.675 9.315 14.965 9.545 ;
      RECT 16.095 8.21 16.385 8.44 ;
      RECT 16.095 8.24 16.555 8.41 ;
      RECT 12.725 4 13.065 4.35 ;
      RECT 12.815 3.32 12.985 4.35 ;
      RECT 15.105 3.26 15.455 3.61 ;
      RECT 12.815 3.32 15.455 3.49 ;
      RECT 15.13 8.945 15.455 9.27 ;
      RECT 9.67 8.895 10.02 9.245 ;
      RECT 15.105 8.945 15.455 9.175 ;
      RECT 9.47 8.945 10.02 9.175 ;
      RECT 9.3 8.975 15.455 9.145 ;
      RECT 14.33 3.66 14.65 3.98 ;
      RECT 14.3 3.66 14.65 3.89 ;
      RECT 14.13 3.69 14.65 3.86 ;
      RECT 14.33 8.545 14.65 8.835 ;
      RECT 14.3 8.575 14.65 8.805 ;
      RECT 14.13 8.605 14.65 8.775 ;
      RECT 10.02 4.28 10.17 4.555 ;
      RECT 10.56 3.36 10.565 3.58 ;
      RECT 11.71 3.56 11.725 3.758 ;
      RECT 11.675 3.552 11.71 3.765 ;
      RECT 11.645 3.545 11.675 3.765 ;
      RECT 11.59 3.51 11.645 3.765 ;
      RECT 11.525 3.447 11.59 3.765 ;
      RECT 11.52 3.412 11.525 3.763 ;
      RECT 11.515 3.407 11.52 3.755 ;
      RECT 11.51 3.402 11.515 3.741 ;
      RECT 11.505 3.399 11.51 3.734 ;
      RECT 11.46 3.389 11.505 3.685 ;
      RECT 11.44 3.376 11.46 3.62 ;
      RECT 11.435 3.371 11.44 3.593 ;
      RECT 11.43 3.37 11.435 3.586 ;
      RECT 11.425 3.369 11.43 3.579 ;
      RECT 11.34 3.354 11.425 3.525 ;
      RECT 11.31 3.335 11.34 3.475 ;
      RECT 11.23 3.318 11.31 3.46 ;
      RECT 11.195 3.305 11.23 3.445 ;
      RECT 11.187 3.305 11.195 3.44 ;
      RECT 11.101 3.306 11.187 3.44 ;
      RECT 11.015 3.308 11.101 3.44 ;
      RECT 10.99 3.309 11.015 3.444 ;
      RECT 10.915 3.315 10.99 3.459 ;
      RECT 10.832 3.327 10.915 3.483 ;
      RECT 10.746 3.34 10.832 3.509 ;
      RECT 10.66 3.353 10.746 3.535 ;
      RECT 10.625 3.362 10.66 3.554 ;
      RECT 10.575 3.362 10.625 3.567 ;
      RECT 10.565 3.36 10.575 3.578 ;
      RECT 10.55 3.357 10.56 3.58 ;
      RECT 10.535 3.349 10.55 3.588 ;
      RECT 10.52 3.341 10.535 3.608 ;
      RECT 10.515 3.336 10.52 3.665 ;
      RECT 10.5 3.331 10.515 3.738 ;
      RECT 10.495 3.326 10.5 3.78 ;
      RECT 10.49 3.324 10.495 3.808 ;
      RECT 10.485 3.322 10.49 3.83 ;
      RECT 10.475 3.318 10.485 3.873 ;
      RECT 10.47 3.315 10.475 3.898 ;
      RECT 10.465 3.313 10.47 3.918 ;
      RECT 10.46 3.311 10.465 3.942 ;
      RECT 10.455 3.307 10.46 3.965 ;
      RECT 10.45 3.303 10.455 3.988 ;
      RECT 10.415 3.293 10.45 4.095 ;
      RECT 10.41 3.283 10.415 4.193 ;
      RECT 10.405 3.281 10.41 4.22 ;
      RECT 10.4 3.28 10.405 4.24 ;
      RECT 10.395 3.272 10.4 4.26 ;
      RECT 10.39 3.267 10.395 4.295 ;
      RECT 10.385 3.265 10.39 4.313 ;
      RECT 10.38 3.265 10.385 4.338 ;
      RECT 10.375 3.265 10.38 4.36 ;
      RECT 10.34 3.265 10.375 4.403 ;
      RECT 10.315 3.265 10.34 4.432 ;
      RECT 10.305 3.265 10.315 3.618 ;
      RECT 10.308 3.675 10.315 4.442 ;
      RECT 10.305 3.732 10.308 4.445 ;
      RECT 10.3 3.265 10.305 3.59 ;
      RECT 10.3 3.782 10.305 4.448 ;
      RECT 10.29 3.265 10.3 3.58 ;
      RECT 10.295 3.835 10.3 4.451 ;
      RECT 10.29 3.92 10.295 4.455 ;
      RECT 10.28 3.265 10.29 3.568 ;
      RECT 10.285 3.967 10.29 4.459 ;
      RECT 10.28 4.042 10.285 4.463 ;
      RECT 10.245 3.265 10.28 3.543 ;
      RECT 10.27 4.125 10.28 4.468 ;
      RECT 10.26 4.192 10.27 4.475 ;
      RECT 10.255 4.22 10.26 4.48 ;
      RECT 10.245 4.233 10.255 4.486 ;
      RECT 10.2 3.265 10.245 3.5 ;
      RECT 10.24 4.238 10.245 4.493 ;
      RECT 10.2 4.255 10.24 4.555 ;
      RECT 10.195 3.267 10.2 3.473 ;
      RECT 10.17 4.275 10.2 4.555 ;
      RECT 10.19 3.272 10.195 3.445 ;
      RECT 9.98 4.284 10.02 4.555 ;
      RECT 9.955 4.292 9.98 4.525 ;
      RECT 9.91 4.3 9.955 4.525 ;
      RECT 9.895 4.305 9.91 4.52 ;
      RECT 9.885 4.305 9.895 4.514 ;
      RECT 9.875 4.312 9.885 4.511 ;
      RECT 9.87 4.35 9.875 4.5 ;
      RECT 9.865 4.412 9.87 4.478 ;
      RECT 11.135 4.287 11.32 4.51 ;
      RECT 11.135 4.302 11.325 4.506 ;
      RECT 11.125 3.575 11.21 4.505 ;
      RECT 11.125 4.302 11.33 4.499 ;
      RECT 11.12 4.31 11.33 4.498 ;
      RECT 11.325 4.03 11.645 4.35 ;
      RECT 11.12 4.202 11.29 4.293 ;
      RECT 11.115 4.202 11.29 4.275 ;
      RECT 11.105 4.01 11.24 4.25 ;
      RECT 11.1 4.01 11.24 4.195 ;
      RECT 11.06 3.59 11.23 4.095 ;
      RECT 11.045 3.59 11.23 3.965 ;
      RECT 11.04 3.59 11.23 3.918 ;
      RECT 11.035 3.59 11.23 3.898 ;
      RECT 11.03 3.59 11.23 3.873 ;
      RECT 11 3.59 11.26 3.85 ;
      RECT 11.01 3.587 11.22 3.85 ;
      RECT 11.135 3.582 11.22 4.51 ;
      RECT 11.02 3.575 11.21 3.85 ;
      RECT 11.015 3.58 11.21 3.85 ;
      RECT 9.845 3.792 10.03 4.005 ;
      RECT 9.845 3.8 10.04 3.998 ;
      RECT 9.825 3.8 10.04 3.995 ;
      RECT 9.82 3.8 10.04 3.98 ;
      RECT 9.75 3.715 10.01 3.975 ;
      RECT 9.75 3.86 10.045 3.888 ;
      RECT 9.405 4.315 9.665 4.575 ;
      RECT 9.43 4.26 9.625 4.575 ;
      RECT 9.425 4.009 9.605 4.303 ;
      RECT 9.425 4.015 9.615 4.303 ;
      RECT 9.405 4.017 9.615 4.248 ;
      RECT 9.4 4.027 9.615 4.115 ;
      RECT 9.43 4.007 9.605 4.575 ;
      RECT 9.516 4.005 9.605 4.575 ;
      RECT 9.375 3.225 9.41 3.595 ;
      RECT 9.165 3.335 9.17 3.595 ;
      RECT 9.41 3.232 9.425 3.595 ;
      RECT 9.3 3.225 9.375 3.673 ;
      RECT 9.29 3.225 9.3 3.758 ;
      RECT 9.265 3.225 9.29 3.793 ;
      RECT 9.225 3.225 9.265 3.861 ;
      RECT 9.215 3.232 9.225 3.913 ;
      RECT 9.185 3.335 9.215 3.954 ;
      RECT 9.18 3.335 9.185 3.993 ;
      RECT 9.17 3.335 9.18 4.013 ;
      RECT 9.165 3.63 9.17 4.05 ;
      RECT 9.16 3.647 9.165 4.07 ;
      RECT 9.145 3.71 9.16 4.11 ;
      RECT 9.14 3.753 9.145 4.145 ;
      RECT 9.135 3.761 9.14 4.158 ;
      RECT 9.125 3.775 9.135 4.18 ;
      RECT 9.1 3.81 9.125 4.245 ;
      RECT 9.09 3.845 9.1 4.308 ;
      RECT 9.07 3.875 9.09 4.369 ;
      RECT 9.055 3.911 9.07 4.436 ;
      RECT 9.045 3.939 9.055 4.475 ;
      RECT 9.035 3.961 9.045 4.495 ;
      RECT 9.03 3.971 9.035 4.506 ;
      RECT 9.025 3.98 9.03 4.509 ;
      RECT 9.015 3.998 9.025 4.513 ;
      RECT 9.005 4.016 9.015 4.514 ;
      RECT 8.98 4.055 9.005 4.511 ;
      RECT 8.96 4.097 8.98 4.508 ;
      RECT 8.945 4.135 8.96 4.507 ;
      RECT 8.91 4.17 8.945 4.504 ;
      RECT 8.905 4.192 8.91 4.502 ;
      RECT 8.84 4.232 8.905 4.499 ;
      RECT 8.835 4.272 8.84 4.495 ;
      RECT 8.82 4.282 8.835 4.486 ;
      RECT 8.81 4.402 8.82 4.471 ;
      RECT 9.29 4.815 9.3 5.075 ;
      RECT 9.29 4.818 9.31 5.074 ;
      RECT 9.28 4.808 9.29 5.073 ;
      RECT 9.27 4.823 9.35 5.069 ;
      RECT 9.255 4.802 9.27 5.067 ;
      RECT 9.23 4.827 9.355 5.063 ;
      RECT 9.215 4.787 9.23 5.058 ;
      RECT 9.215 4.829 9.365 5.057 ;
      RECT 9.215 4.837 9.38 5.05 ;
      RECT 9.155 4.774 9.215 5.04 ;
      RECT 9.145 4.761 9.155 5.022 ;
      RECT 9.12 4.751 9.145 5.012 ;
      RECT 9.115 4.741 9.12 5.004 ;
      RECT 9.05 4.837 9.38 4.986 ;
      RECT 8.965 4.837 9.38 4.948 ;
      RECT 8.855 4.665 9.115 4.925 ;
      RECT 9.23 4.795 9.255 5.063 ;
      RECT 9.27 4.805 9.28 5.069 ;
      RECT 8.855 4.813 9.295 4.925 ;
      RECT 9.04 10.055 9.33 10.285 ;
      RECT 9.1 9.315 9.27 10.285 ;
      RECT 9 9.345 9.37 9.715 ;
      RECT 9.04 9.315 9.33 9.715 ;
      RECT 8.07 4.57 8.1 4.87 ;
      RECT 7.845 4.555 7.85 4.83 ;
      RECT 7.645 4.555 7.8 4.815 ;
      RECT 8.945 3.27 8.975 3.53 ;
      RECT 8.935 3.27 8.945 3.638 ;
      RECT 8.915 3.27 8.935 3.648 ;
      RECT 8.9 3.27 8.915 3.66 ;
      RECT 8.845 3.27 8.9 3.71 ;
      RECT 8.83 3.27 8.845 3.758 ;
      RECT 8.8 3.27 8.83 3.793 ;
      RECT 8.745 3.27 8.8 3.855 ;
      RECT 8.725 3.27 8.745 3.923 ;
      RECT 8.72 3.27 8.725 3.953 ;
      RECT 8.715 3.27 8.72 3.965 ;
      RECT 8.71 3.387 8.715 3.983 ;
      RECT 8.69 3.405 8.71 4.008 ;
      RECT 8.67 3.432 8.69 4.058 ;
      RECT 8.665 3.452 8.67 4.089 ;
      RECT 8.66 3.46 8.665 4.106 ;
      RECT 8.645 3.486 8.66 4.135 ;
      RECT 8.63 3.528 8.645 4.17 ;
      RECT 8.625 3.557 8.63 4.193 ;
      RECT 8.62 3.572 8.625 4.206 ;
      RECT 8.615 3.595 8.62 4.217 ;
      RECT 8.605 3.615 8.615 4.235 ;
      RECT 8.595 3.645 8.605 4.258 ;
      RECT 8.59 3.667 8.595 4.278 ;
      RECT 8.585 3.682 8.59 4.293 ;
      RECT 8.57 3.712 8.585 4.32 ;
      RECT 8.565 3.742 8.57 4.346 ;
      RECT 8.56 3.76 8.565 4.358 ;
      RECT 8.55 3.79 8.56 4.377 ;
      RECT 8.54 3.815 8.55 4.402 ;
      RECT 8.535 3.835 8.54 4.421 ;
      RECT 8.53 3.852 8.535 4.434 ;
      RECT 8.52 3.878 8.53 4.453 ;
      RECT 8.51 3.916 8.52 4.48 ;
      RECT 8.505 3.942 8.51 4.5 ;
      RECT 8.5 3.952 8.505 4.51 ;
      RECT 8.495 3.965 8.5 4.525 ;
      RECT 8.49 3.98 8.495 4.535 ;
      RECT 8.485 4.002 8.49 4.55 ;
      RECT 8.48 4.02 8.485 4.561 ;
      RECT 8.475 4.03 8.48 4.572 ;
      RECT 8.47 4.038 8.475 4.584 ;
      RECT 8.465 4.046 8.47 4.595 ;
      RECT 8.46 4.072 8.465 4.608 ;
      RECT 8.45 4.1 8.46 4.621 ;
      RECT 8.445 4.13 8.45 4.63 ;
      RECT 8.44 4.145 8.445 4.637 ;
      RECT 8.425 4.17 8.44 4.644 ;
      RECT 8.42 4.192 8.425 4.65 ;
      RECT 8.415 4.217 8.42 4.653 ;
      RECT 8.406 4.245 8.415 4.657 ;
      RECT 8.4 4.262 8.406 4.662 ;
      RECT 8.395 4.28 8.4 4.666 ;
      RECT 8.39 4.292 8.395 4.669 ;
      RECT 8.385 4.313 8.39 4.673 ;
      RECT 8.38 4.331 8.385 4.676 ;
      RECT 8.375 4.345 8.38 4.679 ;
      RECT 8.37 4.362 8.375 4.682 ;
      RECT 8.365 4.375 8.37 4.685 ;
      RECT 8.34 4.412 8.365 4.693 ;
      RECT 8.335 4.457 8.34 4.702 ;
      RECT 8.33 4.485 8.335 4.705 ;
      RECT 8.32 4.505 8.33 4.709 ;
      RECT 8.315 4.525 8.32 4.714 ;
      RECT 8.31 4.54 8.315 4.717 ;
      RECT 8.29 4.55 8.31 4.724 ;
      RECT 8.225 4.557 8.29 4.75 ;
      RECT 8.19 4.56 8.225 4.778 ;
      RECT 8.175 4.563 8.19 4.793 ;
      RECT 8.165 4.564 8.175 4.808 ;
      RECT 8.155 4.565 8.165 4.825 ;
      RECT 8.15 4.565 8.155 4.84 ;
      RECT 8.145 4.565 8.15 4.848 ;
      RECT 8.13 4.566 8.145 4.863 ;
      RECT 8.1 4.568 8.13 4.87 ;
      RECT 7.99 4.575 8.07 4.87 ;
      RECT 7.945 4.58 7.99 4.87 ;
      RECT 7.935 4.581 7.945 4.86 ;
      RECT 7.925 4.582 7.935 4.853 ;
      RECT 7.905 4.584 7.925 4.848 ;
      RECT 7.895 4.555 7.905 4.843 ;
      RECT 7.85 4.555 7.895 4.835 ;
      RECT 7.82 4.555 7.845 4.825 ;
      RECT 7.8 4.555 7.82 4.818 ;
      RECT 8.08 3.355 8.34 3.615 ;
      RECT 7.96 3.37 7.97 3.535 ;
      RECT 7.945 3.37 7.95 3.53 ;
      RECT 5.31 3.21 5.495 3.5 ;
      RECT 7.125 3.335 7.14 3.49 ;
      RECT 5.275 3.21 5.3 3.47 ;
      RECT 7.69 3.26 7.695 3.402 ;
      RECT 7.605 3.255 7.63 3.395 ;
      RECT 8.005 3.372 8.08 3.565 ;
      RECT 7.99 3.37 8.005 3.548 ;
      RECT 7.97 3.37 7.99 3.54 ;
      RECT 7.95 3.37 7.96 3.533 ;
      RECT 7.905 3.365 7.945 3.523 ;
      RECT 7.865 3.34 7.905 3.508 ;
      RECT 7.85 3.315 7.865 3.498 ;
      RECT 7.845 3.309 7.85 3.496 ;
      RECT 7.81 3.301 7.845 3.479 ;
      RECT 7.805 3.294 7.81 3.467 ;
      RECT 7.785 3.289 7.805 3.455 ;
      RECT 7.775 3.283 7.785 3.44 ;
      RECT 7.755 3.278 7.775 3.425 ;
      RECT 7.745 3.273 7.755 3.418 ;
      RECT 7.74 3.271 7.745 3.413 ;
      RECT 7.735 3.27 7.74 3.41 ;
      RECT 7.695 3.265 7.735 3.406 ;
      RECT 7.675 3.259 7.69 3.401 ;
      RECT 7.64 3.256 7.675 3.398 ;
      RECT 7.63 3.255 7.64 3.396 ;
      RECT 7.57 3.255 7.605 3.393 ;
      RECT 7.525 3.255 7.57 3.393 ;
      RECT 7.475 3.255 7.525 3.396 ;
      RECT 7.46 3.257 7.475 3.398 ;
      RECT 7.445 3.26 7.46 3.399 ;
      RECT 7.435 3.265 7.445 3.4 ;
      RECT 7.405 3.27 7.435 3.405 ;
      RECT 7.395 3.276 7.405 3.413 ;
      RECT 7.385 3.278 7.395 3.417 ;
      RECT 7.375 3.282 7.385 3.421 ;
      RECT 7.35 3.288 7.375 3.429 ;
      RECT 7.34 3.293 7.35 3.437 ;
      RECT 7.325 3.297 7.34 3.441 ;
      RECT 7.29 3.303 7.325 3.449 ;
      RECT 7.27 3.308 7.29 3.459 ;
      RECT 7.24 3.315 7.27 3.468 ;
      RECT 7.195 3.324 7.24 3.482 ;
      RECT 7.19 3.329 7.195 3.493 ;
      RECT 7.17 3.332 7.19 3.494 ;
      RECT 7.14 3.335 7.17 3.492 ;
      RECT 7.105 3.335 7.125 3.488 ;
      RECT 7.035 3.335 7.105 3.479 ;
      RECT 7.02 3.332 7.035 3.471 ;
      RECT 6.98 3.325 7.02 3.466 ;
      RECT 6.955 3.315 6.98 3.459 ;
      RECT 6.95 3.309 6.955 3.456 ;
      RECT 6.91 3.303 6.95 3.453 ;
      RECT 6.895 3.296 6.91 3.448 ;
      RECT 6.875 3.292 6.895 3.443 ;
      RECT 6.86 3.287 6.875 3.439 ;
      RECT 6.845 3.282 6.86 3.437 ;
      RECT 6.83 3.278 6.845 3.436 ;
      RECT 6.815 3.276 6.83 3.432 ;
      RECT 6.805 3.274 6.815 3.427 ;
      RECT 6.79 3.271 6.805 3.423 ;
      RECT 6.78 3.269 6.79 3.418 ;
      RECT 6.76 3.266 6.78 3.414 ;
      RECT 6.715 3.265 6.76 3.412 ;
      RECT 6.655 3.267 6.715 3.413 ;
      RECT 6.635 3.269 6.655 3.415 ;
      RECT 6.605 3.272 6.635 3.416 ;
      RECT 6.555 3.277 6.605 3.418 ;
      RECT 6.55 3.28 6.555 3.42 ;
      RECT 6.54 3.282 6.55 3.423 ;
      RECT 6.535 3.284 6.54 3.426 ;
      RECT 6.485 3.287 6.535 3.433 ;
      RECT 6.465 3.291 6.485 3.445 ;
      RECT 6.455 3.294 6.465 3.451 ;
      RECT 6.445 3.295 6.455 3.454 ;
      RECT 6.406 3.298 6.445 3.456 ;
      RECT 6.32 3.305 6.406 3.459 ;
      RECT 6.246 3.315 6.32 3.463 ;
      RECT 6.16 3.326 6.246 3.468 ;
      RECT 6.145 3.333 6.16 3.47 ;
      RECT 6.09 3.337 6.145 3.471 ;
      RECT 6.076 3.34 6.09 3.473 ;
      RECT 5.99 3.34 6.076 3.475 ;
      RECT 5.95 3.337 5.99 3.478 ;
      RECT 5.926 3.333 5.95 3.48 ;
      RECT 5.84 3.323 5.926 3.483 ;
      RECT 5.81 3.312 5.84 3.484 ;
      RECT 5.791 3.308 5.81 3.483 ;
      RECT 5.705 3.301 5.791 3.48 ;
      RECT 5.645 3.29 5.705 3.477 ;
      RECT 5.625 3.282 5.645 3.475 ;
      RECT 5.59 3.277 5.625 3.474 ;
      RECT 5.565 3.272 5.59 3.473 ;
      RECT 5.535 3.267 5.565 3.472 ;
      RECT 5.51 3.21 5.535 3.471 ;
      RECT 5.495 3.21 5.51 3.495 ;
      RECT 5.3 3.21 5.31 3.495 ;
      RECT 7.075 4.23 7.08 4.37 ;
      RECT 6.735 4.23 6.77 4.368 ;
      RECT 6.31 4.215 6.325 4.36 ;
      RECT 8.14 3.995 8.23 4.255 ;
      RECT 7.97 3.86 8.07 4.255 ;
      RECT 5.005 3.835 5.085 4.045 ;
      RECT 8.095 3.972 8.14 4.255 ;
      RECT 8.085 3.942 8.095 4.255 ;
      RECT 8.07 3.865 8.085 4.255 ;
      RECT 7.885 3.86 7.97 4.22 ;
      RECT 7.88 3.862 7.885 4.215 ;
      RECT 7.875 3.867 7.88 4.215 ;
      RECT 7.84 3.967 7.875 4.215 ;
      RECT 7.83 3.995 7.84 4.215 ;
      RECT 7.82 4.01 7.83 4.215 ;
      RECT 7.81 4.022 7.82 4.215 ;
      RECT 7.805 4.032 7.81 4.215 ;
      RECT 7.79 4.042 7.805 4.217 ;
      RECT 7.785 4.057 7.79 4.219 ;
      RECT 7.77 4.07 7.785 4.221 ;
      RECT 7.765 4.085 7.77 4.224 ;
      RECT 7.745 4.095 7.765 4.228 ;
      RECT 7.73 4.105 7.745 4.231 ;
      RECT 7.695 4.112 7.73 4.236 ;
      RECT 7.651 4.119 7.695 4.244 ;
      RECT 7.565 4.131 7.651 4.257 ;
      RECT 7.54 4.142 7.565 4.268 ;
      RECT 7.51 4.147 7.54 4.273 ;
      RECT 7.475 4.152 7.51 4.281 ;
      RECT 7.445 4.157 7.475 4.288 ;
      RECT 7.42 4.162 7.445 4.293 ;
      RECT 7.355 4.169 7.42 4.302 ;
      RECT 7.285 4.182 7.355 4.318 ;
      RECT 7.255 4.192 7.285 4.33 ;
      RECT 7.23 4.197 7.255 4.337 ;
      RECT 7.175 4.204 7.23 4.345 ;
      RECT 7.17 4.211 7.175 4.35 ;
      RECT 7.165 4.213 7.17 4.351 ;
      RECT 7.15 4.215 7.165 4.353 ;
      RECT 7.145 4.215 7.15 4.356 ;
      RECT 7.08 4.222 7.145 4.363 ;
      RECT 7.045 4.232 7.075 4.373 ;
      RECT 7.028 4.235 7.045 4.375 ;
      RECT 6.942 4.234 7.028 4.374 ;
      RECT 6.856 4.232 6.942 4.371 ;
      RECT 6.77 4.231 6.856 4.369 ;
      RECT 6.669 4.229 6.735 4.368 ;
      RECT 6.583 4.226 6.669 4.366 ;
      RECT 6.497 4.222 6.583 4.364 ;
      RECT 6.411 4.219 6.497 4.363 ;
      RECT 6.325 4.216 6.411 4.361 ;
      RECT 6.225 4.215 6.31 4.358 ;
      RECT 6.175 4.213 6.225 4.356 ;
      RECT 6.155 4.21 6.175 4.354 ;
      RECT 6.135 4.208 6.155 4.351 ;
      RECT 6.11 4.204 6.135 4.348 ;
      RECT 6.065 4.198 6.11 4.343 ;
      RECT 6.025 4.192 6.065 4.335 ;
      RECT 6 4.187 6.025 4.328 ;
      RECT 5.945 4.18 6 4.32 ;
      RECT 5.921 4.173 5.945 4.313 ;
      RECT 5.835 4.164 5.921 4.303 ;
      RECT 5.805 4.156 5.835 4.293 ;
      RECT 5.775 4.152 5.805 4.288 ;
      RECT 5.77 4.149 5.775 4.285 ;
      RECT 5.765 4.148 5.77 4.285 ;
      RECT 5.69 4.141 5.765 4.278 ;
      RECT 5.651 4.132 5.69 4.267 ;
      RECT 5.565 4.122 5.651 4.255 ;
      RECT 5.525 4.112 5.565 4.243 ;
      RECT 5.486 4.107 5.525 4.236 ;
      RECT 5.4 4.097 5.486 4.225 ;
      RECT 5.36 4.085 5.4 4.214 ;
      RECT 5.325 4.07 5.36 4.207 ;
      RECT 5.315 4.06 5.325 4.204 ;
      RECT 5.295 4.045 5.315 4.202 ;
      RECT 5.265 4.015 5.295 4.198 ;
      RECT 5.255 3.995 5.265 4.193 ;
      RECT 5.25 3.987 5.255 4.19 ;
      RECT 5.245 3.98 5.25 4.188 ;
      RECT 5.23 3.967 5.245 4.181 ;
      RECT 5.225 3.957 5.23 4.173 ;
      RECT 5.22 3.95 5.225 4.168 ;
      RECT 5.215 3.945 5.22 4.164 ;
      RECT 5.2 3.932 5.215 4.156 ;
      RECT 5.195 3.842 5.2 4.145 ;
      RECT 5.19 3.837 5.195 4.138 ;
      RECT 5.115 3.835 5.19 4.098 ;
      RECT 5.085 3.835 5.115 4.053 ;
      RECT 4.99 3.84 5.005 4.04 ;
      RECT 7.475 3.545 7.735 3.805 ;
      RECT 7.46 3.533 7.64 3.77 ;
      RECT 7.455 3.534 7.64 3.768 ;
      RECT 7.44 3.538 7.65 3.758 ;
      RECT 7.435 3.543 7.655 3.728 ;
      RECT 7.44 3.54 7.655 3.758 ;
      RECT 7.455 3.535 7.65 3.768 ;
      RECT 7.475 3.532 7.64 3.805 ;
      RECT 7.475 3.531 7.63 3.805 ;
      RECT 7.5 3.53 7.63 3.805 ;
      RECT 7.06 3.775 7.32 4.035 ;
      RECT 6.935 3.82 7.32 4.03 ;
      RECT 6.925 3.825 7.32 4.025 ;
      RECT 6.94 4.765 6.955 5.075 ;
      RECT 5.535 4.535 5.545 4.665 ;
      RECT 5.315 4.53 5.42 4.665 ;
      RECT 5.23 4.535 5.28 4.665 ;
      RECT 3.78 3.27 3.785 4.375 ;
      RECT 7.035 4.857 7.04 4.993 ;
      RECT 7.03 4.852 7.035 5.053 ;
      RECT 7.025 4.85 7.03 5.066 ;
      RECT 7.01 4.847 7.025 5.068 ;
      RECT 7.005 4.842 7.01 5.07 ;
      RECT 7 4.838 7.005 5.073 ;
      RECT 6.985 4.833 7 5.075 ;
      RECT 6.955 4.825 6.985 5.075 ;
      RECT 6.916 4.765 6.94 5.075 ;
      RECT 6.83 4.765 6.916 5.072 ;
      RECT 6.8 4.765 6.83 5.065 ;
      RECT 6.775 4.765 6.8 5.058 ;
      RECT 6.75 4.765 6.775 5.05 ;
      RECT 6.735 4.765 6.75 5.043 ;
      RECT 6.71 4.765 6.735 5.035 ;
      RECT 6.695 4.765 6.71 5.028 ;
      RECT 6.655 4.775 6.695 5.017 ;
      RECT 6.645 4.77 6.655 5.007 ;
      RECT 6.641 4.769 6.645 5.004 ;
      RECT 6.555 4.761 6.641 4.987 ;
      RECT 6.522 4.75 6.555 4.964 ;
      RECT 6.436 4.739 6.522 4.942 ;
      RECT 6.35 4.723 6.436 4.911 ;
      RECT 6.28 4.708 6.35 4.883 ;
      RECT 6.27 4.701 6.28 4.87 ;
      RECT 6.24 4.698 6.27 4.86 ;
      RECT 6.215 4.694 6.24 4.853 ;
      RECT 6.2 4.691 6.215 4.848 ;
      RECT 6.195 4.69 6.2 4.843 ;
      RECT 6.165 4.685 6.195 4.836 ;
      RECT 6.16 4.68 6.165 4.831 ;
      RECT 6.145 4.677 6.16 4.826 ;
      RECT 6.14 4.672 6.145 4.821 ;
      RECT 6.12 4.667 6.14 4.818 ;
      RECT 6.105 4.662 6.12 4.81 ;
      RECT 6.09 4.656 6.105 4.805 ;
      RECT 6.06 4.647 6.09 4.798 ;
      RECT 6.055 4.64 6.06 4.79 ;
      RECT 6.05 4.638 6.055 4.788 ;
      RECT 6.045 4.637 6.05 4.785 ;
      RECT 6.005 4.63 6.045 4.778 ;
      RECT 5.991 4.62 6.005 4.768 ;
      RECT 5.94 4.609 5.991 4.756 ;
      RECT 5.915 4.595 5.94 4.742 ;
      RECT 5.89 4.584 5.915 4.734 ;
      RECT 5.87 4.573 5.89 4.728 ;
      RECT 5.86 4.567 5.87 4.723 ;
      RECT 5.855 4.565 5.86 4.719 ;
      RECT 5.835 4.56 5.855 4.714 ;
      RECT 5.805 4.55 5.835 4.704 ;
      RECT 5.8 4.542 5.805 4.697 ;
      RECT 5.785 4.54 5.8 4.693 ;
      RECT 5.765 4.54 5.785 4.688 ;
      RECT 5.76 4.539 5.765 4.686 ;
      RECT 5.755 4.539 5.76 4.683 ;
      RECT 5.715 4.538 5.755 4.678 ;
      RECT 5.69 4.537 5.715 4.673 ;
      RECT 5.63 4.536 5.69 4.67 ;
      RECT 5.545 4.535 5.63 4.668 ;
      RECT 5.506 4.534 5.535 4.665 ;
      RECT 5.42 4.532 5.506 4.665 ;
      RECT 5.28 4.532 5.315 4.665 ;
      RECT 5.19 4.536 5.23 4.668 ;
      RECT 5.175 4.539 5.19 4.675 ;
      RECT 5.165 4.54 5.175 4.682 ;
      RECT 5.14 4.543 5.165 4.687 ;
      RECT 5.135 4.545 5.14 4.69 ;
      RECT 5.085 4.547 5.135 4.691 ;
      RECT 5.046 4.551 5.085 4.693 ;
      RECT 4.96 4.553 5.046 4.696 ;
      RECT 4.942 4.555 4.96 4.698 ;
      RECT 4.856 4.558 4.942 4.7 ;
      RECT 4.77 4.562 4.856 4.703 ;
      RECT 4.733 4.566 4.77 4.706 ;
      RECT 4.647 4.569 4.733 4.709 ;
      RECT 4.561 4.573 4.647 4.712 ;
      RECT 4.475 4.578 4.561 4.716 ;
      RECT 4.455 4.58 4.475 4.719 ;
      RECT 4.435 4.579 4.455 4.72 ;
      RECT 4.386 4.576 4.435 4.721 ;
      RECT 4.3 4.571 4.386 4.724 ;
      RECT 4.25 4.566 4.3 4.726 ;
      RECT 4.226 4.564 4.25 4.727 ;
      RECT 4.14 4.559 4.226 4.729 ;
      RECT 4.115 4.555 4.14 4.728 ;
      RECT 4.105 4.552 4.115 4.726 ;
      RECT 4.095 4.545 4.105 4.723 ;
      RECT 4.09 4.525 4.095 4.718 ;
      RECT 4.08 4.495 4.09 4.713 ;
      RECT 4.065 4.365 4.08 4.704 ;
      RECT 4.06 4.357 4.065 4.697 ;
      RECT 4.04 4.35 4.06 4.689 ;
      RECT 4.035 4.332 4.04 4.681 ;
      RECT 4.025 4.312 4.035 4.676 ;
      RECT 4.02 4.285 4.025 4.672 ;
      RECT 4.015 4.262 4.02 4.669 ;
      RECT 3.995 4.22 4.015 4.661 ;
      RECT 3.96 4.135 3.995 4.645 ;
      RECT 3.955 4.067 3.96 4.633 ;
      RECT 3.94 4.037 3.955 4.627 ;
      RECT 3.935 3.282 3.94 3.528 ;
      RECT 3.925 4.007 3.94 4.618 ;
      RECT 3.93 3.277 3.935 3.56 ;
      RECT 3.925 3.272 3.93 3.603 ;
      RECT 3.92 3.27 3.925 3.638 ;
      RECT 3.905 3.97 3.925 4.608 ;
      RECT 3.915 3.27 3.92 3.675 ;
      RECT 3.9 3.27 3.915 3.773 ;
      RECT 3.9 3.943 3.905 4.601 ;
      RECT 3.895 3.27 3.9 3.848 ;
      RECT 3.895 3.931 3.9 4.598 ;
      RECT 3.89 3.27 3.895 3.88 ;
      RECT 3.89 3.91 3.895 4.595 ;
      RECT 3.885 3.27 3.89 4.592 ;
      RECT 3.85 3.27 3.885 4.578 ;
      RECT 3.835 3.27 3.85 4.56 ;
      RECT 3.815 3.27 3.835 4.55 ;
      RECT 3.79 3.27 3.815 4.533 ;
      RECT 3.785 3.27 3.79 4.483 ;
      RECT 3.775 3.27 3.78 4.313 ;
      RECT 3.77 3.27 3.775 4.22 ;
      RECT 3.765 3.27 3.77 4.133 ;
      RECT 3.76 3.27 3.765 4.065 ;
      RECT 3.755 3.27 3.76 4.008 ;
      RECT 3.745 3.27 3.755 3.903 ;
      RECT 3.74 3.27 3.745 3.775 ;
      RECT 3.735 3.27 3.74 3.693 ;
      RECT 3.73 3.272 3.735 3.61 ;
      RECT 3.725 3.277 3.73 3.543 ;
      RECT 3.72 3.282 3.725 3.47 ;
      RECT 6.535 3.6 6.795 3.86 ;
      RECT 6.555 3.567 6.765 3.86 ;
      RECT 6.555 3.565 6.755 3.86 ;
      RECT 6.565 3.552 6.755 3.86 ;
      RECT 6.565 3.55 6.68 3.86 ;
      RECT 6.04 3.675 6.215 3.955 ;
      RECT 6.035 3.675 6.215 3.953 ;
      RECT 6.035 3.675 6.23 3.95 ;
      RECT 6.025 3.675 6.23 3.948 ;
      RECT 5.97 3.675 6.23 3.935 ;
      RECT 5.97 3.75 6.235 3.913 ;
      RECT 5.515 3.687 5.535 3.93 ;
      RECT 5.515 3.687 5.575 3.929 ;
      RECT 5.51 3.689 5.575 3.928 ;
      RECT 5.51 3.689 5.661 3.927 ;
      RECT 5.51 3.689 5.73 3.926 ;
      RECT 5.51 3.689 5.75 3.918 ;
      RECT 5.49 3.692 5.75 3.916 ;
      RECT 5.475 3.702 5.75 3.901 ;
      RECT 5.475 3.702 5.765 3.9 ;
      RECT 5.47 3.711 5.765 3.892 ;
      RECT 5.47 3.711 5.77 3.888 ;
      RECT 5.575 3.625 5.835 3.885 ;
      RECT 5.465 3.713 5.835 3.77 ;
      RECT 5.535 3.68 5.835 3.885 ;
      RECT 5.5 4.873 5.505 5.08 ;
      RECT 5.45 4.867 5.5 5.079 ;
      RECT 5.417 4.881 5.51 5.078 ;
      RECT 5.331 4.881 5.51 5.077 ;
      RECT 5.245 4.881 5.51 5.076 ;
      RECT 5.245 4.98 5.515 5.073 ;
      RECT 5.24 4.98 5.515 5.068 ;
      RECT 5.235 4.98 5.515 5.05 ;
      RECT 5.23 4.98 5.515 5.033 ;
      RECT 5.19 4.765 5.45 5.025 ;
      RECT 4.65 3.915 4.736 4.329 ;
      RECT 4.65 3.915 4.775 4.326 ;
      RECT 4.65 3.915 4.795 4.316 ;
      RECT 4.605 3.915 4.795 4.313 ;
      RECT 4.605 4.067 4.805 4.303 ;
      RECT 4.605 4.088 4.81 4.297 ;
      RECT 4.605 4.106 4.815 4.293 ;
      RECT 4.605 4.126 4.825 4.288 ;
      RECT 4.58 4.126 4.825 4.285 ;
      RECT 4.57 4.126 4.825 4.263 ;
      RECT 4.57 4.142 4.83 4.233 ;
      RECT 4.535 3.915 4.795 4.22 ;
      RECT 4.535 4.154 4.835 4.175 ;
      RECT 1.975 8.945 2.265 9.175 ;
      RECT 1.805 8.975 2.265 9.145 ;
      RECT 1.545 10.055 1.835 10.285 ;
      RECT 1.605 9.315 1.775 10.285 ;
      RECT 1.515 9.315 1.865 9.605 ;
      RECT 1.14 8.575 1.49 8.865 ;
      RECT 1 8.605 1.49 8.775 ;
      RECT 68.16 4.56 68.42 4.82 ;
      RECT 52.9 4.56 53.16 4.82 ;
      RECT 37.64 4.56 37.9 4.82 ;
      RECT 22.38 4.56 22.64 4.82 ;
      RECT 7.12 4.56 7.38 4.82 ;
    LAYER mcon ;
      RECT 78.555 8.61 78.725 8.78 ;
      RECT 78.555 10.09 78.725 10.26 ;
      RECT 78.205 1.395 78.375 1.565 ;
      RECT 78.205 5.455 78.375 5.625 ;
      RECT 78.205 6.84 78.375 7.01 ;
      RECT 78.205 10.9 78.375 11.07 ;
      RECT 78.185 4.055 78.355 4.225 ;
      RECT 78.185 8.24 78.355 8.41 ;
      RECT 77.565 2.205 77.735 2.375 ;
      RECT 77.565 3.685 77.735 3.855 ;
      RECT 77.565 8.61 77.735 8.78 ;
      RECT 77.565 10.09 77.735 10.26 ;
      RECT 77.215 1.395 77.385 1.565 ;
      RECT 77.215 5.455 77.385 5.625 ;
      RECT 77.215 6.84 77.385 7.01 ;
      RECT 77.215 10.9 77.385 11.07 ;
      RECT 77.195 4.055 77.365 4.225 ;
      RECT 77.195 8.24 77.365 8.41 ;
      RECT 76.515 1.4 76.685 1.57 ;
      RECT 76.515 5.46 76.685 5.63 ;
      RECT 76.515 6.835 76.685 7.005 ;
      RECT 76.515 10.895 76.685 11.065 ;
      RECT 76.205 3.32 76.375 3.49 ;
      RECT 76.205 8.975 76.375 9.145 ;
      RECT 75.835 1.4 76.005 1.57 ;
      RECT 75.835 10.895 76.005 11.065 ;
      RECT 75.775 2.21 75.945 2.38 ;
      RECT 75.775 2.95 75.945 3.12 ;
      RECT 75.775 9.345 75.945 9.515 ;
      RECT 75.775 10.085 75.945 10.255 ;
      RECT 75.4 3.69 75.57 3.86 ;
      RECT 75.4 8.605 75.57 8.775 ;
      RECT 75.155 1.4 75.325 1.57 ;
      RECT 75.155 10.895 75.325 11.065 ;
      RECT 74.475 1.4 74.645 1.57 ;
      RECT 74.475 10.895 74.645 11.065 ;
      RECT 73.015 2.71 73.185 2.88 ;
      RECT 73.015 5.43 73.185 5.6 ;
      RECT 72.575 3.575 72.745 3.745 ;
      RECT 72.555 2.71 72.725 2.88 ;
      RECT 72.555 5.43 72.725 5.6 ;
      RECT 72.18 4.32 72.35 4.49 ;
      RECT 72.095 2.71 72.265 2.88 ;
      RECT 72.095 5.43 72.265 5.6 ;
      RECT 72.07 3.595 72.24 3.765 ;
      RECT 71.635 2.71 71.805 2.88 ;
      RECT 71.635 5.43 71.805 5.6 ;
      RECT 71.25 3.285 71.42 3.455 ;
      RECT 71.175 2.71 71.345 2.88 ;
      RECT 71.175 5.43 71.345 5.6 ;
      RECT 70.935 4.325 71.105 4.495 ;
      RECT 70.89 3.815 71.06 3.985 ;
      RECT 70.88 6.835 71.05 7.005 ;
      RECT 70.88 10.895 71.05 11.065 ;
      RECT 70.715 2.71 70.885 2.88 ;
      RECT 70.715 5.43 70.885 5.6 ;
      RECT 70.57 8.975 70.74 9.145 ;
      RECT 70.465 4.025 70.635 4.195 ;
      RECT 70.275 3.245 70.445 3.415 ;
      RECT 70.255 2.71 70.425 2.88 ;
      RECT 70.255 5.43 70.425 5.6 ;
      RECT 70.225 4.855 70.395 5.025 ;
      RECT 70.2 10.895 70.37 11.065 ;
      RECT 70.14 9.345 70.31 9.515 ;
      RECT 70.14 10.085 70.31 10.255 ;
      RECT 69.89 4.295 70.06 4.465 ;
      RECT 69.795 2.71 69.965 2.88 ;
      RECT 69.795 3.455 69.965 3.625 ;
      RECT 69.795 5.43 69.965 5.6 ;
      RECT 69.765 8.605 69.935 8.775 ;
      RECT 69.52 10.895 69.69 11.065 ;
      RECT 69.335 2.71 69.505 2.88 ;
      RECT 69.335 5.43 69.505 5.6 ;
      RECT 68.995 4.68 69.165 4.85 ;
      RECT 68.935 3.88 69.105 4.05 ;
      RECT 68.875 2.71 69.045 2.88 ;
      RECT 68.875 5.43 69.045 5.6 ;
      RECT 68.84 10.895 69.01 11.065 ;
      RECT 68.495 3.55 68.665 3.72 ;
      RECT 68.415 2.71 68.585 2.88 ;
      RECT 68.415 5.43 68.585 5.6 ;
      RECT 68.23 4.6 68.4 4.77 ;
      RECT 67.985 3.84 68.155 4.01 ;
      RECT 67.955 2.71 68.125 2.88 ;
      RECT 67.955 5.43 68.125 5.6 ;
      RECT 67.89 4.87 68.06 5.04 ;
      RECT 67.615 3.565 67.785 3.735 ;
      RECT 67.495 2.71 67.665 2.88 ;
      RECT 67.495 5.43 67.665 5.6 ;
      RECT 67.085 3.765 67.255 3.935 ;
      RECT 67.035 2.71 67.205 2.88 ;
      RECT 67.035 5.43 67.205 5.6 ;
      RECT 66.575 2.71 66.745 2.88 ;
      RECT 66.575 5.43 66.745 5.6 ;
      RECT 66.565 3.71 66.735 3.88 ;
      RECT 66.36 3.31 66.53 3.48 ;
      RECT 66.36 4.89 66.53 5.06 ;
      RECT 66.115 2.71 66.285 2.88 ;
      RECT 66.115 5.43 66.285 5.6 ;
      RECT 66.05 3.855 66.22 4.025 ;
      RECT 65.655 2.71 65.825 2.88 ;
      RECT 65.655 5.43 65.825 5.6 ;
      RECT 65.64 4.08 65.81 4.25 ;
      RECT 65.195 2.71 65.365 2.88 ;
      RECT 65.195 5.43 65.365 5.6 ;
      RECT 64.93 4.38 65.1 4.55 ;
      RECT 64.785 3.29 64.955 3.46 ;
      RECT 64.735 2.71 64.905 2.88 ;
      RECT 64.735 5.43 64.905 5.6 ;
      RECT 63.295 8.61 63.465 8.78 ;
      RECT 63.295 10.09 63.465 10.26 ;
      RECT 62.945 1.395 63.115 1.565 ;
      RECT 62.945 5.455 63.115 5.625 ;
      RECT 62.945 6.84 63.115 7.01 ;
      RECT 62.945 10.9 63.115 11.07 ;
      RECT 62.925 4.055 63.095 4.225 ;
      RECT 62.925 8.24 63.095 8.41 ;
      RECT 62.305 2.205 62.475 2.375 ;
      RECT 62.305 3.685 62.475 3.855 ;
      RECT 62.305 8.61 62.475 8.78 ;
      RECT 62.305 10.09 62.475 10.26 ;
      RECT 61.955 1.395 62.125 1.565 ;
      RECT 61.955 5.455 62.125 5.625 ;
      RECT 61.955 6.84 62.125 7.01 ;
      RECT 61.955 10.9 62.125 11.07 ;
      RECT 61.935 4.055 62.105 4.225 ;
      RECT 61.935 8.24 62.105 8.41 ;
      RECT 61.255 1.4 61.425 1.57 ;
      RECT 61.255 5.46 61.425 5.63 ;
      RECT 61.255 6.835 61.425 7.005 ;
      RECT 61.255 10.895 61.425 11.065 ;
      RECT 60.945 3.32 61.115 3.49 ;
      RECT 60.945 8.975 61.115 9.145 ;
      RECT 60.575 1.4 60.745 1.57 ;
      RECT 60.575 10.895 60.745 11.065 ;
      RECT 60.515 2.21 60.685 2.38 ;
      RECT 60.515 2.95 60.685 3.12 ;
      RECT 60.515 9.345 60.685 9.515 ;
      RECT 60.515 10.085 60.685 10.255 ;
      RECT 60.14 3.69 60.31 3.86 ;
      RECT 60.14 8.605 60.31 8.775 ;
      RECT 59.895 1.4 60.065 1.57 ;
      RECT 59.895 10.895 60.065 11.065 ;
      RECT 59.215 1.4 59.385 1.57 ;
      RECT 59.215 10.895 59.385 11.065 ;
      RECT 57.755 2.71 57.925 2.88 ;
      RECT 57.755 5.43 57.925 5.6 ;
      RECT 57.315 3.575 57.485 3.745 ;
      RECT 57.295 2.71 57.465 2.88 ;
      RECT 57.295 5.43 57.465 5.6 ;
      RECT 56.92 4.32 57.09 4.49 ;
      RECT 56.835 2.71 57.005 2.88 ;
      RECT 56.835 5.43 57.005 5.6 ;
      RECT 56.81 3.595 56.98 3.765 ;
      RECT 56.375 2.71 56.545 2.88 ;
      RECT 56.375 5.43 56.545 5.6 ;
      RECT 55.99 3.285 56.16 3.455 ;
      RECT 55.915 2.71 56.085 2.88 ;
      RECT 55.915 5.43 56.085 5.6 ;
      RECT 55.675 4.325 55.845 4.495 ;
      RECT 55.63 3.815 55.8 3.985 ;
      RECT 55.62 6.835 55.79 7.005 ;
      RECT 55.62 10.895 55.79 11.065 ;
      RECT 55.455 2.71 55.625 2.88 ;
      RECT 55.455 5.43 55.625 5.6 ;
      RECT 55.31 8.975 55.48 9.145 ;
      RECT 55.205 4.025 55.375 4.195 ;
      RECT 55.015 3.245 55.185 3.415 ;
      RECT 54.995 2.71 55.165 2.88 ;
      RECT 54.995 5.43 55.165 5.6 ;
      RECT 54.965 4.855 55.135 5.025 ;
      RECT 54.94 10.895 55.11 11.065 ;
      RECT 54.88 9.345 55.05 9.515 ;
      RECT 54.88 10.085 55.05 10.255 ;
      RECT 54.63 4.295 54.8 4.465 ;
      RECT 54.535 2.71 54.705 2.88 ;
      RECT 54.535 3.455 54.705 3.625 ;
      RECT 54.535 5.43 54.705 5.6 ;
      RECT 54.505 8.605 54.675 8.775 ;
      RECT 54.26 10.895 54.43 11.065 ;
      RECT 54.075 2.71 54.245 2.88 ;
      RECT 54.075 5.43 54.245 5.6 ;
      RECT 53.735 4.68 53.905 4.85 ;
      RECT 53.675 3.88 53.845 4.05 ;
      RECT 53.615 2.71 53.785 2.88 ;
      RECT 53.615 5.43 53.785 5.6 ;
      RECT 53.58 10.895 53.75 11.065 ;
      RECT 53.235 3.55 53.405 3.72 ;
      RECT 53.155 2.71 53.325 2.88 ;
      RECT 53.155 5.43 53.325 5.6 ;
      RECT 52.97 4.6 53.14 4.77 ;
      RECT 52.725 3.84 52.895 4.01 ;
      RECT 52.695 2.71 52.865 2.88 ;
      RECT 52.695 5.43 52.865 5.6 ;
      RECT 52.63 4.87 52.8 5.04 ;
      RECT 52.355 3.565 52.525 3.735 ;
      RECT 52.235 2.71 52.405 2.88 ;
      RECT 52.235 5.43 52.405 5.6 ;
      RECT 51.825 3.765 51.995 3.935 ;
      RECT 51.775 2.71 51.945 2.88 ;
      RECT 51.775 5.43 51.945 5.6 ;
      RECT 51.315 2.71 51.485 2.88 ;
      RECT 51.315 5.43 51.485 5.6 ;
      RECT 51.305 3.71 51.475 3.88 ;
      RECT 51.1 3.31 51.27 3.48 ;
      RECT 51.1 4.89 51.27 5.06 ;
      RECT 50.855 2.71 51.025 2.88 ;
      RECT 50.855 5.43 51.025 5.6 ;
      RECT 50.79 3.855 50.96 4.025 ;
      RECT 50.395 2.71 50.565 2.88 ;
      RECT 50.395 5.43 50.565 5.6 ;
      RECT 50.38 4.08 50.55 4.25 ;
      RECT 49.935 2.71 50.105 2.88 ;
      RECT 49.935 5.43 50.105 5.6 ;
      RECT 49.67 4.38 49.84 4.55 ;
      RECT 49.525 3.29 49.695 3.46 ;
      RECT 49.475 2.71 49.645 2.88 ;
      RECT 49.475 5.43 49.645 5.6 ;
      RECT 48.035 8.61 48.205 8.78 ;
      RECT 48.035 10.09 48.205 10.26 ;
      RECT 47.685 1.395 47.855 1.565 ;
      RECT 47.685 5.455 47.855 5.625 ;
      RECT 47.685 6.84 47.855 7.01 ;
      RECT 47.685 10.9 47.855 11.07 ;
      RECT 47.665 4.055 47.835 4.225 ;
      RECT 47.665 8.24 47.835 8.41 ;
      RECT 47.045 2.205 47.215 2.375 ;
      RECT 47.045 3.685 47.215 3.855 ;
      RECT 47.045 8.61 47.215 8.78 ;
      RECT 47.045 10.09 47.215 10.26 ;
      RECT 46.695 1.395 46.865 1.565 ;
      RECT 46.695 5.455 46.865 5.625 ;
      RECT 46.695 6.84 46.865 7.01 ;
      RECT 46.695 10.9 46.865 11.07 ;
      RECT 46.675 4.055 46.845 4.225 ;
      RECT 46.675 8.24 46.845 8.41 ;
      RECT 45.995 1.4 46.165 1.57 ;
      RECT 45.995 5.46 46.165 5.63 ;
      RECT 45.995 6.835 46.165 7.005 ;
      RECT 45.995 10.895 46.165 11.065 ;
      RECT 45.685 3.32 45.855 3.49 ;
      RECT 45.685 8.975 45.855 9.145 ;
      RECT 45.315 1.4 45.485 1.57 ;
      RECT 45.315 10.895 45.485 11.065 ;
      RECT 45.255 2.21 45.425 2.38 ;
      RECT 45.255 2.95 45.425 3.12 ;
      RECT 45.255 9.345 45.425 9.515 ;
      RECT 45.255 10.085 45.425 10.255 ;
      RECT 44.88 3.69 45.05 3.86 ;
      RECT 44.88 8.605 45.05 8.775 ;
      RECT 44.635 1.4 44.805 1.57 ;
      RECT 44.635 10.895 44.805 11.065 ;
      RECT 43.955 1.4 44.125 1.57 ;
      RECT 43.955 10.895 44.125 11.065 ;
      RECT 42.495 2.71 42.665 2.88 ;
      RECT 42.495 5.43 42.665 5.6 ;
      RECT 42.055 3.575 42.225 3.745 ;
      RECT 42.035 2.71 42.205 2.88 ;
      RECT 42.035 5.43 42.205 5.6 ;
      RECT 41.66 4.32 41.83 4.49 ;
      RECT 41.575 2.71 41.745 2.88 ;
      RECT 41.575 5.43 41.745 5.6 ;
      RECT 41.55 3.595 41.72 3.765 ;
      RECT 41.115 2.71 41.285 2.88 ;
      RECT 41.115 5.43 41.285 5.6 ;
      RECT 40.73 3.285 40.9 3.455 ;
      RECT 40.655 2.71 40.825 2.88 ;
      RECT 40.655 5.43 40.825 5.6 ;
      RECT 40.415 4.325 40.585 4.495 ;
      RECT 40.37 3.815 40.54 3.985 ;
      RECT 40.36 6.835 40.53 7.005 ;
      RECT 40.36 10.895 40.53 11.065 ;
      RECT 40.195 2.71 40.365 2.88 ;
      RECT 40.195 5.43 40.365 5.6 ;
      RECT 40.05 8.975 40.22 9.145 ;
      RECT 39.945 4.025 40.115 4.195 ;
      RECT 39.755 3.245 39.925 3.415 ;
      RECT 39.735 2.71 39.905 2.88 ;
      RECT 39.735 5.43 39.905 5.6 ;
      RECT 39.705 4.855 39.875 5.025 ;
      RECT 39.68 10.895 39.85 11.065 ;
      RECT 39.62 9.345 39.79 9.515 ;
      RECT 39.62 10.085 39.79 10.255 ;
      RECT 39.37 4.295 39.54 4.465 ;
      RECT 39.275 2.71 39.445 2.88 ;
      RECT 39.275 3.455 39.445 3.625 ;
      RECT 39.275 5.43 39.445 5.6 ;
      RECT 39.245 8.605 39.415 8.775 ;
      RECT 39 10.895 39.17 11.065 ;
      RECT 38.815 2.71 38.985 2.88 ;
      RECT 38.815 5.43 38.985 5.6 ;
      RECT 38.475 4.68 38.645 4.85 ;
      RECT 38.415 3.88 38.585 4.05 ;
      RECT 38.355 2.71 38.525 2.88 ;
      RECT 38.355 5.43 38.525 5.6 ;
      RECT 38.32 10.895 38.49 11.065 ;
      RECT 37.975 3.55 38.145 3.72 ;
      RECT 37.895 2.71 38.065 2.88 ;
      RECT 37.895 5.43 38.065 5.6 ;
      RECT 37.71 4.6 37.88 4.77 ;
      RECT 37.465 3.84 37.635 4.01 ;
      RECT 37.435 2.71 37.605 2.88 ;
      RECT 37.435 5.43 37.605 5.6 ;
      RECT 37.37 4.87 37.54 5.04 ;
      RECT 37.095 3.565 37.265 3.735 ;
      RECT 36.975 2.71 37.145 2.88 ;
      RECT 36.975 5.43 37.145 5.6 ;
      RECT 36.565 3.765 36.735 3.935 ;
      RECT 36.515 2.71 36.685 2.88 ;
      RECT 36.515 5.43 36.685 5.6 ;
      RECT 36.055 2.71 36.225 2.88 ;
      RECT 36.055 5.43 36.225 5.6 ;
      RECT 36.045 3.71 36.215 3.88 ;
      RECT 35.84 3.31 36.01 3.48 ;
      RECT 35.84 4.89 36.01 5.06 ;
      RECT 35.595 2.71 35.765 2.88 ;
      RECT 35.595 5.43 35.765 5.6 ;
      RECT 35.53 3.855 35.7 4.025 ;
      RECT 35.135 2.71 35.305 2.88 ;
      RECT 35.135 5.43 35.305 5.6 ;
      RECT 35.12 4.08 35.29 4.25 ;
      RECT 34.675 2.71 34.845 2.88 ;
      RECT 34.675 5.43 34.845 5.6 ;
      RECT 34.41 4.38 34.58 4.55 ;
      RECT 34.265 3.29 34.435 3.46 ;
      RECT 34.215 2.71 34.385 2.88 ;
      RECT 34.215 5.43 34.385 5.6 ;
      RECT 32.775 8.61 32.945 8.78 ;
      RECT 32.775 10.09 32.945 10.26 ;
      RECT 32.425 1.395 32.595 1.565 ;
      RECT 32.425 5.455 32.595 5.625 ;
      RECT 32.425 6.84 32.595 7.01 ;
      RECT 32.425 10.9 32.595 11.07 ;
      RECT 32.405 4.055 32.575 4.225 ;
      RECT 32.405 8.24 32.575 8.41 ;
      RECT 31.785 2.205 31.955 2.375 ;
      RECT 31.785 3.685 31.955 3.855 ;
      RECT 31.785 8.61 31.955 8.78 ;
      RECT 31.785 10.09 31.955 10.26 ;
      RECT 31.435 1.395 31.605 1.565 ;
      RECT 31.435 5.455 31.605 5.625 ;
      RECT 31.435 6.84 31.605 7.01 ;
      RECT 31.435 10.9 31.605 11.07 ;
      RECT 31.415 4.055 31.585 4.225 ;
      RECT 31.415 8.24 31.585 8.41 ;
      RECT 30.735 1.4 30.905 1.57 ;
      RECT 30.735 5.46 30.905 5.63 ;
      RECT 30.735 6.835 30.905 7.005 ;
      RECT 30.735 10.895 30.905 11.065 ;
      RECT 30.425 3.32 30.595 3.49 ;
      RECT 30.425 8.975 30.595 9.145 ;
      RECT 30.055 1.4 30.225 1.57 ;
      RECT 30.055 10.895 30.225 11.065 ;
      RECT 29.995 2.21 30.165 2.38 ;
      RECT 29.995 2.95 30.165 3.12 ;
      RECT 29.995 9.345 30.165 9.515 ;
      RECT 29.995 10.085 30.165 10.255 ;
      RECT 29.62 3.69 29.79 3.86 ;
      RECT 29.62 8.605 29.79 8.775 ;
      RECT 29.375 1.4 29.545 1.57 ;
      RECT 29.375 10.895 29.545 11.065 ;
      RECT 28.695 1.4 28.865 1.57 ;
      RECT 28.695 10.895 28.865 11.065 ;
      RECT 27.235 2.71 27.405 2.88 ;
      RECT 27.235 5.43 27.405 5.6 ;
      RECT 26.795 3.575 26.965 3.745 ;
      RECT 26.775 2.71 26.945 2.88 ;
      RECT 26.775 5.43 26.945 5.6 ;
      RECT 26.4 4.32 26.57 4.49 ;
      RECT 26.315 2.71 26.485 2.88 ;
      RECT 26.315 5.43 26.485 5.6 ;
      RECT 26.29 3.595 26.46 3.765 ;
      RECT 25.855 2.71 26.025 2.88 ;
      RECT 25.855 5.43 26.025 5.6 ;
      RECT 25.47 3.285 25.64 3.455 ;
      RECT 25.395 2.71 25.565 2.88 ;
      RECT 25.395 5.43 25.565 5.6 ;
      RECT 25.155 4.325 25.325 4.495 ;
      RECT 25.11 3.815 25.28 3.985 ;
      RECT 25.1 6.835 25.27 7.005 ;
      RECT 25.1 10.895 25.27 11.065 ;
      RECT 24.935 2.71 25.105 2.88 ;
      RECT 24.935 5.43 25.105 5.6 ;
      RECT 24.79 8.975 24.96 9.145 ;
      RECT 24.685 4.025 24.855 4.195 ;
      RECT 24.495 3.245 24.665 3.415 ;
      RECT 24.475 2.71 24.645 2.88 ;
      RECT 24.475 5.43 24.645 5.6 ;
      RECT 24.445 4.855 24.615 5.025 ;
      RECT 24.42 10.895 24.59 11.065 ;
      RECT 24.36 9.345 24.53 9.515 ;
      RECT 24.36 10.085 24.53 10.255 ;
      RECT 24.11 4.295 24.28 4.465 ;
      RECT 24.015 2.71 24.185 2.88 ;
      RECT 24.015 3.455 24.185 3.625 ;
      RECT 24.015 5.43 24.185 5.6 ;
      RECT 23.985 8.605 24.155 8.775 ;
      RECT 23.74 10.895 23.91 11.065 ;
      RECT 23.555 2.71 23.725 2.88 ;
      RECT 23.555 5.43 23.725 5.6 ;
      RECT 23.215 4.68 23.385 4.85 ;
      RECT 23.155 3.88 23.325 4.05 ;
      RECT 23.095 2.71 23.265 2.88 ;
      RECT 23.095 5.43 23.265 5.6 ;
      RECT 23.06 10.895 23.23 11.065 ;
      RECT 22.715 3.55 22.885 3.72 ;
      RECT 22.635 2.71 22.805 2.88 ;
      RECT 22.635 5.43 22.805 5.6 ;
      RECT 22.45 4.6 22.62 4.77 ;
      RECT 22.205 3.84 22.375 4.01 ;
      RECT 22.175 2.71 22.345 2.88 ;
      RECT 22.175 5.43 22.345 5.6 ;
      RECT 22.11 4.87 22.28 5.04 ;
      RECT 21.835 3.565 22.005 3.735 ;
      RECT 21.715 2.71 21.885 2.88 ;
      RECT 21.715 5.43 21.885 5.6 ;
      RECT 21.305 3.765 21.475 3.935 ;
      RECT 21.255 2.71 21.425 2.88 ;
      RECT 21.255 5.43 21.425 5.6 ;
      RECT 20.795 2.71 20.965 2.88 ;
      RECT 20.795 5.43 20.965 5.6 ;
      RECT 20.785 3.71 20.955 3.88 ;
      RECT 20.58 3.31 20.75 3.48 ;
      RECT 20.58 4.89 20.75 5.06 ;
      RECT 20.335 2.71 20.505 2.88 ;
      RECT 20.335 5.43 20.505 5.6 ;
      RECT 20.27 3.855 20.44 4.025 ;
      RECT 19.875 2.71 20.045 2.88 ;
      RECT 19.875 5.43 20.045 5.6 ;
      RECT 19.86 4.08 20.03 4.25 ;
      RECT 19.415 2.71 19.585 2.88 ;
      RECT 19.415 5.43 19.585 5.6 ;
      RECT 19.15 4.38 19.32 4.55 ;
      RECT 19.005 3.29 19.175 3.46 ;
      RECT 18.955 2.71 19.125 2.88 ;
      RECT 18.955 5.43 19.125 5.6 ;
      RECT 17.515 8.61 17.685 8.78 ;
      RECT 17.515 10.09 17.685 10.26 ;
      RECT 17.165 1.395 17.335 1.565 ;
      RECT 17.165 5.455 17.335 5.625 ;
      RECT 17.165 6.84 17.335 7.01 ;
      RECT 17.165 10.9 17.335 11.07 ;
      RECT 17.145 4.055 17.315 4.225 ;
      RECT 17.145 8.24 17.315 8.41 ;
      RECT 16.525 2.205 16.695 2.375 ;
      RECT 16.525 3.685 16.695 3.855 ;
      RECT 16.525 8.61 16.695 8.78 ;
      RECT 16.525 10.09 16.695 10.26 ;
      RECT 16.175 1.395 16.345 1.565 ;
      RECT 16.175 5.455 16.345 5.625 ;
      RECT 16.175 6.84 16.345 7.01 ;
      RECT 16.175 10.9 16.345 11.07 ;
      RECT 16.155 4.055 16.325 4.225 ;
      RECT 16.155 8.24 16.325 8.41 ;
      RECT 15.475 1.4 15.645 1.57 ;
      RECT 15.475 5.46 15.645 5.63 ;
      RECT 15.475 6.835 15.645 7.005 ;
      RECT 15.475 10.895 15.645 11.065 ;
      RECT 15.165 3.32 15.335 3.49 ;
      RECT 15.165 8.975 15.335 9.145 ;
      RECT 14.795 1.4 14.965 1.57 ;
      RECT 14.795 10.895 14.965 11.065 ;
      RECT 14.735 2.21 14.905 2.38 ;
      RECT 14.735 2.95 14.905 3.12 ;
      RECT 14.735 9.345 14.905 9.515 ;
      RECT 14.735 10.085 14.905 10.255 ;
      RECT 14.36 3.69 14.53 3.86 ;
      RECT 14.36 8.605 14.53 8.775 ;
      RECT 14.115 1.4 14.285 1.57 ;
      RECT 14.115 10.895 14.285 11.065 ;
      RECT 13.435 1.4 13.605 1.57 ;
      RECT 13.435 10.895 13.605 11.065 ;
      RECT 11.975 2.71 12.145 2.88 ;
      RECT 11.975 5.43 12.145 5.6 ;
      RECT 11.535 3.575 11.705 3.745 ;
      RECT 11.515 2.71 11.685 2.88 ;
      RECT 11.515 5.43 11.685 5.6 ;
      RECT 11.14 4.32 11.31 4.49 ;
      RECT 11.055 2.71 11.225 2.88 ;
      RECT 11.055 5.43 11.225 5.6 ;
      RECT 11.03 3.595 11.2 3.765 ;
      RECT 10.595 2.71 10.765 2.88 ;
      RECT 10.595 5.43 10.765 5.6 ;
      RECT 10.21 3.285 10.38 3.455 ;
      RECT 10.135 2.71 10.305 2.88 ;
      RECT 10.135 5.43 10.305 5.6 ;
      RECT 9.895 4.325 10.065 4.495 ;
      RECT 9.85 3.815 10.02 3.985 ;
      RECT 9.84 6.835 10.01 7.005 ;
      RECT 9.84 10.895 10.01 11.065 ;
      RECT 9.675 2.71 9.845 2.88 ;
      RECT 9.675 5.43 9.845 5.6 ;
      RECT 9.53 8.975 9.7 9.145 ;
      RECT 9.425 4.025 9.595 4.195 ;
      RECT 9.235 3.245 9.405 3.415 ;
      RECT 9.215 2.71 9.385 2.88 ;
      RECT 9.215 5.43 9.385 5.6 ;
      RECT 9.185 4.855 9.355 5.025 ;
      RECT 9.16 10.895 9.33 11.065 ;
      RECT 9.1 9.345 9.27 9.515 ;
      RECT 9.1 10.085 9.27 10.255 ;
      RECT 8.85 4.295 9.02 4.465 ;
      RECT 8.755 2.71 8.925 2.88 ;
      RECT 8.755 3.455 8.925 3.625 ;
      RECT 8.755 5.43 8.925 5.6 ;
      RECT 8.725 8.605 8.895 8.775 ;
      RECT 8.48 10.895 8.65 11.065 ;
      RECT 8.295 2.71 8.465 2.88 ;
      RECT 8.295 5.43 8.465 5.6 ;
      RECT 7.955 4.68 8.125 4.85 ;
      RECT 7.895 3.88 8.065 4.05 ;
      RECT 7.835 2.71 8.005 2.88 ;
      RECT 7.835 5.43 8.005 5.6 ;
      RECT 7.8 10.895 7.97 11.065 ;
      RECT 7.455 3.55 7.625 3.72 ;
      RECT 7.375 2.71 7.545 2.88 ;
      RECT 7.375 5.43 7.545 5.6 ;
      RECT 7.19 4.6 7.36 4.77 ;
      RECT 6.945 3.84 7.115 4.01 ;
      RECT 6.915 2.71 7.085 2.88 ;
      RECT 6.915 5.43 7.085 5.6 ;
      RECT 6.85 4.87 7.02 5.04 ;
      RECT 6.575 3.565 6.745 3.735 ;
      RECT 6.455 2.71 6.625 2.88 ;
      RECT 6.455 5.43 6.625 5.6 ;
      RECT 6.045 3.765 6.215 3.935 ;
      RECT 5.995 2.71 6.165 2.88 ;
      RECT 5.995 5.43 6.165 5.6 ;
      RECT 5.535 2.71 5.705 2.88 ;
      RECT 5.535 5.43 5.705 5.6 ;
      RECT 5.525 3.71 5.695 3.88 ;
      RECT 5.32 3.31 5.49 3.48 ;
      RECT 5.32 4.89 5.49 5.06 ;
      RECT 5.075 2.71 5.245 2.88 ;
      RECT 5.075 5.43 5.245 5.6 ;
      RECT 5.01 3.855 5.18 4.025 ;
      RECT 4.615 2.71 4.785 2.88 ;
      RECT 4.615 5.43 4.785 5.6 ;
      RECT 4.6 4.08 4.77 4.25 ;
      RECT 4.155 2.71 4.325 2.88 ;
      RECT 4.155 5.43 4.325 5.6 ;
      RECT 3.89 4.38 4.06 4.55 ;
      RECT 3.745 3.29 3.915 3.46 ;
      RECT 3.695 2.71 3.865 2.88 ;
      RECT 3.695 5.43 3.865 5.6 ;
      RECT 2.345 6.835 2.515 7.005 ;
      RECT 2.345 10.895 2.515 11.065 ;
      RECT 2.035 8.975 2.205 9.145 ;
      RECT 1.665 10.895 1.835 11.065 ;
      RECT 1.605 9.345 1.775 9.515 ;
      RECT 1.605 10.085 1.775 10.255 ;
      RECT 1.23 8.605 1.4 8.775 ;
      RECT 0.985 10.895 1.155 11.065 ;
      RECT 0.305 10.895 0.475 11.065 ;
    LAYER li1 ;
      RECT 72.56 0 72.73 3.38 ;
      RECT 71.62 0 71.79 3.38 ;
      RECT 70.66 0 70.83 3.38 ;
      RECT 68.74 0 68.91 3.38 ;
      RECT 67.78 0 67.95 3.38 ;
      RECT 65.86 0 66.03 3.38 ;
      RECT 57.3 0 57.47 3.38 ;
      RECT 56.36 0 56.53 3.38 ;
      RECT 55.4 0 55.57 3.38 ;
      RECT 53.48 0 53.65 3.38 ;
      RECT 52.52 0 52.69 3.38 ;
      RECT 50.6 0 50.77 3.38 ;
      RECT 42.04 0 42.21 3.38 ;
      RECT 41.1 0 41.27 3.38 ;
      RECT 40.14 0 40.31 3.38 ;
      RECT 38.22 0 38.39 3.38 ;
      RECT 37.26 0 37.43 3.38 ;
      RECT 35.34 0 35.51 3.38 ;
      RECT 26.78 0 26.95 3.38 ;
      RECT 25.84 0 26.01 3.38 ;
      RECT 24.88 0 25.05 3.38 ;
      RECT 22.96 0 23.13 3.38 ;
      RECT 22 0 22.17 3.38 ;
      RECT 20.08 0 20.25 3.38 ;
      RECT 11.52 0 11.69 3.38 ;
      RECT 10.58 0 10.75 3.38 ;
      RECT 9.62 0 9.79 3.38 ;
      RECT 7.7 0 7.87 3.38 ;
      RECT 6.74 0 6.91 3.38 ;
      RECT 4.82 0 4.99 3.38 ;
      RECT 69.615 0 69.81 2.89 ;
      RECT 65.86 0 66.135 2.89 ;
      RECT 54.355 0 54.55 2.89 ;
      RECT 50.6 0 50.875 2.89 ;
      RECT 39.095 0 39.29 2.89 ;
      RECT 35.34 0 35.615 2.89 ;
      RECT 23.835 0 24.03 2.89 ;
      RECT 20.08 0 20.355 2.89 ;
      RECT 8.575 0 8.77 2.89 ;
      RECT 4.82 0 5.095 2.89 ;
      RECT 64.59 0 73.33 2.88 ;
      RECT 49.33 0 58.07 2.88 ;
      RECT 34.07 0 42.81 2.88 ;
      RECT 18.81 0 27.55 2.88 ;
      RECT 3.55 0 12.29 2.88 ;
      RECT 74.395 0 74.565 2.23 ;
      RECT 59.135 0 59.305 2.23 ;
      RECT 43.875 0 44.045 2.23 ;
      RECT 28.615 0 28.785 2.23 ;
      RECT 13.355 0 13.525 2.23 ;
      RECT 78.125 0 78.295 2.225 ;
      RECT 77.135 0 77.305 2.225 ;
      RECT 62.865 0 63.035 2.225 ;
      RECT 61.875 0 62.045 2.225 ;
      RECT 47.605 0 47.775 2.225 ;
      RECT 46.615 0 46.785 2.225 ;
      RECT 32.345 0 32.515 2.225 ;
      RECT 31.355 0 31.525 2.225 ;
      RECT 17.085 0 17.255 2.225 ;
      RECT 16.095 0 16.265 2.225 ;
      RECT 0.005 0 79.1 1.6 ;
      RECT 2.035 5.435 2.205 10.595 ;
      RECT 78.125 4.695 78.295 7.77 ;
      RECT 77.135 4.695 77.305 7.77 ;
      RECT 62.865 4.695 63.035 7.77 ;
      RECT 61.875 4.695 62.045 7.77 ;
      RECT 47.605 4.695 47.775 7.77 ;
      RECT 46.615 4.695 46.785 7.77 ;
      RECT 32.345 4.695 32.515 7.77 ;
      RECT 31.355 4.695 31.525 7.77 ;
      RECT 17.085 4.695 17.255 7.77 ;
      RECT 16.095 4.695 16.265 7.77 ;
      RECT 74.395 4.7 74.565 7.765 ;
      RECT 68.76 4.93 68.93 7.765 ;
      RECT 59.135 4.7 59.305 7.765 ;
      RECT 53.5 4.93 53.67 7.765 ;
      RECT 43.875 4.7 44.045 7.765 ;
      RECT 38.24 4.93 38.41 7.765 ;
      RECT 28.615 4.7 28.785 7.765 ;
      RECT 22.98 4.93 23.15 7.765 ;
      RECT 13.355 4.7 13.525 7.765 ;
      RECT 7.72 4.93 7.89 7.765 ;
      RECT 0.225 5.435 0.395 7.765 ;
      RECT 76.965 5.425 78.945 7.04 ;
      RECT 61.705 5.425 63.685 7.04 ;
      RECT 46.445 5.425 48.425 7.04 ;
      RECT 31.185 5.425 33.165 7.04 ;
      RECT 15.925 5.425 17.905 7.04 ;
      RECT 0 5.435 79.1 7.035 ;
      RECT 64.59 5.43 79.1 7.035 ;
      RECT 49.33 5.43 63.84 7.035 ;
      RECT 34.07 5.43 48.58 7.035 ;
      RECT 18.81 5.43 33.32 7.035 ;
      RECT 3.55 5.43 18.06 7.035 ;
      RECT 71.62 4.93 71.79 7.035 ;
      RECT 69.7 4.93 69.87 7.035 ;
      RECT 67.3 4.93 67.47 7.035 ;
      RECT 65.38 4.93 65.55 7.035 ;
      RECT 56.36 4.93 56.53 7.035 ;
      RECT 54.44 4.93 54.61 7.035 ;
      RECT 52.04 4.93 52.21 7.035 ;
      RECT 50.12 4.93 50.29 7.035 ;
      RECT 41.1 4.93 41.27 7.035 ;
      RECT 39.18 4.93 39.35 7.035 ;
      RECT 36.78 4.93 36.95 7.035 ;
      RECT 34.86 4.93 35.03 7.035 ;
      RECT 25.84 4.93 26.01 7.035 ;
      RECT 23.92 4.93 24.09 7.035 ;
      RECT 21.52 4.93 21.69 7.035 ;
      RECT 19.6 4.93 19.77 7.035 ;
      RECT 10.58 4.93 10.75 7.035 ;
      RECT 8.66 4.93 8.83 7.035 ;
      RECT 6.26 4.93 6.43 7.035 ;
      RECT 4.34 4.93 4.51 7.035 ;
      RECT 0.005 10.865 79.1 12.465 ;
      RECT 78.125 10.24 78.295 12.465 ;
      RECT 77.135 10.24 77.305 12.465 ;
      RECT 74.395 10.235 74.565 12.465 ;
      RECT 68.76 10.235 68.93 12.465 ;
      RECT 62.865 10.24 63.035 12.465 ;
      RECT 61.875 10.24 62.045 12.465 ;
      RECT 59.135 10.235 59.305 12.465 ;
      RECT 53.5 10.235 53.67 12.465 ;
      RECT 47.605 10.24 47.775 12.465 ;
      RECT 46.615 10.24 46.785 12.465 ;
      RECT 43.875 10.235 44.045 12.465 ;
      RECT 38.24 10.235 38.41 12.465 ;
      RECT 32.345 10.24 32.515 12.465 ;
      RECT 31.355 10.24 31.525 12.465 ;
      RECT 28.615 10.235 28.785 12.465 ;
      RECT 22.98 10.235 23.15 12.465 ;
      RECT 17.085 10.24 17.255 12.465 ;
      RECT 16.095 10.24 16.265 12.465 ;
      RECT 13.355 10.235 13.525 12.465 ;
      RECT 7.72 10.235 7.89 12.465 ;
      RECT 0.225 10.235 0.395 12.465 ;
      RECT 78.185 3.035 78.355 4.225 ;
      RECT 78.185 3.035 78.655 3.205 ;
      RECT 78.185 9.26 78.655 9.43 ;
      RECT 78.185 8.24 78.355 9.43 ;
      RECT 77.195 3.035 77.365 4.225 ;
      RECT 77.195 3.035 77.665 3.205 ;
      RECT 77.195 9.26 77.665 9.43 ;
      RECT 77.195 8.24 77.365 9.43 ;
      RECT 75.345 3.93 75.515 5.16 ;
      RECT 75.4 2.15 75.57 4.1 ;
      RECT 75.345 1.87 75.515 2.32 ;
      RECT 75.345 10.145 75.515 10.595 ;
      RECT 75.4 8.365 75.57 10.315 ;
      RECT 75.345 7.305 75.515 8.535 ;
      RECT 74.825 1.87 74.995 5.16 ;
      RECT 74.825 3.37 75.23 3.7 ;
      RECT 74.825 2.53 75.23 2.86 ;
      RECT 74.825 7.305 74.995 10.595 ;
      RECT 74.825 9.605 75.23 9.935 ;
      RECT 74.825 8.765 75.23 9.095 ;
      RECT 72.75 4.421 72.755 4.593 ;
      RECT 72.745 4.414 72.75 4.683 ;
      RECT 72.74 4.408 72.745 4.702 ;
      RECT 72.72 4.402 72.74 4.712 ;
      RECT 72.705 4.397 72.72 4.72 ;
      RECT 72.668 4.391 72.705 4.718 ;
      RECT 72.582 4.377 72.668 4.714 ;
      RECT 72.496 4.359 72.582 4.709 ;
      RECT 72.41 4.34 72.496 4.703 ;
      RECT 72.38 4.328 72.41 4.699 ;
      RECT 72.36 4.322 72.38 4.698 ;
      RECT 72.295 4.32 72.36 4.696 ;
      RECT 72.28 4.32 72.295 4.688 ;
      RECT 72.265 4.32 72.28 4.675 ;
      RECT 72.26 4.32 72.265 4.665 ;
      RECT 72.245 4.32 72.26 4.643 ;
      RECT 72.23 4.32 72.245 4.61 ;
      RECT 72.225 4.32 72.23 4.588 ;
      RECT 72.215 4.32 72.225 4.57 ;
      RECT 72.2 4.32 72.215 4.548 ;
      RECT 72.18 4.32 72.2 4.51 ;
      RECT 72.53 3.605 72.565 4.044 ;
      RECT 72.53 3.605 72.57 4.043 ;
      RECT 72.475 3.665 72.57 4.042 ;
      RECT 72.34 3.837 72.57 4.041 ;
      RECT 72.45 3.715 72.57 4.041 ;
      RECT 72.34 3.837 72.595 4.031 ;
      RECT 72.395 3.782 72.675 3.948 ;
      RECT 72.57 3.576 72.575 4.039 ;
      RECT 72.425 3.752 72.715 3.825 ;
      RECT 72.44 3.735 72.57 4.041 ;
      RECT 72.575 3.575 72.745 3.763 ;
      RECT 72.565 3.578 72.745 3.763 ;
      RECT 72.07 3.455 72.24 3.765 ;
      RECT 72.07 3.455 72.245 3.738 ;
      RECT 72.07 3.455 72.25 3.715 ;
      RECT 72.07 3.455 72.26 3.665 ;
      RECT 72.065 3.56 72.26 3.635 ;
      RECT 72.1 3.13 72.27 3.608 ;
      RECT 72.1 3.13 72.285 3.529 ;
      RECT 72.09 3.34 72.285 3.529 ;
      RECT 72.1 3.14 72.295 3.444 ;
      RECT 72.03 3.882 72.035 4.085 ;
      RECT 72.02 3.87 72.03 4.195 ;
      RECT 71.995 3.87 72.02 4.235 ;
      RECT 71.915 3.87 71.995 4.32 ;
      RECT 71.905 3.87 71.915 4.39 ;
      RECT 71.88 3.87 71.905 4.413 ;
      RECT 71.86 3.87 71.88 4.448 ;
      RECT 71.815 3.88 71.86 4.491 ;
      RECT 71.805 3.892 71.815 4.528 ;
      RECT 71.785 3.906 71.805 4.548 ;
      RECT 71.775 3.924 71.785 4.564 ;
      RECT 71.76 3.95 71.775 4.574 ;
      RECT 71.745 3.991 71.76 4.588 ;
      RECT 71.735 4.026 71.745 4.598 ;
      RECT 71.73 4.042 71.735 4.603 ;
      RECT 71.72 4.057 71.73 4.608 ;
      RECT 71.7 4.1 71.72 4.618 ;
      RECT 71.68 4.137 71.7 4.631 ;
      RECT 71.645 4.16 71.68 4.649 ;
      RECT 71.635 4.174 71.645 4.665 ;
      RECT 71.615 4.184 71.635 4.675 ;
      RECT 71.61 4.193 71.615 4.683 ;
      RECT 71.6 4.2 71.61 4.69 ;
      RECT 71.59 4.207 71.6 4.698 ;
      RECT 71.575 4.217 71.59 4.706 ;
      RECT 71.565 4.231 71.575 4.716 ;
      RECT 71.555 4.243 71.565 4.728 ;
      RECT 71.54 4.265 71.555 4.741 ;
      RECT 71.53 4.287 71.54 4.752 ;
      RECT 71.52 4.307 71.53 4.761 ;
      RECT 71.515 4.322 71.52 4.768 ;
      RECT 71.485 4.355 71.515 4.782 ;
      RECT 71.475 4.39 71.485 4.797 ;
      RECT 71.47 4.397 71.475 4.803 ;
      RECT 71.45 4.412 71.47 4.81 ;
      RECT 71.445 4.427 71.45 4.818 ;
      RECT 71.44 4.436 71.445 4.823 ;
      RECT 71.425 4.442 71.44 4.83 ;
      RECT 71.42 4.448 71.425 4.838 ;
      RECT 71.415 4.452 71.42 4.845 ;
      RECT 71.41 4.456 71.415 4.855 ;
      RECT 71.4 4.461 71.41 4.865 ;
      RECT 71.38 4.472 71.4 4.893 ;
      RECT 71.365 4.484 71.38 4.92 ;
      RECT 71.345 4.497 71.365 4.945 ;
      RECT 71.325 4.512 71.345 4.969 ;
      RECT 71.31 4.527 71.325 4.984 ;
      RECT 71.305 4.538 71.31 4.993 ;
      RECT 71.24 4.583 71.305 5.003 ;
      RECT 71.205 4.642 71.24 5.016 ;
      RECT 71.2 4.665 71.205 5.022 ;
      RECT 71.195 4.672 71.2 5.024 ;
      RECT 71.18 4.682 71.195 5.027 ;
      RECT 71.15 4.707 71.18 5.031 ;
      RECT 71.145 4.725 71.15 5.035 ;
      RECT 71.14 4.732 71.145 5.036 ;
      RECT 71.12 4.74 71.14 5.04 ;
      RECT 71.11 4.747 71.12 5.044 ;
      RECT 71.066 4.758 71.11 5.051 ;
      RECT 70.98 4.786 71.066 5.067 ;
      RECT 70.92 4.81 70.98 5.085 ;
      RECT 70.875 4.82 70.92 5.099 ;
      RECT 70.816 4.828 70.875 5.113 ;
      RECT 70.73 4.835 70.816 5.132 ;
      RECT 70.705 4.84 70.73 5.147 ;
      RECT 70.625 4.843 70.705 5.15 ;
      RECT 70.545 4.847 70.625 5.137 ;
      RECT 70.536 4.85 70.545 5.122 ;
      RECT 70.45 4.85 70.536 5.107 ;
      RECT 70.39 4.852 70.45 5.084 ;
      RECT 70.386 4.855 70.39 5.074 ;
      RECT 70.3 4.855 70.386 5.059 ;
      RECT 70.225 4.855 70.3 5.035 ;
      RECT 71.54 3.864 71.55 4.04 ;
      RECT 71.495 3.831 71.54 4.04 ;
      RECT 71.45 3.782 71.495 4.04 ;
      RECT 71.42 3.752 71.45 4.041 ;
      RECT 71.415 3.735 71.42 4.042 ;
      RECT 71.39 3.715 71.415 4.043 ;
      RECT 71.375 3.69 71.39 4.044 ;
      RECT 71.37 3.677 71.375 4.045 ;
      RECT 71.365 3.671 71.37 4.043 ;
      RECT 71.36 3.663 71.365 4.037 ;
      RECT 71.335 3.655 71.36 4.017 ;
      RECT 71.315 3.644 71.335 3.988 ;
      RECT 71.285 3.629 71.315 3.959 ;
      RECT 71.265 3.615 71.285 3.931 ;
      RECT 71.255 3.609 71.265 3.91 ;
      RECT 71.25 3.606 71.255 3.893 ;
      RECT 71.245 3.603 71.25 3.878 ;
      RECT 71.23 3.598 71.245 3.843 ;
      RECT 71.225 3.594 71.23 3.81 ;
      RECT 71.205 3.589 71.225 3.786 ;
      RECT 71.175 3.581 71.205 3.751 ;
      RECT 71.16 3.575 71.175 3.728 ;
      RECT 71.12 3.568 71.16 3.713 ;
      RECT 71.095 3.56 71.12 3.693 ;
      RECT 71.075 3.555 71.095 3.683 ;
      RECT 71.04 3.549 71.075 3.678 ;
      RECT 70.995 3.54 71.04 3.677 ;
      RECT 70.965 3.536 70.995 3.679 ;
      RECT 70.88 3.544 70.965 3.683 ;
      RECT 70.81 3.555 70.88 3.705 ;
      RECT 70.797 3.561 70.81 3.728 ;
      RECT 70.711 3.568 70.797 3.75 ;
      RECT 70.625 3.58 70.711 3.787 ;
      RECT 70.625 3.957 70.635 4.195 ;
      RECT 70.62 3.586 70.625 3.81 ;
      RECT 70.615 3.842 70.625 4.195 ;
      RECT 70.615 3.587 70.62 3.815 ;
      RECT 70.61 3.588 70.615 4.195 ;
      RECT 70.586 3.59 70.61 4.196 ;
      RECT 70.5 3.598 70.586 4.198 ;
      RECT 70.48 3.612 70.5 4.201 ;
      RECT 70.475 3.64 70.48 4.202 ;
      RECT 70.47 3.652 70.475 4.203 ;
      RECT 70.465 3.667 70.47 4.204 ;
      RECT 70.455 3.697 70.465 4.205 ;
      RECT 70.45 3.735 70.455 4.203 ;
      RECT 70.445 3.755 70.45 4.198 ;
      RECT 70.43 3.79 70.445 4.183 ;
      RECT 70.42 3.842 70.43 4.163 ;
      RECT 70.415 3.872 70.42 4.151 ;
      RECT 70.4 3.885 70.415 4.134 ;
      RECT 70.375 3.889 70.4 4.101 ;
      RECT 70.36 3.887 70.375 4.078 ;
      RECT 70.345 3.886 70.36 4.075 ;
      RECT 70.285 3.884 70.345 4.073 ;
      RECT 70.275 3.882 70.285 4.068 ;
      RECT 70.235 3.881 70.275 4.065 ;
      RECT 70.165 3.878 70.235 4.063 ;
      RECT 70.11 3.876 70.165 4.058 ;
      RECT 70.04 3.87 70.11 4.053 ;
      RECT 70.031 3.87 70.04 4.05 ;
      RECT 69.945 3.87 70.031 4.045 ;
      RECT 69.94 3.87 69.945 4.04 ;
      RECT 71.245 3.105 71.42 3.455 ;
      RECT 71.245 3.12 71.43 3.453 ;
      RECT 71.22 3.07 71.365 3.45 ;
      RECT 71.2 3.071 71.365 3.443 ;
      RECT 71.19 3.072 71.375 3.438 ;
      RECT 71.16 3.073 71.375 3.425 ;
      RECT 71.11 3.074 71.375 3.401 ;
      RECT 71.105 3.076 71.375 3.386 ;
      RECT 71.105 3.142 71.435 3.38 ;
      RECT 71.085 3.083 71.39 3.36 ;
      RECT 71.075 3.092 71.4 3.215 ;
      RECT 71.085 3.087 71.4 3.36 ;
      RECT 71.105 3.077 71.39 3.386 ;
      RECT 70.69 4.402 70.86 4.69 ;
      RECT 70.685 4.42 70.87 4.685 ;
      RECT 70.65 4.428 70.935 4.605 ;
      RECT 70.65 4.428 71.021 4.595 ;
      RECT 70.65 4.428 71.075 4.541 ;
      RECT 70.935 4.325 71.105 4.509 ;
      RECT 70.65 4.48 71.11 4.497 ;
      RECT 70.635 4.45 71.105 4.493 ;
      RECT 70.895 4.332 70.935 4.644 ;
      RECT 70.775 4.369 71.105 4.509 ;
      RECT 70.87 4.344 70.895 4.67 ;
      RECT 70.86 4.351 71.105 4.509 ;
      RECT 70.991 3.815 71.06 4.074 ;
      RECT 70.991 3.87 71.065 4.073 ;
      RECT 70.905 3.87 71.065 4.072 ;
      RECT 70.9 3.87 71.07 4.065 ;
      RECT 70.89 3.815 71.06 4.06 ;
      RECT 70.27 3.114 70.445 3.415 ;
      RECT 70.255 3.102 70.27 3.4 ;
      RECT 70.225 3.101 70.255 3.353 ;
      RECT 70.225 3.119 70.45 3.348 ;
      RECT 70.21 3.103 70.27 3.313 ;
      RECT 70.205 3.125 70.46 3.213 ;
      RECT 70.205 3.108 70.356 3.213 ;
      RECT 70.205 3.11 70.36 3.213 ;
      RECT 70.21 3.106 70.356 3.313 ;
      RECT 70.315 4.342 70.32 4.69 ;
      RECT 70.305 4.332 70.315 4.696 ;
      RECT 70.27 4.322 70.305 4.698 ;
      RECT 70.232 4.317 70.27 4.702 ;
      RECT 70.146 4.31 70.232 4.709 ;
      RECT 70.06 4.3 70.146 4.719 ;
      RECT 70.015 4.295 70.06 4.727 ;
      RECT 70.011 4.295 70.015 4.731 ;
      RECT 69.925 4.295 70.011 4.738 ;
      RECT 69.91 4.295 69.925 4.738 ;
      RECT 69.9 4.293 69.91 4.71 ;
      RECT 69.89 4.289 69.9 4.653 ;
      RECT 69.87 4.283 69.89 4.585 ;
      RECT 69.865 4.279 69.87 4.533 ;
      RECT 69.855 4.278 69.865 4.5 ;
      RECT 69.805 4.276 69.855 4.485 ;
      RECT 69.78 4.274 69.805 4.48 ;
      RECT 69.737 4.272 69.78 4.476 ;
      RECT 69.651 4.268 69.737 4.464 ;
      RECT 69.565 4.263 69.651 4.448 ;
      RECT 69.535 4.26 69.565 4.435 ;
      RECT 69.51 4.259 69.535 4.423 ;
      RECT 69.505 4.259 69.51 4.413 ;
      RECT 69.465 4.258 69.505 4.405 ;
      RECT 69.45 4.257 69.465 4.398 ;
      RECT 69.4 4.256 69.45 4.39 ;
      RECT 69.398 4.255 69.4 4.385 ;
      RECT 69.312 4.253 69.398 4.385 ;
      RECT 69.226 4.248 69.312 4.385 ;
      RECT 69.14 4.244 69.226 4.385 ;
      RECT 69.091 4.24 69.14 4.383 ;
      RECT 69.005 4.237 69.091 4.378 ;
      RECT 68.982 4.234 69.005 4.374 ;
      RECT 68.896 4.231 68.982 4.369 ;
      RECT 68.81 4.227 68.896 4.36 ;
      RECT 68.785 4.22 68.81 4.355 ;
      RECT 68.725 4.185 68.785 4.352 ;
      RECT 68.705 4.11 68.725 4.349 ;
      RECT 68.7 4.052 68.705 4.348 ;
      RECT 68.675 3.992 68.7 4.347 ;
      RECT 68.6 3.87 68.675 4.343 ;
      RECT 68.59 3.87 68.6 4.335 ;
      RECT 68.575 3.87 68.59 4.325 ;
      RECT 68.56 3.87 68.575 4.295 ;
      RECT 68.545 3.87 68.56 4.24 ;
      RECT 68.53 3.87 68.545 4.178 ;
      RECT 68.505 3.87 68.53 4.103 ;
      RECT 68.5 3.87 68.505 4.053 ;
      RECT 69.845 3.415 69.865 3.724 ;
      RECT 69.831 3.417 69.88 3.721 ;
      RECT 69.831 3.422 69.9 3.712 ;
      RECT 69.745 3.42 69.88 3.706 ;
      RECT 69.745 3.428 69.935 3.689 ;
      RECT 69.71 3.43 69.935 3.688 ;
      RECT 69.68 3.438 69.935 3.679 ;
      RECT 69.67 3.443 69.955 3.665 ;
      RECT 69.71 3.433 69.955 3.665 ;
      RECT 69.71 3.436 69.965 3.653 ;
      RECT 69.68 3.438 69.975 3.64 ;
      RECT 69.68 3.442 69.985 3.583 ;
      RECT 69.67 3.447 69.99 3.498 ;
      RECT 69.831 3.415 69.865 3.721 ;
      RECT 69.71 10.145 69.88 10.595 ;
      RECT 69.765 8.365 69.935 10.315 ;
      RECT 69.71 7.305 69.88 8.535 ;
      RECT 69.27 3.518 69.275 3.73 ;
      RECT 69.145 3.515 69.16 3.73 ;
      RECT 68.61 3.545 68.68 3.73 ;
      RECT 68.495 3.545 68.53 3.725 ;
      RECT 69.616 3.847 69.635 4.041 ;
      RECT 69.53 3.802 69.616 4.042 ;
      RECT 69.52 3.755 69.53 4.044 ;
      RECT 69.515 3.735 69.52 4.045 ;
      RECT 69.495 3.7 69.515 4.046 ;
      RECT 69.48 3.65 69.495 4.047 ;
      RECT 69.46 3.587 69.48 4.048 ;
      RECT 69.45 3.55 69.46 4.049 ;
      RECT 69.435 3.539 69.45 4.05 ;
      RECT 69.43 3.531 69.435 4.048 ;
      RECT 69.42 3.53 69.43 4.04 ;
      RECT 69.39 3.527 69.42 4.019 ;
      RECT 69.315 3.522 69.39 3.964 ;
      RECT 69.3 3.518 69.315 3.91 ;
      RECT 69.29 3.518 69.3 3.805 ;
      RECT 69.275 3.518 69.29 3.738 ;
      RECT 69.26 3.518 69.27 3.728 ;
      RECT 69.205 3.517 69.26 3.725 ;
      RECT 69.16 3.515 69.205 3.728 ;
      RECT 69.132 3.515 69.145 3.731 ;
      RECT 69.046 3.519 69.132 3.733 ;
      RECT 68.96 3.525 69.046 3.738 ;
      RECT 68.94 3.529 68.96 3.74 ;
      RECT 68.938 3.53 68.94 3.739 ;
      RECT 68.852 3.532 68.938 3.738 ;
      RECT 68.766 3.537 68.852 3.735 ;
      RECT 68.68 3.542 68.766 3.732 ;
      RECT 68.53 3.545 68.61 3.728 ;
      RECT 69.19 7.305 69.36 10.595 ;
      RECT 69.19 9.605 69.595 9.935 ;
      RECT 69.19 8.765 69.595 9.095 ;
      RECT 69.306 4.52 69.355 4.854 ;
      RECT 69.306 4.52 69.36 4.853 ;
      RECT 69.22 4.52 69.36 4.852 ;
      RECT 68.995 4.628 69.365 4.85 ;
      RECT 69.22 4.52 69.39 4.843 ;
      RECT 69.19 4.532 69.395 4.834 ;
      RECT 69.175 4.55 69.4 4.831 ;
      RECT 68.99 4.634 69.4 4.758 ;
      RECT 68.985 4.641 69.4 4.718 ;
      RECT 69 4.607 69.4 4.831 ;
      RECT 69.161 4.553 69.365 4.85 ;
      RECT 69.075 4.573 69.4 4.831 ;
      RECT 69.175 4.547 69.395 4.834 ;
      RECT 68.945 3.871 69.135 4.065 ;
      RECT 68.94 3.873 69.135 4.064 ;
      RECT 68.935 3.877 69.15 4.061 ;
      RECT 68.95 3.87 69.15 4.061 ;
      RECT 68.935 3.98 69.155 4.056 ;
      RECT 68.23 4.48 68.321 4.778 ;
      RECT 68.225 4.482 68.4 4.773 ;
      RECT 68.23 4.48 68.4 4.773 ;
      RECT 68.225 4.486 68.42 4.771 ;
      RECT 68.225 4.541 68.46 4.77 ;
      RECT 68.225 4.576 68.475 4.764 ;
      RECT 68.225 4.61 68.485 4.754 ;
      RECT 68.215 4.49 68.42 4.605 ;
      RECT 68.215 4.51 68.435 4.605 ;
      RECT 68.215 4.493 68.425 4.605 ;
      RECT 68.44 3.261 68.445 3.323 ;
      RECT 68.435 3.183 68.44 3.346 ;
      RECT 68.43 3.14 68.435 3.357 ;
      RECT 68.425 3.13 68.43 3.369 ;
      RECT 68.42 3.13 68.425 3.378 ;
      RECT 68.395 3.13 68.42 3.41 ;
      RECT 68.39 3.13 68.395 3.443 ;
      RECT 68.375 3.13 68.39 3.468 ;
      RECT 68.365 3.13 68.375 3.495 ;
      RECT 68.36 3.13 68.365 3.508 ;
      RECT 68.355 3.13 68.36 3.523 ;
      RECT 68.345 3.13 68.355 3.538 ;
      RECT 68.34 3.13 68.345 3.558 ;
      RECT 68.315 3.13 68.34 3.593 ;
      RECT 68.27 3.13 68.315 3.638 ;
      RECT 68.26 3.13 68.27 3.651 ;
      RECT 68.175 3.215 68.26 3.658 ;
      RECT 68.14 3.337 68.175 3.667 ;
      RECT 68.135 3.377 68.14 3.671 ;
      RECT 68.115 3.4 68.135 3.673 ;
      RECT 68.11 3.43 68.115 3.676 ;
      RECT 68.1 3.442 68.11 3.677 ;
      RECT 68.055 3.465 68.1 3.682 ;
      RECT 68.015 3.495 68.055 3.69 ;
      RECT 67.98 3.507 68.015 3.696 ;
      RECT 67.975 3.512 67.98 3.7 ;
      RECT 67.905 3.522 67.975 3.707 ;
      RECT 67.865 3.532 67.905 3.717 ;
      RECT 67.845 3.537 67.865 3.723 ;
      RECT 67.835 3.541 67.845 3.728 ;
      RECT 67.83 3.544 67.835 3.731 ;
      RECT 67.82 3.545 67.83 3.732 ;
      RECT 67.795 3.547 67.82 3.736 ;
      RECT 67.785 3.552 67.795 3.739 ;
      RECT 67.74 3.56 67.785 3.74 ;
      RECT 67.615 3.565 67.74 3.74 ;
      RECT 68.17 3.862 68.19 4.044 ;
      RECT 68.121 3.847 68.17 4.043 ;
      RECT 68.035 3.862 68.19 4.041 ;
      RECT 68.02 3.862 68.19 4.04 ;
      RECT 67.985 3.84 68.155 4.025 ;
      RECT 68.055 4.86 68.07 5.069 ;
      RECT 68.055 4.868 68.075 5.068 ;
      RECT 68 4.868 68.075 5.067 ;
      RECT 67.98 4.872 68.08 5.065 ;
      RECT 67.96 4.822 68 5.064 ;
      RECT 67.905 4.88 68.085 5.062 ;
      RECT 67.87 4.837 68 5.06 ;
      RECT 67.866 4.84 68.055 5.059 ;
      RECT 67.78 4.848 68.055 5.057 ;
      RECT 67.78 4.892 68.09 5.05 ;
      RECT 67.77 4.985 68.09 5.048 ;
      RECT 67.78 4.904 68.095 5.033 ;
      RECT 67.78 4.925 68.11 5.003 ;
      RECT 67.78 4.952 68.115 4.973 ;
      RECT 67.905 4.83 68 5.062 ;
      RECT 67.535 3.875 67.54 4.413 ;
      RECT 67.34 4.205 67.345 4.4 ;
      RECT 65.64 3.87 65.655 4.25 ;
      RECT 67.705 3.87 67.71 4.04 ;
      RECT 67.7 3.87 67.705 4.05 ;
      RECT 67.695 3.87 67.7 4.063 ;
      RECT 67.67 3.87 67.695 4.105 ;
      RECT 67.645 3.87 67.67 4.178 ;
      RECT 67.63 3.87 67.645 4.23 ;
      RECT 67.625 3.87 67.63 4.26 ;
      RECT 67.6 3.87 67.625 4.3 ;
      RECT 67.585 3.87 67.6 4.355 ;
      RECT 67.58 3.87 67.585 4.388 ;
      RECT 67.555 3.87 67.58 4.408 ;
      RECT 67.54 3.87 67.555 4.414 ;
      RECT 67.47 3.905 67.535 4.41 ;
      RECT 67.42 3.96 67.47 4.405 ;
      RECT 67.41 3.992 67.42 4.403 ;
      RECT 67.405 4.017 67.41 4.403 ;
      RECT 67.385 4.09 67.405 4.403 ;
      RECT 67.375 4.17 67.385 4.402 ;
      RECT 67.36 4.2 67.375 4.402 ;
      RECT 67.345 4.205 67.36 4.401 ;
      RECT 67.285 4.207 67.34 4.398 ;
      RECT 67.255 4.212 67.285 4.394 ;
      RECT 67.253 4.215 67.255 4.393 ;
      RECT 67.167 4.217 67.253 4.39 ;
      RECT 67.081 4.223 67.167 4.384 ;
      RECT 66.995 4.228 67.081 4.378 ;
      RECT 66.922 4.233 66.995 4.379 ;
      RECT 66.836 4.239 66.922 4.387 ;
      RECT 66.75 4.245 66.836 4.396 ;
      RECT 66.73 4.249 66.75 4.401 ;
      RECT 66.683 4.251 66.73 4.404 ;
      RECT 66.597 4.256 66.683 4.41 ;
      RECT 66.511 4.261 66.597 4.419 ;
      RECT 66.425 4.267 66.511 4.427 ;
      RECT 66.34 4.265 66.425 4.436 ;
      RECT 66.336 4.26 66.34 4.44 ;
      RECT 66.25 4.255 66.336 4.432 ;
      RECT 66.186 4.246 66.25 4.42 ;
      RECT 66.1 4.237 66.186 4.407 ;
      RECT 66.076 4.23 66.1 4.398 ;
      RECT 65.99 4.224 66.076 4.385 ;
      RECT 65.95 4.217 65.99 4.371 ;
      RECT 65.945 4.207 65.95 4.367 ;
      RECT 65.935 4.195 65.945 4.366 ;
      RECT 65.915 4.165 65.935 4.363 ;
      RECT 65.86 4.085 65.915 4.357 ;
      RECT 65.84 4.004 65.86 4.352 ;
      RECT 65.82 3.962 65.84 4.348 ;
      RECT 65.795 3.915 65.82 4.342 ;
      RECT 65.79 3.89 65.795 4.339 ;
      RECT 65.755 3.87 65.79 4.334 ;
      RECT 65.746 3.87 65.755 4.327 ;
      RECT 65.66 3.87 65.746 4.297 ;
      RECT 65.655 3.87 65.66 4.26 ;
      RECT 65.62 3.87 65.64 4.182 ;
      RECT 65.615 3.912 65.62 4.147 ;
      RECT 65.61 3.987 65.615 4.103 ;
      RECT 67.06 3.792 67.235 4.04 ;
      RECT 67.06 3.792 67.24 4.038 ;
      RECT 67.055 3.824 67.24 3.998 ;
      RECT 67.085 3.765 67.255 3.985 ;
      RECT 67.05 3.842 67.255 3.918 ;
      RECT 66.36 3.305 66.53 3.48 ;
      RECT 66.36 3.305 66.702 3.472 ;
      RECT 66.36 3.305 66.785 3.466 ;
      RECT 66.36 3.305 66.82 3.462 ;
      RECT 66.36 3.305 66.84 3.461 ;
      RECT 66.36 3.305 66.926 3.457 ;
      RECT 66.82 3.13 66.99 3.452 ;
      RECT 66.395 3.237 67.02 3.45 ;
      RECT 66.385 3.292 67.025 3.448 ;
      RECT 66.36 3.328 67.035 3.443 ;
      RECT 66.36 3.355 67.04 3.373 ;
      RECT 66.425 3.18 67 3.45 ;
      RECT 66.616 3.165 67 3.45 ;
      RECT 66.45 3.168 67 3.45 ;
      RECT 66.53 3.166 66.616 3.477 ;
      RECT 66.616 3.163 66.995 3.45 ;
      RECT 66.8 3.14 66.995 3.45 ;
      RECT 66.702 3.161 66.995 3.45 ;
      RECT 66.785 3.155 66.8 3.463 ;
      RECT 66.935 4.52 66.94 4.72 ;
      RECT 66.4 4.585 66.445 4.72 ;
      RECT 66.97 4.52 66.99 4.693 ;
      RECT 66.94 4.52 66.97 4.708 ;
      RECT 66.875 4.52 66.935 4.745 ;
      RECT 66.86 4.52 66.875 4.775 ;
      RECT 66.845 4.52 66.86 4.788 ;
      RECT 66.825 4.52 66.845 4.803 ;
      RECT 66.82 4.52 66.825 4.812 ;
      RECT 66.81 4.524 66.82 4.817 ;
      RECT 66.795 4.534 66.81 4.828 ;
      RECT 66.77 4.55 66.795 4.838 ;
      RECT 66.76 4.564 66.77 4.84 ;
      RECT 66.74 4.576 66.76 4.837 ;
      RECT 66.71 4.597 66.74 4.831 ;
      RECT 66.7 4.609 66.71 4.826 ;
      RECT 66.69 4.607 66.7 4.823 ;
      RECT 66.675 4.606 66.69 4.818 ;
      RECT 66.67 4.605 66.675 4.813 ;
      RECT 66.635 4.603 66.67 4.803 ;
      RECT 66.615 4.6 66.635 4.785 ;
      RECT 66.605 4.598 66.615 4.78 ;
      RECT 66.595 4.597 66.605 4.775 ;
      RECT 66.56 4.595 66.595 4.763 ;
      RECT 66.505 4.591 66.56 4.743 ;
      RECT 66.495 4.589 66.505 4.728 ;
      RECT 66.49 4.589 66.495 4.723 ;
      RECT 66.445 4.587 66.49 4.72 ;
      RECT 66.35 4.585 66.4 4.724 ;
      RECT 66.34 4.586 66.35 4.729 ;
      RECT 66.28 4.593 66.34 4.743 ;
      RECT 66.255 4.601 66.28 4.763 ;
      RECT 66.245 4.605 66.255 4.775 ;
      RECT 66.24 4.606 66.245 4.78 ;
      RECT 66.225 4.608 66.24 4.783 ;
      RECT 66.21 4.61 66.225 4.788 ;
      RECT 66.205 4.61 66.21 4.791 ;
      RECT 66.16 4.615 66.205 4.802 ;
      RECT 66.155 4.619 66.16 4.814 ;
      RECT 66.13 4.615 66.155 4.818 ;
      RECT 66.12 4.611 66.13 4.822 ;
      RECT 66.11 4.61 66.12 4.826 ;
      RECT 66.095 4.6 66.11 4.832 ;
      RECT 66.09 4.588 66.095 4.836 ;
      RECT 66.085 4.585 66.09 4.837 ;
      RECT 66.08 4.582 66.085 4.839 ;
      RECT 66.065 4.57 66.08 4.838 ;
      RECT 66.05 4.552 66.065 4.835 ;
      RECT 66.03 4.531 66.05 4.828 ;
      RECT 65.965 4.52 66.03 4.8 ;
      RECT 65.961 4.52 65.965 4.779 ;
      RECT 65.875 4.52 65.961 4.749 ;
      RECT 65.86 4.52 65.875 4.705 ;
      RECT 66.435 3.62 66.44 3.855 ;
      RECT 65.565 3.536 65.57 3.74 ;
      RECT 66.145 3.565 66.15 3.72 ;
      RECT 66.065 3.545 66.07 3.72 ;
      RECT 66.735 3.687 66.75 4.04 ;
      RECT 66.661 3.672 66.735 4.04 ;
      RECT 66.575 3.655 66.661 4.04 ;
      RECT 66.565 3.645 66.575 4.038 ;
      RECT 66.56 3.643 66.565 4.033 ;
      RECT 66.545 3.641 66.56 4.019 ;
      RECT 66.475 3.633 66.545 3.959 ;
      RECT 66.455 3.624 66.475 3.893 ;
      RECT 66.45 3.621 66.455 3.873 ;
      RECT 66.44 3.62 66.45 3.863 ;
      RECT 66.43 3.62 66.435 3.847 ;
      RECT 66.42 3.619 66.43 3.837 ;
      RECT 66.41 3.617 66.42 3.825 ;
      RECT 66.395 3.614 66.41 3.805 ;
      RECT 66.385 3.612 66.395 3.79 ;
      RECT 66.365 3.609 66.385 3.778 ;
      RECT 66.36 3.607 66.365 3.768 ;
      RECT 66.335 3.605 66.36 3.755 ;
      RECT 66.305 3.6 66.335 3.74 ;
      RECT 66.225 3.591 66.305 3.731 ;
      RECT 66.18 3.58 66.225 3.724 ;
      RECT 66.16 3.571 66.18 3.721 ;
      RECT 66.15 3.566 66.16 3.72 ;
      RECT 66.105 3.56 66.145 3.72 ;
      RECT 66.09 3.552 66.105 3.72 ;
      RECT 66.07 3.547 66.09 3.72 ;
      RECT 66.05 3.544 66.065 3.72 ;
      RECT 65.967 3.543 66.05 3.719 ;
      RECT 65.881 3.542 65.967 3.715 ;
      RECT 65.795 3.54 65.881 3.712 ;
      RECT 65.742 3.539 65.795 3.714 ;
      RECT 65.656 3.538 65.742 3.723 ;
      RECT 65.57 3.537 65.656 3.735 ;
      RECT 65.55 3.536 65.565 3.743 ;
      RECT 65.47 3.535 65.55 3.755 ;
      RECT 65.445 3.535 65.47 3.768 ;
      RECT 65.42 3.535 65.445 3.783 ;
      RECT 65.415 3.535 65.42 3.805 ;
      RECT 65.41 3.535 65.415 3.823 ;
      RECT 65.405 3.535 65.41 3.84 ;
      RECT 65.4 3.535 65.405 3.853 ;
      RECT 65.395 3.535 65.4 3.863 ;
      RECT 65.355 3.535 65.395 3.948 ;
      RECT 65.34 3.535 65.355 4.033 ;
      RECT 65.33 3.536 65.34 4.045 ;
      RECT 65.295 3.541 65.33 4.05 ;
      RECT 65.255 3.55 65.295 4.05 ;
      RECT 65.24 3.56 65.255 4.05 ;
      RECT 65.235 3.57 65.24 4.05 ;
      RECT 65.215 3.597 65.235 4.05 ;
      RECT 65.165 3.68 65.215 4.05 ;
      RECT 65.16 3.742 65.165 4.05 ;
      RECT 65.15 3.755 65.16 4.05 ;
      RECT 65.14 3.777 65.15 4.05 ;
      RECT 65.13 3.802 65.14 4.045 ;
      RECT 65.125 3.84 65.13 4.038 ;
      RECT 65.115 3.95 65.125 4.033 ;
      RECT 66.51 4.871 66.525 5.13 ;
      RECT 66.51 4.886 66.53 5.129 ;
      RECT 66.426 4.886 66.53 5.127 ;
      RECT 66.426 4.9 66.535 5.126 ;
      RECT 66.34 4.942 66.54 5.123 ;
      RECT 66.335 4.885 66.525 5.118 ;
      RECT 66.335 4.956 66.545 5.115 ;
      RECT 66.33 4.987 66.545 5.113 ;
      RECT 66.335 4.984 66.56 5.103 ;
      RECT 66.33 5.03 66.575 5.088 ;
      RECT 66.33 5.058 66.58 5.073 ;
      RECT 66.34 4.86 66.51 5.123 ;
      RECT 66.1 3.87 66.27 4.04 ;
      RECT 66.065 3.87 66.27 4.035 ;
      RECT 66.055 3.87 66.27 4.028 ;
      RECT 66.05 3.855 66.22 4.025 ;
      RECT 64.88 4.392 65.145 4.835 ;
      RECT 64.875 4.363 65.09 4.833 ;
      RECT 64.87 4.517 65.15 4.828 ;
      RECT 64.875 4.412 65.15 4.828 ;
      RECT 64.875 4.423 65.16 4.815 ;
      RECT 64.875 4.37 65.12 4.833 ;
      RECT 64.88 4.357 65.09 4.835 ;
      RECT 64.88 4.355 65.04 4.835 ;
      RECT 64.981 4.347 65.04 4.835 ;
      RECT 64.895 4.348 65.04 4.835 ;
      RECT 64.981 4.346 65.03 4.835 ;
      RECT 64.785 3.161 64.96 3.46 ;
      RECT 64.835 3.123 64.96 3.46 ;
      RECT 64.82 3.125 65.046 3.452 ;
      RECT 64.82 3.128 65.085 3.439 ;
      RECT 64.82 3.129 65.095 3.425 ;
      RECT 64.775 3.18 65.095 3.415 ;
      RECT 64.82 3.13 65.1 3.41 ;
      RECT 64.775 3.34 65.105 3.4 ;
      RECT 64.76 3.2 65.1 3.34 ;
      RECT 64.755 3.216 65.1 3.28 ;
      RECT 64.8 3.14 65.1 3.41 ;
      RECT 64.835 3.121 64.921 3.46 ;
      RECT 62.925 3.035 63.095 4.225 ;
      RECT 62.925 3.035 63.395 3.205 ;
      RECT 62.925 9.26 63.395 9.43 ;
      RECT 62.925 8.24 63.095 9.43 ;
      RECT 61.935 3.035 62.105 4.225 ;
      RECT 61.935 3.035 62.405 3.205 ;
      RECT 61.935 9.26 62.405 9.43 ;
      RECT 61.935 8.24 62.105 9.43 ;
      RECT 60.085 3.93 60.255 5.16 ;
      RECT 60.14 2.15 60.31 4.1 ;
      RECT 60.085 1.87 60.255 2.32 ;
      RECT 60.085 10.145 60.255 10.595 ;
      RECT 60.14 8.365 60.31 10.315 ;
      RECT 60.085 7.305 60.255 8.535 ;
      RECT 59.565 1.87 59.735 5.16 ;
      RECT 59.565 3.37 59.97 3.7 ;
      RECT 59.565 2.53 59.97 2.86 ;
      RECT 59.565 7.305 59.735 10.595 ;
      RECT 59.565 9.605 59.97 9.935 ;
      RECT 59.565 8.765 59.97 9.095 ;
      RECT 57.49 4.421 57.495 4.593 ;
      RECT 57.485 4.414 57.49 4.683 ;
      RECT 57.48 4.408 57.485 4.702 ;
      RECT 57.46 4.402 57.48 4.712 ;
      RECT 57.445 4.397 57.46 4.72 ;
      RECT 57.408 4.391 57.445 4.718 ;
      RECT 57.322 4.377 57.408 4.714 ;
      RECT 57.236 4.359 57.322 4.709 ;
      RECT 57.15 4.34 57.236 4.703 ;
      RECT 57.12 4.328 57.15 4.699 ;
      RECT 57.1 4.322 57.12 4.698 ;
      RECT 57.035 4.32 57.1 4.696 ;
      RECT 57.02 4.32 57.035 4.688 ;
      RECT 57.005 4.32 57.02 4.675 ;
      RECT 57 4.32 57.005 4.665 ;
      RECT 56.985 4.32 57 4.643 ;
      RECT 56.97 4.32 56.985 4.61 ;
      RECT 56.965 4.32 56.97 4.588 ;
      RECT 56.955 4.32 56.965 4.57 ;
      RECT 56.94 4.32 56.955 4.548 ;
      RECT 56.92 4.32 56.94 4.51 ;
      RECT 57.27 3.605 57.305 4.044 ;
      RECT 57.27 3.605 57.31 4.043 ;
      RECT 57.215 3.665 57.31 4.042 ;
      RECT 57.08 3.837 57.31 4.041 ;
      RECT 57.19 3.715 57.31 4.041 ;
      RECT 57.08 3.837 57.335 4.031 ;
      RECT 57.135 3.782 57.415 3.948 ;
      RECT 57.31 3.576 57.315 4.039 ;
      RECT 57.165 3.752 57.455 3.825 ;
      RECT 57.18 3.735 57.31 4.041 ;
      RECT 57.315 3.575 57.485 3.763 ;
      RECT 57.305 3.578 57.485 3.763 ;
      RECT 56.81 3.455 56.98 3.765 ;
      RECT 56.81 3.455 56.985 3.738 ;
      RECT 56.81 3.455 56.99 3.715 ;
      RECT 56.81 3.455 57 3.665 ;
      RECT 56.805 3.56 57 3.635 ;
      RECT 56.84 3.13 57.01 3.608 ;
      RECT 56.84 3.13 57.025 3.529 ;
      RECT 56.83 3.34 57.025 3.529 ;
      RECT 56.84 3.14 57.035 3.444 ;
      RECT 56.77 3.882 56.775 4.085 ;
      RECT 56.76 3.87 56.77 4.195 ;
      RECT 56.735 3.87 56.76 4.235 ;
      RECT 56.655 3.87 56.735 4.32 ;
      RECT 56.645 3.87 56.655 4.39 ;
      RECT 56.62 3.87 56.645 4.413 ;
      RECT 56.6 3.87 56.62 4.448 ;
      RECT 56.555 3.88 56.6 4.491 ;
      RECT 56.545 3.892 56.555 4.528 ;
      RECT 56.525 3.906 56.545 4.548 ;
      RECT 56.515 3.924 56.525 4.564 ;
      RECT 56.5 3.95 56.515 4.574 ;
      RECT 56.485 3.991 56.5 4.588 ;
      RECT 56.475 4.026 56.485 4.598 ;
      RECT 56.47 4.042 56.475 4.603 ;
      RECT 56.46 4.057 56.47 4.608 ;
      RECT 56.44 4.1 56.46 4.618 ;
      RECT 56.42 4.137 56.44 4.631 ;
      RECT 56.385 4.16 56.42 4.649 ;
      RECT 56.375 4.174 56.385 4.665 ;
      RECT 56.355 4.184 56.375 4.675 ;
      RECT 56.35 4.193 56.355 4.683 ;
      RECT 56.34 4.2 56.35 4.69 ;
      RECT 56.33 4.207 56.34 4.698 ;
      RECT 56.315 4.217 56.33 4.706 ;
      RECT 56.305 4.231 56.315 4.716 ;
      RECT 56.295 4.243 56.305 4.728 ;
      RECT 56.28 4.265 56.295 4.741 ;
      RECT 56.27 4.287 56.28 4.752 ;
      RECT 56.26 4.307 56.27 4.761 ;
      RECT 56.255 4.322 56.26 4.768 ;
      RECT 56.225 4.355 56.255 4.782 ;
      RECT 56.215 4.39 56.225 4.797 ;
      RECT 56.21 4.397 56.215 4.803 ;
      RECT 56.19 4.412 56.21 4.81 ;
      RECT 56.185 4.427 56.19 4.818 ;
      RECT 56.18 4.436 56.185 4.823 ;
      RECT 56.165 4.442 56.18 4.83 ;
      RECT 56.16 4.448 56.165 4.838 ;
      RECT 56.155 4.452 56.16 4.845 ;
      RECT 56.15 4.456 56.155 4.855 ;
      RECT 56.14 4.461 56.15 4.865 ;
      RECT 56.12 4.472 56.14 4.893 ;
      RECT 56.105 4.484 56.12 4.92 ;
      RECT 56.085 4.497 56.105 4.945 ;
      RECT 56.065 4.512 56.085 4.969 ;
      RECT 56.05 4.527 56.065 4.984 ;
      RECT 56.045 4.538 56.05 4.993 ;
      RECT 55.98 4.583 56.045 5.003 ;
      RECT 55.945 4.642 55.98 5.016 ;
      RECT 55.94 4.665 55.945 5.022 ;
      RECT 55.935 4.672 55.94 5.024 ;
      RECT 55.92 4.682 55.935 5.027 ;
      RECT 55.89 4.707 55.92 5.031 ;
      RECT 55.885 4.725 55.89 5.035 ;
      RECT 55.88 4.732 55.885 5.036 ;
      RECT 55.86 4.74 55.88 5.04 ;
      RECT 55.85 4.747 55.86 5.044 ;
      RECT 55.806 4.758 55.85 5.051 ;
      RECT 55.72 4.786 55.806 5.067 ;
      RECT 55.66 4.81 55.72 5.085 ;
      RECT 55.615 4.82 55.66 5.099 ;
      RECT 55.556 4.828 55.615 5.113 ;
      RECT 55.47 4.835 55.556 5.132 ;
      RECT 55.445 4.84 55.47 5.147 ;
      RECT 55.365 4.843 55.445 5.15 ;
      RECT 55.285 4.847 55.365 5.137 ;
      RECT 55.276 4.85 55.285 5.122 ;
      RECT 55.19 4.85 55.276 5.107 ;
      RECT 55.13 4.852 55.19 5.084 ;
      RECT 55.126 4.855 55.13 5.074 ;
      RECT 55.04 4.855 55.126 5.059 ;
      RECT 54.965 4.855 55.04 5.035 ;
      RECT 56.28 3.864 56.29 4.04 ;
      RECT 56.235 3.831 56.28 4.04 ;
      RECT 56.19 3.782 56.235 4.04 ;
      RECT 56.16 3.752 56.19 4.041 ;
      RECT 56.155 3.735 56.16 4.042 ;
      RECT 56.13 3.715 56.155 4.043 ;
      RECT 56.115 3.69 56.13 4.044 ;
      RECT 56.11 3.677 56.115 4.045 ;
      RECT 56.105 3.671 56.11 4.043 ;
      RECT 56.1 3.663 56.105 4.037 ;
      RECT 56.075 3.655 56.1 4.017 ;
      RECT 56.055 3.644 56.075 3.988 ;
      RECT 56.025 3.629 56.055 3.959 ;
      RECT 56.005 3.615 56.025 3.931 ;
      RECT 55.995 3.609 56.005 3.91 ;
      RECT 55.99 3.606 55.995 3.893 ;
      RECT 55.985 3.603 55.99 3.878 ;
      RECT 55.97 3.598 55.985 3.843 ;
      RECT 55.965 3.594 55.97 3.81 ;
      RECT 55.945 3.589 55.965 3.786 ;
      RECT 55.915 3.581 55.945 3.751 ;
      RECT 55.9 3.575 55.915 3.728 ;
      RECT 55.86 3.568 55.9 3.713 ;
      RECT 55.835 3.56 55.86 3.693 ;
      RECT 55.815 3.555 55.835 3.683 ;
      RECT 55.78 3.549 55.815 3.678 ;
      RECT 55.735 3.54 55.78 3.677 ;
      RECT 55.705 3.536 55.735 3.679 ;
      RECT 55.62 3.544 55.705 3.683 ;
      RECT 55.55 3.555 55.62 3.705 ;
      RECT 55.537 3.561 55.55 3.728 ;
      RECT 55.451 3.568 55.537 3.75 ;
      RECT 55.365 3.58 55.451 3.787 ;
      RECT 55.365 3.957 55.375 4.195 ;
      RECT 55.36 3.586 55.365 3.81 ;
      RECT 55.355 3.842 55.365 4.195 ;
      RECT 55.355 3.587 55.36 3.815 ;
      RECT 55.35 3.588 55.355 4.195 ;
      RECT 55.326 3.59 55.35 4.196 ;
      RECT 55.24 3.598 55.326 4.198 ;
      RECT 55.22 3.612 55.24 4.201 ;
      RECT 55.215 3.64 55.22 4.202 ;
      RECT 55.21 3.652 55.215 4.203 ;
      RECT 55.205 3.667 55.21 4.204 ;
      RECT 55.195 3.697 55.205 4.205 ;
      RECT 55.19 3.735 55.195 4.203 ;
      RECT 55.185 3.755 55.19 4.198 ;
      RECT 55.17 3.79 55.185 4.183 ;
      RECT 55.16 3.842 55.17 4.163 ;
      RECT 55.155 3.872 55.16 4.151 ;
      RECT 55.14 3.885 55.155 4.134 ;
      RECT 55.115 3.889 55.14 4.101 ;
      RECT 55.1 3.887 55.115 4.078 ;
      RECT 55.085 3.886 55.1 4.075 ;
      RECT 55.025 3.884 55.085 4.073 ;
      RECT 55.015 3.882 55.025 4.068 ;
      RECT 54.975 3.881 55.015 4.065 ;
      RECT 54.905 3.878 54.975 4.063 ;
      RECT 54.85 3.876 54.905 4.058 ;
      RECT 54.78 3.87 54.85 4.053 ;
      RECT 54.771 3.87 54.78 4.05 ;
      RECT 54.685 3.87 54.771 4.045 ;
      RECT 54.68 3.87 54.685 4.04 ;
      RECT 55.985 3.105 56.16 3.455 ;
      RECT 55.985 3.12 56.17 3.453 ;
      RECT 55.96 3.07 56.105 3.45 ;
      RECT 55.94 3.071 56.105 3.443 ;
      RECT 55.93 3.072 56.115 3.438 ;
      RECT 55.9 3.073 56.115 3.425 ;
      RECT 55.85 3.074 56.115 3.401 ;
      RECT 55.845 3.076 56.115 3.386 ;
      RECT 55.845 3.142 56.175 3.38 ;
      RECT 55.825 3.083 56.13 3.36 ;
      RECT 55.815 3.092 56.14 3.215 ;
      RECT 55.825 3.087 56.14 3.36 ;
      RECT 55.845 3.077 56.13 3.386 ;
      RECT 55.43 4.402 55.6 4.69 ;
      RECT 55.425 4.42 55.61 4.685 ;
      RECT 55.39 4.428 55.675 4.605 ;
      RECT 55.39 4.428 55.761 4.595 ;
      RECT 55.39 4.428 55.815 4.541 ;
      RECT 55.675 4.325 55.845 4.509 ;
      RECT 55.39 4.48 55.85 4.497 ;
      RECT 55.375 4.45 55.845 4.493 ;
      RECT 55.635 4.332 55.675 4.644 ;
      RECT 55.515 4.369 55.845 4.509 ;
      RECT 55.61 4.344 55.635 4.67 ;
      RECT 55.6 4.351 55.845 4.509 ;
      RECT 55.731 3.815 55.8 4.074 ;
      RECT 55.731 3.87 55.805 4.073 ;
      RECT 55.645 3.87 55.805 4.072 ;
      RECT 55.64 3.87 55.81 4.065 ;
      RECT 55.63 3.815 55.8 4.06 ;
      RECT 55.01 3.114 55.185 3.415 ;
      RECT 54.995 3.102 55.01 3.4 ;
      RECT 54.965 3.101 54.995 3.353 ;
      RECT 54.965 3.119 55.19 3.348 ;
      RECT 54.95 3.103 55.01 3.313 ;
      RECT 54.945 3.125 55.2 3.213 ;
      RECT 54.945 3.108 55.096 3.213 ;
      RECT 54.945 3.11 55.1 3.213 ;
      RECT 54.95 3.106 55.096 3.313 ;
      RECT 55.055 4.342 55.06 4.69 ;
      RECT 55.045 4.332 55.055 4.696 ;
      RECT 55.01 4.322 55.045 4.698 ;
      RECT 54.972 4.317 55.01 4.702 ;
      RECT 54.886 4.31 54.972 4.709 ;
      RECT 54.8 4.3 54.886 4.719 ;
      RECT 54.755 4.295 54.8 4.727 ;
      RECT 54.751 4.295 54.755 4.731 ;
      RECT 54.665 4.295 54.751 4.738 ;
      RECT 54.65 4.295 54.665 4.738 ;
      RECT 54.64 4.293 54.65 4.71 ;
      RECT 54.63 4.289 54.64 4.653 ;
      RECT 54.61 4.283 54.63 4.585 ;
      RECT 54.605 4.279 54.61 4.533 ;
      RECT 54.595 4.278 54.605 4.5 ;
      RECT 54.545 4.276 54.595 4.485 ;
      RECT 54.52 4.274 54.545 4.48 ;
      RECT 54.477 4.272 54.52 4.476 ;
      RECT 54.391 4.268 54.477 4.464 ;
      RECT 54.305 4.263 54.391 4.448 ;
      RECT 54.275 4.26 54.305 4.435 ;
      RECT 54.25 4.259 54.275 4.423 ;
      RECT 54.245 4.259 54.25 4.413 ;
      RECT 54.205 4.258 54.245 4.405 ;
      RECT 54.19 4.257 54.205 4.398 ;
      RECT 54.14 4.256 54.19 4.39 ;
      RECT 54.138 4.255 54.14 4.385 ;
      RECT 54.052 4.253 54.138 4.385 ;
      RECT 53.966 4.248 54.052 4.385 ;
      RECT 53.88 4.244 53.966 4.385 ;
      RECT 53.831 4.24 53.88 4.383 ;
      RECT 53.745 4.237 53.831 4.378 ;
      RECT 53.722 4.234 53.745 4.374 ;
      RECT 53.636 4.231 53.722 4.369 ;
      RECT 53.55 4.227 53.636 4.36 ;
      RECT 53.525 4.22 53.55 4.355 ;
      RECT 53.465 4.185 53.525 4.352 ;
      RECT 53.445 4.11 53.465 4.349 ;
      RECT 53.44 4.052 53.445 4.348 ;
      RECT 53.415 3.992 53.44 4.347 ;
      RECT 53.34 3.87 53.415 4.343 ;
      RECT 53.33 3.87 53.34 4.335 ;
      RECT 53.315 3.87 53.33 4.325 ;
      RECT 53.3 3.87 53.315 4.295 ;
      RECT 53.285 3.87 53.3 4.24 ;
      RECT 53.27 3.87 53.285 4.178 ;
      RECT 53.245 3.87 53.27 4.103 ;
      RECT 53.24 3.87 53.245 4.053 ;
      RECT 54.585 3.415 54.605 3.724 ;
      RECT 54.571 3.417 54.62 3.721 ;
      RECT 54.571 3.422 54.64 3.712 ;
      RECT 54.485 3.42 54.62 3.706 ;
      RECT 54.485 3.428 54.675 3.689 ;
      RECT 54.45 3.43 54.675 3.688 ;
      RECT 54.42 3.438 54.675 3.679 ;
      RECT 54.41 3.443 54.695 3.665 ;
      RECT 54.45 3.433 54.695 3.665 ;
      RECT 54.45 3.436 54.705 3.653 ;
      RECT 54.42 3.438 54.715 3.64 ;
      RECT 54.42 3.442 54.725 3.583 ;
      RECT 54.41 3.447 54.73 3.498 ;
      RECT 54.571 3.415 54.605 3.721 ;
      RECT 54.45 10.145 54.62 10.595 ;
      RECT 54.505 8.365 54.675 10.315 ;
      RECT 54.45 7.305 54.62 8.535 ;
      RECT 54.01 3.518 54.015 3.73 ;
      RECT 53.885 3.515 53.9 3.73 ;
      RECT 53.35 3.545 53.42 3.73 ;
      RECT 53.235 3.545 53.27 3.725 ;
      RECT 54.356 3.847 54.375 4.041 ;
      RECT 54.27 3.802 54.356 4.042 ;
      RECT 54.26 3.755 54.27 4.044 ;
      RECT 54.255 3.735 54.26 4.045 ;
      RECT 54.235 3.7 54.255 4.046 ;
      RECT 54.22 3.65 54.235 4.047 ;
      RECT 54.2 3.587 54.22 4.048 ;
      RECT 54.19 3.55 54.2 4.049 ;
      RECT 54.175 3.539 54.19 4.05 ;
      RECT 54.17 3.531 54.175 4.048 ;
      RECT 54.16 3.53 54.17 4.04 ;
      RECT 54.13 3.527 54.16 4.019 ;
      RECT 54.055 3.522 54.13 3.964 ;
      RECT 54.04 3.518 54.055 3.91 ;
      RECT 54.03 3.518 54.04 3.805 ;
      RECT 54.015 3.518 54.03 3.738 ;
      RECT 54 3.518 54.01 3.728 ;
      RECT 53.945 3.517 54 3.725 ;
      RECT 53.9 3.515 53.945 3.728 ;
      RECT 53.872 3.515 53.885 3.731 ;
      RECT 53.786 3.519 53.872 3.733 ;
      RECT 53.7 3.525 53.786 3.738 ;
      RECT 53.68 3.529 53.7 3.74 ;
      RECT 53.678 3.53 53.68 3.739 ;
      RECT 53.592 3.532 53.678 3.738 ;
      RECT 53.506 3.537 53.592 3.735 ;
      RECT 53.42 3.542 53.506 3.732 ;
      RECT 53.27 3.545 53.35 3.728 ;
      RECT 53.93 7.305 54.1 10.595 ;
      RECT 53.93 9.605 54.335 9.935 ;
      RECT 53.93 8.765 54.335 9.095 ;
      RECT 54.046 4.52 54.095 4.854 ;
      RECT 54.046 4.52 54.1 4.853 ;
      RECT 53.96 4.52 54.1 4.852 ;
      RECT 53.735 4.628 54.105 4.85 ;
      RECT 53.96 4.52 54.13 4.843 ;
      RECT 53.93 4.532 54.135 4.834 ;
      RECT 53.915 4.55 54.14 4.831 ;
      RECT 53.73 4.634 54.14 4.758 ;
      RECT 53.725 4.641 54.14 4.718 ;
      RECT 53.74 4.607 54.14 4.831 ;
      RECT 53.901 4.553 54.105 4.85 ;
      RECT 53.815 4.573 54.14 4.831 ;
      RECT 53.915 4.547 54.135 4.834 ;
      RECT 53.685 3.871 53.875 4.065 ;
      RECT 53.68 3.873 53.875 4.064 ;
      RECT 53.675 3.877 53.89 4.061 ;
      RECT 53.69 3.87 53.89 4.061 ;
      RECT 53.675 3.98 53.895 4.056 ;
      RECT 52.97 4.48 53.061 4.778 ;
      RECT 52.965 4.482 53.14 4.773 ;
      RECT 52.97 4.48 53.14 4.773 ;
      RECT 52.965 4.486 53.16 4.771 ;
      RECT 52.965 4.541 53.2 4.77 ;
      RECT 52.965 4.576 53.215 4.764 ;
      RECT 52.965 4.61 53.225 4.754 ;
      RECT 52.955 4.49 53.16 4.605 ;
      RECT 52.955 4.51 53.175 4.605 ;
      RECT 52.955 4.493 53.165 4.605 ;
      RECT 53.18 3.261 53.185 3.323 ;
      RECT 53.175 3.183 53.18 3.346 ;
      RECT 53.17 3.14 53.175 3.357 ;
      RECT 53.165 3.13 53.17 3.369 ;
      RECT 53.16 3.13 53.165 3.378 ;
      RECT 53.135 3.13 53.16 3.41 ;
      RECT 53.13 3.13 53.135 3.443 ;
      RECT 53.115 3.13 53.13 3.468 ;
      RECT 53.105 3.13 53.115 3.495 ;
      RECT 53.1 3.13 53.105 3.508 ;
      RECT 53.095 3.13 53.1 3.523 ;
      RECT 53.085 3.13 53.095 3.538 ;
      RECT 53.08 3.13 53.085 3.558 ;
      RECT 53.055 3.13 53.08 3.593 ;
      RECT 53.01 3.13 53.055 3.638 ;
      RECT 53 3.13 53.01 3.651 ;
      RECT 52.915 3.215 53 3.658 ;
      RECT 52.88 3.337 52.915 3.667 ;
      RECT 52.875 3.377 52.88 3.671 ;
      RECT 52.855 3.4 52.875 3.673 ;
      RECT 52.85 3.43 52.855 3.676 ;
      RECT 52.84 3.442 52.85 3.677 ;
      RECT 52.795 3.465 52.84 3.682 ;
      RECT 52.755 3.495 52.795 3.69 ;
      RECT 52.72 3.507 52.755 3.696 ;
      RECT 52.715 3.512 52.72 3.7 ;
      RECT 52.645 3.522 52.715 3.707 ;
      RECT 52.605 3.532 52.645 3.717 ;
      RECT 52.585 3.537 52.605 3.723 ;
      RECT 52.575 3.541 52.585 3.728 ;
      RECT 52.57 3.544 52.575 3.731 ;
      RECT 52.56 3.545 52.57 3.732 ;
      RECT 52.535 3.547 52.56 3.736 ;
      RECT 52.525 3.552 52.535 3.739 ;
      RECT 52.48 3.56 52.525 3.74 ;
      RECT 52.355 3.565 52.48 3.74 ;
      RECT 52.91 3.862 52.93 4.044 ;
      RECT 52.861 3.847 52.91 4.043 ;
      RECT 52.775 3.862 52.93 4.041 ;
      RECT 52.76 3.862 52.93 4.04 ;
      RECT 52.725 3.84 52.895 4.025 ;
      RECT 52.795 4.86 52.81 5.069 ;
      RECT 52.795 4.868 52.815 5.068 ;
      RECT 52.74 4.868 52.815 5.067 ;
      RECT 52.72 4.872 52.82 5.065 ;
      RECT 52.7 4.822 52.74 5.064 ;
      RECT 52.645 4.88 52.825 5.062 ;
      RECT 52.61 4.837 52.74 5.06 ;
      RECT 52.606 4.84 52.795 5.059 ;
      RECT 52.52 4.848 52.795 5.057 ;
      RECT 52.52 4.892 52.83 5.05 ;
      RECT 52.51 4.985 52.83 5.048 ;
      RECT 52.52 4.904 52.835 5.033 ;
      RECT 52.52 4.925 52.85 5.003 ;
      RECT 52.52 4.952 52.855 4.973 ;
      RECT 52.645 4.83 52.74 5.062 ;
      RECT 52.275 3.875 52.28 4.413 ;
      RECT 52.08 4.205 52.085 4.4 ;
      RECT 50.38 3.87 50.395 4.25 ;
      RECT 52.445 3.87 52.45 4.04 ;
      RECT 52.44 3.87 52.445 4.05 ;
      RECT 52.435 3.87 52.44 4.063 ;
      RECT 52.41 3.87 52.435 4.105 ;
      RECT 52.385 3.87 52.41 4.178 ;
      RECT 52.37 3.87 52.385 4.23 ;
      RECT 52.365 3.87 52.37 4.26 ;
      RECT 52.34 3.87 52.365 4.3 ;
      RECT 52.325 3.87 52.34 4.355 ;
      RECT 52.32 3.87 52.325 4.388 ;
      RECT 52.295 3.87 52.32 4.408 ;
      RECT 52.28 3.87 52.295 4.414 ;
      RECT 52.21 3.905 52.275 4.41 ;
      RECT 52.16 3.96 52.21 4.405 ;
      RECT 52.15 3.992 52.16 4.403 ;
      RECT 52.145 4.017 52.15 4.403 ;
      RECT 52.125 4.09 52.145 4.403 ;
      RECT 52.115 4.17 52.125 4.402 ;
      RECT 52.1 4.2 52.115 4.402 ;
      RECT 52.085 4.205 52.1 4.401 ;
      RECT 52.025 4.207 52.08 4.398 ;
      RECT 51.995 4.212 52.025 4.394 ;
      RECT 51.993 4.215 51.995 4.393 ;
      RECT 51.907 4.217 51.993 4.39 ;
      RECT 51.821 4.223 51.907 4.384 ;
      RECT 51.735 4.228 51.821 4.378 ;
      RECT 51.662 4.233 51.735 4.379 ;
      RECT 51.576 4.239 51.662 4.387 ;
      RECT 51.49 4.245 51.576 4.396 ;
      RECT 51.47 4.249 51.49 4.401 ;
      RECT 51.423 4.251 51.47 4.404 ;
      RECT 51.337 4.256 51.423 4.41 ;
      RECT 51.251 4.261 51.337 4.419 ;
      RECT 51.165 4.267 51.251 4.427 ;
      RECT 51.08 4.265 51.165 4.436 ;
      RECT 51.076 4.26 51.08 4.44 ;
      RECT 50.99 4.255 51.076 4.432 ;
      RECT 50.926 4.246 50.99 4.42 ;
      RECT 50.84 4.237 50.926 4.407 ;
      RECT 50.816 4.23 50.84 4.398 ;
      RECT 50.73 4.224 50.816 4.385 ;
      RECT 50.69 4.217 50.73 4.371 ;
      RECT 50.685 4.207 50.69 4.367 ;
      RECT 50.675 4.195 50.685 4.366 ;
      RECT 50.655 4.165 50.675 4.363 ;
      RECT 50.6 4.085 50.655 4.357 ;
      RECT 50.58 4.004 50.6 4.352 ;
      RECT 50.56 3.962 50.58 4.348 ;
      RECT 50.535 3.915 50.56 4.342 ;
      RECT 50.53 3.89 50.535 4.339 ;
      RECT 50.495 3.87 50.53 4.334 ;
      RECT 50.486 3.87 50.495 4.327 ;
      RECT 50.4 3.87 50.486 4.297 ;
      RECT 50.395 3.87 50.4 4.26 ;
      RECT 50.36 3.87 50.38 4.182 ;
      RECT 50.355 3.912 50.36 4.147 ;
      RECT 50.35 3.987 50.355 4.103 ;
      RECT 51.8 3.792 51.975 4.04 ;
      RECT 51.8 3.792 51.98 4.038 ;
      RECT 51.795 3.824 51.98 3.998 ;
      RECT 51.825 3.765 51.995 3.985 ;
      RECT 51.79 3.842 51.995 3.918 ;
      RECT 51.1 3.305 51.27 3.48 ;
      RECT 51.1 3.305 51.442 3.472 ;
      RECT 51.1 3.305 51.525 3.466 ;
      RECT 51.1 3.305 51.56 3.462 ;
      RECT 51.1 3.305 51.58 3.461 ;
      RECT 51.1 3.305 51.666 3.457 ;
      RECT 51.56 3.13 51.73 3.452 ;
      RECT 51.135 3.237 51.76 3.45 ;
      RECT 51.125 3.292 51.765 3.448 ;
      RECT 51.1 3.328 51.775 3.443 ;
      RECT 51.1 3.355 51.78 3.373 ;
      RECT 51.165 3.18 51.74 3.45 ;
      RECT 51.356 3.165 51.74 3.45 ;
      RECT 51.19 3.168 51.74 3.45 ;
      RECT 51.27 3.166 51.356 3.477 ;
      RECT 51.356 3.163 51.735 3.45 ;
      RECT 51.54 3.14 51.735 3.45 ;
      RECT 51.442 3.161 51.735 3.45 ;
      RECT 51.525 3.155 51.54 3.463 ;
      RECT 51.675 4.52 51.68 4.72 ;
      RECT 51.14 4.585 51.185 4.72 ;
      RECT 51.71 4.52 51.73 4.693 ;
      RECT 51.68 4.52 51.71 4.708 ;
      RECT 51.615 4.52 51.675 4.745 ;
      RECT 51.6 4.52 51.615 4.775 ;
      RECT 51.585 4.52 51.6 4.788 ;
      RECT 51.565 4.52 51.585 4.803 ;
      RECT 51.56 4.52 51.565 4.812 ;
      RECT 51.55 4.524 51.56 4.817 ;
      RECT 51.535 4.534 51.55 4.828 ;
      RECT 51.51 4.55 51.535 4.838 ;
      RECT 51.5 4.564 51.51 4.84 ;
      RECT 51.48 4.576 51.5 4.837 ;
      RECT 51.45 4.597 51.48 4.831 ;
      RECT 51.44 4.609 51.45 4.826 ;
      RECT 51.43 4.607 51.44 4.823 ;
      RECT 51.415 4.606 51.43 4.818 ;
      RECT 51.41 4.605 51.415 4.813 ;
      RECT 51.375 4.603 51.41 4.803 ;
      RECT 51.355 4.6 51.375 4.785 ;
      RECT 51.345 4.598 51.355 4.78 ;
      RECT 51.335 4.597 51.345 4.775 ;
      RECT 51.3 4.595 51.335 4.763 ;
      RECT 51.245 4.591 51.3 4.743 ;
      RECT 51.235 4.589 51.245 4.728 ;
      RECT 51.23 4.589 51.235 4.723 ;
      RECT 51.185 4.587 51.23 4.72 ;
      RECT 51.09 4.585 51.14 4.724 ;
      RECT 51.08 4.586 51.09 4.729 ;
      RECT 51.02 4.593 51.08 4.743 ;
      RECT 50.995 4.601 51.02 4.763 ;
      RECT 50.985 4.605 50.995 4.775 ;
      RECT 50.98 4.606 50.985 4.78 ;
      RECT 50.965 4.608 50.98 4.783 ;
      RECT 50.95 4.61 50.965 4.788 ;
      RECT 50.945 4.61 50.95 4.791 ;
      RECT 50.9 4.615 50.945 4.802 ;
      RECT 50.895 4.619 50.9 4.814 ;
      RECT 50.87 4.615 50.895 4.818 ;
      RECT 50.86 4.611 50.87 4.822 ;
      RECT 50.85 4.61 50.86 4.826 ;
      RECT 50.835 4.6 50.85 4.832 ;
      RECT 50.83 4.588 50.835 4.836 ;
      RECT 50.825 4.585 50.83 4.837 ;
      RECT 50.82 4.582 50.825 4.839 ;
      RECT 50.805 4.57 50.82 4.838 ;
      RECT 50.79 4.552 50.805 4.835 ;
      RECT 50.77 4.531 50.79 4.828 ;
      RECT 50.705 4.52 50.77 4.8 ;
      RECT 50.701 4.52 50.705 4.779 ;
      RECT 50.615 4.52 50.701 4.749 ;
      RECT 50.6 4.52 50.615 4.705 ;
      RECT 51.175 3.62 51.18 3.855 ;
      RECT 50.305 3.536 50.31 3.74 ;
      RECT 50.885 3.565 50.89 3.72 ;
      RECT 50.805 3.545 50.81 3.72 ;
      RECT 51.475 3.687 51.49 4.04 ;
      RECT 51.401 3.672 51.475 4.04 ;
      RECT 51.315 3.655 51.401 4.04 ;
      RECT 51.305 3.645 51.315 4.038 ;
      RECT 51.3 3.643 51.305 4.033 ;
      RECT 51.285 3.641 51.3 4.019 ;
      RECT 51.215 3.633 51.285 3.959 ;
      RECT 51.195 3.624 51.215 3.893 ;
      RECT 51.19 3.621 51.195 3.873 ;
      RECT 51.18 3.62 51.19 3.863 ;
      RECT 51.17 3.62 51.175 3.847 ;
      RECT 51.16 3.619 51.17 3.837 ;
      RECT 51.15 3.617 51.16 3.825 ;
      RECT 51.135 3.614 51.15 3.805 ;
      RECT 51.125 3.612 51.135 3.79 ;
      RECT 51.105 3.609 51.125 3.778 ;
      RECT 51.1 3.607 51.105 3.768 ;
      RECT 51.075 3.605 51.1 3.755 ;
      RECT 51.045 3.6 51.075 3.74 ;
      RECT 50.965 3.591 51.045 3.731 ;
      RECT 50.92 3.58 50.965 3.724 ;
      RECT 50.9 3.571 50.92 3.721 ;
      RECT 50.89 3.566 50.9 3.72 ;
      RECT 50.845 3.56 50.885 3.72 ;
      RECT 50.83 3.552 50.845 3.72 ;
      RECT 50.81 3.547 50.83 3.72 ;
      RECT 50.79 3.544 50.805 3.72 ;
      RECT 50.707 3.543 50.79 3.719 ;
      RECT 50.621 3.542 50.707 3.715 ;
      RECT 50.535 3.54 50.621 3.712 ;
      RECT 50.482 3.539 50.535 3.714 ;
      RECT 50.396 3.538 50.482 3.723 ;
      RECT 50.31 3.537 50.396 3.735 ;
      RECT 50.29 3.536 50.305 3.743 ;
      RECT 50.21 3.535 50.29 3.755 ;
      RECT 50.185 3.535 50.21 3.768 ;
      RECT 50.16 3.535 50.185 3.783 ;
      RECT 50.155 3.535 50.16 3.805 ;
      RECT 50.15 3.535 50.155 3.823 ;
      RECT 50.145 3.535 50.15 3.84 ;
      RECT 50.14 3.535 50.145 3.853 ;
      RECT 50.135 3.535 50.14 3.863 ;
      RECT 50.095 3.535 50.135 3.948 ;
      RECT 50.08 3.535 50.095 4.033 ;
      RECT 50.07 3.536 50.08 4.045 ;
      RECT 50.035 3.541 50.07 4.05 ;
      RECT 49.995 3.55 50.035 4.05 ;
      RECT 49.98 3.56 49.995 4.05 ;
      RECT 49.975 3.57 49.98 4.05 ;
      RECT 49.955 3.597 49.975 4.05 ;
      RECT 49.905 3.68 49.955 4.05 ;
      RECT 49.9 3.742 49.905 4.05 ;
      RECT 49.89 3.755 49.9 4.05 ;
      RECT 49.88 3.777 49.89 4.05 ;
      RECT 49.87 3.802 49.88 4.045 ;
      RECT 49.865 3.84 49.87 4.038 ;
      RECT 49.855 3.95 49.865 4.033 ;
      RECT 51.25 4.871 51.265 5.13 ;
      RECT 51.25 4.886 51.27 5.129 ;
      RECT 51.166 4.886 51.27 5.127 ;
      RECT 51.166 4.9 51.275 5.126 ;
      RECT 51.08 4.942 51.28 5.123 ;
      RECT 51.075 4.885 51.265 5.118 ;
      RECT 51.075 4.956 51.285 5.115 ;
      RECT 51.07 4.987 51.285 5.113 ;
      RECT 51.075 4.984 51.3 5.103 ;
      RECT 51.07 5.03 51.315 5.088 ;
      RECT 51.07 5.058 51.32 5.073 ;
      RECT 51.08 4.86 51.25 5.123 ;
      RECT 50.84 3.87 51.01 4.04 ;
      RECT 50.805 3.87 51.01 4.035 ;
      RECT 50.795 3.87 51.01 4.028 ;
      RECT 50.79 3.855 50.96 4.025 ;
      RECT 49.62 4.392 49.885 4.835 ;
      RECT 49.615 4.363 49.83 4.833 ;
      RECT 49.61 4.517 49.89 4.828 ;
      RECT 49.615 4.412 49.89 4.828 ;
      RECT 49.615 4.423 49.9 4.815 ;
      RECT 49.615 4.37 49.86 4.833 ;
      RECT 49.62 4.357 49.83 4.835 ;
      RECT 49.62 4.355 49.78 4.835 ;
      RECT 49.721 4.347 49.78 4.835 ;
      RECT 49.635 4.348 49.78 4.835 ;
      RECT 49.721 4.346 49.77 4.835 ;
      RECT 49.525 3.161 49.7 3.46 ;
      RECT 49.575 3.123 49.7 3.46 ;
      RECT 49.56 3.125 49.786 3.452 ;
      RECT 49.56 3.128 49.825 3.439 ;
      RECT 49.56 3.129 49.835 3.425 ;
      RECT 49.515 3.18 49.835 3.415 ;
      RECT 49.56 3.13 49.84 3.41 ;
      RECT 49.515 3.34 49.845 3.4 ;
      RECT 49.5 3.2 49.84 3.34 ;
      RECT 49.495 3.216 49.84 3.28 ;
      RECT 49.54 3.14 49.84 3.41 ;
      RECT 49.575 3.121 49.661 3.46 ;
      RECT 47.665 3.035 47.835 4.225 ;
      RECT 47.665 3.035 48.135 3.205 ;
      RECT 47.665 9.26 48.135 9.43 ;
      RECT 47.665 8.24 47.835 9.43 ;
      RECT 46.675 3.035 46.845 4.225 ;
      RECT 46.675 3.035 47.145 3.205 ;
      RECT 46.675 9.26 47.145 9.43 ;
      RECT 46.675 8.24 46.845 9.43 ;
      RECT 44.825 3.93 44.995 5.16 ;
      RECT 44.88 2.15 45.05 4.1 ;
      RECT 44.825 1.87 44.995 2.32 ;
      RECT 44.825 10.145 44.995 10.595 ;
      RECT 44.88 8.365 45.05 10.315 ;
      RECT 44.825 7.305 44.995 8.535 ;
      RECT 44.305 1.87 44.475 5.16 ;
      RECT 44.305 3.37 44.71 3.7 ;
      RECT 44.305 2.53 44.71 2.86 ;
      RECT 44.305 7.305 44.475 10.595 ;
      RECT 44.305 9.605 44.71 9.935 ;
      RECT 44.305 8.765 44.71 9.095 ;
      RECT 42.23 4.421 42.235 4.593 ;
      RECT 42.225 4.414 42.23 4.683 ;
      RECT 42.22 4.408 42.225 4.702 ;
      RECT 42.2 4.402 42.22 4.712 ;
      RECT 42.185 4.397 42.2 4.72 ;
      RECT 42.148 4.391 42.185 4.718 ;
      RECT 42.062 4.377 42.148 4.714 ;
      RECT 41.976 4.359 42.062 4.709 ;
      RECT 41.89 4.34 41.976 4.703 ;
      RECT 41.86 4.328 41.89 4.699 ;
      RECT 41.84 4.322 41.86 4.698 ;
      RECT 41.775 4.32 41.84 4.696 ;
      RECT 41.76 4.32 41.775 4.688 ;
      RECT 41.745 4.32 41.76 4.675 ;
      RECT 41.74 4.32 41.745 4.665 ;
      RECT 41.725 4.32 41.74 4.643 ;
      RECT 41.71 4.32 41.725 4.61 ;
      RECT 41.705 4.32 41.71 4.588 ;
      RECT 41.695 4.32 41.705 4.57 ;
      RECT 41.68 4.32 41.695 4.548 ;
      RECT 41.66 4.32 41.68 4.51 ;
      RECT 42.01 3.605 42.045 4.044 ;
      RECT 42.01 3.605 42.05 4.043 ;
      RECT 41.955 3.665 42.05 4.042 ;
      RECT 41.82 3.837 42.05 4.041 ;
      RECT 41.93 3.715 42.05 4.041 ;
      RECT 41.82 3.837 42.075 4.031 ;
      RECT 41.875 3.782 42.155 3.948 ;
      RECT 42.05 3.576 42.055 4.039 ;
      RECT 41.905 3.752 42.195 3.825 ;
      RECT 41.92 3.735 42.05 4.041 ;
      RECT 42.055 3.575 42.225 3.763 ;
      RECT 42.045 3.578 42.225 3.763 ;
      RECT 41.55 3.455 41.72 3.765 ;
      RECT 41.55 3.455 41.725 3.738 ;
      RECT 41.55 3.455 41.73 3.715 ;
      RECT 41.55 3.455 41.74 3.665 ;
      RECT 41.545 3.56 41.74 3.635 ;
      RECT 41.58 3.13 41.75 3.608 ;
      RECT 41.58 3.13 41.765 3.529 ;
      RECT 41.57 3.34 41.765 3.529 ;
      RECT 41.58 3.14 41.775 3.444 ;
      RECT 41.51 3.882 41.515 4.085 ;
      RECT 41.5 3.87 41.51 4.195 ;
      RECT 41.475 3.87 41.5 4.235 ;
      RECT 41.395 3.87 41.475 4.32 ;
      RECT 41.385 3.87 41.395 4.39 ;
      RECT 41.36 3.87 41.385 4.413 ;
      RECT 41.34 3.87 41.36 4.448 ;
      RECT 41.295 3.88 41.34 4.491 ;
      RECT 41.285 3.892 41.295 4.528 ;
      RECT 41.265 3.906 41.285 4.548 ;
      RECT 41.255 3.924 41.265 4.564 ;
      RECT 41.24 3.95 41.255 4.574 ;
      RECT 41.225 3.991 41.24 4.588 ;
      RECT 41.215 4.026 41.225 4.598 ;
      RECT 41.21 4.042 41.215 4.603 ;
      RECT 41.2 4.057 41.21 4.608 ;
      RECT 41.18 4.1 41.2 4.618 ;
      RECT 41.16 4.137 41.18 4.631 ;
      RECT 41.125 4.16 41.16 4.649 ;
      RECT 41.115 4.174 41.125 4.665 ;
      RECT 41.095 4.184 41.115 4.675 ;
      RECT 41.09 4.193 41.095 4.683 ;
      RECT 41.08 4.2 41.09 4.69 ;
      RECT 41.07 4.207 41.08 4.698 ;
      RECT 41.055 4.217 41.07 4.706 ;
      RECT 41.045 4.231 41.055 4.716 ;
      RECT 41.035 4.243 41.045 4.728 ;
      RECT 41.02 4.265 41.035 4.741 ;
      RECT 41.01 4.287 41.02 4.752 ;
      RECT 41 4.307 41.01 4.761 ;
      RECT 40.995 4.322 41 4.768 ;
      RECT 40.965 4.355 40.995 4.782 ;
      RECT 40.955 4.39 40.965 4.797 ;
      RECT 40.95 4.397 40.955 4.803 ;
      RECT 40.93 4.412 40.95 4.81 ;
      RECT 40.925 4.427 40.93 4.818 ;
      RECT 40.92 4.436 40.925 4.823 ;
      RECT 40.905 4.442 40.92 4.83 ;
      RECT 40.9 4.448 40.905 4.838 ;
      RECT 40.895 4.452 40.9 4.845 ;
      RECT 40.89 4.456 40.895 4.855 ;
      RECT 40.88 4.461 40.89 4.865 ;
      RECT 40.86 4.472 40.88 4.893 ;
      RECT 40.845 4.484 40.86 4.92 ;
      RECT 40.825 4.497 40.845 4.945 ;
      RECT 40.805 4.512 40.825 4.969 ;
      RECT 40.79 4.527 40.805 4.984 ;
      RECT 40.785 4.538 40.79 4.993 ;
      RECT 40.72 4.583 40.785 5.003 ;
      RECT 40.685 4.642 40.72 5.016 ;
      RECT 40.68 4.665 40.685 5.022 ;
      RECT 40.675 4.672 40.68 5.024 ;
      RECT 40.66 4.682 40.675 5.027 ;
      RECT 40.63 4.707 40.66 5.031 ;
      RECT 40.625 4.725 40.63 5.035 ;
      RECT 40.62 4.732 40.625 5.036 ;
      RECT 40.6 4.74 40.62 5.04 ;
      RECT 40.59 4.747 40.6 5.044 ;
      RECT 40.546 4.758 40.59 5.051 ;
      RECT 40.46 4.786 40.546 5.067 ;
      RECT 40.4 4.81 40.46 5.085 ;
      RECT 40.355 4.82 40.4 5.099 ;
      RECT 40.296 4.828 40.355 5.113 ;
      RECT 40.21 4.835 40.296 5.132 ;
      RECT 40.185 4.84 40.21 5.147 ;
      RECT 40.105 4.843 40.185 5.15 ;
      RECT 40.025 4.847 40.105 5.137 ;
      RECT 40.016 4.85 40.025 5.122 ;
      RECT 39.93 4.85 40.016 5.107 ;
      RECT 39.87 4.852 39.93 5.084 ;
      RECT 39.866 4.855 39.87 5.074 ;
      RECT 39.78 4.855 39.866 5.059 ;
      RECT 39.705 4.855 39.78 5.035 ;
      RECT 41.02 3.864 41.03 4.04 ;
      RECT 40.975 3.831 41.02 4.04 ;
      RECT 40.93 3.782 40.975 4.04 ;
      RECT 40.9 3.752 40.93 4.041 ;
      RECT 40.895 3.735 40.9 4.042 ;
      RECT 40.87 3.715 40.895 4.043 ;
      RECT 40.855 3.69 40.87 4.044 ;
      RECT 40.85 3.677 40.855 4.045 ;
      RECT 40.845 3.671 40.85 4.043 ;
      RECT 40.84 3.663 40.845 4.037 ;
      RECT 40.815 3.655 40.84 4.017 ;
      RECT 40.795 3.644 40.815 3.988 ;
      RECT 40.765 3.629 40.795 3.959 ;
      RECT 40.745 3.615 40.765 3.931 ;
      RECT 40.735 3.609 40.745 3.91 ;
      RECT 40.73 3.606 40.735 3.893 ;
      RECT 40.725 3.603 40.73 3.878 ;
      RECT 40.71 3.598 40.725 3.843 ;
      RECT 40.705 3.594 40.71 3.81 ;
      RECT 40.685 3.589 40.705 3.786 ;
      RECT 40.655 3.581 40.685 3.751 ;
      RECT 40.64 3.575 40.655 3.728 ;
      RECT 40.6 3.568 40.64 3.713 ;
      RECT 40.575 3.56 40.6 3.693 ;
      RECT 40.555 3.555 40.575 3.683 ;
      RECT 40.52 3.549 40.555 3.678 ;
      RECT 40.475 3.54 40.52 3.677 ;
      RECT 40.445 3.536 40.475 3.679 ;
      RECT 40.36 3.544 40.445 3.683 ;
      RECT 40.29 3.555 40.36 3.705 ;
      RECT 40.277 3.561 40.29 3.728 ;
      RECT 40.191 3.568 40.277 3.75 ;
      RECT 40.105 3.58 40.191 3.787 ;
      RECT 40.105 3.957 40.115 4.195 ;
      RECT 40.1 3.586 40.105 3.81 ;
      RECT 40.095 3.842 40.105 4.195 ;
      RECT 40.095 3.587 40.1 3.815 ;
      RECT 40.09 3.588 40.095 4.195 ;
      RECT 40.066 3.59 40.09 4.196 ;
      RECT 39.98 3.598 40.066 4.198 ;
      RECT 39.96 3.612 39.98 4.201 ;
      RECT 39.955 3.64 39.96 4.202 ;
      RECT 39.95 3.652 39.955 4.203 ;
      RECT 39.945 3.667 39.95 4.204 ;
      RECT 39.935 3.697 39.945 4.205 ;
      RECT 39.93 3.735 39.935 4.203 ;
      RECT 39.925 3.755 39.93 4.198 ;
      RECT 39.91 3.79 39.925 4.183 ;
      RECT 39.9 3.842 39.91 4.163 ;
      RECT 39.895 3.872 39.9 4.151 ;
      RECT 39.88 3.885 39.895 4.134 ;
      RECT 39.855 3.889 39.88 4.101 ;
      RECT 39.84 3.887 39.855 4.078 ;
      RECT 39.825 3.886 39.84 4.075 ;
      RECT 39.765 3.884 39.825 4.073 ;
      RECT 39.755 3.882 39.765 4.068 ;
      RECT 39.715 3.881 39.755 4.065 ;
      RECT 39.645 3.878 39.715 4.063 ;
      RECT 39.59 3.876 39.645 4.058 ;
      RECT 39.52 3.87 39.59 4.053 ;
      RECT 39.511 3.87 39.52 4.05 ;
      RECT 39.425 3.87 39.511 4.045 ;
      RECT 39.42 3.87 39.425 4.04 ;
      RECT 40.725 3.105 40.9 3.455 ;
      RECT 40.725 3.12 40.91 3.453 ;
      RECT 40.7 3.07 40.845 3.45 ;
      RECT 40.68 3.071 40.845 3.443 ;
      RECT 40.67 3.072 40.855 3.438 ;
      RECT 40.64 3.073 40.855 3.425 ;
      RECT 40.59 3.074 40.855 3.401 ;
      RECT 40.585 3.076 40.855 3.386 ;
      RECT 40.585 3.142 40.915 3.38 ;
      RECT 40.565 3.083 40.87 3.36 ;
      RECT 40.555 3.092 40.88 3.215 ;
      RECT 40.565 3.087 40.88 3.36 ;
      RECT 40.585 3.077 40.87 3.386 ;
      RECT 40.17 4.402 40.34 4.69 ;
      RECT 40.165 4.42 40.35 4.685 ;
      RECT 40.13 4.428 40.415 4.605 ;
      RECT 40.13 4.428 40.501 4.595 ;
      RECT 40.13 4.428 40.555 4.541 ;
      RECT 40.415 4.325 40.585 4.509 ;
      RECT 40.13 4.48 40.59 4.497 ;
      RECT 40.115 4.45 40.585 4.493 ;
      RECT 40.375 4.332 40.415 4.644 ;
      RECT 40.255 4.369 40.585 4.509 ;
      RECT 40.35 4.344 40.375 4.67 ;
      RECT 40.34 4.351 40.585 4.509 ;
      RECT 40.471 3.815 40.54 4.074 ;
      RECT 40.471 3.87 40.545 4.073 ;
      RECT 40.385 3.87 40.545 4.072 ;
      RECT 40.38 3.87 40.55 4.065 ;
      RECT 40.37 3.815 40.54 4.06 ;
      RECT 39.75 3.114 39.925 3.415 ;
      RECT 39.735 3.102 39.75 3.4 ;
      RECT 39.705 3.101 39.735 3.353 ;
      RECT 39.705 3.119 39.93 3.348 ;
      RECT 39.69 3.103 39.75 3.313 ;
      RECT 39.685 3.125 39.94 3.213 ;
      RECT 39.685 3.108 39.836 3.213 ;
      RECT 39.685 3.11 39.84 3.213 ;
      RECT 39.69 3.106 39.836 3.313 ;
      RECT 39.795 4.342 39.8 4.69 ;
      RECT 39.785 4.332 39.795 4.696 ;
      RECT 39.75 4.322 39.785 4.698 ;
      RECT 39.712 4.317 39.75 4.702 ;
      RECT 39.626 4.31 39.712 4.709 ;
      RECT 39.54 4.3 39.626 4.719 ;
      RECT 39.495 4.295 39.54 4.727 ;
      RECT 39.491 4.295 39.495 4.731 ;
      RECT 39.405 4.295 39.491 4.738 ;
      RECT 39.39 4.295 39.405 4.738 ;
      RECT 39.38 4.293 39.39 4.71 ;
      RECT 39.37 4.289 39.38 4.653 ;
      RECT 39.35 4.283 39.37 4.585 ;
      RECT 39.345 4.279 39.35 4.533 ;
      RECT 39.335 4.278 39.345 4.5 ;
      RECT 39.285 4.276 39.335 4.485 ;
      RECT 39.26 4.274 39.285 4.48 ;
      RECT 39.217 4.272 39.26 4.476 ;
      RECT 39.131 4.268 39.217 4.464 ;
      RECT 39.045 4.263 39.131 4.448 ;
      RECT 39.015 4.26 39.045 4.435 ;
      RECT 38.99 4.259 39.015 4.423 ;
      RECT 38.985 4.259 38.99 4.413 ;
      RECT 38.945 4.258 38.985 4.405 ;
      RECT 38.93 4.257 38.945 4.398 ;
      RECT 38.88 4.256 38.93 4.39 ;
      RECT 38.878 4.255 38.88 4.385 ;
      RECT 38.792 4.253 38.878 4.385 ;
      RECT 38.706 4.248 38.792 4.385 ;
      RECT 38.62 4.244 38.706 4.385 ;
      RECT 38.571 4.24 38.62 4.383 ;
      RECT 38.485 4.237 38.571 4.378 ;
      RECT 38.462 4.234 38.485 4.374 ;
      RECT 38.376 4.231 38.462 4.369 ;
      RECT 38.29 4.227 38.376 4.36 ;
      RECT 38.265 4.22 38.29 4.355 ;
      RECT 38.205 4.185 38.265 4.352 ;
      RECT 38.185 4.11 38.205 4.349 ;
      RECT 38.18 4.052 38.185 4.348 ;
      RECT 38.155 3.992 38.18 4.347 ;
      RECT 38.08 3.87 38.155 4.343 ;
      RECT 38.07 3.87 38.08 4.335 ;
      RECT 38.055 3.87 38.07 4.325 ;
      RECT 38.04 3.87 38.055 4.295 ;
      RECT 38.025 3.87 38.04 4.24 ;
      RECT 38.01 3.87 38.025 4.178 ;
      RECT 37.985 3.87 38.01 4.103 ;
      RECT 37.98 3.87 37.985 4.053 ;
      RECT 39.325 3.415 39.345 3.724 ;
      RECT 39.311 3.417 39.36 3.721 ;
      RECT 39.311 3.422 39.38 3.712 ;
      RECT 39.225 3.42 39.36 3.706 ;
      RECT 39.225 3.428 39.415 3.689 ;
      RECT 39.19 3.43 39.415 3.688 ;
      RECT 39.16 3.438 39.415 3.679 ;
      RECT 39.15 3.443 39.435 3.665 ;
      RECT 39.19 3.433 39.435 3.665 ;
      RECT 39.19 3.436 39.445 3.653 ;
      RECT 39.16 3.438 39.455 3.64 ;
      RECT 39.16 3.442 39.465 3.583 ;
      RECT 39.15 3.447 39.47 3.498 ;
      RECT 39.311 3.415 39.345 3.721 ;
      RECT 39.19 10.145 39.36 10.595 ;
      RECT 39.245 8.365 39.415 10.315 ;
      RECT 39.19 7.305 39.36 8.535 ;
      RECT 38.75 3.518 38.755 3.73 ;
      RECT 38.625 3.515 38.64 3.73 ;
      RECT 38.09 3.545 38.16 3.73 ;
      RECT 37.975 3.545 38.01 3.725 ;
      RECT 39.096 3.847 39.115 4.041 ;
      RECT 39.01 3.802 39.096 4.042 ;
      RECT 39 3.755 39.01 4.044 ;
      RECT 38.995 3.735 39 4.045 ;
      RECT 38.975 3.7 38.995 4.046 ;
      RECT 38.96 3.65 38.975 4.047 ;
      RECT 38.94 3.587 38.96 4.048 ;
      RECT 38.93 3.55 38.94 4.049 ;
      RECT 38.915 3.539 38.93 4.05 ;
      RECT 38.91 3.531 38.915 4.048 ;
      RECT 38.9 3.53 38.91 4.04 ;
      RECT 38.87 3.527 38.9 4.019 ;
      RECT 38.795 3.522 38.87 3.964 ;
      RECT 38.78 3.518 38.795 3.91 ;
      RECT 38.77 3.518 38.78 3.805 ;
      RECT 38.755 3.518 38.77 3.738 ;
      RECT 38.74 3.518 38.75 3.728 ;
      RECT 38.685 3.517 38.74 3.725 ;
      RECT 38.64 3.515 38.685 3.728 ;
      RECT 38.612 3.515 38.625 3.731 ;
      RECT 38.526 3.519 38.612 3.733 ;
      RECT 38.44 3.525 38.526 3.738 ;
      RECT 38.42 3.529 38.44 3.74 ;
      RECT 38.418 3.53 38.42 3.739 ;
      RECT 38.332 3.532 38.418 3.738 ;
      RECT 38.246 3.537 38.332 3.735 ;
      RECT 38.16 3.542 38.246 3.732 ;
      RECT 38.01 3.545 38.09 3.728 ;
      RECT 38.67 7.305 38.84 10.595 ;
      RECT 38.67 9.605 39.075 9.935 ;
      RECT 38.67 8.765 39.075 9.095 ;
      RECT 38.786 4.52 38.835 4.854 ;
      RECT 38.786 4.52 38.84 4.853 ;
      RECT 38.7 4.52 38.84 4.852 ;
      RECT 38.475 4.628 38.845 4.85 ;
      RECT 38.7 4.52 38.87 4.843 ;
      RECT 38.67 4.532 38.875 4.834 ;
      RECT 38.655 4.55 38.88 4.831 ;
      RECT 38.47 4.634 38.88 4.758 ;
      RECT 38.465 4.641 38.88 4.718 ;
      RECT 38.48 4.607 38.88 4.831 ;
      RECT 38.641 4.553 38.845 4.85 ;
      RECT 38.555 4.573 38.88 4.831 ;
      RECT 38.655 4.547 38.875 4.834 ;
      RECT 38.425 3.871 38.615 4.065 ;
      RECT 38.42 3.873 38.615 4.064 ;
      RECT 38.415 3.877 38.63 4.061 ;
      RECT 38.43 3.87 38.63 4.061 ;
      RECT 38.415 3.98 38.635 4.056 ;
      RECT 37.71 4.48 37.801 4.778 ;
      RECT 37.705 4.482 37.88 4.773 ;
      RECT 37.71 4.48 37.88 4.773 ;
      RECT 37.705 4.486 37.9 4.771 ;
      RECT 37.705 4.541 37.94 4.77 ;
      RECT 37.705 4.576 37.955 4.764 ;
      RECT 37.705 4.61 37.965 4.754 ;
      RECT 37.695 4.49 37.9 4.605 ;
      RECT 37.695 4.51 37.915 4.605 ;
      RECT 37.695 4.493 37.905 4.605 ;
      RECT 37.92 3.261 37.925 3.323 ;
      RECT 37.915 3.183 37.92 3.346 ;
      RECT 37.91 3.14 37.915 3.357 ;
      RECT 37.905 3.13 37.91 3.369 ;
      RECT 37.9 3.13 37.905 3.378 ;
      RECT 37.875 3.13 37.9 3.41 ;
      RECT 37.87 3.13 37.875 3.443 ;
      RECT 37.855 3.13 37.87 3.468 ;
      RECT 37.845 3.13 37.855 3.495 ;
      RECT 37.84 3.13 37.845 3.508 ;
      RECT 37.835 3.13 37.84 3.523 ;
      RECT 37.825 3.13 37.835 3.538 ;
      RECT 37.82 3.13 37.825 3.558 ;
      RECT 37.795 3.13 37.82 3.593 ;
      RECT 37.75 3.13 37.795 3.638 ;
      RECT 37.74 3.13 37.75 3.651 ;
      RECT 37.655 3.215 37.74 3.658 ;
      RECT 37.62 3.337 37.655 3.667 ;
      RECT 37.615 3.377 37.62 3.671 ;
      RECT 37.595 3.4 37.615 3.673 ;
      RECT 37.59 3.43 37.595 3.676 ;
      RECT 37.58 3.442 37.59 3.677 ;
      RECT 37.535 3.465 37.58 3.682 ;
      RECT 37.495 3.495 37.535 3.69 ;
      RECT 37.46 3.507 37.495 3.696 ;
      RECT 37.455 3.512 37.46 3.7 ;
      RECT 37.385 3.522 37.455 3.707 ;
      RECT 37.345 3.532 37.385 3.717 ;
      RECT 37.325 3.537 37.345 3.723 ;
      RECT 37.315 3.541 37.325 3.728 ;
      RECT 37.31 3.544 37.315 3.731 ;
      RECT 37.3 3.545 37.31 3.732 ;
      RECT 37.275 3.547 37.3 3.736 ;
      RECT 37.265 3.552 37.275 3.739 ;
      RECT 37.22 3.56 37.265 3.74 ;
      RECT 37.095 3.565 37.22 3.74 ;
      RECT 37.65 3.862 37.67 4.044 ;
      RECT 37.601 3.847 37.65 4.043 ;
      RECT 37.515 3.862 37.67 4.041 ;
      RECT 37.5 3.862 37.67 4.04 ;
      RECT 37.465 3.84 37.635 4.025 ;
      RECT 37.535 4.86 37.55 5.069 ;
      RECT 37.535 4.868 37.555 5.068 ;
      RECT 37.48 4.868 37.555 5.067 ;
      RECT 37.46 4.872 37.56 5.065 ;
      RECT 37.44 4.822 37.48 5.064 ;
      RECT 37.385 4.88 37.565 5.062 ;
      RECT 37.35 4.837 37.48 5.06 ;
      RECT 37.346 4.84 37.535 5.059 ;
      RECT 37.26 4.848 37.535 5.057 ;
      RECT 37.26 4.892 37.57 5.05 ;
      RECT 37.25 4.985 37.57 5.048 ;
      RECT 37.26 4.904 37.575 5.033 ;
      RECT 37.26 4.925 37.59 5.003 ;
      RECT 37.26 4.952 37.595 4.973 ;
      RECT 37.385 4.83 37.48 5.062 ;
      RECT 37.015 3.875 37.02 4.413 ;
      RECT 36.82 4.205 36.825 4.4 ;
      RECT 35.12 3.87 35.135 4.25 ;
      RECT 37.185 3.87 37.19 4.04 ;
      RECT 37.18 3.87 37.185 4.05 ;
      RECT 37.175 3.87 37.18 4.063 ;
      RECT 37.15 3.87 37.175 4.105 ;
      RECT 37.125 3.87 37.15 4.178 ;
      RECT 37.11 3.87 37.125 4.23 ;
      RECT 37.105 3.87 37.11 4.26 ;
      RECT 37.08 3.87 37.105 4.3 ;
      RECT 37.065 3.87 37.08 4.355 ;
      RECT 37.06 3.87 37.065 4.388 ;
      RECT 37.035 3.87 37.06 4.408 ;
      RECT 37.02 3.87 37.035 4.414 ;
      RECT 36.95 3.905 37.015 4.41 ;
      RECT 36.9 3.96 36.95 4.405 ;
      RECT 36.89 3.992 36.9 4.403 ;
      RECT 36.885 4.017 36.89 4.403 ;
      RECT 36.865 4.09 36.885 4.403 ;
      RECT 36.855 4.17 36.865 4.402 ;
      RECT 36.84 4.2 36.855 4.402 ;
      RECT 36.825 4.205 36.84 4.401 ;
      RECT 36.765 4.207 36.82 4.398 ;
      RECT 36.735 4.212 36.765 4.394 ;
      RECT 36.733 4.215 36.735 4.393 ;
      RECT 36.647 4.217 36.733 4.39 ;
      RECT 36.561 4.223 36.647 4.384 ;
      RECT 36.475 4.228 36.561 4.378 ;
      RECT 36.402 4.233 36.475 4.379 ;
      RECT 36.316 4.239 36.402 4.387 ;
      RECT 36.23 4.245 36.316 4.396 ;
      RECT 36.21 4.249 36.23 4.401 ;
      RECT 36.163 4.251 36.21 4.404 ;
      RECT 36.077 4.256 36.163 4.41 ;
      RECT 35.991 4.261 36.077 4.419 ;
      RECT 35.905 4.267 35.991 4.427 ;
      RECT 35.82 4.265 35.905 4.436 ;
      RECT 35.816 4.26 35.82 4.44 ;
      RECT 35.73 4.255 35.816 4.432 ;
      RECT 35.666 4.246 35.73 4.42 ;
      RECT 35.58 4.237 35.666 4.407 ;
      RECT 35.556 4.23 35.58 4.398 ;
      RECT 35.47 4.224 35.556 4.385 ;
      RECT 35.43 4.217 35.47 4.371 ;
      RECT 35.425 4.207 35.43 4.367 ;
      RECT 35.415 4.195 35.425 4.366 ;
      RECT 35.395 4.165 35.415 4.363 ;
      RECT 35.34 4.085 35.395 4.357 ;
      RECT 35.32 4.004 35.34 4.352 ;
      RECT 35.3 3.962 35.32 4.348 ;
      RECT 35.275 3.915 35.3 4.342 ;
      RECT 35.27 3.89 35.275 4.339 ;
      RECT 35.235 3.87 35.27 4.334 ;
      RECT 35.226 3.87 35.235 4.327 ;
      RECT 35.14 3.87 35.226 4.297 ;
      RECT 35.135 3.87 35.14 4.26 ;
      RECT 35.1 3.87 35.12 4.182 ;
      RECT 35.095 3.912 35.1 4.147 ;
      RECT 35.09 3.987 35.095 4.103 ;
      RECT 36.54 3.792 36.715 4.04 ;
      RECT 36.54 3.792 36.72 4.038 ;
      RECT 36.535 3.824 36.72 3.998 ;
      RECT 36.565 3.765 36.735 3.985 ;
      RECT 36.53 3.842 36.735 3.918 ;
      RECT 35.84 3.305 36.01 3.48 ;
      RECT 35.84 3.305 36.182 3.472 ;
      RECT 35.84 3.305 36.265 3.466 ;
      RECT 35.84 3.305 36.3 3.462 ;
      RECT 35.84 3.305 36.32 3.461 ;
      RECT 35.84 3.305 36.406 3.457 ;
      RECT 36.3 3.13 36.47 3.452 ;
      RECT 35.875 3.237 36.5 3.45 ;
      RECT 35.865 3.292 36.505 3.448 ;
      RECT 35.84 3.328 36.515 3.443 ;
      RECT 35.84 3.355 36.52 3.373 ;
      RECT 35.905 3.18 36.48 3.45 ;
      RECT 36.096 3.165 36.48 3.45 ;
      RECT 35.93 3.168 36.48 3.45 ;
      RECT 36.01 3.166 36.096 3.477 ;
      RECT 36.096 3.163 36.475 3.45 ;
      RECT 36.28 3.14 36.475 3.45 ;
      RECT 36.182 3.161 36.475 3.45 ;
      RECT 36.265 3.155 36.28 3.463 ;
      RECT 36.415 4.52 36.42 4.72 ;
      RECT 35.88 4.585 35.925 4.72 ;
      RECT 36.45 4.52 36.47 4.693 ;
      RECT 36.42 4.52 36.45 4.708 ;
      RECT 36.355 4.52 36.415 4.745 ;
      RECT 36.34 4.52 36.355 4.775 ;
      RECT 36.325 4.52 36.34 4.788 ;
      RECT 36.305 4.52 36.325 4.803 ;
      RECT 36.3 4.52 36.305 4.812 ;
      RECT 36.29 4.524 36.3 4.817 ;
      RECT 36.275 4.534 36.29 4.828 ;
      RECT 36.25 4.55 36.275 4.838 ;
      RECT 36.24 4.564 36.25 4.84 ;
      RECT 36.22 4.576 36.24 4.837 ;
      RECT 36.19 4.597 36.22 4.831 ;
      RECT 36.18 4.609 36.19 4.826 ;
      RECT 36.17 4.607 36.18 4.823 ;
      RECT 36.155 4.606 36.17 4.818 ;
      RECT 36.15 4.605 36.155 4.813 ;
      RECT 36.115 4.603 36.15 4.803 ;
      RECT 36.095 4.6 36.115 4.785 ;
      RECT 36.085 4.598 36.095 4.78 ;
      RECT 36.075 4.597 36.085 4.775 ;
      RECT 36.04 4.595 36.075 4.763 ;
      RECT 35.985 4.591 36.04 4.743 ;
      RECT 35.975 4.589 35.985 4.728 ;
      RECT 35.97 4.589 35.975 4.723 ;
      RECT 35.925 4.587 35.97 4.72 ;
      RECT 35.83 4.585 35.88 4.724 ;
      RECT 35.82 4.586 35.83 4.729 ;
      RECT 35.76 4.593 35.82 4.743 ;
      RECT 35.735 4.601 35.76 4.763 ;
      RECT 35.725 4.605 35.735 4.775 ;
      RECT 35.72 4.606 35.725 4.78 ;
      RECT 35.705 4.608 35.72 4.783 ;
      RECT 35.69 4.61 35.705 4.788 ;
      RECT 35.685 4.61 35.69 4.791 ;
      RECT 35.64 4.615 35.685 4.802 ;
      RECT 35.635 4.619 35.64 4.814 ;
      RECT 35.61 4.615 35.635 4.818 ;
      RECT 35.6 4.611 35.61 4.822 ;
      RECT 35.59 4.61 35.6 4.826 ;
      RECT 35.575 4.6 35.59 4.832 ;
      RECT 35.57 4.588 35.575 4.836 ;
      RECT 35.565 4.585 35.57 4.837 ;
      RECT 35.56 4.582 35.565 4.839 ;
      RECT 35.545 4.57 35.56 4.838 ;
      RECT 35.53 4.552 35.545 4.835 ;
      RECT 35.51 4.531 35.53 4.828 ;
      RECT 35.445 4.52 35.51 4.8 ;
      RECT 35.441 4.52 35.445 4.779 ;
      RECT 35.355 4.52 35.441 4.749 ;
      RECT 35.34 4.52 35.355 4.705 ;
      RECT 35.915 3.62 35.92 3.855 ;
      RECT 35.045 3.536 35.05 3.74 ;
      RECT 35.625 3.565 35.63 3.72 ;
      RECT 35.545 3.545 35.55 3.72 ;
      RECT 36.215 3.687 36.23 4.04 ;
      RECT 36.141 3.672 36.215 4.04 ;
      RECT 36.055 3.655 36.141 4.04 ;
      RECT 36.045 3.645 36.055 4.038 ;
      RECT 36.04 3.643 36.045 4.033 ;
      RECT 36.025 3.641 36.04 4.019 ;
      RECT 35.955 3.633 36.025 3.959 ;
      RECT 35.935 3.624 35.955 3.893 ;
      RECT 35.93 3.621 35.935 3.873 ;
      RECT 35.92 3.62 35.93 3.863 ;
      RECT 35.91 3.62 35.915 3.847 ;
      RECT 35.9 3.619 35.91 3.837 ;
      RECT 35.89 3.617 35.9 3.825 ;
      RECT 35.875 3.614 35.89 3.805 ;
      RECT 35.865 3.612 35.875 3.79 ;
      RECT 35.845 3.609 35.865 3.778 ;
      RECT 35.84 3.607 35.845 3.768 ;
      RECT 35.815 3.605 35.84 3.755 ;
      RECT 35.785 3.6 35.815 3.74 ;
      RECT 35.705 3.591 35.785 3.731 ;
      RECT 35.66 3.58 35.705 3.724 ;
      RECT 35.64 3.571 35.66 3.721 ;
      RECT 35.63 3.566 35.64 3.72 ;
      RECT 35.585 3.56 35.625 3.72 ;
      RECT 35.57 3.552 35.585 3.72 ;
      RECT 35.55 3.547 35.57 3.72 ;
      RECT 35.53 3.544 35.545 3.72 ;
      RECT 35.447 3.543 35.53 3.719 ;
      RECT 35.361 3.542 35.447 3.715 ;
      RECT 35.275 3.54 35.361 3.712 ;
      RECT 35.222 3.539 35.275 3.714 ;
      RECT 35.136 3.538 35.222 3.723 ;
      RECT 35.05 3.537 35.136 3.735 ;
      RECT 35.03 3.536 35.045 3.743 ;
      RECT 34.95 3.535 35.03 3.755 ;
      RECT 34.925 3.535 34.95 3.768 ;
      RECT 34.9 3.535 34.925 3.783 ;
      RECT 34.895 3.535 34.9 3.805 ;
      RECT 34.89 3.535 34.895 3.823 ;
      RECT 34.885 3.535 34.89 3.84 ;
      RECT 34.88 3.535 34.885 3.853 ;
      RECT 34.875 3.535 34.88 3.863 ;
      RECT 34.835 3.535 34.875 3.948 ;
      RECT 34.82 3.535 34.835 4.033 ;
      RECT 34.81 3.536 34.82 4.045 ;
      RECT 34.775 3.541 34.81 4.05 ;
      RECT 34.735 3.55 34.775 4.05 ;
      RECT 34.72 3.56 34.735 4.05 ;
      RECT 34.715 3.57 34.72 4.05 ;
      RECT 34.695 3.597 34.715 4.05 ;
      RECT 34.645 3.68 34.695 4.05 ;
      RECT 34.64 3.742 34.645 4.05 ;
      RECT 34.63 3.755 34.64 4.05 ;
      RECT 34.62 3.777 34.63 4.05 ;
      RECT 34.61 3.802 34.62 4.045 ;
      RECT 34.605 3.84 34.61 4.038 ;
      RECT 34.595 3.95 34.605 4.033 ;
      RECT 35.99 4.871 36.005 5.13 ;
      RECT 35.99 4.886 36.01 5.129 ;
      RECT 35.906 4.886 36.01 5.127 ;
      RECT 35.906 4.9 36.015 5.126 ;
      RECT 35.82 4.942 36.02 5.123 ;
      RECT 35.815 4.885 36.005 5.118 ;
      RECT 35.815 4.956 36.025 5.115 ;
      RECT 35.81 4.987 36.025 5.113 ;
      RECT 35.815 4.984 36.04 5.103 ;
      RECT 35.81 5.03 36.055 5.088 ;
      RECT 35.81 5.058 36.06 5.073 ;
      RECT 35.82 4.86 35.99 5.123 ;
      RECT 35.58 3.87 35.75 4.04 ;
      RECT 35.545 3.87 35.75 4.035 ;
      RECT 35.535 3.87 35.75 4.028 ;
      RECT 35.53 3.855 35.7 4.025 ;
      RECT 34.36 4.392 34.625 4.835 ;
      RECT 34.355 4.363 34.57 4.833 ;
      RECT 34.35 4.517 34.63 4.828 ;
      RECT 34.355 4.412 34.63 4.828 ;
      RECT 34.355 4.423 34.64 4.815 ;
      RECT 34.355 4.37 34.6 4.833 ;
      RECT 34.36 4.357 34.57 4.835 ;
      RECT 34.36 4.355 34.52 4.835 ;
      RECT 34.461 4.347 34.52 4.835 ;
      RECT 34.375 4.348 34.52 4.835 ;
      RECT 34.461 4.346 34.51 4.835 ;
      RECT 34.265 3.161 34.44 3.46 ;
      RECT 34.315 3.123 34.44 3.46 ;
      RECT 34.3 3.125 34.526 3.452 ;
      RECT 34.3 3.128 34.565 3.439 ;
      RECT 34.3 3.129 34.575 3.425 ;
      RECT 34.255 3.18 34.575 3.415 ;
      RECT 34.3 3.13 34.58 3.41 ;
      RECT 34.255 3.34 34.585 3.4 ;
      RECT 34.24 3.2 34.58 3.34 ;
      RECT 34.235 3.216 34.58 3.28 ;
      RECT 34.28 3.14 34.58 3.41 ;
      RECT 34.315 3.121 34.401 3.46 ;
      RECT 32.405 3.035 32.575 4.225 ;
      RECT 32.405 3.035 32.875 3.205 ;
      RECT 32.405 9.26 32.875 9.43 ;
      RECT 32.405 8.24 32.575 9.43 ;
      RECT 31.415 3.035 31.585 4.225 ;
      RECT 31.415 3.035 31.885 3.205 ;
      RECT 31.415 9.26 31.885 9.43 ;
      RECT 31.415 8.24 31.585 9.43 ;
      RECT 29.565 3.93 29.735 5.16 ;
      RECT 29.62 2.15 29.79 4.1 ;
      RECT 29.565 1.87 29.735 2.32 ;
      RECT 29.565 10.145 29.735 10.595 ;
      RECT 29.62 8.365 29.79 10.315 ;
      RECT 29.565 7.305 29.735 8.535 ;
      RECT 29.045 1.87 29.215 5.16 ;
      RECT 29.045 3.37 29.45 3.7 ;
      RECT 29.045 2.53 29.45 2.86 ;
      RECT 29.045 7.305 29.215 10.595 ;
      RECT 29.045 9.605 29.45 9.935 ;
      RECT 29.045 8.765 29.45 9.095 ;
      RECT 26.97 4.421 26.975 4.593 ;
      RECT 26.965 4.414 26.97 4.683 ;
      RECT 26.96 4.408 26.965 4.702 ;
      RECT 26.94 4.402 26.96 4.712 ;
      RECT 26.925 4.397 26.94 4.72 ;
      RECT 26.888 4.391 26.925 4.718 ;
      RECT 26.802 4.377 26.888 4.714 ;
      RECT 26.716 4.359 26.802 4.709 ;
      RECT 26.63 4.34 26.716 4.703 ;
      RECT 26.6 4.328 26.63 4.699 ;
      RECT 26.58 4.322 26.6 4.698 ;
      RECT 26.515 4.32 26.58 4.696 ;
      RECT 26.5 4.32 26.515 4.688 ;
      RECT 26.485 4.32 26.5 4.675 ;
      RECT 26.48 4.32 26.485 4.665 ;
      RECT 26.465 4.32 26.48 4.643 ;
      RECT 26.45 4.32 26.465 4.61 ;
      RECT 26.445 4.32 26.45 4.588 ;
      RECT 26.435 4.32 26.445 4.57 ;
      RECT 26.42 4.32 26.435 4.548 ;
      RECT 26.4 4.32 26.42 4.51 ;
      RECT 26.75 3.605 26.785 4.044 ;
      RECT 26.75 3.605 26.79 4.043 ;
      RECT 26.695 3.665 26.79 4.042 ;
      RECT 26.56 3.837 26.79 4.041 ;
      RECT 26.67 3.715 26.79 4.041 ;
      RECT 26.56 3.837 26.815 4.031 ;
      RECT 26.615 3.782 26.895 3.948 ;
      RECT 26.79 3.576 26.795 4.039 ;
      RECT 26.645 3.752 26.935 3.825 ;
      RECT 26.66 3.735 26.79 4.041 ;
      RECT 26.795 3.575 26.965 3.763 ;
      RECT 26.785 3.578 26.965 3.763 ;
      RECT 26.29 3.455 26.46 3.765 ;
      RECT 26.29 3.455 26.465 3.738 ;
      RECT 26.29 3.455 26.47 3.715 ;
      RECT 26.29 3.455 26.48 3.665 ;
      RECT 26.285 3.56 26.48 3.635 ;
      RECT 26.32 3.13 26.49 3.608 ;
      RECT 26.32 3.13 26.505 3.529 ;
      RECT 26.31 3.34 26.505 3.529 ;
      RECT 26.32 3.14 26.515 3.444 ;
      RECT 26.25 3.882 26.255 4.085 ;
      RECT 26.24 3.87 26.25 4.195 ;
      RECT 26.215 3.87 26.24 4.235 ;
      RECT 26.135 3.87 26.215 4.32 ;
      RECT 26.125 3.87 26.135 4.39 ;
      RECT 26.1 3.87 26.125 4.413 ;
      RECT 26.08 3.87 26.1 4.448 ;
      RECT 26.035 3.88 26.08 4.491 ;
      RECT 26.025 3.892 26.035 4.528 ;
      RECT 26.005 3.906 26.025 4.548 ;
      RECT 25.995 3.924 26.005 4.564 ;
      RECT 25.98 3.95 25.995 4.574 ;
      RECT 25.965 3.991 25.98 4.588 ;
      RECT 25.955 4.026 25.965 4.598 ;
      RECT 25.95 4.042 25.955 4.603 ;
      RECT 25.94 4.057 25.95 4.608 ;
      RECT 25.92 4.1 25.94 4.618 ;
      RECT 25.9 4.137 25.92 4.631 ;
      RECT 25.865 4.16 25.9 4.649 ;
      RECT 25.855 4.174 25.865 4.665 ;
      RECT 25.835 4.184 25.855 4.675 ;
      RECT 25.83 4.193 25.835 4.683 ;
      RECT 25.82 4.2 25.83 4.69 ;
      RECT 25.81 4.207 25.82 4.698 ;
      RECT 25.795 4.217 25.81 4.706 ;
      RECT 25.785 4.231 25.795 4.716 ;
      RECT 25.775 4.243 25.785 4.728 ;
      RECT 25.76 4.265 25.775 4.741 ;
      RECT 25.75 4.287 25.76 4.752 ;
      RECT 25.74 4.307 25.75 4.761 ;
      RECT 25.735 4.322 25.74 4.768 ;
      RECT 25.705 4.355 25.735 4.782 ;
      RECT 25.695 4.39 25.705 4.797 ;
      RECT 25.69 4.397 25.695 4.803 ;
      RECT 25.67 4.412 25.69 4.81 ;
      RECT 25.665 4.427 25.67 4.818 ;
      RECT 25.66 4.436 25.665 4.823 ;
      RECT 25.645 4.442 25.66 4.83 ;
      RECT 25.64 4.448 25.645 4.838 ;
      RECT 25.635 4.452 25.64 4.845 ;
      RECT 25.63 4.456 25.635 4.855 ;
      RECT 25.62 4.461 25.63 4.865 ;
      RECT 25.6 4.472 25.62 4.893 ;
      RECT 25.585 4.484 25.6 4.92 ;
      RECT 25.565 4.497 25.585 4.945 ;
      RECT 25.545 4.512 25.565 4.969 ;
      RECT 25.53 4.527 25.545 4.984 ;
      RECT 25.525 4.538 25.53 4.993 ;
      RECT 25.46 4.583 25.525 5.003 ;
      RECT 25.425 4.642 25.46 5.016 ;
      RECT 25.42 4.665 25.425 5.022 ;
      RECT 25.415 4.672 25.42 5.024 ;
      RECT 25.4 4.682 25.415 5.027 ;
      RECT 25.37 4.707 25.4 5.031 ;
      RECT 25.365 4.725 25.37 5.035 ;
      RECT 25.36 4.732 25.365 5.036 ;
      RECT 25.34 4.74 25.36 5.04 ;
      RECT 25.33 4.747 25.34 5.044 ;
      RECT 25.286 4.758 25.33 5.051 ;
      RECT 25.2 4.786 25.286 5.067 ;
      RECT 25.14 4.81 25.2 5.085 ;
      RECT 25.095 4.82 25.14 5.099 ;
      RECT 25.036 4.828 25.095 5.113 ;
      RECT 24.95 4.835 25.036 5.132 ;
      RECT 24.925 4.84 24.95 5.147 ;
      RECT 24.845 4.843 24.925 5.15 ;
      RECT 24.765 4.847 24.845 5.137 ;
      RECT 24.756 4.85 24.765 5.122 ;
      RECT 24.67 4.85 24.756 5.107 ;
      RECT 24.61 4.852 24.67 5.084 ;
      RECT 24.606 4.855 24.61 5.074 ;
      RECT 24.52 4.855 24.606 5.059 ;
      RECT 24.445 4.855 24.52 5.035 ;
      RECT 25.76 3.864 25.77 4.04 ;
      RECT 25.715 3.831 25.76 4.04 ;
      RECT 25.67 3.782 25.715 4.04 ;
      RECT 25.64 3.752 25.67 4.041 ;
      RECT 25.635 3.735 25.64 4.042 ;
      RECT 25.61 3.715 25.635 4.043 ;
      RECT 25.595 3.69 25.61 4.044 ;
      RECT 25.59 3.677 25.595 4.045 ;
      RECT 25.585 3.671 25.59 4.043 ;
      RECT 25.58 3.663 25.585 4.037 ;
      RECT 25.555 3.655 25.58 4.017 ;
      RECT 25.535 3.644 25.555 3.988 ;
      RECT 25.505 3.629 25.535 3.959 ;
      RECT 25.485 3.615 25.505 3.931 ;
      RECT 25.475 3.609 25.485 3.91 ;
      RECT 25.47 3.606 25.475 3.893 ;
      RECT 25.465 3.603 25.47 3.878 ;
      RECT 25.45 3.598 25.465 3.843 ;
      RECT 25.445 3.594 25.45 3.81 ;
      RECT 25.425 3.589 25.445 3.786 ;
      RECT 25.395 3.581 25.425 3.751 ;
      RECT 25.38 3.575 25.395 3.728 ;
      RECT 25.34 3.568 25.38 3.713 ;
      RECT 25.315 3.56 25.34 3.693 ;
      RECT 25.295 3.555 25.315 3.683 ;
      RECT 25.26 3.549 25.295 3.678 ;
      RECT 25.215 3.54 25.26 3.677 ;
      RECT 25.185 3.536 25.215 3.679 ;
      RECT 25.1 3.544 25.185 3.683 ;
      RECT 25.03 3.555 25.1 3.705 ;
      RECT 25.017 3.561 25.03 3.728 ;
      RECT 24.931 3.568 25.017 3.75 ;
      RECT 24.845 3.58 24.931 3.787 ;
      RECT 24.845 3.957 24.855 4.195 ;
      RECT 24.84 3.586 24.845 3.81 ;
      RECT 24.835 3.842 24.845 4.195 ;
      RECT 24.835 3.587 24.84 3.815 ;
      RECT 24.83 3.588 24.835 4.195 ;
      RECT 24.806 3.59 24.83 4.196 ;
      RECT 24.72 3.598 24.806 4.198 ;
      RECT 24.7 3.612 24.72 4.201 ;
      RECT 24.695 3.64 24.7 4.202 ;
      RECT 24.69 3.652 24.695 4.203 ;
      RECT 24.685 3.667 24.69 4.204 ;
      RECT 24.675 3.697 24.685 4.205 ;
      RECT 24.67 3.735 24.675 4.203 ;
      RECT 24.665 3.755 24.67 4.198 ;
      RECT 24.65 3.79 24.665 4.183 ;
      RECT 24.64 3.842 24.65 4.163 ;
      RECT 24.635 3.872 24.64 4.151 ;
      RECT 24.62 3.885 24.635 4.134 ;
      RECT 24.595 3.889 24.62 4.101 ;
      RECT 24.58 3.887 24.595 4.078 ;
      RECT 24.565 3.886 24.58 4.075 ;
      RECT 24.505 3.884 24.565 4.073 ;
      RECT 24.495 3.882 24.505 4.068 ;
      RECT 24.455 3.881 24.495 4.065 ;
      RECT 24.385 3.878 24.455 4.063 ;
      RECT 24.33 3.876 24.385 4.058 ;
      RECT 24.26 3.87 24.33 4.053 ;
      RECT 24.251 3.87 24.26 4.05 ;
      RECT 24.165 3.87 24.251 4.045 ;
      RECT 24.16 3.87 24.165 4.04 ;
      RECT 25.465 3.105 25.64 3.455 ;
      RECT 25.465 3.12 25.65 3.453 ;
      RECT 25.44 3.07 25.585 3.45 ;
      RECT 25.42 3.071 25.585 3.443 ;
      RECT 25.41 3.072 25.595 3.438 ;
      RECT 25.38 3.073 25.595 3.425 ;
      RECT 25.33 3.074 25.595 3.401 ;
      RECT 25.325 3.076 25.595 3.386 ;
      RECT 25.325 3.142 25.655 3.38 ;
      RECT 25.305 3.083 25.61 3.36 ;
      RECT 25.295 3.092 25.62 3.215 ;
      RECT 25.305 3.087 25.62 3.36 ;
      RECT 25.325 3.077 25.61 3.386 ;
      RECT 24.91 4.402 25.08 4.69 ;
      RECT 24.905 4.42 25.09 4.685 ;
      RECT 24.87 4.428 25.155 4.605 ;
      RECT 24.87 4.428 25.241 4.595 ;
      RECT 24.87 4.428 25.295 4.541 ;
      RECT 25.155 4.325 25.325 4.509 ;
      RECT 24.87 4.48 25.33 4.497 ;
      RECT 24.855 4.45 25.325 4.493 ;
      RECT 25.115 4.332 25.155 4.644 ;
      RECT 24.995 4.369 25.325 4.509 ;
      RECT 25.09 4.344 25.115 4.67 ;
      RECT 25.08 4.351 25.325 4.509 ;
      RECT 25.211 3.815 25.28 4.074 ;
      RECT 25.211 3.87 25.285 4.073 ;
      RECT 25.125 3.87 25.285 4.072 ;
      RECT 25.12 3.87 25.29 4.065 ;
      RECT 25.11 3.815 25.28 4.06 ;
      RECT 24.49 3.114 24.665 3.415 ;
      RECT 24.475 3.102 24.49 3.4 ;
      RECT 24.445 3.101 24.475 3.353 ;
      RECT 24.445 3.119 24.67 3.348 ;
      RECT 24.43 3.103 24.49 3.313 ;
      RECT 24.425 3.125 24.68 3.213 ;
      RECT 24.425 3.108 24.576 3.213 ;
      RECT 24.425 3.11 24.58 3.213 ;
      RECT 24.43 3.106 24.576 3.313 ;
      RECT 24.535 4.342 24.54 4.69 ;
      RECT 24.525 4.332 24.535 4.696 ;
      RECT 24.49 4.322 24.525 4.698 ;
      RECT 24.452 4.317 24.49 4.702 ;
      RECT 24.366 4.31 24.452 4.709 ;
      RECT 24.28 4.3 24.366 4.719 ;
      RECT 24.235 4.295 24.28 4.727 ;
      RECT 24.231 4.295 24.235 4.731 ;
      RECT 24.145 4.295 24.231 4.738 ;
      RECT 24.13 4.295 24.145 4.738 ;
      RECT 24.12 4.293 24.13 4.71 ;
      RECT 24.11 4.289 24.12 4.653 ;
      RECT 24.09 4.283 24.11 4.585 ;
      RECT 24.085 4.279 24.09 4.533 ;
      RECT 24.075 4.278 24.085 4.5 ;
      RECT 24.025 4.276 24.075 4.485 ;
      RECT 24 4.274 24.025 4.48 ;
      RECT 23.957 4.272 24 4.476 ;
      RECT 23.871 4.268 23.957 4.464 ;
      RECT 23.785 4.263 23.871 4.448 ;
      RECT 23.755 4.26 23.785 4.435 ;
      RECT 23.73 4.259 23.755 4.423 ;
      RECT 23.725 4.259 23.73 4.413 ;
      RECT 23.685 4.258 23.725 4.405 ;
      RECT 23.67 4.257 23.685 4.398 ;
      RECT 23.62 4.256 23.67 4.39 ;
      RECT 23.618 4.255 23.62 4.385 ;
      RECT 23.532 4.253 23.618 4.385 ;
      RECT 23.446 4.248 23.532 4.385 ;
      RECT 23.36 4.244 23.446 4.385 ;
      RECT 23.311 4.24 23.36 4.383 ;
      RECT 23.225 4.237 23.311 4.378 ;
      RECT 23.202 4.234 23.225 4.374 ;
      RECT 23.116 4.231 23.202 4.369 ;
      RECT 23.03 4.227 23.116 4.36 ;
      RECT 23.005 4.22 23.03 4.355 ;
      RECT 22.945 4.185 23.005 4.352 ;
      RECT 22.925 4.11 22.945 4.349 ;
      RECT 22.92 4.052 22.925 4.348 ;
      RECT 22.895 3.992 22.92 4.347 ;
      RECT 22.82 3.87 22.895 4.343 ;
      RECT 22.81 3.87 22.82 4.335 ;
      RECT 22.795 3.87 22.81 4.325 ;
      RECT 22.78 3.87 22.795 4.295 ;
      RECT 22.765 3.87 22.78 4.24 ;
      RECT 22.75 3.87 22.765 4.178 ;
      RECT 22.725 3.87 22.75 4.103 ;
      RECT 22.72 3.87 22.725 4.053 ;
      RECT 24.065 3.415 24.085 3.724 ;
      RECT 24.051 3.417 24.1 3.721 ;
      RECT 24.051 3.422 24.12 3.712 ;
      RECT 23.965 3.42 24.1 3.706 ;
      RECT 23.965 3.428 24.155 3.689 ;
      RECT 23.93 3.43 24.155 3.688 ;
      RECT 23.9 3.438 24.155 3.679 ;
      RECT 23.89 3.443 24.175 3.665 ;
      RECT 23.93 3.433 24.175 3.665 ;
      RECT 23.93 3.436 24.185 3.653 ;
      RECT 23.9 3.438 24.195 3.64 ;
      RECT 23.9 3.442 24.205 3.583 ;
      RECT 23.89 3.447 24.21 3.498 ;
      RECT 24.051 3.415 24.085 3.721 ;
      RECT 23.93 10.145 24.1 10.595 ;
      RECT 23.985 8.365 24.155 10.315 ;
      RECT 23.93 7.305 24.1 8.535 ;
      RECT 23.49 3.518 23.495 3.73 ;
      RECT 23.365 3.515 23.38 3.73 ;
      RECT 22.83 3.545 22.9 3.73 ;
      RECT 22.715 3.545 22.75 3.725 ;
      RECT 23.836 3.847 23.855 4.041 ;
      RECT 23.75 3.802 23.836 4.042 ;
      RECT 23.74 3.755 23.75 4.044 ;
      RECT 23.735 3.735 23.74 4.045 ;
      RECT 23.715 3.7 23.735 4.046 ;
      RECT 23.7 3.65 23.715 4.047 ;
      RECT 23.68 3.587 23.7 4.048 ;
      RECT 23.67 3.55 23.68 4.049 ;
      RECT 23.655 3.539 23.67 4.05 ;
      RECT 23.65 3.531 23.655 4.048 ;
      RECT 23.64 3.53 23.65 4.04 ;
      RECT 23.61 3.527 23.64 4.019 ;
      RECT 23.535 3.522 23.61 3.964 ;
      RECT 23.52 3.518 23.535 3.91 ;
      RECT 23.51 3.518 23.52 3.805 ;
      RECT 23.495 3.518 23.51 3.738 ;
      RECT 23.48 3.518 23.49 3.728 ;
      RECT 23.425 3.517 23.48 3.725 ;
      RECT 23.38 3.515 23.425 3.728 ;
      RECT 23.352 3.515 23.365 3.731 ;
      RECT 23.266 3.519 23.352 3.733 ;
      RECT 23.18 3.525 23.266 3.738 ;
      RECT 23.16 3.529 23.18 3.74 ;
      RECT 23.158 3.53 23.16 3.739 ;
      RECT 23.072 3.532 23.158 3.738 ;
      RECT 22.986 3.537 23.072 3.735 ;
      RECT 22.9 3.542 22.986 3.732 ;
      RECT 22.75 3.545 22.83 3.728 ;
      RECT 23.41 7.305 23.58 10.595 ;
      RECT 23.41 9.605 23.815 9.935 ;
      RECT 23.41 8.765 23.815 9.095 ;
      RECT 23.526 4.52 23.575 4.854 ;
      RECT 23.526 4.52 23.58 4.853 ;
      RECT 23.44 4.52 23.58 4.852 ;
      RECT 23.215 4.628 23.585 4.85 ;
      RECT 23.44 4.52 23.61 4.843 ;
      RECT 23.41 4.532 23.615 4.834 ;
      RECT 23.395 4.55 23.62 4.831 ;
      RECT 23.21 4.634 23.62 4.758 ;
      RECT 23.205 4.641 23.62 4.718 ;
      RECT 23.22 4.607 23.62 4.831 ;
      RECT 23.381 4.553 23.585 4.85 ;
      RECT 23.295 4.573 23.62 4.831 ;
      RECT 23.395 4.547 23.615 4.834 ;
      RECT 23.165 3.871 23.355 4.065 ;
      RECT 23.16 3.873 23.355 4.064 ;
      RECT 23.155 3.877 23.37 4.061 ;
      RECT 23.17 3.87 23.37 4.061 ;
      RECT 23.155 3.98 23.375 4.056 ;
      RECT 22.45 4.48 22.541 4.778 ;
      RECT 22.445 4.482 22.62 4.773 ;
      RECT 22.45 4.48 22.62 4.773 ;
      RECT 22.445 4.486 22.64 4.771 ;
      RECT 22.445 4.541 22.68 4.77 ;
      RECT 22.445 4.576 22.695 4.764 ;
      RECT 22.445 4.61 22.705 4.754 ;
      RECT 22.435 4.49 22.64 4.605 ;
      RECT 22.435 4.51 22.655 4.605 ;
      RECT 22.435 4.493 22.645 4.605 ;
      RECT 22.66 3.261 22.665 3.323 ;
      RECT 22.655 3.183 22.66 3.346 ;
      RECT 22.65 3.14 22.655 3.357 ;
      RECT 22.645 3.13 22.65 3.369 ;
      RECT 22.64 3.13 22.645 3.378 ;
      RECT 22.615 3.13 22.64 3.41 ;
      RECT 22.61 3.13 22.615 3.443 ;
      RECT 22.595 3.13 22.61 3.468 ;
      RECT 22.585 3.13 22.595 3.495 ;
      RECT 22.58 3.13 22.585 3.508 ;
      RECT 22.575 3.13 22.58 3.523 ;
      RECT 22.565 3.13 22.575 3.538 ;
      RECT 22.56 3.13 22.565 3.558 ;
      RECT 22.535 3.13 22.56 3.593 ;
      RECT 22.49 3.13 22.535 3.638 ;
      RECT 22.48 3.13 22.49 3.651 ;
      RECT 22.395 3.215 22.48 3.658 ;
      RECT 22.36 3.337 22.395 3.667 ;
      RECT 22.355 3.377 22.36 3.671 ;
      RECT 22.335 3.4 22.355 3.673 ;
      RECT 22.33 3.43 22.335 3.676 ;
      RECT 22.32 3.442 22.33 3.677 ;
      RECT 22.275 3.465 22.32 3.682 ;
      RECT 22.235 3.495 22.275 3.69 ;
      RECT 22.2 3.507 22.235 3.696 ;
      RECT 22.195 3.512 22.2 3.7 ;
      RECT 22.125 3.522 22.195 3.707 ;
      RECT 22.085 3.532 22.125 3.717 ;
      RECT 22.065 3.537 22.085 3.723 ;
      RECT 22.055 3.541 22.065 3.728 ;
      RECT 22.05 3.544 22.055 3.731 ;
      RECT 22.04 3.545 22.05 3.732 ;
      RECT 22.015 3.547 22.04 3.736 ;
      RECT 22.005 3.552 22.015 3.739 ;
      RECT 21.96 3.56 22.005 3.74 ;
      RECT 21.835 3.565 21.96 3.74 ;
      RECT 22.39 3.862 22.41 4.044 ;
      RECT 22.341 3.847 22.39 4.043 ;
      RECT 22.255 3.862 22.41 4.041 ;
      RECT 22.24 3.862 22.41 4.04 ;
      RECT 22.205 3.84 22.375 4.025 ;
      RECT 22.275 4.86 22.29 5.069 ;
      RECT 22.275 4.868 22.295 5.068 ;
      RECT 22.22 4.868 22.295 5.067 ;
      RECT 22.2 4.872 22.3 5.065 ;
      RECT 22.18 4.822 22.22 5.064 ;
      RECT 22.125 4.88 22.305 5.062 ;
      RECT 22.09 4.837 22.22 5.06 ;
      RECT 22.086 4.84 22.275 5.059 ;
      RECT 22 4.848 22.275 5.057 ;
      RECT 22 4.892 22.31 5.05 ;
      RECT 21.99 4.985 22.31 5.048 ;
      RECT 22 4.904 22.315 5.033 ;
      RECT 22 4.925 22.33 5.003 ;
      RECT 22 4.952 22.335 4.973 ;
      RECT 22.125 4.83 22.22 5.062 ;
      RECT 21.755 3.875 21.76 4.413 ;
      RECT 21.56 4.205 21.565 4.4 ;
      RECT 19.86 3.87 19.875 4.25 ;
      RECT 21.925 3.87 21.93 4.04 ;
      RECT 21.92 3.87 21.925 4.05 ;
      RECT 21.915 3.87 21.92 4.063 ;
      RECT 21.89 3.87 21.915 4.105 ;
      RECT 21.865 3.87 21.89 4.178 ;
      RECT 21.85 3.87 21.865 4.23 ;
      RECT 21.845 3.87 21.85 4.26 ;
      RECT 21.82 3.87 21.845 4.3 ;
      RECT 21.805 3.87 21.82 4.355 ;
      RECT 21.8 3.87 21.805 4.388 ;
      RECT 21.775 3.87 21.8 4.408 ;
      RECT 21.76 3.87 21.775 4.414 ;
      RECT 21.69 3.905 21.755 4.41 ;
      RECT 21.64 3.96 21.69 4.405 ;
      RECT 21.63 3.992 21.64 4.403 ;
      RECT 21.625 4.017 21.63 4.403 ;
      RECT 21.605 4.09 21.625 4.403 ;
      RECT 21.595 4.17 21.605 4.402 ;
      RECT 21.58 4.2 21.595 4.402 ;
      RECT 21.565 4.205 21.58 4.401 ;
      RECT 21.505 4.207 21.56 4.398 ;
      RECT 21.475 4.212 21.505 4.394 ;
      RECT 21.473 4.215 21.475 4.393 ;
      RECT 21.387 4.217 21.473 4.39 ;
      RECT 21.301 4.223 21.387 4.384 ;
      RECT 21.215 4.228 21.301 4.378 ;
      RECT 21.142 4.233 21.215 4.379 ;
      RECT 21.056 4.239 21.142 4.387 ;
      RECT 20.97 4.245 21.056 4.396 ;
      RECT 20.95 4.249 20.97 4.401 ;
      RECT 20.903 4.251 20.95 4.404 ;
      RECT 20.817 4.256 20.903 4.41 ;
      RECT 20.731 4.261 20.817 4.419 ;
      RECT 20.645 4.267 20.731 4.427 ;
      RECT 20.56 4.265 20.645 4.436 ;
      RECT 20.556 4.26 20.56 4.44 ;
      RECT 20.47 4.255 20.556 4.432 ;
      RECT 20.406 4.246 20.47 4.42 ;
      RECT 20.32 4.237 20.406 4.407 ;
      RECT 20.296 4.23 20.32 4.398 ;
      RECT 20.21 4.224 20.296 4.385 ;
      RECT 20.17 4.217 20.21 4.371 ;
      RECT 20.165 4.207 20.17 4.367 ;
      RECT 20.155 4.195 20.165 4.366 ;
      RECT 20.135 4.165 20.155 4.363 ;
      RECT 20.08 4.085 20.135 4.357 ;
      RECT 20.06 4.004 20.08 4.352 ;
      RECT 20.04 3.962 20.06 4.348 ;
      RECT 20.015 3.915 20.04 4.342 ;
      RECT 20.01 3.89 20.015 4.339 ;
      RECT 19.975 3.87 20.01 4.334 ;
      RECT 19.966 3.87 19.975 4.327 ;
      RECT 19.88 3.87 19.966 4.297 ;
      RECT 19.875 3.87 19.88 4.26 ;
      RECT 19.84 3.87 19.86 4.182 ;
      RECT 19.835 3.912 19.84 4.147 ;
      RECT 19.83 3.987 19.835 4.103 ;
      RECT 21.28 3.792 21.455 4.04 ;
      RECT 21.28 3.792 21.46 4.038 ;
      RECT 21.275 3.824 21.46 3.998 ;
      RECT 21.305 3.765 21.475 3.985 ;
      RECT 21.27 3.842 21.475 3.918 ;
      RECT 20.58 3.305 20.75 3.48 ;
      RECT 20.58 3.305 20.922 3.472 ;
      RECT 20.58 3.305 21.005 3.466 ;
      RECT 20.58 3.305 21.04 3.462 ;
      RECT 20.58 3.305 21.06 3.461 ;
      RECT 20.58 3.305 21.146 3.457 ;
      RECT 21.04 3.13 21.21 3.452 ;
      RECT 20.615 3.237 21.24 3.45 ;
      RECT 20.605 3.292 21.245 3.448 ;
      RECT 20.58 3.328 21.255 3.443 ;
      RECT 20.58 3.355 21.26 3.373 ;
      RECT 20.645 3.18 21.22 3.45 ;
      RECT 20.836 3.165 21.22 3.45 ;
      RECT 20.67 3.168 21.22 3.45 ;
      RECT 20.75 3.166 20.836 3.477 ;
      RECT 20.836 3.163 21.215 3.45 ;
      RECT 21.02 3.14 21.215 3.45 ;
      RECT 20.922 3.161 21.215 3.45 ;
      RECT 21.005 3.155 21.02 3.463 ;
      RECT 21.155 4.52 21.16 4.72 ;
      RECT 20.62 4.585 20.665 4.72 ;
      RECT 21.19 4.52 21.21 4.693 ;
      RECT 21.16 4.52 21.19 4.708 ;
      RECT 21.095 4.52 21.155 4.745 ;
      RECT 21.08 4.52 21.095 4.775 ;
      RECT 21.065 4.52 21.08 4.788 ;
      RECT 21.045 4.52 21.065 4.803 ;
      RECT 21.04 4.52 21.045 4.812 ;
      RECT 21.03 4.524 21.04 4.817 ;
      RECT 21.015 4.534 21.03 4.828 ;
      RECT 20.99 4.55 21.015 4.838 ;
      RECT 20.98 4.564 20.99 4.84 ;
      RECT 20.96 4.576 20.98 4.837 ;
      RECT 20.93 4.597 20.96 4.831 ;
      RECT 20.92 4.609 20.93 4.826 ;
      RECT 20.91 4.607 20.92 4.823 ;
      RECT 20.895 4.606 20.91 4.818 ;
      RECT 20.89 4.605 20.895 4.813 ;
      RECT 20.855 4.603 20.89 4.803 ;
      RECT 20.835 4.6 20.855 4.785 ;
      RECT 20.825 4.598 20.835 4.78 ;
      RECT 20.815 4.597 20.825 4.775 ;
      RECT 20.78 4.595 20.815 4.763 ;
      RECT 20.725 4.591 20.78 4.743 ;
      RECT 20.715 4.589 20.725 4.728 ;
      RECT 20.71 4.589 20.715 4.723 ;
      RECT 20.665 4.587 20.71 4.72 ;
      RECT 20.57 4.585 20.62 4.724 ;
      RECT 20.56 4.586 20.57 4.729 ;
      RECT 20.5 4.593 20.56 4.743 ;
      RECT 20.475 4.601 20.5 4.763 ;
      RECT 20.465 4.605 20.475 4.775 ;
      RECT 20.46 4.606 20.465 4.78 ;
      RECT 20.445 4.608 20.46 4.783 ;
      RECT 20.43 4.61 20.445 4.788 ;
      RECT 20.425 4.61 20.43 4.791 ;
      RECT 20.38 4.615 20.425 4.802 ;
      RECT 20.375 4.619 20.38 4.814 ;
      RECT 20.35 4.615 20.375 4.818 ;
      RECT 20.34 4.611 20.35 4.822 ;
      RECT 20.33 4.61 20.34 4.826 ;
      RECT 20.315 4.6 20.33 4.832 ;
      RECT 20.31 4.588 20.315 4.836 ;
      RECT 20.305 4.585 20.31 4.837 ;
      RECT 20.3 4.582 20.305 4.839 ;
      RECT 20.285 4.57 20.3 4.838 ;
      RECT 20.27 4.552 20.285 4.835 ;
      RECT 20.25 4.531 20.27 4.828 ;
      RECT 20.185 4.52 20.25 4.8 ;
      RECT 20.181 4.52 20.185 4.779 ;
      RECT 20.095 4.52 20.181 4.749 ;
      RECT 20.08 4.52 20.095 4.705 ;
      RECT 20.655 3.62 20.66 3.855 ;
      RECT 19.785 3.536 19.79 3.74 ;
      RECT 20.365 3.565 20.37 3.72 ;
      RECT 20.285 3.545 20.29 3.72 ;
      RECT 20.955 3.687 20.97 4.04 ;
      RECT 20.881 3.672 20.955 4.04 ;
      RECT 20.795 3.655 20.881 4.04 ;
      RECT 20.785 3.645 20.795 4.038 ;
      RECT 20.78 3.643 20.785 4.033 ;
      RECT 20.765 3.641 20.78 4.019 ;
      RECT 20.695 3.633 20.765 3.959 ;
      RECT 20.675 3.624 20.695 3.893 ;
      RECT 20.67 3.621 20.675 3.873 ;
      RECT 20.66 3.62 20.67 3.863 ;
      RECT 20.65 3.62 20.655 3.847 ;
      RECT 20.64 3.619 20.65 3.837 ;
      RECT 20.63 3.617 20.64 3.825 ;
      RECT 20.615 3.614 20.63 3.805 ;
      RECT 20.605 3.612 20.615 3.79 ;
      RECT 20.585 3.609 20.605 3.778 ;
      RECT 20.58 3.607 20.585 3.768 ;
      RECT 20.555 3.605 20.58 3.755 ;
      RECT 20.525 3.6 20.555 3.74 ;
      RECT 20.445 3.591 20.525 3.731 ;
      RECT 20.4 3.58 20.445 3.724 ;
      RECT 20.38 3.571 20.4 3.721 ;
      RECT 20.37 3.566 20.38 3.72 ;
      RECT 20.325 3.56 20.365 3.72 ;
      RECT 20.31 3.552 20.325 3.72 ;
      RECT 20.29 3.547 20.31 3.72 ;
      RECT 20.27 3.544 20.285 3.72 ;
      RECT 20.187 3.543 20.27 3.719 ;
      RECT 20.101 3.542 20.187 3.715 ;
      RECT 20.015 3.54 20.101 3.712 ;
      RECT 19.962 3.539 20.015 3.714 ;
      RECT 19.876 3.538 19.962 3.723 ;
      RECT 19.79 3.537 19.876 3.735 ;
      RECT 19.77 3.536 19.785 3.743 ;
      RECT 19.69 3.535 19.77 3.755 ;
      RECT 19.665 3.535 19.69 3.768 ;
      RECT 19.64 3.535 19.665 3.783 ;
      RECT 19.635 3.535 19.64 3.805 ;
      RECT 19.63 3.535 19.635 3.823 ;
      RECT 19.625 3.535 19.63 3.84 ;
      RECT 19.62 3.535 19.625 3.853 ;
      RECT 19.615 3.535 19.62 3.863 ;
      RECT 19.575 3.535 19.615 3.948 ;
      RECT 19.56 3.535 19.575 4.033 ;
      RECT 19.55 3.536 19.56 4.045 ;
      RECT 19.515 3.541 19.55 4.05 ;
      RECT 19.475 3.55 19.515 4.05 ;
      RECT 19.46 3.56 19.475 4.05 ;
      RECT 19.455 3.57 19.46 4.05 ;
      RECT 19.435 3.597 19.455 4.05 ;
      RECT 19.385 3.68 19.435 4.05 ;
      RECT 19.38 3.742 19.385 4.05 ;
      RECT 19.37 3.755 19.38 4.05 ;
      RECT 19.36 3.777 19.37 4.05 ;
      RECT 19.35 3.802 19.36 4.045 ;
      RECT 19.345 3.84 19.35 4.038 ;
      RECT 19.335 3.95 19.345 4.033 ;
      RECT 20.73 4.871 20.745 5.13 ;
      RECT 20.73 4.886 20.75 5.129 ;
      RECT 20.646 4.886 20.75 5.127 ;
      RECT 20.646 4.9 20.755 5.126 ;
      RECT 20.56 4.942 20.76 5.123 ;
      RECT 20.555 4.885 20.745 5.118 ;
      RECT 20.555 4.956 20.765 5.115 ;
      RECT 20.55 4.987 20.765 5.113 ;
      RECT 20.555 4.984 20.78 5.103 ;
      RECT 20.55 5.03 20.795 5.088 ;
      RECT 20.55 5.058 20.8 5.073 ;
      RECT 20.56 4.86 20.73 5.123 ;
      RECT 20.32 3.87 20.49 4.04 ;
      RECT 20.285 3.87 20.49 4.035 ;
      RECT 20.275 3.87 20.49 4.028 ;
      RECT 20.27 3.855 20.44 4.025 ;
      RECT 19.1 4.392 19.365 4.835 ;
      RECT 19.095 4.363 19.31 4.833 ;
      RECT 19.09 4.517 19.37 4.828 ;
      RECT 19.095 4.412 19.37 4.828 ;
      RECT 19.095 4.423 19.38 4.815 ;
      RECT 19.095 4.37 19.34 4.833 ;
      RECT 19.1 4.357 19.31 4.835 ;
      RECT 19.1 4.355 19.26 4.835 ;
      RECT 19.201 4.347 19.26 4.835 ;
      RECT 19.115 4.348 19.26 4.835 ;
      RECT 19.201 4.346 19.25 4.835 ;
      RECT 19.005 3.161 19.18 3.46 ;
      RECT 19.055 3.123 19.18 3.46 ;
      RECT 19.04 3.125 19.266 3.452 ;
      RECT 19.04 3.128 19.305 3.439 ;
      RECT 19.04 3.129 19.315 3.425 ;
      RECT 18.995 3.18 19.315 3.415 ;
      RECT 19.04 3.13 19.32 3.41 ;
      RECT 18.995 3.34 19.325 3.4 ;
      RECT 18.98 3.2 19.32 3.34 ;
      RECT 18.975 3.216 19.32 3.28 ;
      RECT 19.02 3.14 19.32 3.41 ;
      RECT 19.055 3.121 19.141 3.46 ;
      RECT 17.145 3.035 17.315 4.225 ;
      RECT 17.145 3.035 17.615 3.205 ;
      RECT 17.145 9.26 17.615 9.43 ;
      RECT 17.145 8.24 17.315 9.43 ;
      RECT 16.155 3.035 16.325 4.225 ;
      RECT 16.155 3.035 16.625 3.205 ;
      RECT 16.155 9.26 16.625 9.43 ;
      RECT 16.155 8.24 16.325 9.43 ;
      RECT 14.305 3.93 14.475 5.16 ;
      RECT 14.36 2.15 14.53 4.1 ;
      RECT 14.305 1.87 14.475 2.32 ;
      RECT 14.305 10.145 14.475 10.595 ;
      RECT 14.36 8.365 14.53 10.315 ;
      RECT 14.305 7.305 14.475 8.535 ;
      RECT 13.785 1.87 13.955 5.16 ;
      RECT 13.785 3.37 14.19 3.7 ;
      RECT 13.785 2.53 14.19 2.86 ;
      RECT 13.785 7.305 13.955 10.595 ;
      RECT 13.785 9.605 14.19 9.935 ;
      RECT 13.785 8.765 14.19 9.095 ;
      RECT 11.71 4.421 11.715 4.593 ;
      RECT 11.705 4.414 11.71 4.683 ;
      RECT 11.7 4.408 11.705 4.702 ;
      RECT 11.68 4.402 11.7 4.712 ;
      RECT 11.665 4.397 11.68 4.72 ;
      RECT 11.628 4.391 11.665 4.718 ;
      RECT 11.542 4.377 11.628 4.714 ;
      RECT 11.456 4.359 11.542 4.709 ;
      RECT 11.37 4.34 11.456 4.703 ;
      RECT 11.34 4.328 11.37 4.699 ;
      RECT 11.32 4.322 11.34 4.698 ;
      RECT 11.255 4.32 11.32 4.696 ;
      RECT 11.24 4.32 11.255 4.688 ;
      RECT 11.225 4.32 11.24 4.675 ;
      RECT 11.22 4.32 11.225 4.665 ;
      RECT 11.205 4.32 11.22 4.643 ;
      RECT 11.19 4.32 11.205 4.61 ;
      RECT 11.185 4.32 11.19 4.588 ;
      RECT 11.175 4.32 11.185 4.57 ;
      RECT 11.16 4.32 11.175 4.548 ;
      RECT 11.14 4.32 11.16 4.51 ;
      RECT 11.49 3.605 11.525 4.044 ;
      RECT 11.49 3.605 11.53 4.043 ;
      RECT 11.435 3.665 11.53 4.042 ;
      RECT 11.3 3.837 11.53 4.041 ;
      RECT 11.41 3.715 11.53 4.041 ;
      RECT 11.3 3.837 11.555 4.031 ;
      RECT 11.355 3.782 11.635 3.948 ;
      RECT 11.53 3.576 11.535 4.039 ;
      RECT 11.385 3.752 11.675 3.825 ;
      RECT 11.4 3.735 11.53 4.041 ;
      RECT 11.535 3.575 11.705 3.763 ;
      RECT 11.525 3.578 11.705 3.763 ;
      RECT 11.03 3.455 11.2 3.765 ;
      RECT 11.03 3.455 11.205 3.738 ;
      RECT 11.03 3.455 11.21 3.715 ;
      RECT 11.03 3.455 11.22 3.665 ;
      RECT 11.025 3.56 11.22 3.635 ;
      RECT 11.06 3.13 11.23 3.608 ;
      RECT 11.06 3.13 11.245 3.529 ;
      RECT 11.05 3.34 11.245 3.529 ;
      RECT 11.06 3.14 11.255 3.444 ;
      RECT 10.99 3.882 10.995 4.085 ;
      RECT 10.98 3.87 10.99 4.195 ;
      RECT 10.955 3.87 10.98 4.235 ;
      RECT 10.875 3.87 10.955 4.32 ;
      RECT 10.865 3.87 10.875 4.39 ;
      RECT 10.84 3.87 10.865 4.413 ;
      RECT 10.82 3.87 10.84 4.448 ;
      RECT 10.775 3.88 10.82 4.491 ;
      RECT 10.765 3.892 10.775 4.528 ;
      RECT 10.745 3.906 10.765 4.548 ;
      RECT 10.735 3.924 10.745 4.564 ;
      RECT 10.72 3.95 10.735 4.574 ;
      RECT 10.705 3.991 10.72 4.588 ;
      RECT 10.695 4.026 10.705 4.598 ;
      RECT 10.69 4.042 10.695 4.603 ;
      RECT 10.68 4.057 10.69 4.608 ;
      RECT 10.66 4.1 10.68 4.618 ;
      RECT 10.64 4.137 10.66 4.631 ;
      RECT 10.605 4.16 10.64 4.649 ;
      RECT 10.595 4.174 10.605 4.665 ;
      RECT 10.575 4.184 10.595 4.675 ;
      RECT 10.57 4.193 10.575 4.683 ;
      RECT 10.56 4.2 10.57 4.69 ;
      RECT 10.55 4.207 10.56 4.698 ;
      RECT 10.535 4.217 10.55 4.706 ;
      RECT 10.525 4.231 10.535 4.716 ;
      RECT 10.515 4.243 10.525 4.728 ;
      RECT 10.5 4.265 10.515 4.741 ;
      RECT 10.49 4.287 10.5 4.752 ;
      RECT 10.48 4.307 10.49 4.761 ;
      RECT 10.475 4.322 10.48 4.768 ;
      RECT 10.445 4.355 10.475 4.782 ;
      RECT 10.435 4.39 10.445 4.797 ;
      RECT 10.43 4.397 10.435 4.803 ;
      RECT 10.41 4.412 10.43 4.81 ;
      RECT 10.405 4.427 10.41 4.818 ;
      RECT 10.4 4.436 10.405 4.823 ;
      RECT 10.385 4.442 10.4 4.83 ;
      RECT 10.38 4.448 10.385 4.838 ;
      RECT 10.375 4.452 10.38 4.845 ;
      RECT 10.37 4.456 10.375 4.855 ;
      RECT 10.36 4.461 10.37 4.865 ;
      RECT 10.34 4.472 10.36 4.893 ;
      RECT 10.325 4.484 10.34 4.92 ;
      RECT 10.305 4.497 10.325 4.945 ;
      RECT 10.285 4.512 10.305 4.969 ;
      RECT 10.27 4.527 10.285 4.984 ;
      RECT 10.265 4.538 10.27 4.993 ;
      RECT 10.2 4.583 10.265 5.003 ;
      RECT 10.165 4.642 10.2 5.016 ;
      RECT 10.16 4.665 10.165 5.022 ;
      RECT 10.155 4.672 10.16 5.024 ;
      RECT 10.14 4.682 10.155 5.027 ;
      RECT 10.11 4.707 10.14 5.031 ;
      RECT 10.105 4.725 10.11 5.035 ;
      RECT 10.1 4.732 10.105 5.036 ;
      RECT 10.08 4.74 10.1 5.04 ;
      RECT 10.07 4.747 10.08 5.044 ;
      RECT 10.026 4.758 10.07 5.051 ;
      RECT 9.94 4.786 10.026 5.067 ;
      RECT 9.88 4.81 9.94 5.085 ;
      RECT 9.835 4.82 9.88 5.099 ;
      RECT 9.776 4.828 9.835 5.113 ;
      RECT 9.69 4.835 9.776 5.132 ;
      RECT 9.665 4.84 9.69 5.147 ;
      RECT 9.585 4.843 9.665 5.15 ;
      RECT 9.505 4.847 9.585 5.137 ;
      RECT 9.496 4.85 9.505 5.122 ;
      RECT 9.41 4.85 9.496 5.107 ;
      RECT 9.35 4.852 9.41 5.084 ;
      RECT 9.346 4.855 9.35 5.074 ;
      RECT 9.26 4.855 9.346 5.059 ;
      RECT 9.185 4.855 9.26 5.035 ;
      RECT 10.5 3.864 10.51 4.04 ;
      RECT 10.455 3.831 10.5 4.04 ;
      RECT 10.41 3.782 10.455 4.04 ;
      RECT 10.38 3.752 10.41 4.041 ;
      RECT 10.375 3.735 10.38 4.042 ;
      RECT 10.35 3.715 10.375 4.043 ;
      RECT 10.335 3.69 10.35 4.044 ;
      RECT 10.33 3.677 10.335 4.045 ;
      RECT 10.325 3.671 10.33 4.043 ;
      RECT 10.32 3.663 10.325 4.037 ;
      RECT 10.295 3.655 10.32 4.017 ;
      RECT 10.275 3.644 10.295 3.988 ;
      RECT 10.245 3.629 10.275 3.959 ;
      RECT 10.225 3.615 10.245 3.931 ;
      RECT 10.215 3.609 10.225 3.91 ;
      RECT 10.21 3.606 10.215 3.893 ;
      RECT 10.205 3.603 10.21 3.878 ;
      RECT 10.19 3.598 10.205 3.843 ;
      RECT 10.185 3.594 10.19 3.81 ;
      RECT 10.165 3.589 10.185 3.786 ;
      RECT 10.135 3.581 10.165 3.751 ;
      RECT 10.12 3.575 10.135 3.728 ;
      RECT 10.08 3.568 10.12 3.713 ;
      RECT 10.055 3.56 10.08 3.693 ;
      RECT 10.035 3.555 10.055 3.683 ;
      RECT 10 3.549 10.035 3.678 ;
      RECT 9.955 3.54 10 3.677 ;
      RECT 9.925 3.536 9.955 3.679 ;
      RECT 9.84 3.544 9.925 3.683 ;
      RECT 9.77 3.555 9.84 3.705 ;
      RECT 9.757 3.561 9.77 3.728 ;
      RECT 9.671 3.568 9.757 3.75 ;
      RECT 9.585 3.58 9.671 3.787 ;
      RECT 9.585 3.957 9.595 4.195 ;
      RECT 9.58 3.586 9.585 3.81 ;
      RECT 9.575 3.842 9.585 4.195 ;
      RECT 9.575 3.587 9.58 3.815 ;
      RECT 9.57 3.588 9.575 4.195 ;
      RECT 9.546 3.59 9.57 4.196 ;
      RECT 9.46 3.598 9.546 4.198 ;
      RECT 9.44 3.612 9.46 4.201 ;
      RECT 9.435 3.64 9.44 4.202 ;
      RECT 9.43 3.652 9.435 4.203 ;
      RECT 9.425 3.667 9.43 4.204 ;
      RECT 9.415 3.697 9.425 4.205 ;
      RECT 9.41 3.735 9.415 4.203 ;
      RECT 9.405 3.755 9.41 4.198 ;
      RECT 9.39 3.79 9.405 4.183 ;
      RECT 9.38 3.842 9.39 4.163 ;
      RECT 9.375 3.872 9.38 4.151 ;
      RECT 9.36 3.885 9.375 4.134 ;
      RECT 9.335 3.889 9.36 4.101 ;
      RECT 9.32 3.887 9.335 4.078 ;
      RECT 9.305 3.886 9.32 4.075 ;
      RECT 9.245 3.884 9.305 4.073 ;
      RECT 9.235 3.882 9.245 4.068 ;
      RECT 9.195 3.881 9.235 4.065 ;
      RECT 9.125 3.878 9.195 4.063 ;
      RECT 9.07 3.876 9.125 4.058 ;
      RECT 9 3.87 9.07 4.053 ;
      RECT 8.991 3.87 9 4.05 ;
      RECT 8.905 3.87 8.991 4.045 ;
      RECT 8.9 3.87 8.905 4.04 ;
      RECT 10.205 3.105 10.38 3.455 ;
      RECT 10.205 3.12 10.39 3.453 ;
      RECT 10.18 3.07 10.325 3.45 ;
      RECT 10.16 3.071 10.325 3.443 ;
      RECT 10.15 3.072 10.335 3.438 ;
      RECT 10.12 3.073 10.335 3.425 ;
      RECT 10.07 3.074 10.335 3.401 ;
      RECT 10.065 3.076 10.335 3.386 ;
      RECT 10.065 3.142 10.395 3.38 ;
      RECT 10.045 3.083 10.35 3.36 ;
      RECT 10.035 3.092 10.36 3.215 ;
      RECT 10.045 3.087 10.36 3.36 ;
      RECT 10.065 3.077 10.35 3.386 ;
      RECT 9.65 4.402 9.82 4.69 ;
      RECT 9.645 4.42 9.83 4.685 ;
      RECT 9.61 4.428 9.895 4.605 ;
      RECT 9.61 4.428 9.981 4.595 ;
      RECT 9.61 4.428 10.035 4.541 ;
      RECT 9.895 4.325 10.065 4.509 ;
      RECT 9.61 4.48 10.07 4.497 ;
      RECT 9.595 4.45 10.065 4.493 ;
      RECT 9.855 4.332 9.895 4.644 ;
      RECT 9.735 4.369 10.065 4.509 ;
      RECT 9.83 4.344 9.855 4.67 ;
      RECT 9.82 4.351 10.065 4.509 ;
      RECT 9.951 3.815 10.02 4.074 ;
      RECT 9.951 3.87 10.025 4.073 ;
      RECT 9.865 3.87 10.025 4.072 ;
      RECT 9.86 3.87 10.03 4.065 ;
      RECT 9.85 3.815 10.02 4.06 ;
      RECT 9.23 3.114 9.405 3.415 ;
      RECT 9.215 3.102 9.23 3.4 ;
      RECT 9.185 3.101 9.215 3.353 ;
      RECT 9.185 3.119 9.41 3.348 ;
      RECT 9.17 3.103 9.23 3.313 ;
      RECT 9.165 3.125 9.42 3.213 ;
      RECT 9.165 3.108 9.316 3.213 ;
      RECT 9.165 3.11 9.32 3.213 ;
      RECT 9.17 3.106 9.316 3.313 ;
      RECT 9.275 4.342 9.28 4.69 ;
      RECT 9.265 4.332 9.275 4.696 ;
      RECT 9.23 4.322 9.265 4.698 ;
      RECT 9.192 4.317 9.23 4.702 ;
      RECT 9.106 4.31 9.192 4.709 ;
      RECT 9.02 4.3 9.106 4.719 ;
      RECT 8.975 4.295 9.02 4.727 ;
      RECT 8.971 4.295 8.975 4.731 ;
      RECT 8.885 4.295 8.971 4.738 ;
      RECT 8.87 4.295 8.885 4.738 ;
      RECT 8.86 4.293 8.87 4.71 ;
      RECT 8.85 4.289 8.86 4.653 ;
      RECT 8.83 4.283 8.85 4.585 ;
      RECT 8.825 4.279 8.83 4.533 ;
      RECT 8.815 4.278 8.825 4.5 ;
      RECT 8.765 4.276 8.815 4.485 ;
      RECT 8.74 4.274 8.765 4.48 ;
      RECT 8.697 4.272 8.74 4.476 ;
      RECT 8.611 4.268 8.697 4.464 ;
      RECT 8.525 4.263 8.611 4.448 ;
      RECT 8.495 4.26 8.525 4.435 ;
      RECT 8.47 4.259 8.495 4.423 ;
      RECT 8.465 4.259 8.47 4.413 ;
      RECT 8.425 4.258 8.465 4.405 ;
      RECT 8.41 4.257 8.425 4.398 ;
      RECT 8.36 4.256 8.41 4.39 ;
      RECT 8.358 4.255 8.36 4.385 ;
      RECT 8.272 4.253 8.358 4.385 ;
      RECT 8.186 4.248 8.272 4.385 ;
      RECT 8.1 4.244 8.186 4.385 ;
      RECT 8.051 4.24 8.1 4.383 ;
      RECT 7.965 4.237 8.051 4.378 ;
      RECT 7.942 4.234 7.965 4.374 ;
      RECT 7.856 4.231 7.942 4.369 ;
      RECT 7.77 4.227 7.856 4.36 ;
      RECT 7.745 4.22 7.77 4.355 ;
      RECT 7.685 4.185 7.745 4.352 ;
      RECT 7.665 4.11 7.685 4.349 ;
      RECT 7.66 4.052 7.665 4.348 ;
      RECT 7.635 3.992 7.66 4.347 ;
      RECT 7.56 3.87 7.635 4.343 ;
      RECT 7.55 3.87 7.56 4.335 ;
      RECT 7.535 3.87 7.55 4.325 ;
      RECT 7.52 3.87 7.535 4.295 ;
      RECT 7.505 3.87 7.52 4.24 ;
      RECT 7.49 3.87 7.505 4.178 ;
      RECT 7.465 3.87 7.49 4.103 ;
      RECT 7.46 3.87 7.465 4.053 ;
      RECT 8.805 3.415 8.825 3.724 ;
      RECT 8.791 3.417 8.84 3.721 ;
      RECT 8.791 3.422 8.86 3.712 ;
      RECT 8.705 3.42 8.84 3.706 ;
      RECT 8.705 3.428 8.895 3.689 ;
      RECT 8.67 3.43 8.895 3.688 ;
      RECT 8.64 3.438 8.895 3.679 ;
      RECT 8.63 3.443 8.915 3.665 ;
      RECT 8.67 3.433 8.915 3.665 ;
      RECT 8.67 3.436 8.925 3.653 ;
      RECT 8.64 3.438 8.935 3.64 ;
      RECT 8.64 3.442 8.945 3.583 ;
      RECT 8.63 3.447 8.95 3.498 ;
      RECT 8.791 3.415 8.825 3.721 ;
      RECT 8.67 10.145 8.84 10.595 ;
      RECT 8.725 8.365 8.895 10.315 ;
      RECT 8.67 7.305 8.84 8.535 ;
      RECT 8.23 3.518 8.235 3.73 ;
      RECT 8.105 3.515 8.12 3.73 ;
      RECT 7.57 3.545 7.64 3.73 ;
      RECT 7.455 3.545 7.49 3.725 ;
      RECT 8.576 3.847 8.595 4.041 ;
      RECT 8.49 3.802 8.576 4.042 ;
      RECT 8.48 3.755 8.49 4.044 ;
      RECT 8.475 3.735 8.48 4.045 ;
      RECT 8.455 3.7 8.475 4.046 ;
      RECT 8.44 3.65 8.455 4.047 ;
      RECT 8.42 3.587 8.44 4.048 ;
      RECT 8.41 3.55 8.42 4.049 ;
      RECT 8.395 3.539 8.41 4.05 ;
      RECT 8.39 3.531 8.395 4.048 ;
      RECT 8.38 3.53 8.39 4.04 ;
      RECT 8.35 3.527 8.38 4.019 ;
      RECT 8.275 3.522 8.35 3.964 ;
      RECT 8.26 3.518 8.275 3.91 ;
      RECT 8.25 3.518 8.26 3.805 ;
      RECT 8.235 3.518 8.25 3.738 ;
      RECT 8.22 3.518 8.23 3.728 ;
      RECT 8.165 3.517 8.22 3.725 ;
      RECT 8.12 3.515 8.165 3.728 ;
      RECT 8.092 3.515 8.105 3.731 ;
      RECT 8.006 3.519 8.092 3.733 ;
      RECT 7.92 3.525 8.006 3.738 ;
      RECT 7.9 3.529 7.92 3.74 ;
      RECT 7.898 3.53 7.9 3.739 ;
      RECT 7.812 3.532 7.898 3.738 ;
      RECT 7.726 3.537 7.812 3.735 ;
      RECT 7.64 3.542 7.726 3.732 ;
      RECT 7.49 3.545 7.57 3.728 ;
      RECT 8.15 7.305 8.32 10.595 ;
      RECT 8.15 9.605 8.555 9.935 ;
      RECT 8.15 8.765 8.555 9.095 ;
      RECT 8.266 4.52 8.315 4.854 ;
      RECT 8.266 4.52 8.32 4.853 ;
      RECT 8.18 4.52 8.32 4.852 ;
      RECT 7.955 4.628 8.325 4.85 ;
      RECT 8.18 4.52 8.35 4.843 ;
      RECT 8.15 4.532 8.355 4.834 ;
      RECT 8.135 4.55 8.36 4.831 ;
      RECT 7.95 4.634 8.36 4.758 ;
      RECT 7.945 4.641 8.36 4.718 ;
      RECT 7.96 4.607 8.36 4.831 ;
      RECT 8.121 4.553 8.325 4.85 ;
      RECT 8.035 4.573 8.36 4.831 ;
      RECT 8.135 4.547 8.355 4.834 ;
      RECT 7.905 3.871 8.095 4.065 ;
      RECT 7.9 3.873 8.095 4.064 ;
      RECT 7.895 3.877 8.11 4.061 ;
      RECT 7.91 3.87 8.11 4.061 ;
      RECT 7.895 3.98 8.115 4.056 ;
      RECT 7.19 4.48 7.281 4.778 ;
      RECT 7.185 4.482 7.36 4.773 ;
      RECT 7.19 4.48 7.36 4.773 ;
      RECT 7.185 4.486 7.38 4.771 ;
      RECT 7.185 4.541 7.42 4.77 ;
      RECT 7.185 4.576 7.435 4.764 ;
      RECT 7.185 4.61 7.445 4.754 ;
      RECT 7.175 4.49 7.38 4.605 ;
      RECT 7.175 4.51 7.395 4.605 ;
      RECT 7.175 4.493 7.385 4.605 ;
      RECT 7.4 3.261 7.405 3.323 ;
      RECT 7.395 3.183 7.4 3.346 ;
      RECT 7.39 3.14 7.395 3.357 ;
      RECT 7.385 3.13 7.39 3.369 ;
      RECT 7.38 3.13 7.385 3.378 ;
      RECT 7.355 3.13 7.38 3.41 ;
      RECT 7.35 3.13 7.355 3.443 ;
      RECT 7.335 3.13 7.35 3.468 ;
      RECT 7.325 3.13 7.335 3.495 ;
      RECT 7.32 3.13 7.325 3.508 ;
      RECT 7.315 3.13 7.32 3.523 ;
      RECT 7.305 3.13 7.315 3.538 ;
      RECT 7.3 3.13 7.305 3.558 ;
      RECT 7.275 3.13 7.3 3.593 ;
      RECT 7.23 3.13 7.275 3.638 ;
      RECT 7.22 3.13 7.23 3.651 ;
      RECT 7.135 3.215 7.22 3.658 ;
      RECT 7.1 3.337 7.135 3.667 ;
      RECT 7.095 3.377 7.1 3.671 ;
      RECT 7.075 3.4 7.095 3.673 ;
      RECT 7.07 3.43 7.075 3.676 ;
      RECT 7.06 3.442 7.07 3.677 ;
      RECT 7.015 3.465 7.06 3.682 ;
      RECT 6.975 3.495 7.015 3.69 ;
      RECT 6.94 3.507 6.975 3.696 ;
      RECT 6.935 3.512 6.94 3.7 ;
      RECT 6.865 3.522 6.935 3.707 ;
      RECT 6.825 3.532 6.865 3.717 ;
      RECT 6.805 3.537 6.825 3.723 ;
      RECT 6.795 3.541 6.805 3.728 ;
      RECT 6.79 3.544 6.795 3.731 ;
      RECT 6.78 3.545 6.79 3.732 ;
      RECT 6.755 3.547 6.78 3.736 ;
      RECT 6.745 3.552 6.755 3.739 ;
      RECT 6.7 3.56 6.745 3.74 ;
      RECT 6.575 3.565 6.7 3.74 ;
      RECT 7.13 3.862 7.15 4.044 ;
      RECT 7.081 3.847 7.13 4.043 ;
      RECT 6.995 3.862 7.15 4.041 ;
      RECT 6.98 3.862 7.15 4.04 ;
      RECT 6.945 3.84 7.115 4.025 ;
      RECT 7.015 4.86 7.03 5.069 ;
      RECT 7.015 4.868 7.035 5.068 ;
      RECT 6.96 4.868 7.035 5.067 ;
      RECT 6.94 4.872 7.04 5.065 ;
      RECT 6.92 4.822 6.96 5.064 ;
      RECT 6.865 4.88 7.045 5.062 ;
      RECT 6.83 4.837 6.96 5.06 ;
      RECT 6.826 4.84 7.015 5.059 ;
      RECT 6.74 4.848 7.015 5.057 ;
      RECT 6.74 4.892 7.05 5.05 ;
      RECT 6.73 4.985 7.05 5.048 ;
      RECT 6.74 4.904 7.055 5.033 ;
      RECT 6.74 4.925 7.07 5.003 ;
      RECT 6.74 4.952 7.075 4.973 ;
      RECT 6.865 4.83 6.96 5.062 ;
      RECT 6.495 3.875 6.5 4.413 ;
      RECT 6.3 4.205 6.305 4.4 ;
      RECT 4.6 3.87 4.615 4.25 ;
      RECT 6.665 3.87 6.67 4.04 ;
      RECT 6.66 3.87 6.665 4.05 ;
      RECT 6.655 3.87 6.66 4.063 ;
      RECT 6.63 3.87 6.655 4.105 ;
      RECT 6.605 3.87 6.63 4.178 ;
      RECT 6.59 3.87 6.605 4.23 ;
      RECT 6.585 3.87 6.59 4.26 ;
      RECT 6.56 3.87 6.585 4.3 ;
      RECT 6.545 3.87 6.56 4.355 ;
      RECT 6.54 3.87 6.545 4.388 ;
      RECT 6.515 3.87 6.54 4.408 ;
      RECT 6.5 3.87 6.515 4.414 ;
      RECT 6.43 3.905 6.495 4.41 ;
      RECT 6.38 3.96 6.43 4.405 ;
      RECT 6.37 3.992 6.38 4.403 ;
      RECT 6.365 4.017 6.37 4.403 ;
      RECT 6.345 4.09 6.365 4.403 ;
      RECT 6.335 4.17 6.345 4.402 ;
      RECT 6.32 4.2 6.335 4.402 ;
      RECT 6.305 4.205 6.32 4.401 ;
      RECT 6.245 4.207 6.3 4.398 ;
      RECT 6.215 4.212 6.245 4.394 ;
      RECT 6.213 4.215 6.215 4.393 ;
      RECT 6.127 4.217 6.213 4.39 ;
      RECT 6.041 4.223 6.127 4.384 ;
      RECT 5.955 4.228 6.041 4.378 ;
      RECT 5.882 4.233 5.955 4.379 ;
      RECT 5.796 4.239 5.882 4.387 ;
      RECT 5.71 4.245 5.796 4.396 ;
      RECT 5.69 4.249 5.71 4.401 ;
      RECT 5.643 4.251 5.69 4.404 ;
      RECT 5.557 4.256 5.643 4.41 ;
      RECT 5.471 4.261 5.557 4.419 ;
      RECT 5.385 4.267 5.471 4.427 ;
      RECT 5.3 4.265 5.385 4.436 ;
      RECT 5.296 4.26 5.3 4.44 ;
      RECT 5.21 4.255 5.296 4.432 ;
      RECT 5.146 4.246 5.21 4.42 ;
      RECT 5.06 4.237 5.146 4.407 ;
      RECT 5.036 4.23 5.06 4.398 ;
      RECT 4.95 4.224 5.036 4.385 ;
      RECT 4.91 4.217 4.95 4.371 ;
      RECT 4.905 4.207 4.91 4.367 ;
      RECT 4.895 4.195 4.905 4.366 ;
      RECT 4.875 4.165 4.895 4.363 ;
      RECT 4.82 4.085 4.875 4.357 ;
      RECT 4.8 4.004 4.82 4.352 ;
      RECT 4.78 3.962 4.8 4.348 ;
      RECT 4.755 3.915 4.78 4.342 ;
      RECT 4.75 3.89 4.755 4.339 ;
      RECT 4.715 3.87 4.75 4.334 ;
      RECT 4.706 3.87 4.715 4.327 ;
      RECT 4.62 3.87 4.706 4.297 ;
      RECT 4.615 3.87 4.62 4.26 ;
      RECT 4.58 3.87 4.6 4.182 ;
      RECT 4.575 3.912 4.58 4.147 ;
      RECT 4.57 3.987 4.575 4.103 ;
      RECT 6.02 3.792 6.195 4.04 ;
      RECT 6.02 3.792 6.2 4.038 ;
      RECT 6.015 3.824 6.2 3.998 ;
      RECT 6.045 3.765 6.215 3.985 ;
      RECT 6.01 3.842 6.215 3.918 ;
      RECT 5.32 3.305 5.49 3.48 ;
      RECT 5.32 3.305 5.662 3.472 ;
      RECT 5.32 3.305 5.745 3.466 ;
      RECT 5.32 3.305 5.78 3.462 ;
      RECT 5.32 3.305 5.8 3.461 ;
      RECT 5.32 3.305 5.886 3.457 ;
      RECT 5.78 3.13 5.95 3.452 ;
      RECT 5.355 3.237 5.98 3.45 ;
      RECT 5.345 3.292 5.985 3.448 ;
      RECT 5.32 3.328 5.995 3.443 ;
      RECT 5.32 3.355 6 3.373 ;
      RECT 5.385 3.18 5.96 3.45 ;
      RECT 5.576 3.165 5.96 3.45 ;
      RECT 5.41 3.168 5.96 3.45 ;
      RECT 5.49 3.166 5.576 3.477 ;
      RECT 5.576 3.163 5.955 3.45 ;
      RECT 5.76 3.14 5.955 3.45 ;
      RECT 5.662 3.161 5.955 3.45 ;
      RECT 5.745 3.155 5.76 3.463 ;
      RECT 5.895 4.52 5.9 4.72 ;
      RECT 5.36 4.585 5.405 4.72 ;
      RECT 5.93 4.52 5.95 4.693 ;
      RECT 5.9 4.52 5.93 4.708 ;
      RECT 5.835 4.52 5.895 4.745 ;
      RECT 5.82 4.52 5.835 4.775 ;
      RECT 5.805 4.52 5.82 4.788 ;
      RECT 5.785 4.52 5.805 4.803 ;
      RECT 5.78 4.52 5.785 4.812 ;
      RECT 5.77 4.524 5.78 4.817 ;
      RECT 5.755 4.534 5.77 4.828 ;
      RECT 5.73 4.55 5.755 4.838 ;
      RECT 5.72 4.564 5.73 4.84 ;
      RECT 5.7 4.576 5.72 4.837 ;
      RECT 5.67 4.597 5.7 4.831 ;
      RECT 5.66 4.609 5.67 4.826 ;
      RECT 5.65 4.607 5.66 4.823 ;
      RECT 5.635 4.606 5.65 4.818 ;
      RECT 5.63 4.605 5.635 4.813 ;
      RECT 5.595 4.603 5.63 4.803 ;
      RECT 5.575 4.6 5.595 4.785 ;
      RECT 5.565 4.598 5.575 4.78 ;
      RECT 5.555 4.597 5.565 4.775 ;
      RECT 5.52 4.595 5.555 4.763 ;
      RECT 5.465 4.591 5.52 4.743 ;
      RECT 5.455 4.589 5.465 4.728 ;
      RECT 5.45 4.589 5.455 4.723 ;
      RECT 5.405 4.587 5.45 4.72 ;
      RECT 5.31 4.585 5.36 4.724 ;
      RECT 5.3 4.586 5.31 4.729 ;
      RECT 5.24 4.593 5.3 4.743 ;
      RECT 5.215 4.601 5.24 4.763 ;
      RECT 5.205 4.605 5.215 4.775 ;
      RECT 5.2 4.606 5.205 4.78 ;
      RECT 5.185 4.608 5.2 4.783 ;
      RECT 5.17 4.61 5.185 4.788 ;
      RECT 5.165 4.61 5.17 4.791 ;
      RECT 5.12 4.615 5.165 4.802 ;
      RECT 5.115 4.619 5.12 4.814 ;
      RECT 5.09 4.615 5.115 4.818 ;
      RECT 5.08 4.611 5.09 4.822 ;
      RECT 5.07 4.61 5.08 4.826 ;
      RECT 5.055 4.6 5.07 4.832 ;
      RECT 5.05 4.588 5.055 4.836 ;
      RECT 5.045 4.585 5.05 4.837 ;
      RECT 5.04 4.582 5.045 4.839 ;
      RECT 5.025 4.57 5.04 4.838 ;
      RECT 5.01 4.552 5.025 4.835 ;
      RECT 4.99 4.531 5.01 4.828 ;
      RECT 4.925 4.52 4.99 4.8 ;
      RECT 4.921 4.52 4.925 4.779 ;
      RECT 4.835 4.52 4.921 4.749 ;
      RECT 4.82 4.52 4.835 4.705 ;
      RECT 5.395 3.62 5.4 3.855 ;
      RECT 4.525 3.536 4.53 3.74 ;
      RECT 5.105 3.565 5.11 3.72 ;
      RECT 5.025 3.545 5.03 3.72 ;
      RECT 5.695 3.687 5.71 4.04 ;
      RECT 5.621 3.672 5.695 4.04 ;
      RECT 5.535 3.655 5.621 4.04 ;
      RECT 5.525 3.645 5.535 4.038 ;
      RECT 5.52 3.643 5.525 4.033 ;
      RECT 5.505 3.641 5.52 4.019 ;
      RECT 5.435 3.633 5.505 3.959 ;
      RECT 5.415 3.624 5.435 3.893 ;
      RECT 5.41 3.621 5.415 3.873 ;
      RECT 5.4 3.62 5.41 3.863 ;
      RECT 5.39 3.62 5.395 3.847 ;
      RECT 5.38 3.619 5.39 3.837 ;
      RECT 5.37 3.617 5.38 3.825 ;
      RECT 5.355 3.614 5.37 3.805 ;
      RECT 5.345 3.612 5.355 3.79 ;
      RECT 5.325 3.609 5.345 3.778 ;
      RECT 5.32 3.607 5.325 3.768 ;
      RECT 5.295 3.605 5.32 3.755 ;
      RECT 5.265 3.6 5.295 3.74 ;
      RECT 5.185 3.591 5.265 3.731 ;
      RECT 5.14 3.58 5.185 3.724 ;
      RECT 5.12 3.571 5.14 3.721 ;
      RECT 5.11 3.566 5.12 3.72 ;
      RECT 5.065 3.56 5.105 3.72 ;
      RECT 5.05 3.552 5.065 3.72 ;
      RECT 5.03 3.547 5.05 3.72 ;
      RECT 5.01 3.544 5.025 3.72 ;
      RECT 4.927 3.543 5.01 3.719 ;
      RECT 4.841 3.542 4.927 3.715 ;
      RECT 4.755 3.54 4.841 3.712 ;
      RECT 4.702 3.539 4.755 3.714 ;
      RECT 4.616 3.538 4.702 3.723 ;
      RECT 4.53 3.537 4.616 3.735 ;
      RECT 4.51 3.536 4.525 3.743 ;
      RECT 4.43 3.535 4.51 3.755 ;
      RECT 4.405 3.535 4.43 3.768 ;
      RECT 4.38 3.535 4.405 3.783 ;
      RECT 4.375 3.535 4.38 3.805 ;
      RECT 4.37 3.535 4.375 3.823 ;
      RECT 4.365 3.535 4.37 3.84 ;
      RECT 4.36 3.535 4.365 3.853 ;
      RECT 4.355 3.535 4.36 3.863 ;
      RECT 4.315 3.535 4.355 3.948 ;
      RECT 4.3 3.535 4.315 4.033 ;
      RECT 4.29 3.536 4.3 4.045 ;
      RECT 4.255 3.541 4.29 4.05 ;
      RECT 4.215 3.55 4.255 4.05 ;
      RECT 4.2 3.56 4.215 4.05 ;
      RECT 4.195 3.57 4.2 4.05 ;
      RECT 4.175 3.597 4.195 4.05 ;
      RECT 4.125 3.68 4.175 4.05 ;
      RECT 4.12 3.742 4.125 4.05 ;
      RECT 4.11 3.755 4.12 4.05 ;
      RECT 4.1 3.777 4.11 4.05 ;
      RECT 4.09 3.802 4.1 4.045 ;
      RECT 4.085 3.84 4.09 4.038 ;
      RECT 4.075 3.95 4.085 4.033 ;
      RECT 5.47 4.871 5.485 5.13 ;
      RECT 5.47 4.886 5.49 5.129 ;
      RECT 5.386 4.886 5.49 5.127 ;
      RECT 5.386 4.9 5.495 5.126 ;
      RECT 5.3 4.942 5.5 5.123 ;
      RECT 5.295 4.885 5.485 5.118 ;
      RECT 5.295 4.956 5.505 5.115 ;
      RECT 5.29 4.987 5.505 5.113 ;
      RECT 5.295 4.984 5.52 5.103 ;
      RECT 5.29 5.03 5.535 5.088 ;
      RECT 5.29 5.058 5.54 5.073 ;
      RECT 5.3 4.86 5.47 5.123 ;
      RECT 5.06 3.87 5.23 4.04 ;
      RECT 5.025 3.87 5.23 4.035 ;
      RECT 5.015 3.87 5.23 4.028 ;
      RECT 5.01 3.855 5.18 4.025 ;
      RECT 3.84 4.392 4.105 4.835 ;
      RECT 3.835 4.363 4.05 4.833 ;
      RECT 3.83 4.517 4.11 4.828 ;
      RECT 3.835 4.412 4.11 4.828 ;
      RECT 3.835 4.423 4.12 4.815 ;
      RECT 3.835 4.37 4.08 4.833 ;
      RECT 3.84 4.357 4.05 4.835 ;
      RECT 3.84 4.355 4 4.835 ;
      RECT 3.941 4.347 4 4.835 ;
      RECT 3.855 4.348 4 4.835 ;
      RECT 3.941 4.346 3.99 4.835 ;
      RECT 3.745 3.161 3.92 3.46 ;
      RECT 3.795 3.123 3.92 3.46 ;
      RECT 3.78 3.125 4.006 3.452 ;
      RECT 3.78 3.128 4.045 3.439 ;
      RECT 3.78 3.129 4.055 3.425 ;
      RECT 3.735 3.18 4.055 3.415 ;
      RECT 3.78 3.13 4.06 3.41 ;
      RECT 3.735 3.34 4.065 3.4 ;
      RECT 3.72 3.2 4.06 3.34 ;
      RECT 3.715 3.216 4.06 3.28 ;
      RECT 3.76 3.14 4.06 3.41 ;
      RECT 3.795 3.121 3.881 3.46 ;
      RECT 1.175 10.145 1.345 10.595 ;
      RECT 1.23 8.365 1.4 10.315 ;
      RECT 1.175 7.305 1.345 8.535 ;
      RECT 0.655 7.305 0.825 10.595 ;
      RECT 0.655 9.605 1.06 9.935 ;
      RECT 0.655 8.765 1.06 9.095 ;
      RECT 78.555 7.31 78.725 8.78 ;
      RECT 78.555 10.09 78.725 10.6 ;
      RECT 77.565 1.865 77.735 2.375 ;
      RECT 77.565 3.685 77.735 5.155 ;
      RECT 77.565 7.31 77.735 8.78 ;
      RECT 77.565 10.09 77.735 10.6 ;
      RECT 76.205 1.87 76.375 5.16 ;
      RECT 76.205 7.305 76.375 10.595 ;
      RECT 75.775 1.87 75.945 2.38 ;
      RECT 75.775 2.95 75.945 5.16 ;
      RECT 75.775 7.305 75.945 9.515 ;
      RECT 75.775 10.085 75.945 10.595 ;
      RECT 70.57 7.305 70.74 10.595 ;
      RECT 70.14 7.305 70.31 9.515 ;
      RECT 70.14 10.085 70.31 10.595 ;
      RECT 63.295 7.31 63.465 8.78 ;
      RECT 63.295 10.09 63.465 10.6 ;
      RECT 62.305 1.865 62.475 2.375 ;
      RECT 62.305 3.685 62.475 5.155 ;
      RECT 62.305 7.31 62.475 8.78 ;
      RECT 62.305 10.09 62.475 10.6 ;
      RECT 60.945 1.87 61.115 5.16 ;
      RECT 60.945 7.305 61.115 10.595 ;
      RECT 60.515 1.87 60.685 2.38 ;
      RECT 60.515 2.95 60.685 5.16 ;
      RECT 60.515 7.305 60.685 9.515 ;
      RECT 60.515 10.085 60.685 10.595 ;
      RECT 55.31 7.305 55.48 10.595 ;
      RECT 54.88 7.305 55.05 9.515 ;
      RECT 54.88 10.085 55.05 10.595 ;
      RECT 48.035 7.31 48.205 8.78 ;
      RECT 48.035 10.09 48.205 10.6 ;
      RECT 47.045 1.865 47.215 2.375 ;
      RECT 47.045 3.685 47.215 5.155 ;
      RECT 47.045 7.31 47.215 8.78 ;
      RECT 47.045 10.09 47.215 10.6 ;
      RECT 45.685 1.87 45.855 5.16 ;
      RECT 45.685 7.305 45.855 10.595 ;
      RECT 45.255 1.87 45.425 2.38 ;
      RECT 45.255 2.95 45.425 5.16 ;
      RECT 45.255 7.305 45.425 9.515 ;
      RECT 45.255 10.085 45.425 10.595 ;
      RECT 40.05 7.305 40.22 10.595 ;
      RECT 39.62 7.305 39.79 9.515 ;
      RECT 39.62 10.085 39.79 10.595 ;
      RECT 32.775 7.31 32.945 8.78 ;
      RECT 32.775 10.09 32.945 10.6 ;
      RECT 31.785 1.865 31.955 2.375 ;
      RECT 31.785 3.685 31.955 5.155 ;
      RECT 31.785 7.31 31.955 8.78 ;
      RECT 31.785 10.09 31.955 10.6 ;
      RECT 30.425 1.87 30.595 5.16 ;
      RECT 30.425 7.305 30.595 10.595 ;
      RECT 29.995 1.87 30.165 2.38 ;
      RECT 29.995 2.95 30.165 5.16 ;
      RECT 29.995 7.305 30.165 9.515 ;
      RECT 29.995 10.085 30.165 10.595 ;
      RECT 24.79 7.305 24.96 10.595 ;
      RECT 24.36 7.305 24.53 9.515 ;
      RECT 24.36 10.085 24.53 10.595 ;
      RECT 17.515 7.31 17.685 8.78 ;
      RECT 17.515 10.09 17.685 10.6 ;
      RECT 16.525 1.865 16.695 2.375 ;
      RECT 16.525 3.685 16.695 5.155 ;
      RECT 16.525 7.31 16.695 8.78 ;
      RECT 16.525 10.09 16.695 10.6 ;
      RECT 15.165 1.87 15.335 5.16 ;
      RECT 15.165 7.305 15.335 10.595 ;
      RECT 14.735 1.87 14.905 2.38 ;
      RECT 14.735 2.95 14.905 5.16 ;
      RECT 14.735 7.305 14.905 9.515 ;
      RECT 14.735 10.085 14.905 10.595 ;
      RECT 9.53 7.305 9.7 10.595 ;
      RECT 9.1 7.305 9.27 9.515 ;
      RECT 9.1 10.085 9.27 10.595 ;
      RECT 1.605 7.305 1.775 9.515 ;
      RECT 1.605 10.085 1.775 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r2

END LIBRARY
