magic
tech sky130A
magscale 1 2
timestamp 1708003897
<< error_s >>
rect 1058 2104 1059 2115
rect 1248 2104 1249 2115
rect 1334 2104 1335 2115
rect 2185 2104 2186 2115
rect 2375 2104 2376 2115
rect 2461 2104 2462 2115
rect 2734 2104 2735 2115
rect 2932 2104 2933 2115
rect 1069 2064 1070 2104
rect 1259 2064 1260 2104
rect 1345 2064 1346 2104
rect 2196 2064 2197 2104
rect 2386 2064 2387 2104
rect 2472 2064 2473 2104
rect 2745 2064 2746 2104
rect 2943 2064 2944 2104
rect 2393 1937 2420 1944
rect 2393 1916 2461 1937
rect 2393 1910 2448 1916
rect 2432 1909 2433 1910
rect 2405 1903 2460 1909
rect 2432 1881 2433 1903
rect 1058 1674 1059 1685
rect 1248 1674 1249 1685
rect 1334 1674 1335 1685
rect 2185 1674 2186 1685
rect 2375 1674 2376 1685
rect 2461 1674 2462 1685
rect 2734 1674 2735 1685
rect 2932 1674 2933 1685
rect 1069 1478 1070 1674
rect 1259 1478 1260 1674
rect 1345 1478 1346 1674
rect 2196 1478 2197 1674
rect 2386 1478 2387 1674
rect 2472 1478 2473 1674
rect 2745 1478 2746 1674
rect 2943 1478 2944 1674
rect 1383 1374 1407 1408
rect 2510 1374 2534 1408
rect 2510 1085 2534 1119
rect 1230 1054 1239 1055
rect 1150 1049 1230 1054
rect 1239 1050 1275 1054
rect 1275 1049 1277 1050
rect 882 1041 1150 1049
rect 1277 1041 1294 1049
rect 871 1040 882 1041
rect 851 1038 882 1040
rect 1295 1038 1299 1041
rect 833 1027 871 1038
rect 1301 1030 1307 1036
rect 500 1025 539 1026
rect 500 1024 537 1025
rect 539 1024 540 1025
rect 498 1022 500 1024
rect 526 1016 538 1024
rect 540 1022 541 1024
rect 800 1022 833 1027
rect 1205 1025 1261 1027
rect 541 1016 547 1022
rect 788 1020 833 1022
rect 1100 1021 1205 1025
rect 1261 1021 1271 1025
rect 788 1016 844 1020
rect 489 1015 541 1016
rect 488 1012 489 1015
rect 547 1013 548 1016
rect 544 1012 548 1013
rect 788 1014 804 1016
rect 832 1015 844 1016
rect 806 1014 828 1015
rect 840 1014 844 1015
rect 788 1012 849 1014
rect 880 1012 1100 1021
rect 1271 1017 1282 1021
rect 1271 1014 1289 1017
rect 1292 1014 1357 1030
rect 1271 1012 1357 1014
rect 478 1005 484 1011
rect 487 1008 488 1012
rect 486 1005 487 1008
rect 524 1005 530 1011
rect 472 999 478 1005
rect 530 999 536 1005
rect 498 990 499 997
rect 537 995 538 1012
rect 543 1001 550 1012
rect 788 1011 846 1012
rect 779 1008 785 1011
rect 786 1009 788 1011
rect 790 1010 795 1011
rect 789 1009 795 1010
rect 849 1009 850 1011
rect 871 1010 879 1012
rect 1277 1011 1286 1012
rect 1271 1010 1284 1011
rect 1292 1010 1357 1012
rect 786 1008 793 1009
rect 851 1008 871 1010
rect 779 1006 787 1008
rect 772 1005 787 1006
rect 789 1005 793 1008
rect 769 1001 787 1005
rect 841 1001 844 1008
rect 543 998 544 1001
rect 542 997 543 998
rect 536 990 538 994
rect 539 990 543 997
rect 751 994 769 1001
rect 772 997 787 1001
rect 498 989 515 990
rect 499 988 515 989
rect 484 978 515 988
rect 519 978 550 990
rect 726 985 751 994
rect 772 990 788 997
rect 842 996 843 1000
rect 847 998 871 1008
rect 1271 1009 1283 1010
rect 1284 1009 1357 1010
rect 1373 1009 1454 1030
rect 2185 1015 2186 1026
rect 2375 1015 2376 1026
rect 2461 1015 2462 1026
rect 2734 1015 2735 1026
rect 2931 1015 2932 1026
rect 1271 1005 1292 1009
rect 847 996 856 998
rect 842 995 844 996
rect 847 995 851 996
rect 787 988 788 990
rect 710 979 726 985
rect 484 972 550 978
rect 696 974 710 979
rect 445 967 451 968
rect 206 965 208 967
rect 261 964 262 967
rect 438 964 442 967
rect 451 964 458 967
rect 262 962 264 964
rect 425 956 438 964
rect 458 963 463 964
rect 463 959 474 963
rect 500 961 516 972
rect 518 966 538 972
rect 688 971 694 973
rect 772 972 788 988
rect 832 992 847 995
rect 853 993 855 996
rect 832 986 848 992
rect 854 988 855 993
rect 851 986 854 988
rect 997 986 1018 1002
rect 1264 1001 1271 1005
rect 1277 1001 1292 1005
rect 1250 994 1264 1001
rect 1284 998 1292 1001
rect 1310 1005 1320 1009
rect 1454 1005 1471 1009
rect 1310 1003 1323 1005
rect 1292 995 1293 998
rect 832 985 856 986
rect 1211 985 1217 991
rect 1233 985 1250 994
rect 1257 985 1263 991
rect 1293 985 1300 995
rect 831 983 832 985
rect 836 974 856 985
rect 1031 974 1043 982
rect 1053 974 1065 982
rect 1205 979 1211 985
rect 1263 979 1269 985
rect 1295 980 1303 985
rect 1295 979 1304 980
rect 1295 978 1305 979
rect 1295 975 1307 978
rect 836 971 848 974
rect 1295 973 1309 975
rect 1310 973 1311 1003
rect 1316 993 1337 1003
rect 1471 999 1493 1005
rect 1493 997 1495 999
rect 1320 983 1337 993
rect 1495 992 1501 997
rect 1501 986 1505 992
rect 1295 971 1311 973
rect 1316 972 1337 983
rect 1505 982 1508 986
rect 1508 975 1512 982
rect 1316 971 1438 972
rect 1512 971 1514 975
rect 683 970 688 971
rect 680 969 683 970
rect 788 968 806 971
rect 832 970 848 971
rect 1025 970 1027 971
rect 1067 970 1104 971
rect 832 969 845 970
rect 580 967 584 968
rect 586 967 591 968
rect 518 961 534 966
rect 572 965 580 967
rect 570 964 572 965
rect 591 964 594 967
rect 672 966 679 968
rect 668 964 672 966
rect 567 963 570 964
rect 566 962 567 963
rect 594 962 597 964
rect 664 963 668 964
rect 486 959 534 961
rect 463 958 478 959
rect 486 958 536 959
rect 559 958 568 962
rect 597 959 601 962
rect 644 961 664 963
rect 466 956 480 958
rect 481 957 536 958
rect 422 954 425 956
rect 466 954 483 956
rect 486 954 536 957
rect 555 956 568 958
rect 601 956 604 959
rect 652 958 658 961
rect 551 954 568 956
rect 604 954 607 956
rect 641 954 649 957
rect 773 956 779 959
rect 788 956 804 968
rect 806 967 813 968
rect 813 965 824 967
rect 832 966 844 969
rect 831 965 844 966
rect 824 964 844 965
rect 864 964 870 970
rect 910 966 916 970
rect 1019 969 1025 970
rect 900 964 916 966
rect 832 962 844 964
rect 751 954 779 956
rect 262 946 263 949
rect 261 945 300 946
rect 259 944 261 945
rect 244 934 259 944
rect 220 920 244 934
rect 217 918 220 920
rect 210 913 217 918
rect 262 913 263 945
rect 300 944 327 945
rect 404 944 422 954
rect 466 953 536 954
rect 466 951 488 953
rect 517 951 518 953
rect 524 951 530 953
rect 544 951 568 954
rect 466 948 568 951
rect 466 947 521 948
rect 524 947 530 948
rect 466 946 500 947
rect 502 946 521 947
rect 533 946 568 948
rect 466 944 521 946
rect 531 945 568 946
rect 530 944 568 945
rect 607 953 630 954
rect 638 953 641 954
rect 607 946 638 953
rect 607 944 630 946
rect 327 938 568 944
rect 597 938 612 944
rect 620 939 630 944
rect 626 938 630 939
rect 679 938 769 954
rect 773 953 799 954
rect 831 953 837 959
rect 858 958 922 964
rect 969 963 975 969
rect 1015 968 1021 969
rect 1010 966 1021 968
rect 1004 964 1009 966
rect 1000 963 1004 964
rect 1015 963 1021 966
rect 1031 968 1065 970
rect 1069 969 1077 970
rect 864 954 916 958
rect 963 957 969 963
rect 1021 957 1027 963
rect 779 947 785 953
rect 825 947 831 953
rect 864 938 878 954
rect 388 922 404 938
rect 450 937 473 938
rect 450 934 478 937
rect 450 933 486 934
rect 488 933 496 935
rect 517 934 518 938
rect 592 937 597 938
rect 583 935 591 936
rect 519 934 566 935
rect 578 934 583 935
rect 503 933 566 934
rect 630 933 646 938
rect 673 936 679 938
rect 864 936 879 938
rect 669 935 672 936
rect 664 933 668 934
rect 450 925 558 933
rect 517 924 518 925
rect 456 922 473 924
rect 388 916 404 920
rect 439 917 454 922
rect 477 920 502 922
rect 290 913 331 916
rect 335 913 404 916
rect 207 911 210 913
rect 262 911 290 913
rect 388 911 432 913
rect 438 911 454 917
rect 475 917 502 920
rect 521 918 580 922
rect 628 920 664 933
rect 862 931 879 936
rect 858 928 862 931
rect 851 924 858 928
rect 843 920 851 924
rect 864 920 879 931
rect 910 920 912 954
rect 916 950 929 954
rect 1031 953 1052 968
rect 1062 967 1065 968
rect 1070 963 1077 969
rect 1105 966 1112 970
rect 1295 969 1309 971
rect 1310 970 1438 971
rect 1320 969 1337 970
rect 1341 969 1438 970
rect 1073 960 1075 963
rect 1291 960 1294 961
rect 1078 954 1085 957
rect 1030 952 1052 953
rect 1030 950 1031 952
rect 916 942 924 950
rect 1029 938 1030 949
rect 1085 940 1108 954
rect 1210 953 1211 957
rect 1269 954 1291 960
rect 1295 957 1314 969
rect 1269 952 1296 954
rect 916 920 924 932
rect 623 918 628 920
rect 503 917 580 918
rect 475 915 487 917
rect 547 916 558 917
rect 495 914 507 916
rect 546 915 548 916
rect 203 909 207 911
rect 261 910 263 911
rect 259 906 264 910
rect 206 903 207 904
rect 197 894 198 899
rect 251 896 252 904
rect 258 903 264 906
rect 388 904 404 911
rect 432 910 457 911
rect 423 908 454 910
rect 457 909 468 910
rect 468 908 475 909
rect 413 906 454 908
rect 475 907 488 908
rect 496 906 503 907
rect 423 905 454 906
rect 438 904 454 905
rect 256 899 264 903
rect 256 895 258 899
rect 250 876 252 895
rect 404 888 420 904
rect 422 888 438 904
rect 515 888 517 911
rect 580 909 596 917
rect 612 913 623 918
rect 607 911 611 913
rect 601 909 607 911
rect 630 909 646 920
rect 830 912 843 920
rect 862 918 916 920
rect 927 918 929 926
rect 966 920 969 937
rect 1108 935 1117 940
rect 1204 939 1210 952
rect 1214 946 1235 949
rect 1251 946 1252 949
rect 1263 948 1269 952
rect 1280 946 1296 952
rect 1204 936 1211 939
rect 1212 938 1214 946
rect 1235 939 1296 946
rect 1309 942 1314 957
rect 1337 968 1438 969
rect 1515 968 1516 970
rect 1243 938 1296 939
rect 1262 937 1312 938
rect 1029 925 1032 929
rect 1117 928 1128 935
rect 1204 933 1212 936
rect 1262 933 1269 937
rect 858 912 928 918
rect 963 917 965 919
rect 1032 918 1047 925
rect 1128 923 1132 928
rect 1132 920 1133 923
rect 1047 917 1070 918
rect 963 916 969 917
rect 961 912 969 916
rect 828 911 830 912
rect 862 911 877 912
rect 878 911 879 912
rect 580 908 646 909
rect 566 907 646 908
rect 822 907 828 911
rect 862 907 883 911
rect 900 908 916 912
rect 524 906 547 907
rect 580 904 646 907
rect 614 888 630 904
rect 808 900 822 907
rect 862 904 877 907
rect 878 904 879 907
rect 910 906 916 908
rect 919 904 928 912
rect 963 911 969 912
rect 1021 916 1070 917
rect 1021 911 1027 916
rect 1038 914 1070 916
rect 1047 913 1071 914
rect 1047 911 1070 913
rect 1073 911 1098 913
rect 1112 911 1126 920
rect 1133 918 1134 920
rect 1199 918 1204 933
rect 1210 927 1217 933
rect 1210 925 1212 927
rect 1134 911 1137 918
rect 1197 911 1199 915
rect 958 907 960 911
rect 863 900 876 904
rect 917 900 919 904
rect 954 900 958 907
rect 969 905 975 911
rect 788 888 811 900
rect 858 897 863 900
rect 842 888 858 897
rect 875 896 878 899
rect 912 896 917 899
rect 952 897 954 900
rect 878 888 894 896
rect 896 888 912 896
rect 946 888 952 897
rect 256 875 264 888
rect 452 880 582 888
rect 785 883 788 888
rect 834 883 842 888
rect 943 883 946 888
rect 700 880 748 883
rect 430 875 472 880
rect 250 873 256 875
rect 419 873 472 875
rect 207 870 211 873
rect 240 871 250 873
rect 253 872 256 873
rect 240 870 252 871
rect 400 870 472 873
rect 515 870 517 880
rect 559 879 700 880
rect 562 875 700 879
rect 748 875 749 880
rect 781 875 785 883
rect 820 876 834 883
rect 938 876 943 883
rect 814 875 820 876
rect 981 875 1005 910
rect 1015 905 1021 911
rect 1047 909 1126 911
rect 1137 909 1138 911
rect 1060 904 1126 909
rect 1138 904 1140 908
rect 1076 888 1092 904
rect 1094 893 1110 904
rect 1140 899 1142 903
rect 1142 893 1144 899
rect 1185 898 1197 910
rect 1206 909 1210 925
rect 1243 916 1251 933
rect 1257 927 1263 933
rect 1205 904 1206 909
rect 1223 905 1243 915
rect 1210 903 1222 905
rect 1223 903 1244 905
rect 1262 904 1263 927
rect 1296 922 1312 937
rect 1314 936 1315 941
rect 1337 938 1358 968
rect 1378 965 1438 968
rect 1516 967 1517 968
rect 1517 965 1520 967
rect 1407 963 1438 965
rect 1520 963 1522 965
rect 1416 961 1438 963
rect 1522 961 1526 963
rect 1370 938 1386 954
rect 1388 938 1404 954
rect 1428 949 1456 961
rect 1526 954 1535 961
rect 1414 938 1415 949
rect 1456 947 1460 949
rect 1535 947 1543 954
rect 1460 946 1461 947
rect 1461 944 1462 946
rect 1543 944 1545 947
rect 1731 944 1732 949
rect 1760 944 1776 954
rect 1462 939 1468 944
rect 1545 940 1550 944
rect 1714 940 1781 944
rect 1550 939 1552 940
rect 1691 939 1714 940
rect 1337 936 1370 938
rect 1375 936 1420 938
rect 1468 936 1470 938
rect 1552 936 1555 939
rect 1688 936 1691 939
rect 1731 938 1732 940
rect 1781 938 1782 939
rect 1315 916 1320 933
rect 1337 922 1369 936
rect 1406 934 1420 936
rect 1470 934 1472 936
rect 1555 934 1559 936
rect 1685 934 1688 936
rect 1400 932 1420 934
rect 1472 932 1473 934
rect 1559 932 1561 934
rect 1684 932 1685 934
rect 1321 915 1327 921
rect 1337 919 1358 922
rect 1362 921 1369 922
rect 1358 915 1361 919
rect 1362 915 1373 921
rect 1315 909 1321 915
rect 1320 908 1321 909
rect 1362 906 1369 915
rect 1373 909 1379 915
rect 1411 904 1447 932
rect 1473 925 1480 932
rect 1561 925 1572 932
rect 1681 925 1684 932
rect 1480 924 1494 925
rect 1472 915 1494 924
rect 1572 919 1581 925
rect 1678 919 1681 925
rect 1581 916 1584 919
rect 1677 916 1678 919
rect 1480 907 1494 915
rect 1584 912 1589 916
rect 1675 912 1677 916
rect 1589 907 1593 912
rect 1672 910 1675 912
rect 1488 905 1497 907
rect 1494 904 1497 905
rect 1593 904 1595 907
rect 1207 901 1247 903
rect 1204 900 1205 901
rect 1203 899 1204 900
rect 1207 899 1243 901
rect 1202 898 1207 899
rect 1185 896 1207 898
rect 1145 893 1197 896
rect 1202 893 1207 896
rect 1094 888 1113 893
rect 1144 888 1197 893
rect 1041 877 1050 881
rect 1088 877 1097 881
rect 1107 879 1113 888
rect 1139 886 1153 888
rect 1134 883 1139 886
rect 1144 883 1153 886
rect 1133 882 1153 883
rect 1125 880 1153 882
rect 1122 879 1153 880
rect 1107 877 1153 879
rect 1033 875 1153 877
rect 562 870 664 875
rect 702 874 856 875
rect 702 872 849 874
rect 675 871 702 872
rect 667 870 675 871
rect 211 869 240 870
rect 248 867 252 870
rect 396 869 400 870
rect 662 869 667 870
rect 247 866 252 867
rect 383 866 396 869
rect 653 868 662 869
rect 645 866 653 868
rect 749 867 752 872
rect 781 871 785 872
rect 814 871 820 872
rect 856 871 870 874
rect 936 871 938 875
rect 952 872 1033 875
rect 1041 872 1153 875
rect 1185 872 1197 888
rect 1198 881 1203 893
rect 1202 880 1203 881
rect 870 870 874 871
rect 195 859 196 866
rect 245 864 252 866
rect 361 865 395 866
rect 640 865 645 866
rect 245 859 247 864
rect 361 862 383 865
rect 360 859 383 862
rect 395 859 402 865
rect 607 859 640 865
rect 244 855 245 859
rect 356 855 361 859
rect 364 854 383 859
rect 402 857 405 859
rect 601 858 607 859
rect 594 857 601 858
rect 578 854 593 857
rect 752 854 757 866
rect 779 863 781 870
rect 811 863 814 870
rect 874 868 886 870
rect 778 860 779 863
rect 810 860 811 863
rect 886 859 924 868
rect 929 863 934 870
rect 952 868 1041 872
rect 1042 870 1153 872
rect 1223 871 1243 899
rect 1247 893 1251 901
rect 1251 873 1256 893
rect 1359 887 1362 904
rect 1419 903 1422 904
rect 1415 902 1419 903
rect 1414 899 1415 901
rect 1447 899 1454 904
rect 1407 887 1414 899
rect 1419 897 1420 899
rect 1453 893 1454 899
rect 1489 893 1496 898
rect 1497 893 1512 904
rect 1362 877 1387 887
rect 1413 877 1414 887
rect 1496 885 1508 893
rect 1512 887 1521 893
rect 1595 887 1608 904
rect 1668 902 1680 910
rect 1690 902 1702 910
rect 1742 904 1743 938
rect 1781 934 1792 938
rect 1782 922 1792 934
rect 1782 903 1783 922
rect 1668 898 1671 902
rect 1704 899 1706 902
rect 1656 886 1664 898
rect 1668 896 1702 898
rect 1668 895 1671 896
rect 1387 870 1414 877
rect 1508 876 1515 885
rect 1521 879 1527 886
rect 1608 879 1613 886
rect 1527 877 1529 879
rect 1613 877 1615 879
rect 1419 870 1420 872
rect 950 866 952 868
rect 947 864 950 866
rect 977 864 980 868
rect 927 860 929 863
rect 243 851 244 854
rect 354 851 356 854
rect 363 850 364 854
rect 194 838 195 850
rect 239 838 243 850
rect 347 838 354 850
rect 193 816 194 837
rect 232 816 239 838
rect 347 835 353 838
rect 341 829 347 835
rect 355 828 360 842
rect 393 835 399 841
rect 405 839 406 854
rect 482 850 578 854
rect 757 850 758 854
rect 776 853 778 859
rect 807 853 810 859
rect 919 858 929 859
rect 919 853 926 858
rect 929 857 935 858
rect 944 857 947 864
rect 1032 863 1041 868
rect 1097 863 1106 870
rect 1115 868 1116 870
rect 1153 868 1154 870
rect 975 860 977 863
rect 1116 861 1118 868
rect 1154 860 1157 868
rect 1183 864 1184 866
rect 1182 861 1183 863
rect 1198 859 1204 870
rect 1220 864 1223 870
rect 1256 866 1258 870
rect 1295 868 1296 869
rect 1293 865 1295 868
rect 1286 864 1293 865
rect 1210 859 1212 861
rect 935 855 958 857
rect 973 856 975 859
rect 1034 856 1040 857
rect 1080 856 1086 857
rect 1119 856 1120 857
rect 1158 856 1159 857
rect 1180 856 1181 859
rect 1206 856 1214 859
rect 935 854 948 855
rect 968 854 973 856
rect 919 852 922 853
rect 919 851 921 852
rect 943 851 944 854
rect 948 851 989 854
rect 422 843 483 850
rect 421 841 422 842
rect 399 832 405 835
rect 406 832 407 838
rect 399 829 407 832
rect 415 829 421 841
rect 425 840 436 842
rect 482 840 483 843
rect 493 843 683 850
rect 758 846 761 850
rect 768 846 776 851
rect 799 847 807 851
rect 794 846 855 847
rect 705 843 787 846
rect 493 839 578 843
rect 671 842 689 843
rect 758 842 761 843
rect 653 839 671 842
rect 689 841 701 842
rect 704 839 707 841
rect 491 838 493 839
rect 486 835 490 838
rect 480 830 486 835
rect 513 831 515 839
rect 645 838 653 839
rect 629 835 645 838
rect 403 828 407 829
rect 479 828 480 830
rect 192 810 193 816
rect 231 811 232 816
rect 260 810 276 824
rect 354 813 355 828
rect 399 826 401 827
rect 403 826 415 828
rect 401 816 422 826
rect 452 817 468 824
rect 399 813 422 816
rect 399 811 401 813
rect 229 807 231 810
rect 405 808 415 813
rect 244 805 255 808
rect 404 806 405 808
rect 422 807 432 813
rect 442 812 468 817
rect 440 809 468 812
rect 438 808 449 809
rect 452 808 468 809
rect 470 808 486 824
rect 509 818 515 831
rect 595 830 629 835
rect 553 824 595 830
rect 707 829 709 839
rect 761 829 766 842
rect 768 828 776 843
rect 548 823 595 824
rect 545 822 564 823
rect 520 818 545 822
rect 509 816 520 818
rect 505 813 515 816
rect 505 812 513 813
rect 436 807 452 808
rect 432 806 452 807
rect 432 805 449 806
rect 486 805 502 808
rect 191 800 192 805
rect 226 800 228 805
rect 225 798 226 800
rect 221 790 225 798
rect 244 792 257 805
rect 400 797 404 805
rect 430 803 463 805
rect 485 804 502 805
rect 190 782 191 789
rect 219 785 221 789
rect 189 771 190 781
rect 218 773 219 782
rect 255 775 257 792
rect 354 790 355 796
rect 340 787 355 790
rect 396 789 400 796
rect 430 794 458 803
rect 482 800 502 804
rect 479 797 502 800
rect 430 793 452 794
rect 436 792 452 793
rect 442 789 452 792
rect 476 792 502 797
rect 476 790 486 792
rect 476 789 502 790
rect 396 788 406 789
rect 340 783 376 787
rect 340 782 379 783
rect 393 782 406 788
rect 436 783 452 789
rect 468 786 502 789
rect 465 783 502 786
rect 340 778 390 782
rect 391 778 406 782
rect 340 774 406 778
rect 430 781 452 783
rect 458 781 502 783
rect 430 774 502 781
rect 509 777 513 812
rect 532 803 533 808
rect 537 803 546 812
rect 548 808 564 822
rect 566 808 582 823
rect 584 808 593 812
rect 644 808 660 824
rect 662 808 678 824
rect 709 808 713 828
rect 766 825 776 828
rect 799 825 807 846
rect 856 843 869 846
rect 873 842 875 843
rect 877 842 919 851
rect 875 839 919 842
rect 877 835 919 839
rect 935 846 989 851
rect 994 853 1206 856
rect 1216 855 1220 863
rect 1244 859 1286 864
rect 1315 863 1321 869
rect 1373 863 1379 869
rect 1387 868 1415 870
rect 1515 868 1516 870
rect 1407 867 1425 868
rect 1407 865 1428 867
rect 1488 865 1490 868
rect 1529 865 1535 877
rect 1416 863 1425 865
rect 1215 854 1216 855
rect 1208 853 1221 854
rect 994 846 1221 853
rect 935 835 965 846
rect 989 845 1221 846
rect 989 843 1001 845
rect 1016 843 1034 845
rect 877 830 965 835
rect 977 831 989 843
rect 1123 842 1124 845
rect 1159 840 1165 845
rect 877 825 919 830
rect 929 828 953 830
rect 973 828 977 831
rect 1125 830 1128 838
rect 1166 830 1169 838
rect 1172 830 1178 845
rect 1199 839 1221 845
rect 1260 840 1265 858
rect 1321 857 1327 863
rect 1321 841 1326 857
rect 1363 841 1365 863
rect 1367 857 1373 863
rect 1415 862 1425 863
rect 1416 861 1425 862
rect 1416 859 1431 861
rect 1488 859 1494 865
rect 1535 864 1536 865
rect 1419 856 1444 859
rect 1419 853 1434 856
rect 1436 853 1442 856
rect 1472 854 1481 859
rect 1482 854 1488 859
rect 1518 857 1519 861
rect 1536 859 1538 864
rect 1538 856 1540 859
rect 1425 850 1434 853
rect 1472 850 1491 854
rect 1480 846 1491 850
rect 1491 842 1492 846
rect 1519 842 1522 854
rect 1540 850 1543 856
rect 1615 851 1631 877
rect 1668 868 1670 895
rect 1668 864 1671 868
rect 1700 864 1702 896
rect 1706 889 1714 898
rect 1706 879 1733 889
rect 1780 881 1783 885
rect 1773 879 1780 881
rect 1706 870 1773 879
rect 1708 865 1773 870
rect 1704 864 1708 865
rect 1664 856 1665 861
rect 1663 854 1665 856
rect 1543 845 1547 850
rect 1547 843 1549 845
rect 1631 844 1636 850
rect 1549 842 1550 843
rect 1550 841 1552 842
rect 1321 839 1354 841
rect 1128 828 1129 830
rect 929 825 938 828
rect 765 824 771 825
rect 765 814 774 824
rect 584 803 598 808
rect 528 794 541 803
rect 537 787 541 794
rect 587 794 602 803
rect 587 792 598 794
rect 628 792 644 808
rect 679 807 694 808
rect 763 807 765 813
rect 771 812 774 814
rect 796 813 798 824
rect 836 814 852 824
rect 829 813 852 814
rect 854 813 877 824
rect 921 820 929 825
rect 933 824 938 825
rect 912 813 921 820
rect 932 813 938 824
rect 953 823 979 828
rect 943 822 986 823
rect 943 821 984 822
rect 973 813 977 821
rect 986 818 993 822
rect 993 816 994 818
rect 772 808 774 812
rect 678 802 694 807
rect 680 799 694 802
rect 713 800 714 807
rect 762 804 763 807
rect 761 800 762 803
rect 774 800 790 808
rect 795 807 796 813
rect 829 808 870 813
rect 820 806 841 808
rect 852 807 858 808
rect 794 800 795 806
rect 820 802 836 806
rect 846 802 852 807
rect 817 801 863 802
rect 817 800 858 801
rect 634 790 640 792
rect 643 791 644 792
rect 671 792 694 799
rect 714 797 716 800
rect 671 791 686 792
rect 642 790 644 791
rect 628 787 644 790
rect 645 789 647 790
rect 680 789 686 791
rect 645 787 686 789
rect 716 787 726 797
rect 759 790 761 797
rect 774 792 794 800
rect 789 790 794 792
rect 817 792 836 800
rect 870 792 886 808
rect 898 807 904 813
rect 905 807 912 813
rect 932 809 933 813
rect 994 812 997 816
rect 1028 813 1044 824
rect 1046 813 1062 824
rect 1097 816 1106 825
rect 1129 824 1130 828
rect 1086 815 1097 816
rect 1019 812 1021 813
rect 1059 812 1063 813
rect 972 809 973 812
rect 1019 810 1063 812
rect 1019 808 1053 810
rect 904 801 910 807
rect 916 792 932 808
rect 817 790 827 792
rect 829 790 836 792
rect 758 787 759 789
rect 628 785 683 787
rect 539 777 540 785
rect 601 777 607 783
rect 628 781 651 785
rect 219 768 220 771
rect 356 767 372 774
rect 374 767 390 774
rect 430 771 438 774
rect 442 771 488 774
rect 438 767 441 769
rect 452 767 468 771
rect 470 767 486 771
rect 188 743 189 767
rect 220 742 223 767
rect 356 759 390 767
rect 442 759 486 767
rect 356 758 372 759
rect 374 758 393 759
rect 452 758 468 759
rect 470 758 486 759
rect 509 763 512 777
rect 519 770 520 771
rect 516 766 520 770
rect 513 763 520 766
rect 322 749 342 753
rect 378 752 393 758
rect 509 757 520 763
rect 322 748 345 749
rect 322 746 368 748
rect 384 747 393 752
rect 449 751 458 756
rect 485 755 520 757
rect 537 756 540 777
rect 502 754 520 755
rect 485 751 520 754
rect 445 747 520 751
rect 528 747 540 756
rect 606 771 613 777
rect 628 774 649 781
rect 322 744 376 746
rect 322 743 383 744
rect 393 743 402 747
rect 427 745 520 747
rect 414 743 520 745
rect 322 740 520 743
rect 393 738 402 740
rect 408 737 514 740
rect 537 738 546 747
rect 548 741 555 747
rect 223 733 224 737
rect 486 730 488 737
rect 509 730 515 737
rect 606 731 607 771
rect 634 753 649 774
rect 681 778 682 785
rect 686 778 695 787
rect 681 756 683 778
rect 687 775 695 778
rect 724 782 739 787
rect 756 782 758 787
rect 774 782 794 790
rect 724 778 794 782
rect 820 780 836 790
rect 724 774 799 778
rect 740 772 756 774
rect 758 772 774 774
rect 789 772 799 774
rect 817 774 836 780
rect 870 774 886 790
rect 916 780 932 790
rect 967 789 972 808
rect 1002 803 1004 806
rect 1012 805 1028 808
rect 1063 807 1078 808
rect 1088 807 1097 815
rect 1124 810 1140 824
rect 1142 810 1158 824
rect 1169 823 1172 830
rect 1169 818 1174 823
rect 1168 816 1169 818
rect 1172 816 1174 818
rect 1199 816 1215 839
rect 1222 830 1229 838
rect 1265 830 1268 839
rect 1316 835 1327 839
rect 1316 831 1321 835
rect 1229 824 1232 830
rect 1268 828 1269 830
rect 1220 816 1236 824
rect 1164 813 1167 815
rect 1116 808 1159 810
rect 1174 808 1178 816
rect 1198 814 1199 816
rect 1108 807 1119 808
rect 1133 807 1135 808
rect 1159 807 1178 808
rect 1012 799 1034 805
rect 1012 798 1028 799
rect 1008 792 1028 798
rect 1034 793 1040 799
rect 1008 789 1015 792
rect 1019 789 1028 792
rect 1062 792 1078 807
rect 1086 799 1092 805
rect 1080 793 1086 799
rect 1062 790 1063 792
rect 967 780 982 789
rect 1012 788 1028 789
rect 916 774 982 780
rect 1007 778 1028 788
rect 1057 787 1059 790
rect 1062 787 1078 790
rect 1051 778 1053 787
rect 1007 776 1053 778
rect 1057 776 1078 787
rect 1095 785 1116 807
rect 1136 803 1137 805
rect 1150 800 1155 804
rect 1138 795 1139 797
rect 1159 795 1174 807
rect 1194 806 1198 813
rect 1220 812 1241 816
rect 1269 813 1274 828
rect 1307 817 1316 831
rect 1325 828 1327 835
rect 1320 818 1321 828
rect 1307 816 1320 817
rect 1304 815 1307 816
rect 1289 814 1301 815
rect 1287 813 1289 814
rect 1265 812 1279 813
rect 1220 810 1265 812
rect 1220 808 1241 810
rect 1269 808 1274 812
rect 1178 801 1180 805
rect 1189 800 1194 806
rect 1185 795 1188 799
rect 1129 787 1145 795
rect 1159 792 1185 795
rect 1204 792 1220 808
rect 1236 806 1241 808
rect 1313 806 1320 816
rect 1325 809 1326 828
rect 1325 806 1328 809
rect 1357 807 1359 839
rect 1492 836 1494 841
rect 1522 836 1523 841
rect 1552 839 1576 841
rect 1313 805 1321 806
rect 1349 805 1359 807
rect 1363 805 1371 817
rect 1412 815 1428 824
rect 1430 815 1446 824
rect 1412 814 1446 815
rect 1494 814 1496 836
rect 1523 824 1529 836
rect 1554 830 1568 839
rect 1636 836 1638 842
rect 1661 841 1665 854
rect 1660 836 1665 841
rect 1653 834 1665 836
rect 1677 860 1705 861
rect 1677 855 1704 860
rect 1568 825 1572 830
rect 1412 813 1447 814
rect 1410 811 1412 813
rect 1445 812 1446 813
rect 1410 808 1446 811
rect 1508 809 1542 824
rect 1572 815 1576 825
rect 1576 809 1578 814
rect 1638 809 1639 825
rect 1505 808 1542 809
rect 1578 808 1579 809
rect 1241 801 1243 805
rect 1274 800 1276 805
rect 1321 802 1325 805
rect 1325 801 1349 802
rect 1357 801 1359 805
rect 1396 801 1422 808
rect 1432 801 1444 808
rect 1276 797 1277 800
rect 1245 795 1246 797
rect 1173 790 1185 792
rect 1246 791 1249 795
rect 1012 774 1023 776
rect 1058 774 1078 776
rect 740 766 805 772
rect 817 768 827 774
rect 829 771 863 774
rect 866 771 870 774
rect 829 768 870 771
rect 740 758 799 766
rect 825 764 827 768
rect 836 764 852 768
rect 680 753 683 756
rect 686 753 689 754
rect 634 744 689 753
rect 747 749 799 758
rect 829 758 852 764
rect 854 758 870 768
rect 932 761 948 774
rect 829 756 841 758
rect 846 755 852 758
rect 904 755 910 761
rect 929 758 948 761
rect 950 758 966 774
rect 1028 772 1044 774
rect 1046 772 1062 774
rect 981 761 987 767
rect 1019 764 1062 772
rect 1092 768 1096 785
rect 1129 780 1146 787
rect 1116 768 1122 773
rect 1142 772 1146 780
rect 1159 780 1189 790
rect 1159 774 1174 780
rect 1185 779 1189 780
rect 1168 773 1173 774
rect 1146 771 1147 772
rect 929 755 935 758
rect 987 755 993 761
rect 1028 758 1044 764
rect 1046 758 1062 764
rect 852 749 858 755
rect 898 749 904 755
rect 931 754 935 755
rect 1090 754 1096 768
rect 1138 767 1159 771
rect 1163 767 1168 773
rect 1104 757 1106 758
rect 1103 755 1104 757
rect 928 750 932 754
rect 1099 752 1103 755
rect 1138 753 1163 767
rect 1189 763 1200 779
rect 1204 774 1220 790
rect 1249 779 1254 790
rect 1254 776 1262 779
rect 1277 778 1293 797
rect 1325 793 1337 801
rect 1347 793 1359 801
rect 1390 797 1412 801
rect 1436 797 1442 801
rect 1390 795 1444 797
rect 1446 795 1462 808
rect 1492 795 1505 808
rect 1523 806 1529 808
rect 1529 802 1530 806
rect 1355 778 1359 793
rect 1384 789 1412 795
rect 1277 776 1315 778
rect 1254 775 1293 776
rect 1254 774 1270 775
rect 1200 754 1206 763
rect 1220 758 1236 774
rect 1238 763 1262 774
rect 1277 764 1293 775
rect 1300 775 1315 776
rect 1300 774 1316 775
rect 1316 763 1318 774
rect 1355 763 1357 778
rect 1238 758 1254 763
rect 1262 753 1267 763
rect 1293 754 1298 763
rect 1316 758 1321 763
rect 1356 761 1357 763
rect 1390 774 1412 789
rect 1442 792 1462 795
rect 1442 790 1456 792
rect 1442 789 1462 790
rect 1442 781 1444 789
rect 1443 774 1444 781
rect 1446 774 1462 789
rect 1485 784 1495 795
rect 1497 787 1498 795
rect 1530 786 1533 800
rect 1542 792 1558 808
rect 1483 780 1485 784
rect 1498 782 1499 786
rect 1533 781 1534 786
rect 1481 774 1483 780
rect 1534 778 1535 781
rect 1535 774 1537 778
rect 1542 774 1558 790
rect 1579 786 1587 808
rect 1653 806 1660 834
rect 1677 826 1698 855
rect 1652 802 1653 806
rect 1665 803 1674 812
rect 1677 808 1688 826
rect 1714 824 1724 847
rect 1700 818 1734 824
rect 2196 819 2197 1015
rect 2386 819 2387 1015
rect 2472 819 2473 1015
rect 2745 819 2746 1015
rect 2942 819 2943 1015
rect 1700 812 1716 818
rect 1718 812 1734 818
rect 1700 809 1734 812
rect 1700 808 1746 809
rect 1649 790 1652 800
rect 1656 794 1665 803
rect 1677 792 1700 808
rect 1712 803 1721 808
rect 1746 805 1751 808
rect 1721 794 1730 803
rect 1639 787 1654 790
rect 1587 779 1593 786
rect 1612 780 1654 787
rect 1660 786 1664 792
rect 1677 790 1687 792
rect 1677 787 1700 790
rect 1656 780 1658 784
rect 1677 781 1714 787
rect 1588 774 1604 779
rect 1612 774 1656 780
rect 1684 774 1714 781
rect 1751 774 1767 805
rect 1390 761 1446 774
rect 1448 763 1456 774
rect 1478 763 1481 774
rect 1499 764 1500 770
rect 1318 753 1321 758
rect 1357 758 1446 761
rect 1477 760 1480 763
rect 1531 760 1542 774
rect 747 745 806 749
rect 928 746 935 750
rect 1089 748 1099 752
rect 1136 749 1138 753
rect 967 746 1064 748
rect 1087 746 1099 748
rect 1135 746 1136 748
rect 927 745 935 746
rect 938 745 1073 746
rect 1084 745 1086 746
rect 1089 745 1099 746
rect 634 741 686 744
rect 689 742 690 744
rect 628 736 692 741
rect 747 740 886 745
rect 927 744 1099 745
rect 628 735 694 736
rect 549 730 555 731
rect 470 727 572 730
rect 470 726 588 727
rect 186 713 187 726
rect 224 717 226 726
rect 470 724 530 726
rect 549 725 555 726
rect 606 725 613 731
rect 634 729 640 735
rect 649 727 652 732
rect 680 729 686 735
rect 691 727 694 735
rect 653 725 654 727
rect 694 725 695 727
rect 747 726 755 740
rect 799 736 886 740
rect 801 730 886 736
rect 919 743 1099 744
rect 1131 743 1135 745
rect 1145 744 1163 753
rect 1267 750 1269 753
rect 1298 750 1300 753
rect 1168 744 1208 745
rect 1209 744 1220 750
rect 919 740 1096 743
rect 919 732 933 740
rect 1131 735 1145 743
rect 808 729 809 730
rect 809 727 810 729
rect 470 720 519 724
rect 470 717 526 720
rect 555 719 561 725
rect 470 713 479 717
rect 226 711 227 713
rect 489 712 491 717
rect 519 710 526 717
rect 185 707 186 710
rect 370 709 450 710
rect 370 707 445 709
rect 491 696 494 709
rect 526 708 536 709
rect 504 700 516 708
rect 526 700 538 708
rect 495 696 500 700
rect 502 698 547 700
rect 526 696 536 698
rect 541 697 547 698
rect 573 697 575 722
rect 601 719 607 725
rect 654 723 655 725
rect 695 720 696 722
rect 741 720 757 726
rect 657 715 659 719
rect 696 716 697 719
rect 743 716 757 720
rect 761 716 764 719
rect 787 718 789 726
rect 799 720 805 726
rect 886 725 895 730
rect 811 723 812 725
rect 786 716 789 718
rect 793 716 801 720
rect 659 709 663 715
rect 697 710 699 715
rect 743 714 753 716
rect 743 713 752 714
rect 755 713 776 716
rect 786 713 788 716
rect 791 713 801 716
rect 752 710 753 713
rect 764 710 767 713
rect 780 711 789 713
rect 791 711 793 713
rect 776 710 791 711
rect 812 710 819 722
rect 895 713 900 724
rect 927 722 933 732
rect 1056 723 1062 729
rect 1072 727 1078 732
rect 1067 723 1072 727
rect 1102 723 1108 729
rect 1128 727 1131 735
rect 1132 727 1145 735
rect 1128 725 1132 727
rect 1153 726 1161 744
rect 1168 740 1220 744
rect 1166 735 1202 740
rect 1208 737 1220 740
rect 1269 747 1272 750
rect 1208 735 1225 737
rect 1166 731 1168 735
rect 1209 734 1225 735
rect 1269 734 1274 747
rect 1219 731 1225 734
rect 1220 730 1225 731
rect 1223 729 1227 730
rect 1272 729 1274 734
rect 1225 726 1229 729
rect 919 719 933 722
rect 919 716 935 719
rect 987 716 988 719
rect 1050 717 1056 723
rect 1108 717 1114 723
rect 1124 722 1128 724
rect 1129 723 1132 725
rect 1155 724 1156 726
rect 1227 725 1229 726
rect 1273 725 1274 729
rect 1161 724 1162 725
rect 664 698 670 708
rect 700 698 702 708
rect 755 701 767 710
rect 768 698 774 708
rect 777 701 789 710
rect 791 709 856 710
rect 798 707 856 709
rect 805 706 856 707
rect 813 703 856 706
rect 819 700 825 703
rect 827 702 856 703
rect 828 701 856 702
rect 819 698 833 700
rect 670 697 674 698
rect 541 696 674 697
rect 184 692 185 696
rect 491 695 500 696
rect 492 694 500 695
rect 504 694 674 696
rect 702 694 706 698
rect 189 690 190 692
rect 187 676 190 690
rect 184 670 187 676
rect 177 663 187 670
rect 189 663 190 676
rect 222 687 223 692
rect 224 687 249 692
rect 489 688 495 694
rect 222 673 253 687
rect 492 684 495 688
rect 504 692 600 694
rect 504 690 564 692
rect 504 688 553 690
rect 504 683 538 688
rect 504 679 513 683
rect 404 673 438 676
rect 222 663 223 673
rect 228 663 235 670
rect 177 658 235 663
rect 252 660 253 673
rect 183 657 228 658
rect 183 653 184 657
rect 187 654 225 657
rect 189 646 201 654
rect 211 646 223 654
rect 183 630 192 644
rect 262 642 263 671
rect 545 663 547 688
rect 573 663 575 692
rect 600 690 632 692
rect 670 691 729 694
rect 670 690 674 691
rect 702 690 706 691
rect 729 690 733 691
rect 774 690 775 696
rect 825 695 833 698
rect 835 697 856 701
rect 897 709 901 713
rect 919 712 937 716
rect 962 712 965 713
rect 919 711 935 712
rect 919 710 933 711
rect 940 710 965 712
rect 980 710 982 712
rect 987 710 993 715
rect 1041 710 1056 716
rect 1123 715 1128 722
rect 1116 711 1122 714
rect 1124 711 1128 715
rect 1150 716 1167 724
rect 927 709 935 710
rect 938 709 941 710
rect 946 709 1048 710
rect 897 706 903 709
rect 927 707 933 709
rect 968 707 1048 709
rect 930 706 1048 707
rect 1116 709 1124 711
rect 1116 706 1122 709
rect 1150 708 1172 716
rect 1164 706 1172 708
rect 1183 706 1189 712
rect 897 702 904 706
rect 897 701 905 702
rect 868 698 878 699
rect 897 698 907 701
rect 930 698 943 706
rect 981 703 987 706
rect 992 705 1061 706
rect 1108 705 1116 706
rect 992 703 1116 705
rect 992 700 1029 703
rect 861 697 865 698
rect 879 697 907 698
rect 843 695 861 697
rect 819 694 861 695
rect 825 692 856 694
rect 825 691 844 692
rect 822 690 830 691
rect 636 688 639 690
rect 675 687 676 690
rect 733 688 737 690
rect 815 688 822 690
rect 676 678 682 687
rect 709 678 716 687
rect 725 685 748 688
rect 806 687 815 688
rect 725 684 750 685
rect 725 683 771 684
rect 775 683 777 687
rect 801 685 806 687
rect 798 684 801 685
rect 796 683 798 684
rect 725 682 796 683
rect 833 682 842 691
rect 849 690 856 692
rect 879 691 910 697
rect 928 691 930 698
rect 992 691 1025 700
rect 1108 695 1116 703
rect 1150 693 1172 706
rect 1177 700 1183 706
rect 1223 700 1225 725
rect 1227 713 1237 725
rect 1273 719 1279 725
rect 1300 719 1315 750
rect 1321 749 1322 753
rect 1357 751 1444 758
rect 1472 753 1478 760
rect 1522 758 1542 760
rect 1604 758 1620 774
rect 1622 770 1638 774
rect 1640 771 1647 774
rect 1651 773 1656 774
rect 1640 770 1646 771
rect 1649 770 1651 773
rect 1686 770 1692 774
rect 1622 764 1640 770
rect 1692 764 1698 770
rect 1622 758 1638 764
rect 1700 760 1714 774
rect 1767 761 1775 774
rect 1700 758 1717 760
rect 1522 753 1531 758
rect 1539 755 1540 757
rect 1711 753 1717 758
rect 1357 749 1442 751
rect 1467 750 1480 753
rect 1322 746 1323 748
rect 1357 745 1448 749
rect 1460 748 1480 750
rect 1516 748 1522 753
rect 1460 746 1478 748
rect 1515 746 1516 748
rect 1464 745 1478 746
rect 1323 735 1325 744
rect 1376 743 1478 745
rect 1376 740 1408 743
rect 1424 740 1478 743
rect 1325 732 1326 735
rect 1326 730 1327 731
rect 1327 726 1328 730
rect 1376 729 1478 740
rect 1501 732 1503 743
rect 1510 740 1515 746
rect 1540 742 1543 753
rect 1507 736 1510 740
rect 1506 735 1507 736
rect 1504 732 1506 735
rect 1499 730 1504 732
rect 1387 727 1391 729
rect 1428 728 1432 729
rect 1386 725 1391 727
rect 1427 725 1428 727
rect 1489 725 1499 730
rect 1319 719 1325 725
rect 1328 721 1332 724
rect 1385 722 1391 725
rect 1447 724 1499 725
rect 1384 721 1391 722
rect 1425 721 1426 722
rect 1447 721 1489 724
rect 1267 713 1273 719
rect 1325 713 1331 719
rect 1332 717 1431 721
rect 1447 717 1482 721
rect 1501 720 1503 730
rect 1543 724 1544 742
rect 1646 740 1672 753
rect 1675 748 1680 753
rect 1717 748 1720 753
rect 1721 748 1730 756
rect 1747 753 1759 761
rect 1767 756 1781 761
rect 1769 753 1781 756
rect 1743 750 1744 752
rect 1775 749 1781 753
rect 1675 747 1681 748
rect 1720 747 1730 748
rect 1675 740 1680 747
rect 1711 746 1722 747
rect 1735 746 1743 749
rect 1747 747 1781 749
rect 1778 746 1781 747
rect 1681 740 1682 746
rect 1544 719 1547 724
rect 1500 717 1501 719
rect 1634 718 1640 731
rect 1645 724 1646 730
rect 1682 726 1684 740
rect 1711 738 1721 746
rect 1722 740 1727 746
rect 1728 740 1741 746
rect 1708 732 1711 738
rect 1705 727 1708 732
rect 1646 722 1648 724
rect 1646 721 1650 722
rect 1678 721 1680 724
rect 1646 719 1680 721
rect 1684 719 1686 726
rect 1704 725 1705 727
rect 1727 726 1741 740
rect 1692 722 1698 724
rect 1692 719 1702 722
rect 1728 720 1745 726
rect 1672 718 1702 719
rect 1227 712 1229 713
rect 1227 707 1235 712
rect 1332 707 1473 717
rect 1474 712 1482 717
rect 1640 716 1646 718
rect 1682 717 1692 718
rect 1682 716 1684 717
rect 1553 715 1555 716
rect 1640 715 1684 716
rect 1496 712 1498 715
rect 1229 706 1235 707
rect 1229 700 1241 706
rect 852 687 856 690
rect 854 685 856 687
rect 855 683 856 685
rect 897 690 910 691
rect 897 687 911 690
rect 897 683 919 687
rect 775 678 777 682
rect 639 673 640 676
rect 637 668 640 673
rect 682 671 686 678
rect 716 671 721 678
rect 855 677 859 683
rect 897 679 916 683
rect 919 682 921 683
rect 924 682 928 690
rect 995 686 1015 691
rect 989 683 1015 686
rect 988 682 1015 683
rect 1025 682 1034 691
rect 1150 690 1167 693
rect 1172 691 1173 693
rect 1174 689 1178 690
rect 1229 689 1235 700
rect 1257 698 1266 700
rect 1257 691 1270 698
rect 1166 687 1178 689
rect 1227 688 1235 689
rect 1223 687 1227 688
rect 1166 685 1181 687
rect 1212 685 1223 687
rect 1166 683 1201 685
rect 1205 683 1212 685
rect 921 681 928 682
rect 975 681 1015 682
rect 921 680 957 681
rect 975 680 987 681
rect 924 679 945 680
rect 966 679 998 680
rect 897 678 994 679
rect 897 677 916 678
rect 788 675 798 676
rect 859 675 860 676
rect 916 675 918 676
rect 801 674 809 675
rect 806 671 820 674
rect 686 668 688 671
rect 630 667 640 668
rect 658 667 669 668
rect 613 664 630 667
rect 602 663 613 664
rect 495 662 613 663
rect 637 662 640 667
rect 669 666 690 667
rect 669 664 692 666
rect 689 663 704 664
rect 724 663 729 668
rect 820 667 822 671
rect 836 664 847 667
rect 831 663 836 664
rect 689 662 836 663
rect 495 659 602 662
rect 495 657 581 659
rect 636 657 637 660
rect 495 656 569 657
rect 495 655 565 656
rect 495 654 558 655
rect 495 653 553 654
rect 495 648 547 653
rect 489 642 553 648
rect 192 626 196 630
rect 252 626 268 642
rect 495 636 501 642
rect 511 638 517 642
rect 517 634 522 638
rect 541 636 547 642
rect 573 634 575 657
rect 632 642 636 657
rect 692 655 696 660
rect 704 659 831 662
rect 860 660 867 675
rect 917 671 920 675
rect 924 674 928 678
rect 1050 675 1056 677
rect 1028 674 1056 675
rect 923 672 924 674
rect 1021 672 1029 674
rect 1050 671 1058 674
rect 1108 671 1114 677
rect 1166 674 1182 683
rect 906 668 923 671
rect 874 664 888 667
rect 888 663 894 664
rect 901 663 921 668
rect 1056 665 1062 671
rect 1102 665 1108 671
rect 1010 663 1013 664
rect 1229 663 1235 688
rect 1248 682 1263 691
rect 1376 689 1382 707
rect 1409 706 1424 707
rect 1409 705 1438 706
rect 888 662 1013 663
rect 894 660 1010 662
rect 1183 660 1235 663
rect 730 657 819 659
rect 730 654 734 657
rect 747 656 812 657
rect 751 655 809 656
rect 761 654 803 655
rect 696 652 697 654
rect 734 652 735 654
rect 767 653 803 654
rect 697 649 699 652
rect 700 642 705 648
rect 735 642 744 652
rect 777 644 778 646
rect 768 642 783 644
rect 632 634 646 642
rect 744 639 746 642
rect 768 639 784 642
rect 746 637 747 639
rect 768 637 795 639
rect 522 632 589 634
rect 196 624 252 626
rect 236 610 252 624
rect 573 614 575 632
rect 580 630 592 632
rect 631 630 646 634
rect 748 633 751 637
rect 768 635 777 637
rect 781 635 826 637
rect 833 635 842 644
rect 867 642 884 660
rect 901 659 1010 660
rect 904 657 1002 659
rect 904 655 910 657
rect 915 656 997 657
rect 917 655 997 656
rect 919 652 991 655
rect 1177 654 1241 660
rect 898 650 901 652
rect 919 651 978 652
rect 919 650 934 651
rect 944 650 950 651
rect 891 645 897 649
rect 919 645 942 650
rect 953 645 972 650
rect 1183 648 1189 654
rect 1198 652 1199 654
rect 1199 650 1200 652
rect 919 644 939 645
rect 919 642 921 644
rect 923 642 939 644
rect 963 642 972 645
rect 1200 644 1202 649
rect 1229 648 1235 654
rect 867 639 888 642
rect 580 626 596 630
rect 630 626 646 630
rect 596 610 612 626
rect 614 610 630 626
rect 714 615 731 633
rect 749 625 771 633
rect 777 626 786 635
rect 824 626 833 635
rect 867 630 884 639
rect 919 634 934 642
rect 960 635 972 642
rect 1025 635 1034 644
rect 1229 643 1232 648
rect 1257 645 1263 682
rect 1283 677 1286 683
rect 1319 676 1321 683
rect 1267 667 1273 673
rect 1274 667 1283 676
rect 1273 663 1283 667
rect 1287 663 1289 673
rect 1319 671 1322 676
rect 1371 674 1376 689
rect 1318 667 1322 671
rect 1325 667 1331 673
rect 1409 672 1424 705
rect 1455 704 1459 705
rect 1479 694 1489 705
rect 1555 694 1623 715
rect 1640 712 1658 715
rect 1645 708 1658 712
rect 1646 707 1658 708
rect 1686 712 1692 717
rect 1725 715 1727 718
rect 1738 716 1745 720
rect 1745 715 1747 716
rect 1779 715 1781 746
rect 1785 737 1793 749
rect 1785 715 1793 727
rect 1470 689 1481 691
rect 1470 688 1479 689
rect 1470 687 1480 688
rect 1483 687 1484 690
rect 1486 688 1495 691
rect 1516 690 1518 691
rect 1623 688 1643 694
rect 1646 691 1648 706
rect 1686 694 1691 712
rect 1708 696 1725 714
rect 1782 711 1785 713
rect 1775 710 1782 711
rect 1769 708 1781 710
rect 1758 703 1781 708
rect 1758 696 1769 703
rect 1702 694 1720 696
rect 1648 688 1650 691
rect 1679 690 1720 694
rect 1679 688 1702 690
rect 1616 687 1710 688
rect 1467 685 1480 687
rect 1464 683 1467 685
rect 1453 677 1464 683
rect 1470 679 1478 685
rect 1369 667 1371 671
rect 1318 663 1325 667
rect 1273 661 1325 663
rect 1274 660 1333 661
rect 1257 644 1265 645
rect 1203 637 1205 641
rect 1229 637 1239 643
rect 1248 642 1265 644
rect 1273 642 1274 659
rect 1275 649 1333 660
rect 1366 655 1369 667
rect 1365 652 1366 654
rect 1402 652 1409 672
rect 1449 668 1453 676
rect 1470 663 1478 669
rect 1482 663 1484 687
rect 1648 676 1650 687
rect 1686 682 1691 687
rect 1732 676 1742 680
rect 1552 672 1572 673
rect 1536 664 1552 672
rect 1572 664 1624 672
rect 1532 663 1536 664
rect 1470 662 1536 663
rect 1624 663 1638 664
rect 1650 663 1652 676
rect 1726 674 1732 676
rect 1695 664 1726 674
rect 1686 663 1695 664
rect 1624 662 1695 663
rect 1283 648 1325 649
rect 1283 645 1324 648
rect 1229 635 1236 637
rect 1248 635 1274 642
rect 1287 637 1299 645
rect 1309 644 1321 645
rect 1322 644 1324 645
rect 1309 641 1324 644
rect 1362 643 1364 647
rect 1400 645 1402 651
rect 1399 643 1400 645
rect 1359 641 1362 643
rect 1306 639 1324 641
rect 1309 637 1324 639
rect 1354 637 1359 641
rect 1311 636 1324 637
rect 1301 635 1307 636
rect 1313 635 1324 636
rect 866 626 884 630
rect 897 626 934 634
rect 969 626 978 635
rect 1016 626 1025 635
rect 866 625 872 626
rect 749 621 764 625
rect 861 621 866 625
rect 749 618 771 621
rect 857 618 861 621
rect 749 615 772 618
rect 853 615 857 618
rect 897 615 921 626
rect 1206 615 1213 634
rect 1229 629 1239 635
rect 731 614 772 615
rect 731 609 786 614
rect 847 610 852 614
rect 891 610 897 615
rect 902 610 918 615
rect 1213 610 1217 615
rect 1229 614 1253 629
rect 1257 626 1274 635
rect 1304 626 1313 635
rect 1318 626 1319 635
rect 1322 624 1324 635
rect 1334 635 1354 637
rect 1396 635 1399 643
rect 1447 642 1449 660
rect 1470 657 1531 662
rect 1638 661 1695 662
rect 1650 660 1652 661
rect 1478 656 1531 657
rect 1478 655 1520 656
rect 1480 653 1518 655
rect 1482 645 1494 653
rect 1504 645 1516 653
rect 1334 632 1351 635
rect 1329 627 1351 632
rect 1391 628 1396 635
rect 1389 627 1391 628
rect 1329 625 1341 627
rect 1304 622 1322 624
rect 1273 620 1308 622
rect 1328 620 1341 625
rect 1229 612 1257 614
rect 1229 611 1271 612
rect 1274 611 1290 620
rect 1292 614 1308 620
rect 1310 615 1341 620
rect 1372 616 1389 627
rect 1444 626 1449 642
rect 1518 626 1519 631
rect 1636 626 1652 642
rect 1691 630 1702 642
rect 1689 626 1702 630
rect 1512 619 1518 625
rect 1322 614 1341 615
rect 1291 612 1341 614
rect 1292 611 1341 612
rect 826 609 847 610
rect 1229 609 1341 611
rect 1363 610 1372 616
rect 1447 615 1454 619
rect 1510 616 1512 619
rect 1507 615 1510 616
rect 1454 614 1507 615
rect 1460 610 1476 614
rect 1652 610 1668 626
rect 1670 610 1686 626
rect 2405 623 2432 629
rect 2433 623 2460 624
rect 731 607 861 609
rect 731 606 751 607
rect 871 606 890 609
rect 1218 607 1341 609
rect 212 557 262 606
rect 292 557 358 606
rect 388 557 454 606
rect 484 557 550 606
rect 580 557 646 606
rect 676 594 751 606
rect 676 557 742 594
rect 751 588 758 594
rect 758 586 767 588
rect 772 585 838 606
rect 868 594 918 606
rect 865 589 918 594
rect 861 586 864 588
rect 767 584 838 585
rect 859 584 861 585
rect 772 557 838 584
rect 852 581 858 584
rect 868 557 918 589
rect 980 557 1030 606
rect 1060 557 1126 606
rect 1156 557 1206 606
rect 1218 594 1234 607
rect 1344 598 1362 610
rect 1229 593 1232 594
rect 1234 589 1240 594
rect 1240 586 1243 588
rect 1323 586 1344 598
rect 1345 596 1356 598
rect 1243 585 1247 586
rect 1247 584 1294 585
rect 1314 584 1319 585
rect 1364 557 1414 606
rect 1444 557 1510 606
rect 1540 557 1606 606
rect 1636 557 1702 606
rect 1732 557 1782 606
rect 2976 481 2977 487
rect 2942 441 2977 475
rect 2988 463 2989 475
rect 2988 441 2989 453
rect 2185 429 2186 440
rect 2375 429 2376 440
rect 2461 429 2462 440
rect 2734 429 2735 440
rect 2931 429 2932 440
rect 2965 429 2977 435
rect 2196 389 2197 429
rect 2386 389 2387 429
rect 2472 389 2473 429
rect 2745 389 2746 429
rect 2942 389 2943 429
<< nwell >>
rect 2941 1749 2977 1750
rect 0 1748 2977 1749
rect 2978 1748 3052 1749
rect 0 1087 3052 1748
rect 0 820 109 1087
rect 1860 1086 2086 1087
rect 1862 744 2076 1086
rect 2097 800 2165 870
rect 2858 772 2888 807
rect 3007 744 3052 1087
<< ndiff >>
rect 2943 441 2977 475
<< locali >>
rect 0 2173 3052 2493
rect 0 1087 3052 1407
rect 1860 1086 2086 1087
rect 3016 1086 3052 1087
rect 255 805 264 810
rect 297 805 311 810
rect 303 774 311 805
rect 533 796 587 808
rect 532 789 587 796
rect 527 782 587 789
rect 523 776 587 782
rect 523 775 588 776
rect 522 774 588 775
rect 303 773 312 774
rect 257 771 312 773
rect 520 771 588 774
rect 257 770 313 771
rect 519 770 588 771
rect 257 766 314 770
rect 516 766 588 770
rect 257 763 315 766
rect 513 763 588 766
rect 257 759 316 763
rect 257 754 321 759
rect 509 757 588 763
rect 506 755 588 757
rect 257 753 326 754
rect 257 749 342 753
rect 502 752 588 755
rect 499 749 588 752
rect 257 748 345 749
rect 257 746 368 748
rect 492 747 588 749
rect 257 744 376 746
rect 473 745 588 747
rect 257 743 383 744
rect 414 743 588 745
rect 257 726 588 743
rect 257 724 530 726
rect 257 717 519 724
rect 257 713 479 717
rect 257 711 461 713
rect 257 710 453 711
rect 257 709 450 710
rect 257 707 445 709
rect 420 555 459 578
rect 787 555 826 572
rect 1155 555 1194 578
rect 1525 555 1565 576
rect 1859 555 1898 576
rect 182 544 1898 555
rect 150 320 1898 544
rect 0 0 3052 320
<< viali >>
rect 2943 1722 2977 1756
rect 2944 1462 2978 1496
rect 2943 997 2977 1031
rect 2943 441 2977 475
<< metal1 >>
rect 0 2173 3052 2493
rect 1139 1721 1173 2173
rect 1240 1934 1314 1943
rect 1240 1878 1249 1934
rect 1305 1878 1314 1934
rect 2421 1909 2705 1916
rect 2433 1903 2705 1909
rect 1240 1869 1314 1878
rect 2387 1882 2705 1903
rect 2387 1869 2433 1882
rect 2466 1847 2531 1854
rect 2466 1829 2473 1847
rect 1310 1795 2473 1829
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2096 1694 2164 1700
rect 2096 1681 2102 1694
rect 1020 1647 2102 1681
rect 2096 1636 2102 1647
rect 2160 1636 2164 1694
rect 2671 1646 2705 1882
rect 2780 1723 2903 1755
rect 2780 1722 2812 1723
rect 2870 1688 2903 1723
rect 2870 1687 2904 1688
rect 2872 1647 2904 1687
rect 2096 1630 2164 1636
rect 2926 1450 2932 1508
rect 2990 1450 2996 1508
rect 1484 1406 1528 1407
rect 1 1086 3053 1406
rect 2925 985 2931 1043
rect 2989 985 2995 1043
rect 1705 806 1769 870
rect 1985 864 2053 870
rect 1985 806 1991 864
rect 2049 806 2053 864
rect 1985 800 2053 806
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2672 819 2706 846
rect 2672 812 2707 819
rect 2673 809 2707 812
rect 2097 800 2165 806
rect 2672 806 2707 809
rect 527 786 587 789
rect 527 782 596 786
rect 523 728 596 782
rect 523 726 587 728
rect 2003 698 2037 800
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 2300 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2461 716 2531 722
rect 2461 698 2467 716
rect 2003 664 2467 698
rect 2461 658 2467 664
rect 2525 658 2531 716
rect 2461 652 2531 658
rect 2672 624 2705 806
rect 2850 801 2914 852
rect 2850 772 2888 801
rect 2779 738 2888 772
rect 2387 623 2421 624
rect 2433 623 2705 624
rect 2387 590 2705 623
rect 420 555 459 578
rect 787 555 826 572
rect 1155 555 1194 578
rect 1859 576 1884 584
rect 1525 568 1565 576
rect 1859 555 1898 576
rect 182 544 1898 555
rect 150 513 1898 544
rect 150 457 562 513
rect 618 457 1898 513
rect 150 320 1898 457
rect 0 0 3052 320
<< via1 >>
rect 1249 1878 1305 1934
rect 2473 1795 2525 1847
rect 2312 1709 2364 1767
rect 2102 1636 2160 1694
rect 2932 1496 2990 1508
rect 2932 1462 2944 1496
rect 2944 1462 2978 1496
rect 2978 1462 2990 1496
rect 2932 1450 2990 1462
rect 2931 1031 2989 1043
rect 2931 997 2943 1031
rect 2943 997 2977 1031
rect 2977 997 2989 1031
rect 2931 985 2989 997
rect 1991 806 2049 864
rect 2103 806 2161 864
rect 2312 738 2364 790
rect 2467 658 2525 716
rect 562 457 618 513
<< metal2 >>
rect 1240 1934 1314 1943
rect 1240 1878 1249 1934
rect 1305 1878 1314 1934
rect 1240 1869 1314 1878
rect 2466 1847 2531 1854
rect 2466 1841 2473 1847
rect 2243 1807 2473 1841
rect 2096 1694 2164 1700
rect 2096 1636 2102 1694
rect 2160 1636 2164 1694
rect 2096 1630 2164 1636
rect 2112 870 2147 1630
rect 1976 864 2053 870
rect 1976 853 1985 864
rect 1974 813 1985 853
rect 1976 806 1985 813
rect 2049 806 2053 864
rect 1976 800 2053 806
rect 2097 864 2165 870
rect 2097 806 2103 864
rect 2161 806 2165 864
rect 2097 800 2165 806
rect 2003 799 2037 800
rect 592 777 598 789
rect 2243 772 2275 1807
rect 2466 1795 2473 1807
rect 2525 1795 2531 1847
rect 2466 1789 2531 1795
rect 2306 1709 2312 1767
rect 2364 1709 2370 1767
rect 2306 1702 2370 1709
rect 2312 1667 2346 1702
rect 2312 1632 2347 1667
rect 2312 1597 2507 1632
rect 2306 790 2370 796
rect 2306 772 2312 790
rect 573 522 606 737
rect 1675 727 1693 767
rect 2243 738 2312 772
rect 2364 738 2370 790
rect 2306 732 2370 738
rect 2472 722 2507 1597
rect 2923 1508 2999 1517
rect 2923 1450 2932 1508
rect 2990 1450 2999 1508
rect 2923 1441 2999 1450
rect 2922 1043 2998 1052
rect 2922 985 2931 1043
rect 2989 985 2998 1043
rect 2922 976 2998 985
rect 2461 716 2531 722
rect 2461 658 2467 716
rect 2525 658 2531 716
rect 2461 652 2531 658
rect 553 513 627 522
rect 553 457 562 513
rect 618 457 627 513
rect 553 448 627 457
<< via2 >>
rect 1249 1878 1305 1934
rect 1985 806 1991 864
rect 1991 806 2043 864
rect 2932 1450 2990 1508
rect 2931 985 2989 1043
<< metal3 >>
rect 1240 1934 1314 1943
rect 1240 1878 1249 1934
rect 1305 1878 1314 1934
rect 1240 1869 1314 1878
rect 1247 1372 1307 1869
rect 2923 1508 2999 2493
rect 2923 1450 2932 1508
rect 2990 1450 2999 1508
rect 2923 1441 2999 1450
rect 409 1305 1307 1372
rect 409 1087 470 1305
rect 1037 1113 1307 1305
rect 409 746 469 1087
rect 772 515 838 657
rect 1045 631 1105 1113
rect 2922 1043 2998 1052
rect 2922 985 2931 1043
rect 2989 985 2998 1043
rect 1973 864 2053 871
rect 1973 806 1985 864
rect 2043 806 2053 864
rect 1973 794 2053 806
rect 1974 515 2040 794
rect 772 449 2040 515
rect 2922 0 2998 985
use scs130hd_mpr2ya_8  scs130hd_mpr2ya_8_0
timestamp 1696006315
transform 1 0 150 0 1 559
box -48 -48 1796 592
use sky130_osu_sc_12T_hs__fill_2  sky130_osu_sc_12T_hs__fill_2_0
timestamp 1604095901
transform 1 0 1513 0 -1 2234
box -7 0 161 1341
use sky130_osu_sc_12T_hs__fill_8  sky130_osu_sc_12T_hs__fill_8_0
timestamp 1604095905
transform 1 0 1684 0 -1 2234
box -9 0 179 897
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1706264206
transform 1 0 2625 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1706264206
transform 1 0 2822 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1706264206
transform 1 0 2823 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1706264206
transform 1 0 2625 0 -1 2234
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 2076 0 1 259
box -8 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1698882961
transform 1 0 949 0 -1 2234
box -8 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1698882961
transform 1 0 2076 0 -1 2234
box -8 0 552 902
<< labels >>
rlabel metal1 36 290 36 290 1 vssd1
port 5 n
rlabel metal2 2128 836 2128 836 1 sel
port 7 n
rlabel metal1 31 2204 31 2204 1 vssd1
port 5 n
rlabel metal1 1310 1795 1332 1829 1 in
port 10 n
rlabel metal1 46 1146 46 1146 1 vccd1
port 6 n
rlabel viali 2943 441 2977 475 1 Y1
port 9 n
rlabel viali 2943 1722 2977 1756 1 Y0
port 8 n
<< end >>
