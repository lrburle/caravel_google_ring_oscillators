magic
tech sky130A
magscale 1 2
timestamp 1714057206
<< nwell >>
rect -48 260 1796 582
<< pwell >>
rect 76 -16 110 16
<< nmos >>
rect 112 46 142 176
rect 208 46 238 176
rect 304 46 334 176
rect 400 46 430 176
rect 496 46 526 176
rect 592 46 622 176
rect 688 46 718 176
rect 784 46 814 176
rect 880 46 910 176
rect 976 46 1006 176
rect 1168 46 1198 176
rect 1264 46 1294 176
rect 1360 46 1390 176
rect 1456 46 1486 176
rect 1552 46 1582 176
<< pmos >>
rect 112 296 142 496
rect 208 296 238 496
rect 304 296 334 496
rect 400 296 430 496
rect 496 296 526 496
rect 592 296 622 496
rect 688 296 718 496
rect 880 296 910 496
rect 976 296 1006 496
rect 1072 296 1102 496
rect 1264 296 1294 496
rect 1360 296 1390 496
rect 1456 296 1486 496
rect 1552 296 1582 496
<< ndiff >>
rect 58 142 112 176
rect 56 100 112 142
rect 56 66 66 100
rect 100 66 112 100
rect 56 48 112 66
rect 58 46 112 48
rect 142 46 208 176
rect 238 100 304 176
rect 238 66 254 100
rect 288 66 304 100
rect 238 46 304 66
rect 334 46 400 176
rect 430 100 496 176
rect 430 66 446 100
rect 480 66 496 100
rect 430 46 496 66
rect 526 46 592 176
rect 622 100 688 176
rect 622 66 638 100
rect 672 66 688 100
rect 622 46 688 66
rect 718 100 784 176
rect 718 66 734 100
rect 768 66 784 100
rect 718 46 784 66
rect 814 100 880 176
rect 814 66 830 100
rect 864 66 880 100
rect 814 46 880 66
rect 910 46 976 176
rect 1006 164 1060 176
rect 1006 130 1017 164
rect 1051 130 1060 164
rect 1006 46 1060 130
rect 1114 96 1168 176
rect 1114 62 1122 96
rect 1156 62 1168 96
rect 1114 46 1168 62
rect 1198 100 1264 176
rect 1198 66 1214 100
rect 1248 66 1264 100
rect 1198 46 1264 66
rect 1294 100 1360 176
rect 1294 66 1310 100
rect 1344 66 1360 100
rect 1294 46 1360 66
rect 1390 100 1456 176
rect 1390 66 1406 100
rect 1440 66 1456 100
rect 1390 46 1456 66
rect 1486 100 1552 176
rect 1486 66 1502 100
rect 1536 66 1552 100
rect 1486 46 1552 66
rect 1582 100 1636 176
rect 1582 66 1594 100
rect 1628 66 1636 100
rect 1582 46 1636 66
<< pdiff >>
rect 58 378 112 496
rect 58 344 66 378
rect 100 344 112 378
rect 58 296 112 344
rect 142 476 208 496
rect 142 442 158 476
rect 192 442 208 476
rect 142 296 208 442
rect 238 378 304 496
rect 238 344 254 378
rect 288 344 304 378
rect 238 296 304 344
rect 334 378 400 496
rect 334 344 350 378
rect 384 344 400 378
rect 334 296 400 344
rect 430 378 496 496
rect 430 344 446 378
rect 480 344 496 378
rect 430 296 496 344
rect 526 476 592 496
rect 526 442 542 476
rect 576 442 592 476
rect 526 296 592 442
rect 622 446 688 496
rect 622 412 638 446
rect 672 412 688 446
rect 622 296 688 412
rect 718 378 772 496
rect 718 344 729 378
rect 763 344 772 378
rect 718 296 772 344
rect 826 476 880 496
rect 826 442 834 476
rect 868 442 880 476
rect 826 296 880 442
rect 910 378 976 496
rect 910 344 926 378
rect 960 344 976 378
rect 910 296 976 344
rect 1006 476 1072 496
rect 1006 442 1022 476
rect 1056 442 1072 476
rect 1006 296 1072 442
rect 1102 446 1156 496
rect 1102 412 1113 446
rect 1147 412 1156 446
rect 1102 296 1156 412
rect 1210 378 1264 496
rect 1210 344 1218 378
rect 1252 344 1264 378
rect 1210 296 1264 344
rect 1294 296 1360 496
rect 1390 476 1456 496
rect 1390 442 1406 476
rect 1440 442 1456 476
rect 1390 296 1456 442
rect 1486 296 1552 496
rect 1582 378 1636 496
rect 1582 344 1593 378
rect 1627 344 1636 378
rect 1582 296 1636 344
<< ndiffc >>
rect 66 66 100 100
rect 254 66 288 100
rect 446 66 480 100
rect 638 66 672 100
rect 734 66 768 100
rect 830 66 864 100
rect 1017 130 1051 164
rect 1122 62 1156 96
rect 1214 66 1248 100
rect 1310 66 1344 100
rect 1406 66 1440 100
rect 1502 66 1536 100
rect 1594 66 1628 100
<< pdiffc >>
rect 66 344 100 378
rect 158 442 192 476
rect 254 344 288 378
rect 350 344 384 378
rect 446 344 480 378
rect 542 442 576 476
rect 638 412 672 446
rect 729 344 763 378
rect 834 442 868 476
rect 926 344 960 378
rect 1022 442 1056 476
rect 1113 412 1147 446
rect 1218 344 1252 378
rect 1406 442 1440 476
rect 1593 344 1627 378
<< poly >>
rect 112 496 142 522
rect 208 496 238 522
rect 304 496 334 522
rect 400 496 430 522
rect 496 496 526 522
rect 592 496 622 522
rect 688 496 718 522
rect 880 496 910 522
rect 976 496 1006 522
rect 1072 496 1102 522
rect 1264 496 1294 522
rect 1360 496 1390 522
rect 1456 496 1486 522
rect 1552 496 1582 522
rect 112 264 142 296
rect 208 264 238 296
rect 304 264 334 296
rect 400 264 430 296
rect 496 264 526 296
rect 592 264 622 296
rect 688 264 718 296
rect 880 264 910 296
rect 976 264 1006 296
rect 1072 264 1102 296
rect 1264 264 1294 296
rect 1360 264 1390 296
rect 1456 264 1486 296
rect 1552 264 1582 296
rect 100 248 154 264
rect 100 214 110 248
rect 144 214 154 248
rect 100 198 154 214
rect 196 248 250 264
rect 196 214 206 248
rect 240 214 250 248
rect 196 198 250 214
rect 292 248 346 264
rect 292 214 302 248
rect 336 214 346 248
rect 292 198 346 214
rect 388 248 442 264
rect 388 214 398 248
rect 432 214 442 248
rect 388 198 442 214
rect 484 248 538 264
rect 484 214 494 248
rect 528 214 538 248
rect 484 198 538 214
rect 580 248 634 264
rect 580 214 590 248
rect 624 214 634 248
rect 580 198 634 214
rect 676 248 730 264
rect 676 214 686 248
rect 720 214 730 248
rect 676 198 730 214
rect 772 248 826 264
rect 772 214 782 248
rect 816 214 826 248
rect 772 198 826 214
rect 868 248 922 264
rect 868 214 878 248
rect 912 214 922 248
rect 868 198 922 214
rect 964 248 1018 264
rect 964 214 974 248
rect 1008 214 1018 248
rect 964 198 1018 214
rect 1060 248 1114 264
rect 1060 214 1070 248
rect 1104 214 1114 248
rect 1060 198 1114 214
rect 1156 248 1210 264
rect 1156 214 1166 248
rect 1200 214 1210 248
rect 1156 198 1210 214
rect 1252 248 1306 264
rect 1252 214 1262 248
rect 1296 214 1306 248
rect 1252 198 1306 214
rect 1348 248 1402 264
rect 1348 214 1358 248
rect 1392 214 1402 248
rect 1348 198 1402 214
rect 1444 248 1498 264
rect 1444 214 1454 248
rect 1488 214 1498 248
rect 1444 198 1498 214
rect 1540 248 1594 264
rect 1540 214 1550 248
rect 1584 214 1594 248
rect 1540 198 1594 214
rect 112 176 142 198
rect 208 176 238 198
rect 304 176 334 198
rect 400 176 430 198
rect 496 176 526 198
rect 592 176 622 198
rect 688 176 718 198
rect 784 176 814 198
rect 880 176 910 198
rect 976 176 1006 198
rect 1168 176 1198 198
rect 1264 176 1294 198
rect 1360 176 1390 198
rect 1456 176 1486 198
rect 1552 176 1582 198
rect 112 20 142 46
rect 208 20 238 46
rect 304 20 334 46
rect 400 20 430 46
rect 496 20 526 46
rect 592 20 622 46
rect 688 20 718 46
rect 784 20 814 46
rect 880 20 910 46
rect 976 20 1006 46
rect 1168 20 1198 46
rect 1264 20 1294 46
rect 1360 20 1390 46
rect 1456 20 1486 46
rect 1552 20 1582 46
<< polycont >>
rect 110 214 144 248
rect 206 214 240 248
rect 302 214 336 248
rect 398 214 432 248
rect 494 214 528 248
rect 590 214 624 248
rect 686 214 720 248
rect 782 214 816 248
rect 878 214 912 248
rect 974 214 1008 248
rect 1070 214 1104 248
rect 1166 214 1200 248
rect 1262 214 1296 248
rect 1358 214 1392 248
rect 1454 214 1488 248
rect 1550 214 1584 248
<< locali >>
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1748 560
rect 158 476 192 526
rect 542 476 576 526
rect 158 426 192 442
rect 422 422 446 456
rect 834 476 868 526
rect 542 426 576 442
rect 638 456 672 462
rect 66 328 100 344
rect 254 328 288 344
rect 350 378 384 394
rect 422 378 480 422
rect 638 396 672 412
rect 834 426 868 442
rect 1022 476 1056 526
rect 1406 476 1440 526
rect 1022 426 1056 442
rect 1113 456 1148 462
rect 734 378 768 422
rect 1147 412 1148 456
rect 1406 426 1440 442
rect 1536 422 1604 456
rect 1113 396 1148 412
rect 1218 378 1220 400
rect 1570 394 1604 422
rect 1570 378 1627 394
rect 422 344 446 378
rect 712 344 729 378
rect 763 344 779 378
rect 878 344 926 378
rect 960 344 976 378
rect 1254 366 1488 378
rect 1252 344 1488 366
rect 1570 344 1593 378
rect 446 328 480 344
rect 1218 328 1254 344
rect 1592 328 1627 344
rect 110 248 144 254
rect 110 198 144 214
rect 206 248 240 254
rect 206 198 240 214
rect 302 248 336 264
rect 494 248 528 264
rect 374 214 398 248
rect 432 214 448 248
rect 374 120 408 214
rect 590 248 624 310
rect 590 198 624 214
rect 686 248 720 254
rect 686 198 720 214
rect 782 248 816 264
rect 878 248 912 264
rect 974 248 1008 254
rect 1070 254 1166 268
rect 1070 248 1200 254
rect 1262 248 1296 264
rect 1054 214 1070 248
rect 1104 214 1166 248
rect 1200 214 1216 248
rect 974 198 1008 214
rect 1358 248 1392 254
rect 1358 198 1392 214
rect 1454 248 1488 264
rect 1584 254 1604 288
rect 1550 248 1604 254
rect 1526 214 1550 248
rect 1584 214 1604 248
rect 1526 206 1604 214
rect 998 130 1017 164
rect 1051 138 1070 164
rect 1051 130 1104 138
rect 66 50 100 66
rect 254 100 288 116
rect 384 86 408 120
rect 254 16 288 66
rect 446 50 480 66
rect 638 100 672 116
rect 706 86 726 110
rect 760 100 768 116
rect 706 66 734 86
rect 638 16 672 66
rect 734 50 768 66
rect 830 100 864 116
rect 830 16 864 66
rect 1214 100 1248 116
rect 960 86 1122 96
rect 926 62 1122 86
rect 1156 62 1174 96
rect 1214 16 1248 66
rect 1310 50 1344 66
rect 1406 100 1440 116
rect 1406 16 1440 66
rect 1502 50 1536 66
rect 1594 100 1628 116
rect 1594 16 1628 66
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1748 16
<< viali >>
rect 28 526 62 560
rect 120 526 154 560
rect 212 526 246 560
rect 304 526 338 560
rect 396 526 430 560
rect 488 526 522 560
rect 580 526 614 560
rect 672 526 706 560
rect 764 526 798 560
rect 856 526 890 560
rect 948 526 982 560
rect 1040 526 1074 560
rect 1132 526 1166 560
rect 1224 526 1258 560
rect 1316 526 1350 560
rect 1408 526 1442 560
rect 1500 526 1534 560
rect 1592 526 1626 560
rect 1684 526 1718 560
rect 446 422 480 456
rect 638 446 672 456
rect 66 378 100 400
rect 66 366 100 378
rect 254 378 288 400
rect 254 366 288 378
rect 638 422 672 446
rect 734 422 768 456
rect 1113 446 1147 456
rect 1113 422 1147 446
rect 1502 422 1536 456
rect 1220 378 1254 400
rect 1220 366 1252 378
rect 1252 366 1254 378
rect 350 310 384 344
rect 590 310 624 344
rect 878 310 912 344
rect 1454 310 1488 344
rect 110 254 144 288
rect 206 254 240 288
rect 302 214 336 232
rect 302 198 336 214
rect 494 214 528 232
rect 494 198 528 214
rect 686 254 720 288
rect 782 214 816 232
rect 782 198 816 214
rect 878 214 912 232
rect 878 198 912 214
rect 974 254 1008 288
rect 1166 254 1200 288
rect 1262 214 1296 232
rect 1262 198 1296 214
rect 1358 254 1392 288
rect 1550 254 1584 288
rect 1454 214 1488 232
rect 1454 198 1488 214
rect 1070 138 1104 172
rect 66 100 100 120
rect 66 86 100 100
rect 350 86 384 120
rect 446 100 480 120
rect 446 86 480 100
rect 726 100 760 120
rect 726 86 734 100
rect 734 86 760 100
rect 926 86 960 120
rect 1310 100 1344 120
rect 1310 86 1344 100
rect 1502 100 1536 120
rect 1502 86 1536 100
rect 28 -18 62 16
rect 120 -18 154 16
rect 212 -18 246 16
rect 304 -18 338 16
rect 396 -18 430 16
rect 488 -18 522 16
rect 580 -18 614 16
rect 672 -18 706 16
rect 764 -18 798 16
rect 856 -18 890 16
rect 948 -18 982 16
rect 1040 -18 1074 16
rect 1132 -18 1166 16
rect 1224 -18 1258 16
rect 1316 -18 1350 16
rect 1408 -18 1442 16
rect 1500 -18 1534 16
rect 1592 -18 1626 16
rect 1684 -18 1718 16
<< metal1 >>
rect 0 560 1748 592
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1748 560
rect 0 520 1748 526
rect 434 456 492 462
rect 434 422 446 456
rect 480 422 492 456
rect 434 420 492 422
rect 256 416 492 420
rect 52 358 58 410
rect 110 358 116 410
rect 256 406 476 416
rect 622 414 628 466
rect 680 414 686 466
rect 742 462 748 466
rect 722 456 748 462
rect 722 422 734 456
rect 722 416 748 422
rect 742 414 748 416
rect 800 414 806 466
rect 1054 414 1060 466
rect 1115 462 1121 466
rect 1115 456 1159 462
rect 1147 422 1159 456
rect 1115 416 1159 422
rect 1490 456 1548 462
rect 1490 422 1502 456
rect 1536 454 1548 456
rect 1576 454 1582 466
rect 1536 426 1582 454
rect 1536 422 1548 426
rect 1490 416 1548 422
rect 1115 414 1121 416
rect 1576 414 1582 426
rect 1634 414 1640 466
rect 242 400 476 406
rect 242 366 254 400
rect 288 392 476 400
rect 288 366 300 392
rect 242 360 300 366
rect 728 358 762 378
rect 1204 358 1210 410
rect 1262 358 1268 410
rect 338 344 396 350
rect 338 310 350 344
rect 384 342 396 344
rect 384 310 428 342
rect 338 304 428 310
rect 98 288 156 294
rect 98 254 110 288
rect 144 254 156 288
rect 98 248 156 254
rect 112 202 140 248
rect 190 246 196 298
rect 248 246 254 298
rect 112 174 236 202
rect 286 190 292 242
rect 344 190 350 242
rect 400 238 428 304
rect 526 302 532 354
rect 584 350 590 354
rect 584 344 636 350
rect 584 310 590 344
rect 624 310 636 344
rect 584 304 636 310
rect 664 344 1100 358
rect 664 314 878 344
rect 584 302 590 304
rect 664 288 732 314
rect 866 310 878 314
rect 912 330 1100 344
rect 912 310 924 330
rect 866 304 924 310
rect 664 258 686 288
rect 674 254 686 258
rect 720 254 732 288
rect 674 248 732 254
rect 958 246 964 298
rect 1016 246 1022 298
rect 400 210 452 238
rect 208 142 236 174
rect 160 130 236 142
rect 52 78 58 130
rect 110 78 116 130
rect 160 90 220 130
rect 214 78 220 90
rect 272 118 278 130
rect 424 126 452 210
rect 482 232 540 238
rect 482 198 494 232
rect 528 230 540 232
rect 574 230 580 242
rect 528 202 580 230
rect 528 198 540 202
rect 482 192 540 198
rect 574 190 580 202
rect 632 190 638 242
rect 770 232 828 238
rect 770 198 782 232
rect 816 198 828 232
rect 770 192 828 198
rect 800 142 828 192
rect 862 190 868 242
rect 920 190 926 242
rect 1072 202 1100 330
rect 1442 344 1500 350
rect 1168 298 1388 314
rect 1442 310 1454 344
rect 1488 342 1500 344
rect 1488 314 1556 342
rect 1488 310 1500 314
rect 1442 304 1500 310
rect 1130 246 1136 298
rect 1188 294 1388 298
rect 1528 294 1580 314
rect 1188 288 1404 294
rect 1200 286 1358 288
rect 1200 254 1212 286
rect 1188 248 1212 254
rect 1346 254 1358 286
rect 1392 254 1404 288
rect 1528 288 1596 294
rect 1528 286 1550 288
rect 1346 248 1404 254
rect 1538 254 1550 286
rect 1584 254 1596 288
rect 1538 248 1596 254
rect 1188 246 1194 248
rect 1250 232 1308 238
rect 1250 202 1262 232
rect 1072 198 1262 202
rect 1296 198 1308 232
rect 1072 192 1308 198
rect 1072 182 1292 192
rect 1438 190 1444 242
rect 1496 190 1502 242
rect 1058 174 1292 182
rect 1058 172 1116 174
rect 800 130 860 142
rect 1058 138 1070 172
rect 1104 138 1116 172
rect 1058 132 1116 138
rect 338 120 396 126
rect 338 118 350 120
rect 272 90 350 118
rect 272 78 278 90
rect 338 86 350 90
rect 384 86 396 120
rect 424 120 492 126
rect 424 90 446 120
rect 338 80 396 86
rect 434 86 446 90
rect 480 118 492 120
rect 598 118 604 130
rect 480 90 604 118
rect 480 86 492 90
rect 434 80 492 86
rect 598 78 604 90
rect 656 78 662 130
rect 692 78 698 130
rect 750 120 772 130
rect 760 86 772 120
rect 800 114 820 130
rect 750 78 772 86
rect 814 78 820 114
rect 872 118 878 130
rect 958 126 964 130
rect 914 120 964 126
rect 914 118 926 120
rect 872 90 926 118
rect 872 78 878 90
rect 914 86 926 90
rect 960 86 964 120
rect 914 80 964 86
rect 958 78 964 80
rect 1016 78 1022 130
rect 1204 78 1210 130
rect 1262 118 1268 130
rect 1298 120 1356 126
rect 1298 118 1310 120
rect 1262 90 1310 118
rect 1262 78 1268 90
rect 1298 86 1310 90
rect 1344 86 1356 120
rect 1298 80 1356 86
rect 1490 120 1548 126
rect 1490 86 1502 120
rect 1536 118 1548 120
rect 1576 118 1582 130
rect 1536 90 1582 118
rect 1536 86 1548 90
rect 1490 80 1548 86
rect 1576 78 1582 90
rect 1634 78 1640 130
rect 0 16 1748 24
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1748 16
rect 0 -48 1748 -18
<< via1 >>
rect 58 400 110 410
rect 58 366 66 400
rect 66 366 100 400
rect 100 366 110 400
rect 58 358 110 366
rect 628 456 680 466
rect 628 422 638 456
rect 638 422 672 456
rect 672 422 680 456
rect 628 414 680 422
rect 748 456 800 466
rect 748 422 768 456
rect 768 422 800 456
rect 748 414 800 422
rect 1060 456 1115 466
rect 1060 422 1113 456
rect 1113 422 1115 456
rect 1060 414 1115 422
rect 1582 414 1634 466
rect 1210 400 1262 410
rect 1210 366 1220 400
rect 1220 366 1254 400
rect 1254 366 1262 400
rect 1210 358 1262 366
rect 196 288 248 298
rect 196 254 206 288
rect 206 254 240 288
rect 240 254 248 288
rect 196 246 248 254
rect 292 232 344 242
rect 292 198 302 232
rect 302 198 336 232
rect 336 198 344 232
rect 292 190 344 198
rect 532 302 584 354
rect 964 288 1016 298
rect 964 254 974 288
rect 974 254 1008 288
rect 1008 254 1016 288
rect 964 246 1016 254
rect 58 120 110 130
rect 58 86 66 120
rect 66 86 100 120
rect 100 86 110 120
rect 58 78 110 86
rect 220 78 272 130
rect 580 190 632 242
rect 868 232 920 242
rect 868 198 878 232
rect 878 198 912 232
rect 912 198 920 232
rect 868 190 920 198
rect 1136 288 1188 298
rect 1136 254 1166 288
rect 1166 254 1188 288
rect 1136 246 1188 254
rect 1444 232 1496 242
rect 1444 198 1454 232
rect 1454 198 1488 232
rect 1488 198 1496 232
rect 1444 190 1496 198
rect 604 78 656 130
rect 698 120 750 130
rect 698 86 726 120
rect 726 86 750 120
rect 698 78 750 86
rect 820 78 872 130
rect 964 78 1016 130
rect 1210 78 1262 130
rect 1582 78 1634 130
<< metal2 >>
rect 688 502 1176 530
rect 688 472 716 502
rect 628 466 716 472
rect 160 426 628 454
rect 58 410 110 416
rect 160 398 188 426
rect 680 426 716 466
rect 748 466 800 472
rect 628 408 680 414
rect 748 408 800 414
rect 962 462 1018 472
rect 748 398 788 408
rect 110 370 188 398
rect 710 370 788 398
rect 1060 466 1115 472
rect 1060 408 1115 414
rect 962 396 1018 406
rect 58 352 110 358
rect 242 356 298 365
rect 70 136 98 352
rect 208 304 242 342
rect 196 300 242 304
rect 532 354 584 360
rect 298 314 532 342
rect 196 298 298 300
rect 194 246 196 252
rect 248 290 298 298
rect 532 296 584 302
rect 431 252 492 253
rect 248 246 250 252
rect 194 178 250 246
rect 292 242 344 248
rect 410 244 492 252
rect 410 230 436 244
rect 344 202 436 230
rect 292 184 344 190
rect 410 188 436 202
rect 410 178 492 188
rect 578 244 634 253
rect 578 178 634 188
rect 710 146 738 370
rect 976 304 1004 396
rect 964 298 1016 304
rect 866 262 922 272
rect 866 190 868 206
rect 920 190 922 206
rect 866 178 922 190
rect 962 246 964 252
rect 1016 246 1018 252
rect 962 178 1018 246
rect 194 136 250 141
rect 710 136 772 146
rect 1072 144 1100 408
rect 1148 304 1176 502
rect 1582 466 1634 472
rect 1210 410 1262 416
rect 1582 408 1634 414
rect 1210 352 1262 358
rect 1136 298 1188 304
rect 1136 240 1188 246
rect 1222 144 1250 352
rect 1594 252 1622 408
rect 1444 242 1496 248
rect 1312 202 1444 230
rect 1004 140 1100 144
rect 58 130 110 136
rect 58 72 110 78
rect 194 132 272 136
rect 250 130 272 132
rect 250 76 272 78
rect 194 72 272 76
rect 604 130 656 136
rect 698 130 716 136
rect 818 130 874 140
rect 656 78 668 118
rect 604 72 668 78
rect 194 66 250 72
rect 640 42 668 72
rect 772 80 780 130
rect 750 78 780 80
rect 698 71 780 78
rect 818 78 820 130
rect 872 78 874 130
rect 818 72 874 78
rect 964 136 1100 140
rect 964 130 1004 136
rect 1060 90 1100 136
rect 1208 134 1264 144
rect 1016 78 1060 80
rect 1198 78 1208 130
rect 1264 78 1273 130
rect 964 70 1060 78
rect 1208 70 1264 78
rect 1312 42 1340 202
rect 1444 184 1496 190
rect 1560 178 1622 252
rect 1574 141 1622 178
rect 1574 132 1636 141
rect 1574 90 1580 132
rect 1580 66 1636 76
rect 640 14 1340 42
<< via2 >>
rect 962 406 1018 462
rect 242 300 298 356
rect 436 188 492 244
rect 578 242 634 244
rect 578 190 580 242
rect 580 190 632 242
rect 632 190 634 242
rect 578 188 634 190
rect 866 242 922 262
rect 866 206 868 242
rect 868 206 920 242
rect 920 206 922 242
rect 194 130 250 132
rect 194 78 220 130
rect 220 78 250 130
rect 194 76 250 78
rect 716 130 772 136
rect 716 80 750 130
rect 750 80 772 130
rect 1004 130 1060 136
rect 1004 80 1016 130
rect 1016 80 1060 130
rect 1208 130 1264 134
rect 1208 78 1210 130
rect 1210 78 1262 130
rect 1262 78 1264 130
rect 1580 130 1636 132
rect 1580 78 1582 130
rect 1582 78 1634 130
rect 1634 78 1636 130
rect 1580 76 1636 78
<< metal3 >>
rect 958 470 1024 472
rect 576 462 1024 470
rect 576 410 962 462
rect 238 360 301 361
rect 430 360 494 366
rect 192 356 338 360
rect 192 300 242 356
rect 298 300 338 356
rect 192 294 338 300
rect 430 290 494 296
rect 430 252 496 290
rect 576 252 636 410
rect 956 406 962 410
rect 1018 406 1024 462
rect 956 400 1024 406
rect 430 244 497 252
rect 430 188 436 244
rect 492 188 497 244
rect 430 182 497 188
rect 572 249 636 252
rect 772 266 928 272
rect 572 244 640 249
rect 572 188 578 244
rect 634 188 640 244
rect 772 204 862 266
rect 860 202 862 204
rect 926 202 928 266
rect 862 196 928 202
rect 572 182 640 188
rect 186 136 257 137
rect 686 136 832 142
rect 166 132 312 136
rect 166 76 194 132
rect 250 76 312 132
rect 166 70 312 76
rect 686 80 716 136
rect 772 80 832 136
rect 686 76 832 80
rect 995 140 1065 141
rect 995 136 1142 140
rect 995 80 1004 136
rect 1060 80 1142 136
rect 686 74 782 76
rect 995 70 1142 80
rect 1202 134 1350 140
rect 1574 136 1646 137
rect 1202 78 1208 134
rect 1264 78 1350 134
rect 1202 74 1350 78
rect 1542 132 1688 136
rect 1542 76 1580 132
rect 1636 76 1688 132
rect 1202 72 1268 74
rect 1542 70 1688 76
rect 995 69 1065 70
rect 1574 69 1646 70
<< via3 >>
rect 430 296 494 360
rect 862 262 926 266
rect 862 206 866 262
rect 866 206 922 262
rect 922 206 926 262
rect 862 202 926 206
<< metal4 >>
rect 428 360 496 361
rect 428 296 430 360
rect 494 296 496 360
rect 428 294 496 296
rect 432 260 496 294
rect 860 266 928 268
rect 860 260 862 266
rect 432 202 862 260
rect 926 202 928 266
rect 432 200 928 202
rect 862 196 928 200
<< labels >>
flabel nwell s 76 526 110 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 76 -16 110 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 0 0 0 0 FreeSans 100 0 0 0 scs130hd_mpr2xa_8
rlabel metal3 s 996 70 1142 140 4 R0
port 3 nsew
rlabel metal3 s 1542 70 1688 136 4 R1
port 4 nsew
rlabel metal3 s 686 76 832 142 4 R2
port 5 nsew
rlabel metal3 s 1204 74 1350 140 4 R3
port 6 nsew
rlabel metal3 s 958 470 1024 472 4 B1
port 7 nsew
rlabel metal3 s 166 70 312 136 4 B0
port 8 nsew
rlabel metal3 s 192 294 338 360 4 A0
port 9 nsew
flabel metal1 s 30 -16 64 16 0 FreeSans 100 0 0 0 vgnd
port 10 nsew
flabel metal1 s 30 526 64 560 0 FreeSans 100 0 0 0 vpwr
port 11 nsew
rlabel metal4 s 928 248 928 248 4 A1
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 1748 544
<< end >>
