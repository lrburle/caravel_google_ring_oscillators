magic
tech sky130A
magscale 1 2
timestamp 1716047795
<< error_s >>
rect 295 1755 311 1785
rect 323 1755 339 1757
rect 193 1630 219 1646
rect 221 1640 247 1646
<< nwell >>
rect 0 1428 714 1748
rect 2307 1645 2465 1748
rect 2507 1645 2539 1681
rect 2307 1626 2470 1645
rect 0 1401 728 1428
rect 2268 1406 2470 1626
rect 3401 1406 3446 1748
rect 0 1128 831 1401
rect 2249 1391 3446 1406
rect 2231 1360 3446 1391
rect 2229 1128 3446 1360
rect 0 1084 830 1128
rect 2231 1097 3446 1128
rect 2248 1086 3446 1097
rect 0 862 834 1084
rect 2248 1055 2470 1086
rect 1886 1022 2470 1055
rect 2248 862 2470 1022
rect 0 742 719 862
rect 2307 744 2470 862
rect 3252 772 3282 807
rect 3401 744 3446 1086
<< ndiff >>
rect 3336 441 3371 475
<< psubdiff >>
rect 2477 2206 2499 2213
rect 2477 2173 2507 2206
rect 2633 2173 2708 2206
<< locali >>
rect 1 2176 3449 2492
rect 1 2172 824 2176
rect 759 1706 824 2172
rect 889 1706 954 2176
rect 1019 1706 1084 2176
rect 1149 1706 1214 2176
rect 1195 1702 1214 1706
rect 1279 1702 1344 2176
rect 1409 1702 1474 2176
rect 1539 1702 1604 2176
rect 1669 1702 1734 2176
rect 1799 1702 1864 2176
rect 1929 1706 1994 2176
rect 2059 1706 2124 2176
rect 2189 2172 3449 2176
rect 2189 1706 2231 2172
rect 3171 1721 3279 1756
rect 1929 1702 1934 1706
rect 1195 1695 1934 1702
rect 1254 1465 1288 1680
rect 2505 1645 2541 1693
rect 3171 1690 3174 1721
rect 3338 1461 3372 1495
rect 1 1401 714 1405
rect 1 1360 715 1401
rect 2249 1360 3446 1406
rect 1 1128 831 1360
rect 2229 1128 3446 1360
rect 1 1085 830 1128
rect 2248 1086 3446 1128
rect 3337 997 3371 1031
rect 3173 725 3272 761
rect 758 586 765 618
rect 2229 591 2307 618
rect 933 586 962 590
rect 758 320 827 586
rect 896 320 962 586
rect 1031 321 1100 590
rect 1169 321 1238 590
rect 1307 321 1376 590
rect 1445 321 1514 590
rect 1583 321 1652 590
rect 1721 321 1790 590
rect 1859 321 1928 590
rect 1997 321 2066 590
rect 2135 321 2204 590
rect 2230 584 2307 591
rect 2273 321 2307 584
rect 1031 320 2307 321
rect 1 0 3449 320
<< viali >>
rect 3053 1877 3099 1923
rect 3337 1743 3371 1777
rect 3048 589 3094 635
rect 3337 441 3371 475
<< metal1 >>
rect 1 2176 3449 2492
rect 1 2172 824 2176
rect 277 1755 311 2172
rect 425 1929 499 1938
rect 425 1873 434 1929
rect 490 1873 499 1929
rect 425 1864 499 1873
rect 514 1772 520 1828
rect 576 1772 582 1828
rect 277 1754 344 1755
rect 277 1729 357 1754
rect 277 1720 369 1729
rect 759 1706 824 2172
rect 889 1706 954 2176
rect 1019 1706 1084 2176
rect 1149 1706 1214 2176
rect 1195 1702 1214 1706
rect 1279 1702 1344 2176
rect 1409 1702 1474 2176
rect 1539 1702 1604 2176
rect 1669 1702 1734 2176
rect 1799 1702 1864 2176
rect 1929 1706 1994 2176
rect 2059 1706 2124 2176
rect 2189 2172 3449 2176
rect 2189 1706 2231 2172
rect 3053 1930 3099 1935
rect 3047 1923 3105 1930
rect 3047 1915 3053 1923
rect 2815 1908 3053 1915
rect 2827 1902 3053 1908
rect 2781 1881 3053 1902
rect 2781 1868 2827 1881
rect 3047 1877 3053 1881
rect 3099 1877 3105 1923
rect 3047 1871 3105 1877
rect 3053 1865 3099 1871
rect 2860 1846 2925 1853
rect 2860 1794 2867 1846
rect 2919 1794 2925 1846
rect 2860 1788 2925 1794
rect 2700 1772 2764 1778
rect 2700 1720 2706 1772
rect 2758 1720 2764 1772
rect 2700 1713 2764 1720
rect 1929 1702 1934 1706
rect 151 1692 219 1698
rect 1195 1695 1934 1702
rect 151 1636 157 1692
rect 213 1680 219 1692
rect 213 1675 222 1680
rect 614 1675 620 1691
rect 213 1646 620 1675
rect 213 1636 219 1646
rect 221 1640 620 1646
rect 151 1630 219 1636
rect 614 1635 620 1640
rect 676 1635 682 1691
rect 2491 1686 2556 1693
rect 2491 1634 2498 1686
rect 2550 1634 2556 1686
rect 2491 1628 2556 1634
rect 1 1401 714 1405
rect 1 1360 715 1401
rect 2249 1391 3446 1406
rect 2231 1360 3446 1391
rect 1 1128 831 1360
rect 2229 1128 3446 1360
rect 1 1085 830 1128
rect 2231 1097 3446 1128
rect 2248 1086 3446 1097
rect 2491 1016 2556 1023
rect 2491 964 2498 1016
rect 2550 964 2556 1016
rect 2491 958 2556 964
rect 2507 845 2541 958
rect 2700 790 2764 796
rect 2700 772 2706 790
rect 2637 738 2706 772
rect 2758 738 2764 790
rect 2700 732 2764 738
rect 2366 716 2431 723
rect 2366 664 2373 716
rect 2425 664 2431 716
rect 2366 658 2431 664
rect 2855 716 2925 722
rect 2855 658 2861 716
rect 2919 658 2925 716
rect 2855 652 2925 658
rect 3048 641 3094 647
rect 3042 635 3100 641
rect 3042 624 3048 635
rect 758 586 766 624
rect 2230 618 2307 624
rect 2229 591 2307 618
rect 2230 590 2307 591
rect 2781 623 2815 624
rect 2827 623 3048 624
rect 2781 590 3048 623
rect 933 586 962 590
rect 758 320 827 586
rect 896 320 962 586
rect 1031 321 1100 590
rect 1169 321 1238 590
rect 1307 321 1376 590
rect 1445 321 1514 590
rect 1583 321 1652 590
rect 1721 321 1790 590
rect 1859 321 1928 590
rect 1997 321 2066 590
rect 2135 553 2307 590
rect 3042 589 3048 590
rect 3094 589 3100 635
rect 3042 582 3100 589
rect 3048 577 3094 582
rect 2135 321 2204 553
rect 2273 321 2307 553
rect 1031 320 2307 321
rect 1 0 3449 320
<< via1 >>
rect 434 1873 490 1929
rect 520 1772 576 1828
rect 2867 1794 2919 1846
rect 2706 1720 2758 1772
rect 157 1636 213 1692
rect 620 1635 676 1691
rect 2498 1634 2550 1686
rect 2498 964 2550 1016
rect 2706 738 2758 790
rect 2373 664 2425 716
rect 2861 658 2919 716
<< metal2 >>
rect 425 1929 499 1938
rect 425 1873 434 1929
rect 490 1873 499 1929
rect 425 1864 499 1873
rect 530 1910 2669 1944
rect 530 1834 564 1910
rect 631 1848 2541 1882
rect 520 1828 576 1834
rect 520 1766 576 1772
rect 147 1692 222 1701
rect 631 1697 665 1848
rect 147 1636 157 1692
rect 213 1636 222 1692
rect 147 1627 222 1636
rect 620 1691 676 1697
rect 2507 1693 2541 1848
rect 2637 1840 2669 1910
rect 2860 1846 2925 1853
rect 2860 1840 2867 1846
rect 2637 1806 2867 1840
rect 620 1629 676 1635
rect 2491 1686 2556 1693
rect 2491 1634 2498 1686
rect 2550 1634 2556 1686
rect 2491 1628 2556 1634
rect 2505 1023 2539 1628
rect 2491 1016 2556 1023
rect 2491 964 2498 1016
rect 2550 964 2556 1016
rect 2491 958 2556 964
rect 1663 874 1698 895
rect 2637 772 2669 1806
rect 2860 1794 2867 1806
rect 2919 1794 2925 1846
rect 2860 1788 2925 1794
rect 2700 1772 2764 1778
rect 2700 1720 2706 1772
rect 2758 1720 2764 1772
rect 2700 1713 2764 1720
rect 2706 1666 2740 1713
rect 2706 1631 2741 1666
rect 2706 1596 2901 1631
rect 2700 790 2764 796
rect 2700 772 2706 790
rect 1379 728 2307 763
rect 2637 738 2706 772
rect 2758 738 2764 790
rect 2700 732 2764 738
rect 2272 698 2307 728
rect 2366 716 2431 723
rect 2866 722 2901 1596
rect 2366 698 2373 716
rect 2272 664 2373 698
rect 2425 698 2431 716
rect 2855 716 2925 722
rect 2855 698 2861 716
rect 2425 664 2861 698
rect 2366 658 2431 664
rect 2855 658 2861 664
rect 2919 658 2925 716
rect 2855 652 2925 658
<< via2 >>
rect 434 1873 490 1929
rect 157 1636 213 1692
<< metal3 >>
rect 151 1701 218 2477
rect 425 1929 499 1938
rect 425 1873 434 1929
rect 490 1924 499 1929
rect 490 1873 1855 1924
rect 425 1864 1855 1873
rect 147 1692 222 1701
rect 147 1636 157 1692
rect 213 1636 222 1692
rect 147 1627 222 1636
rect 1378 1557 1438 1864
rect 1584 1620 1645 1864
rect 1584 1486 1644 1620
rect 1795 1493 1855 1864
rect 1576 1416 1644 1486
rect 1780 1420 1855 1493
use scs130hd_mpr2ct_8  scs130hd_mpr2ct_8_1
timestamp 1710282110
transform 1 0 759 0 1 601
box -43 -60 1510 1148
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1714057206
transform 1 0 3019 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1714057206
transform 1 0 3216 0 1 259
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1714057206
transform 1 0 3217 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1714057206
transform 1 0 3019 0 -1 2233
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 2470 0 1 259
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1714057206
transform 1 0 133 0 -1 2233
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1714057206
transform 1 0 2470 0 -1 2233
box -10 0 552 902
<< labels >>
rlabel metal2 2523 992 2523 992 1 sel
port 8 n
rlabel metal1 53 285 53 285 1 vssd1
port 5 n
rlabel metal1 62 1347 62 1347 1 vccd1
port 6 n
rlabel metal2 547 1796 547 1796 1 in
port 11 n
rlabel metal1 57 2203 57 2203 1 vssd1
port 5 n
rlabel viali 3337 441 3371 475 1 Y1
port 10 n
rlabel viali 3337 1743 3371 1777 1 Y0
port 9 n
<< end >>
