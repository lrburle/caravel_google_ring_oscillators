magic
tech sky130A
magscale 1 2
timestamp 1701971135
<< locali >>
rect 59 63 93 67
rect 0 49 161 63
rect 0 15 59 49
rect 93 15 161 49
rect 0 0 161 15
<< viali >>
rect 59 15 93 49
<< metal1 >>
rect 41 63 47 67
rect 0 9 47 63
rect 105 63 111 67
rect 105 9 161 63
rect 0 0 161 9
<< via1 >>
rect 47 49 105 67
rect 47 15 59 49
rect 59 15 93 49
rect 93 15 105 49
rect 47 9 105 15
<< metal2 >>
rect 38 67 114 76
rect 38 9 47 67
rect 105 9 114 67
rect 38 0 114 9
<< via2 >>
rect 47 9 105 67
<< metal3 >>
rect 0 67 161 76
rect 0 9 47 67
rect 105 9 161 67
rect 0 0 161 9
<< end >>
