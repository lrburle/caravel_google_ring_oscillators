// This is the unpowered netlist.
module mux16x1_project (io_out,
    io_in);
 output io_out;
 input [19:0] io_in;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__13__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__14__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__15__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__15__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__16__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__16__D1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__17__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__17__S (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__18__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__19__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__19__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__19__C (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__20__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__20__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__21__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__22__S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__22__S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__23__S0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__23__S1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__24__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__25__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__26__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_1481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__mux2_1 _13_ (.A0(net5),
    .A1(net7),
    .S(net12),
    .X(_00_));
 sky130_fd_sc_hd__and3b_1 _14_ (.A_N(net1),
    .B(net12),
    .C(net6),
    .X(_01_));
 sky130_fd_sc_hd__nor3b_1 _15_ (.A(net1),
    .B(net12),
    .C_N(net4),
    .Y(_02_));
 sky130_fd_sc_hd__a2111oi_1 _16_ (.A1(net1),
    .A2(_00_),
    .B1(_01_),
    .C1(_02_),
    .D1(net13),
    .Y(_03_));
 sky130_fd_sc_hd__mux2_1 _17_ (.A0(net9),
    .A1(net11),
    .S(net12),
    .X(_04_));
 sky130_fd_sc_hd__nand2_1 _18_ (.A(net1),
    .B(_04_),
    .Y(_05_));
 sky130_fd_sc_hd__nand3b_1 _19_ (.A_N(net1),
    .B(net12),
    .C(net10),
    .Y(_06_));
 sky130_fd_sc_hd__or3b_1 _20_ (.A(net1),
    .B(net12),
    .C_N(net8),
    .X(_07_));
 sky130_fd_sc_hd__a41o_1 _21_ (.A1(net13),
    .A2(_05_),
    .A3(_06_),
    .A4(_07_),
    .B1(_03_),
    .X(_08_));
 sky130_fd_sc_hd__mux4_1 _22_ (.A0(net16),
    .A1(net18),
    .A2(net20),
    .A3(net3),
    .S0(net12),
    .S1(net13),
    .X(_09_));
 sky130_fd_sc_hd__mux4_1 _23_ (.A0(net15),
    .A1(net17),
    .A2(net19),
    .A3(net2),
    .S0(net12),
    .S1(net13),
    .X(_10_));
 sky130_fd_sc_hd__mux2_1 _24_ (.A0(_10_),
    .A1(_09_),
    .S(net1),
    .X(_11_));
 sky130_fd_sc_hd__nor2_1 _25_ (.A(net14),
    .B(_11_),
    .Y(_12_));
 sky130_fd_sc_hd__a21oi_4 _26_ (.A1(net14),
    .A2(_08_),
    .B1(_12_),
    .Y(net21));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(io_in[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(io_in[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(io_in[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(io_in[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(io_in[3]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(io_in[4]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(io_in[5]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(io_in[6]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(io_in[7]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(io_in[8]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(io_in[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(io_in[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(io_in[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(io_in[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_out));
endmodule

