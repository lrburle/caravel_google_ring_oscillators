magic
tech sky130A
magscale 1 2
timestamp 1714141509
<< viali >>
rect 478943 431409 478977 431443
rect 485831 431409 485865 431443
rect 478581 410397 478615 410431
rect 485111 410397 485145 410431
rect 479474 389453 479508 389487
rect 490610 389453 490644 389487
rect 426541 373405 426575 373439
rect 477091 356813 477125 356847
rect 480143 356813 480177 356847
rect 482075 340833 482109 340867
rect 475442 340357 475476 340391
rect 478759 340357 478793 340391
rect 478939 320365 478973 320399
rect 485827 320365 485861 320399
rect 478580 305405 478614 305439
rect 485110 305405 485144 305439
rect 490610 285957 490644 285991
rect 479474 285821 479508 285855
rect 477101 265829 477135 265863
<< metal1 >>
rect 470234 451485 470854 451491
rect 470234 451433 470262 451485
rect 470314 451433 470326 451485
rect 470378 451433 470390 451485
rect 470442 451433 470454 451485
rect 470506 451433 470518 451485
rect 470570 451433 470582 451485
rect 470634 451433 470646 451485
rect 470698 451433 470710 451485
rect 470762 451433 470774 451485
rect 470826 451433 470854 451485
rect 470234 451421 470854 451433
rect 470234 451369 470262 451421
rect 470314 451369 470326 451421
rect 470378 451369 470390 451421
rect 470442 451369 470454 451421
rect 470506 451369 470518 451421
rect 470570 451369 470582 451421
rect 470634 451369 470646 451421
rect 470698 451369 470710 451421
rect 470762 451369 470774 451421
rect 470826 451369 470854 451421
rect 470234 451357 470854 451369
rect 470234 451305 470262 451357
rect 470314 451305 470326 451357
rect 470378 451305 470390 451357
rect 470442 451305 470454 451357
rect 470506 451305 470518 451357
rect 470570 451305 470582 451357
rect 470634 451305 470646 451357
rect 470698 451305 470710 451357
rect 470762 451305 470774 451357
rect 470826 451305 470854 451357
rect 470234 451293 470854 451305
rect 470234 451241 470262 451293
rect 470314 451241 470326 451293
rect 470378 451241 470390 451293
rect 470442 451241 470454 451293
rect 470506 451241 470518 451293
rect 470570 451241 470582 451293
rect 470634 451241 470646 451293
rect 470698 451241 470710 451293
rect 470762 451241 470774 451293
rect 470826 451241 470854 451293
rect 470234 451229 470854 451241
rect 470234 451177 470262 451229
rect 470314 451177 470326 451229
rect 470378 451177 470390 451229
rect 470442 451177 470454 451229
rect 470506 451177 470518 451229
rect 470570 451177 470582 451229
rect 470634 451177 470646 451229
rect 470698 451177 470710 451229
rect 470762 451177 470774 451229
rect 470826 451177 470854 451229
rect 470234 451171 470854 451177
rect 471330 450644 471336 450696
rect 471388 450684 471394 450696
rect 471388 450656 471652 450684
rect 471388 450644 471394 450656
rect 468994 450399 469614 450405
rect 468994 450347 469022 450399
rect 469074 450347 469086 450399
rect 469138 450347 469150 450399
rect 469202 450347 469214 450399
rect 469266 450347 469278 450399
rect 469330 450347 469342 450399
rect 469394 450347 469406 450399
rect 469458 450347 469470 450399
rect 469522 450347 469534 450399
rect 469586 450347 469614 450399
rect 468994 450335 469614 450347
rect 468994 450283 469022 450335
rect 469074 450283 469086 450335
rect 469138 450283 469150 450335
rect 469202 450283 469214 450335
rect 469266 450283 469278 450335
rect 469330 450283 469342 450335
rect 469394 450283 469406 450335
rect 469458 450283 469470 450335
rect 469522 450283 469534 450335
rect 469586 450283 469614 450335
rect 468994 450271 469614 450283
rect 468994 450219 469022 450271
rect 469074 450219 469086 450271
rect 469138 450219 469150 450271
rect 469202 450219 469214 450271
rect 469266 450219 469278 450271
rect 469330 450219 469342 450271
rect 469394 450219 469406 450271
rect 469458 450219 469470 450271
rect 469522 450219 469534 450271
rect 469586 450219 469614 450271
rect 468994 450207 469614 450219
rect 468994 450155 469022 450207
rect 469074 450155 469086 450207
rect 469138 450155 469150 450207
rect 469202 450155 469214 450207
rect 469266 450155 469278 450207
rect 469330 450155 469342 450207
rect 469394 450155 469406 450207
rect 469458 450155 469470 450207
rect 469522 450155 469534 450207
rect 469586 450155 469614 450207
rect 468994 450143 469614 450155
rect 468994 450091 469022 450143
rect 469074 450091 469086 450143
rect 469138 450091 469150 450143
rect 469202 450091 469214 450143
rect 469266 450091 469278 450143
rect 469330 450091 469342 450143
rect 469394 450091 469406 450143
rect 469458 450091 469470 450143
rect 469522 450091 469534 450143
rect 469586 450091 469614 450143
rect 468994 450085 469614 450091
rect 475378 449436 475384 449488
rect 475436 449436 475442 449488
rect 478690 449436 478696 449488
rect 478748 449436 478754 449488
rect 482002 449436 482008 449488
rect 482060 449436 482066 449488
rect 485314 449436 485320 449488
rect 485372 449436 485378 449488
rect 488644 449392 488672 449462
rect 491938 449392 491944 449404
rect 488644 449364 491944 449392
rect 491938 449352 491944 449364
rect 491996 449352 492002 449404
rect 470234 449314 470854 449320
rect 470234 449262 470262 449314
rect 470314 449262 470326 449314
rect 470378 449262 470390 449314
rect 470442 449262 470454 449314
rect 470506 449262 470518 449314
rect 470570 449262 470582 449314
rect 470634 449262 470646 449314
rect 470698 449262 470710 449314
rect 470762 449262 470774 449314
rect 470826 449262 470854 449314
rect 470234 449250 470854 449262
rect 470234 449198 470262 449250
rect 470314 449198 470326 449250
rect 470378 449198 470390 449250
rect 470442 449198 470454 449250
rect 470506 449198 470518 449250
rect 470570 449198 470582 449250
rect 470634 449198 470646 449250
rect 470698 449198 470710 449250
rect 470762 449198 470774 449250
rect 470826 449198 470854 449250
rect 470234 449186 470854 449198
rect 470234 449134 470262 449186
rect 470314 449134 470326 449186
rect 470378 449134 470390 449186
rect 470442 449134 470454 449186
rect 470506 449134 470518 449186
rect 470570 449134 470582 449186
rect 470634 449134 470646 449186
rect 470698 449134 470710 449186
rect 470762 449134 470774 449186
rect 470826 449134 470854 449186
rect 470234 449122 470854 449134
rect 470234 449070 470262 449122
rect 470314 449070 470326 449122
rect 470378 449070 470390 449122
rect 470442 449070 470454 449122
rect 470506 449070 470518 449122
rect 470570 449070 470582 449122
rect 470634 449070 470646 449122
rect 470698 449070 470710 449122
rect 470762 449070 470774 449122
rect 470826 449070 470854 449122
rect 470234 449058 470854 449070
rect 470234 449006 470262 449058
rect 470314 449006 470326 449058
rect 470378 449006 470390 449058
rect 470442 449006 470454 449058
rect 470506 449006 470518 449058
rect 470570 449006 470582 449058
rect 470634 449006 470646 449058
rect 470698 449006 470710 449058
rect 470762 449006 470774 449058
rect 470826 449006 470854 449058
rect 470234 449000 470854 449006
rect 478690 446224 478696 446276
rect 478748 446264 478754 446276
rect 478748 446236 480254 446264
rect 478748 446224 478754 446236
rect 480226 445924 480254 446236
rect 515398 445924 515404 445936
rect 480226 445896 515404 445924
rect 515398 445884 515404 445896
rect 515456 445884 515462 445936
rect 482002 445816 482008 445868
rect 482060 445816 482066 445868
rect 485314 445816 485320 445868
rect 485372 445856 485378 445868
rect 523678 445856 523684 445868
rect 485372 445828 523684 445856
rect 485372 445816 485378 445828
rect 523678 445816 523684 445828
rect 523736 445816 523742 445868
rect 482020 445788 482048 445816
rect 520918 445788 520924 445800
rect 482020 445760 520924 445788
rect 520918 445748 520924 445760
rect 520976 445748 520982 445800
rect 475378 445680 475384 445732
rect 475436 445720 475442 445732
rect 535454 445720 535460 445732
rect 475436 445692 535460 445720
rect 475436 445680 475442 445692
rect 535454 445680 535460 445692
rect 535512 445680 535518 445732
rect 490558 442960 490564 443012
rect 490616 443000 490622 443012
rect 535454 443000 535460 443012
rect 490616 442972 535460 443000
rect 490616 442960 490622 442972
rect 535454 442960 535460 442972
rect 535512 442960 535518 443012
rect 493318 441600 493324 441652
rect 493376 441640 493382 441652
rect 535454 441640 535460 441652
rect 493376 441612 535460 441640
rect 493376 441600 493382 441612
rect 535454 441600 535460 441612
rect 535512 441600 535518 441652
rect 494698 440240 494704 440292
rect 494756 440280 494762 440292
rect 535454 440280 535460 440292
rect 494756 440252 535460 440280
rect 494756 440240 494762 440252
rect 535454 440240 535460 440252
rect 535512 440240 535518 440292
rect 496078 438880 496084 438932
rect 496136 438920 496142 438932
rect 535454 438920 535460 438932
rect 496136 438892 535460 438920
rect 496136 438880 496142 438892
rect 535454 438880 535460 438892
rect 535512 438880 535518 438932
rect 497458 437452 497464 437504
rect 497516 437492 497522 437504
rect 535454 437492 535460 437504
rect 497516 437464 535460 437492
rect 497516 437452 497522 437464
rect 535454 437452 535460 437464
rect 535512 437452 535518 437504
rect 498838 436092 498844 436144
rect 498896 436132 498902 436144
rect 535454 436132 535460 436144
rect 498896 436104 535460 436132
rect 498896 436092 498902 436104
rect 535454 436092 535460 436104
rect 535512 436092 535518 436144
rect 500218 434732 500224 434784
rect 500276 434772 500282 434784
rect 535454 434772 535460 434784
rect 500276 434744 535460 434772
rect 500276 434732 500282 434744
rect 535454 434732 535460 434744
rect 535512 434732 535518 434784
rect 501598 433304 501604 433356
rect 501656 433344 501662 433356
rect 535454 433344 535460 433356
rect 501656 433316 535460 433344
rect 501656 433304 501662 433316
rect 535454 433304 535460 433316
rect 535512 433304 535518 433356
rect 470234 433086 470854 433092
rect 470234 433034 470262 433086
rect 470314 433034 470326 433086
rect 470378 433034 470390 433086
rect 470442 433034 470454 433086
rect 470506 433034 470518 433086
rect 470570 433034 470582 433086
rect 470634 433034 470646 433086
rect 470698 433034 470710 433086
rect 470762 433034 470774 433086
rect 470826 433034 470854 433086
rect 470234 433022 470854 433034
rect 470234 432970 470262 433022
rect 470314 432970 470326 433022
rect 470378 432970 470390 433022
rect 470442 432970 470454 433022
rect 470506 432970 470518 433022
rect 470570 432970 470582 433022
rect 470634 432970 470646 433022
rect 470698 432970 470710 433022
rect 470762 432970 470774 433022
rect 470826 432970 470854 433022
rect 470234 432958 470854 432970
rect 470234 432906 470262 432958
rect 470314 432906 470326 432958
rect 470378 432906 470390 432958
rect 470442 432906 470454 432958
rect 470506 432906 470518 432958
rect 470570 432906 470582 432958
rect 470634 432906 470646 432958
rect 470698 432906 470710 432958
rect 470762 432906 470774 432958
rect 470826 432906 470854 432958
rect 470234 432894 470854 432906
rect 470234 432842 470262 432894
rect 470314 432842 470326 432894
rect 470378 432842 470390 432894
rect 470442 432842 470454 432894
rect 470506 432842 470518 432894
rect 470570 432842 470582 432894
rect 470634 432842 470646 432894
rect 470698 432842 470710 432894
rect 470762 432842 470774 432894
rect 470826 432842 470854 432894
rect 470234 432830 470854 432842
rect 470234 432778 470262 432830
rect 470314 432778 470326 432830
rect 470378 432778 470390 432830
rect 470442 432778 470454 432830
rect 470506 432778 470518 432830
rect 470570 432778 470582 432830
rect 470634 432778 470646 432830
rect 470698 432778 470710 432830
rect 470762 432778 470774 432830
rect 470826 432778 470854 432830
rect 470234 432772 470854 432778
rect 471612 432290 471664 432296
rect 471612 432232 471664 432238
rect 468994 431999 469614 432005
rect 468994 431947 469022 431999
rect 469074 431947 469086 431999
rect 469138 431947 469150 431999
rect 469202 431947 469214 431999
rect 469266 431947 469278 431999
rect 469330 431947 469342 431999
rect 469394 431947 469406 431999
rect 469458 431947 469470 431999
rect 469522 431947 469534 431999
rect 469586 431947 469614 431999
rect 468994 431935 469614 431947
rect 502978 431944 502984 431996
rect 503036 431984 503042 431996
rect 535454 431984 535460 431996
rect 503036 431956 535460 431984
rect 503036 431944 503042 431956
rect 535454 431944 535460 431956
rect 535512 431944 535518 431996
rect 468994 431883 469022 431935
rect 469074 431883 469086 431935
rect 469138 431883 469150 431935
rect 469202 431883 469214 431935
rect 469266 431883 469278 431935
rect 469330 431883 469342 431935
rect 469394 431883 469406 431935
rect 469458 431883 469470 431935
rect 469522 431883 469534 431935
rect 469586 431883 469614 431935
rect 468994 431871 469614 431883
rect 468994 431819 469022 431871
rect 469074 431819 469086 431871
rect 469138 431819 469150 431871
rect 469202 431819 469214 431871
rect 469266 431819 469278 431871
rect 469330 431819 469342 431871
rect 469394 431819 469406 431871
rect 469458 431819 469470 431871
rect 469522 431819 469534 431871
rect 469586 431819 469614 431871
rect 468994 431807 469614 431819
rect 468994 431755 469022 431807
rect 469074 431755 469086 431807
rect 469138 431755 469150 431807
rect 469202 431755 469214 431807
rect 469266 431755 469278 431807
rect 469330 431755 469342 431807
rect 469394 431755 469406 431807
rect 469458 431755 469470 431807
rect 469522 431755 469534 431807
rect 469586 431755 469614 431807
rect 468994 431743 469614 431755
rect 468994 431691 469022 431743
rect 469074 431691 469086 431743
rect 469138 431691 469150 431743
rect 469202 431691 469214 431743
rect 469266 431691 469278 431743
rect 469330 431691 469342 431743
rect 469394 431691 469406 431743
rect 469458 431691 469470 431743
rect 469522 431691 469534 431743
rect 469586 431691 469614 431743
rect 468994 431685 469614 431691
rect 478966 431449 478972 431452
rect 478931 431443 478972 431449
rect 478931 431409 478943 431443
rect 478931 431403 478972 431409
rect 478966 431400 478972 431403
rect 479024 431400 479030 431452
rect 485774 431400 485780 431452
rect 485832 431449 485838 431452
rect 485832 431443 485877 431449
rect 485865 431409 485877 431443
rect 485832 431403 485877 431409
rect 485832 431400 485838 431403
rect 475470 431035 475476 431087
rect 475528 431035 475534 431087
rect 482370 431035 482376 431087
rect 482428 431035 482434 431087
rect 489302 431047 489592 431075
rect 489564 431032 489592 431047
rect 492030 431032 492036 431044
rect 489564 431004 492036 431032
rect 492030 430992 492036 431004
rect 492088 430992 492094 431044
rect 470234 430914 470854 430920
rect 470234 430862 470262 430914
rect 470314 430862 470326 430914
rect 470378 430862 470390 430914
rect 470442 430862 470454 430914
rect 470506 430862 470518 430914
rect 470570 430862 470582 430914
rect 470634 430862 470646 430914
rect 470698 430862 470710 430914
rect 470762 430862 470774 430914
rect 470826 430862 470854 430914
rect 470234 430850 470854 430862
rect 470234 430798 470262 430850
rect 470314 430798 470326 430850
rect 470378 430798 470390 430850
rect 470442 430798 470454 430850
rect 470506 430798 470518 430850
rect 470570 430798 470582 430850
rect 470634 430798 470646 430850
rect 470698 430798 470710 430850
rect 470762 430798 470774 430850
rect 470826 430798 470854 430850
rect 470234 430786 470854 430798
rect 470234 430734 470262 430786
rect 470314 430734 470326 430786
rect 470378 430734 470390 430786
rect 470442 430734 470454 430786
rect 470506 430734 470518 430786
rect 470570 430734 470582 430786
rect 470634 430734 470646 430786
rect 470698 430734 470710 430786
rect 470762 430734 470774 430786
rect 470826 430734 470854 430786
rect 470234 430722 470854 430734
rect 470234 430670 470262 430722
rect 470314 430670 470326 430722
rect 470378 430670 470390 430722
rect 470442 430670 470454 430722
rect 470506 430670 470518 430722
rect 470570 430670 470582 430722
rect 470634 430670 470646 430722
rect 470698 430670 470710 430722
rect 470762 430670 470774 430722
rect 470826 430670 470854 430722
rect 470234 430658 470854 430670
rect 470234 430606 470262 430658
rect 470314 430606 470326 430658
rect 470378 430606 470390 430658
rect 470442 430606 470454 430658
rect 470506 430606 470518 430658
rect 470570 430606 470582 430658
rect 470634 430606 470646 430658
rect 470698 430606 470710 430658
rect 470762 430606 470774 430658
rect 470826 430606 470854 430658
rect 470234 430600 470854 430606
rect 475470 429088 475476 429140
rect 475528 429128 475534 429140
rect 490558 429128 490564 429140
rect 475528 429100 490564 429128
rect 475528 429088 475534 429100
rect 490558 429088 490564 429100
rect 490616 429088 490622 429140
rect 482370 427796 482376 427848
rect 482428 427836 482434 427848
rect 522298 427836 522304 427848
rect 482428 427808 522304 427836
rect 482428 427796 482434 427808
rect 522298 427796 522304 427808
rect 522356 427796 522362 427848
rect 470234 412086 470854 412092
rect 470234 412034 470262 412086
rect 470314 412034 470326 412086
rect 470378 412034 470390 412086
rect 470442 412034 470454 412086
rect 470506 412034 470518 412086
rect 470570 412034 470582 412086
rect 470634 412034 470646 412086
rect 470698 412034 470710 412086
rect 470762 412034 470774 412086
rect 470826 412034 470854 412086
rect 470234 412022 470854 412034
rect 470234 411970 470262 412022
rect 470314 411970 470326 412022
rect 470378 411970 470390 412022
rect 470442 411970 470454 412022
rect 470506 411970 470518 412022
rect 470570 411970 470582 412022
rect 470634 411970 470646 412022
rect 470698 411970 470710 412022
rect 470762 411970 470774 412022
rect 470826 411970 470854 412022
rect 470234 411958 470854 411970
rect 470234 411906 470262 411958
rect 470314 411906 470326 411958
rect 470378 411906 470390 411958
rect 470442 411906 470454 411958
rect 470506 411906 470518 411958
rect 470570 411906 470582 411958
rect 470634 411906 470646 411958
rect 470698 411906 470710 411958
rect 470762 411906 470774 411958
rect 470826 411906 470854 411958
rect 470234 411894 470854 411906
rect 470234 411842 470262 411894
rect 470314 411842 470326 411894
rect 470378 411842 470390 411894
rect 470442 411842 470454 411894
rect 470506 411842 470518 411894
rect 470570 411842 470582 411894
rect 470634 411842 470646 411894
rect 470698 411842 470710 411894
rect 470762 411842 470774 411894
rect 470826 411842 470854 411894
rect 470234 411830 470854 411842
rect 470234 411778 470262 411830
rect 470314 411778 470326 411830
rect 470378 411778 470390 411830
rect 470442 411778 470454 411830
rect 470506 411778 470518 411830
rect 470570 411778 470582 411830
rect 470634 411778 470646 411830
rect 470698 411778 470710 411830
rect 470762 411778 470774 411830
rect 470826 411778 470854 411830
rect 470234 411772 470854 411778
rect 471238 411204 471244 411256
rect 471296 411244 471302 411256
rect 471624 411244 471652 411263
rect 471296 411216 471652 411244
rect 473722 411232 473728 411284
rect 473780 411232 473786 411284
rect 471296 411204 471302 411216
rect 468994 411000 469614 411006
rect 468994 410948 469022 411000
rect 469074 410948 469086 411000
rect 469138 410948 469150 411000
rect 469202 410948 469214 411000
rect 469266 410948 469278 411000
rect 469330 410948 469342 411000
rect 469394 410948 469406 411000
rect 469458 410948 469470 411000
rect 469522 410948 469534 411000
rect 469586 410948 469614 411000
rect 468994 410936 469614 410948
rect 468994 410884 469022 410936
rect 469074 410884 469086 410936
rect 469138 410884 469150 410936
rect 469202 410884 469214 410936
rect 469266 410884 469278 410936
rect 469330 410884 469342 410936
rect 469394 410884 469406 410936
rect 469458 410884 469470 410936
rect 469522 410884 469534 410936
rect 469586 410884 469614 410936
rect 468994 410872 469614 410884
rect 468994 410820 469022 410872
rect 469074 410820 469086 410872
rect 469138 410820 469150 410872
rect 469202 410820 469214 410872
rect 469266 410820 469278 410872
rect 469330 410820 469342 410872
rect 469394 410820 469406 410872
rect 469458 410820 469470 410872
rect 469522 410820 469534 410872
rect 469586 410820 469614 410872
rect 468994 410808 469614 410820
rect 468994 410756 469022 410808
rect 469074 410756 469086 410808
rect 469138 410756 469150 410808
rect 469202 410756 469214 410808
rect 469266 410756 469278 410808
rect 469330 410756 469342 410808
rect 469394 410756 469406 410808
rect 469458 410756 469470 410808
rect 469522 410756 469534 410808
rect 469586 410756 469614 410808
rect 468994 410744 469614 410756
rect 468994 410692 469022 410744
rect 469074 410692 469086 410744
rect 469138 410692 469150 410744
rect 469202 410692 469214 410744
rect 469266 410692 469278 410744
rect 469330 410692 469342 410744
rect 469394 410692 469406 410744
rect 469458 410692 469470 410744
rect 469522 410692 469534 410744
rect 469586 410692 469614 410744
rect 468994 410686 469614 410692
rect 478414 410428 478420 410440
rect 477788 410400 478420 410428
rect 478414 410388 478420 410400
rect 478472 410388 478478 410440
rect 478598 410437 478604 410440
rect 478569 410431 478604 410437
rect 478569 410397 478581 410431
rect 478569 410391 478604 410397
rect 478598 410388 478604 410391
rect 478656 410388 478662 410440
rect 485130 410437 485136 410440
rect 485099 410431 485136 410437
rect 485099 410397 485111 410431
rect 485099 410391 485136 410397
rect 485130 410388 485136 410391
rect 485188 410388 485194 410440
rect 475286 410036 475292 410088
rect 475344 410036 475350 410088
rect 481818 410036 481824 410088
rect 481876 410036 481882 410088
rect 488382 410048 488672 410076
rect 488644 410020 488672 410048
rect 490742 410020 490748 410032
rect 488644 409992 490748 410020
rect 490742 409980 490748 409992
rect 490800 409980 490806 410032
rect 470234 409914 470854 409920
rect 470234 409862 470262 409914
rect 470314 409862 470326 409914
rect 470378 409862 470390 409914
rect 470442 409862 470454 409914
rect 470506 409862 470518 409914
rect 470570 409862 470582 409914
rect 470634 409862 470646 409914
rect 470698 409862 470710 409914
rect 470762 409862 470774 409914
rect 470826 409862 470854 409914
rect 470234 409850 470854 409862
rect 470234 409798 470262 409850
rect 470314 409798 470326 409850
rect 470378 409798 470390 409850
rect 470442 409798 470454 409850
rect 470506 409798 470518 409850
rect 470570 409798 470582 409850
rect 470634 409798 470646 409850
rect 470698 409798 470710 409850
rect 470762 409798 470774 409850
rect 470826 409798 470854 409850
rect 470234 409786 470854 409798
rect 470234 409734 470262 409786
rect 470314 409734 470326 409786
rect 470378 409734 470390 409786
rect 470442 409734 470454 409786
rect 470506 409734 470518 409786
rect 470570 409734 470582 409786
rect 470634 409734 470646 409786
rect 470698 409734 470710 409786
rect 470762 409734 470774 409786
rect 470826 409734 470854 409786
rect 515398 409776 515404 409828
rect 515456 409816 515462 409828
rect 535454 409816 535460 409828
rect 515456 409788 535460 409816
rect 515456 409776 515462 409788
rect 535454 409776 535460 409788
rect 535512 409776 535518 409828
rect 470234 409722 470854 409734
rect 470234 409670 470262 409722
rect 470314 409670 470326 409722
rect 470378 409670 470390 409722
rect 470442 409670 470454 409722
rect 470506 409670 470518 409722
rect 470570 409670 470582 409722
rect 470634 409670 470646 409722
rect 470698 409670 470710 409722
rect 470762 409670 470774 409722
rect 470826 409670 470854 409722
rect 470234 409658 470854 409670
rect 470234 409606 470262 409658
rect 470314 409606 470326 409658
rect 470378 409606 470390 409658
rect 470442 409606 470454 409658
rect 470506 409606 470518 409658
rect 470570 409606 470582 409658
rect 470634 409606 470646 409658
rect 470698 409606 470710 409658
rect 470762 409606 470774 409658
rect 470826 409606 470854 409658
rect 470234 409600 470854 409606
rect 475286 408416 475292 408468
rect 475344 408456 475350 408468
rect 493318 408456 493324 408468
rect 475344 408428 493324 408456
rect 475344 408416 475350 408428
rect 493318 408416 493324 408428
rect 493376 408416 493382 408468
rect 478598 407056 478604 407108
rect 478656 407096 478662 407108
rect 535454 407096 535460 407108
rect 478656 407068 535460 407096
rect 478656 407056 478662 407068
rect 535454 407056 535460 407068
rect 535512 407056 535518 407108
rect 515398 404336 515404 404388
rect 515456 404376 515462 404388
rect 535454 404376 535460 404388
rect 515456 404348 535460 404376
rect 515456 404336 515462 404348
rect 535454 404336 535460 404348
rect 535512 404336 535518 404388
rect 516778 402976 516784 403028
rect 516836 403016 516842 403028
rect 535454 403016 535460 403028
rect 516836 402988 535460 403016
rect 516836 402976 516842 402988
rect 535454 402976 535460 402988
rect 535512 402976 535518 403028
rect 518158 398828 518164 398880
rect 518216 398868 518222 398880
rect 535454 398868 535460 398880
rect 518216 398840 535460 398868
rect 518216 398828 518222 398840
rect 535454 398828 535460 398840
rect 535512 398828 535518 398880
rect 519538 396040 519544 396092
rect 519596 396080 519602 396092
rect 535454 396080 535460 396092
rect 519596 396052 535460 396080
rect 519596 396040 519602 396052
rect 535454 396040 535460 396052
rect 535512 396040 535518 396092
rect 470234 391087 470854 391093
rect 470234 391035 470262 391087
rect 470314 391035 470326 391087
rect 470378 391035 470390 391087
rect 470442 391035 470454 391087
rect 470506 391035 470518 391087
rect 470570 391035 470582 391087
rect 470634 391035 470646 391087
rect 470698 391035 470710 391087
rect 470762 391035 470774 391087
rect 470826 391035 470854 391087
rect 470234 391023 470854 391035
rect 470234 390971 470262 391023
rect 470314 390971 470326 391023
rect 470378 390971 470390 391023
rect 470442 390971 470454 391023
rect 470506 390971 470518 391023
rect 470570 390971 470582 391023
rect 470634 390971 470646 391023
rect 470698 390971 470710 391023
rect 470762 390971 470774 391023
rect 470826 390971 470854 391023
rect 470234 390959 470854 390971
rect 470234 390907 470262 390959
rect 470314 390907 470326 390959
rect 470378 390907 470390 390959
rect 470442 390907 470454 390959
rect 470506 390907 470518 390959
rect 470570 390907 470582 390959
rect 470634 390907 470646 390959
rect 470698 390907 470710 390959
rect 470762 390907 470774 390959
rect 470826 390907 470854 390959
rect 470234 390895 470854 390907
rect 470234 390843 470262 390895
rect 470314 390843 470326 390895
rect 470378 390843 470390 390895
rect 470442 390843 470454 390895
rect 470506 390843 470518 390895
rect 470570 390843 470582 390895
rect 470634 390843 470646 390895
rect 470698 390843 470710 390895
rect 470762 390843 470774 390895
rect 470826 390843 470854 390895
rect 470234 390831 470854 390843
rect 470234 390779 470262 390831
rect 470314 390779 470326 390831
rect 470378 390779 470390 390831
rect 470442 390779 470454 390831
rect 470506 390779 470518 390831
rect 470570 390779 470582 390831
rect 470634 390779 470646 390831
rect 470698 390779 470710 390831
rect 470762 390779 470774 390831
rect 470826 390779 470854 390831
rect 470234 390773 470854 390779
rect 471238 390260 471244 390312
rect 471296 390300 471302 390312
rect 471296 390272 471652 390300
rect 471296 390260 471302 390272
rect 471624 390096 471652 390272
rect 471698 390096 471704 390108
rect 471624 390068 471704 390096
rect 471698 390056 471704 390068
rect 471756 390056 471762 390108
rect 468994 390004 469614 390010
rect 468994 389952 469022 390004
rect 469074 389952 469086 390004
rect 469138 389952 469150 390004
rect 469202 389952 469214 390004
rect 469266 389952 469278 390004
rect 469330 389952 469342 390004
rect 469394 389952 469406 390004
rect 469458 389952 469470 390004
rect 469522 389952 469534 390004
rect 469586 389952 469614 390004
rect 468994 389940 469614 389952
rect 468994 389888 469022 389940
rect 469074 389888 469086 389940
rect 469138 389888 469150 389940
rect 469202 389888 469214 389940
rect 469266 389888 469278 389940
rect 469330 389888 469342 389940
rect 469394 389888 469406 389940
rect 469458 389888 469470 389940
rect 469522 389888 469534 389940
rect 469586 389888 469614 389940
rect 468994 389876 469614 389888
rect 468994 389824 469022 389876
rect 469074 389824 469086 389876
rect 469138 389824 469150 389876
rect 469202 389824 469214 389876
rect 469266 389824 469278 389876
rect 469330 389824 469342 389876
rect 469394 389824 469406 389876
rect 469458 389824 469470 389876
rect 469522 389824 469534 389876
rect 469586 389824 469614 389876
rect 468994 389812 469614 389824
rect 468994 389760 469022 389812
rect 469074 389760 469086 389812
rect 469138 389760 469150 389812
rect 469202 389760 469214 389812
rect 469266 389760 469278 389812
rect 469330 389760 469342 389812
rect 469394 389760 469406 389812
rect 469458 389760 469470 389812
rect 469522 389760 469534 389812
rect 469586 389760 469614 389812
rect 468994 389748 469614 389760
rect 468994 389696 469022 389748
rect 469074 389696 469086 389748
rect 469138 389696 469150 389748
rect 469202 389696 469214 389748
rect 469266 389696 469278 389748
rect 469330 389696 469342 389748
rect 469394 389696 469406 389748
rect 469458 389696 469470 389748
rect 469522 389696 469534 389748
rect 469586 389696 469614 389748
rect 468994 389690 469614 389696
rect 479426 389444 479432 389496
rect 479484 389493 479490 389496
rect 479484 389487 479520 389493
rect 479508 389453 479520 389487
rect 479484 389447 479520 389453
rect 490598 389487 490656 389493
rect 490598 389453 490610 389487
rect 490644 389484 490656 389487
rect 493318 389484 493324 389496
rect 490644 389456 493324 389484
rect 490644 389453 490656 389456
rect 490598 389447 490656 389453
rect 479484 389444 479490 389447
rect 493318 389444 493324 389456
rect 493376 389444 493382 389496
rect 475746 389036 475752 389088
rect 475804 389036 475810 389088
rect 483198 389036 483204 389088
rect 483256 389036 483262 389088
rect 486878 389036 486884 389088
rect 486936 389036 486942 389088
rect 470234 388914 470854 388920
rect 470234 388862 470262 388914
rect 470314 388862 470326 388914
rect 470378 388862 470390 388914
rect 470442 388862 470454 388914
rect 470506 388862 470518 388914
rect 470570 388862 470582 388914
rect 470634 388862 470646 388914
rect 470698 388862 470710 388914
rect 470762 388862 470774 388914
rect 470826 388862 470854 388914
rect 470234 388850 470854 388862
rect 470234 388798 470262 388850
rect 470314 388798 470326 388850
rect 470378 388798 470390 388850
rect 470442 388798 470454 388850
rect 470506 388798 470518 388850
rect 470570 388798 470582 388850
rect 470634 388798 470646 388850
rect 470698 388798 470710 388850
rect 470762 388798 470774 388850
rect 470826 388798 470854 388850
rect 470234 388786 470854 388798
rect 470234 388734 470262 388786
rect 470314 388734 470326 388786
rect 470378 388734 470390 388786
rect 470442 388734 470454 388786
rect 470506 388734 470518 388786
rect 470570 388734 470582 388786
rect 470634 388734 470646 388786
rect 470698 388734 470710 388786
rect 470762 388734 470774 388786
rect 470826 388734 470854 388786
rect 470234 388722 470854 388734
rect 470234 388670 470262 388722
rect 470314 388670 470326 388722
rect 470378 388670 470390 388722
rect 470442 388670 470454 388722
rect 470506 388670 470518 388722
rect 470570 388670 470582 388722
rect 470634 388670 470646 388722
rect 470698 388670 470710 388722
rect 470762 388670 470774 388722
rect 470826 388670 470854 388722
rect 470234 388658 470854 388670
rect 470234 388606 470262 388658
rect 470314 388606 470326 388658
rect 470378 388606 470390 388658
rect 470442 388606 470454 388658
rect 470506 388606 470518 388658
rect 470570 388606 470582 388658
rect 470634 388606 470646 388658
rect 470698 388606 470710 388658
rect 470762 388606 470774 388658
rect 470826 388606 470854 388658
rect 470234 388600 470854 388606
rect 475746 387744 475752 387796
rect 475804 387744 475810 387796
rect 479426 387744 479432 387796
rect 479484 387784 479490 387796
rect 515398 387784 515404 387796
rect 479484 387756 515404 387784
rect 479484 387744 479490 387756
rect 515398 387744 515404 387756
rect 515456 387744 515462 387796
rect 475764 387716 475792 387744
rect 494698 387716 494704 387728
rect 475764 387688 494704 387716
rect 494698 387676 494704 387688
rect 494756 387676 494762 387728
rect 483198 386384 483204 386436
rect 483256 386424 483262 386436
rect 484302 386424 484308 386436
rect 483256 386396 484308 386424
rect 483256 386384 483262 386396
rect 484302 386384 484308 386396
rect 484360 386384 484366 386436
rect 520918 373940 520924 373992
rect 520976 373980 520982 373992
rect 535454 373980 535460 373992
rect 520976 373952 535460 373980
rect 520976 373940 520982 373952
rect 535454 373940 535460 373952
rect 535512 373940 535518 373992
rect 426529 373439 426587 373445
rect 426529 373405 426541 373439
rect 426575 373436 426587 373439
rect 536190 373436 536196 373448
rect 426575 373408 536196 373436
rect 426575 373405 426587 373408
rect 426529 373399 426587 373405
rect 536190 373396 536196 373408
rect 536248 373396 536254 373448
rect 522298 372512 522304 372564
rect 522356 372552 522362 372564
rect 535454 372552 535460 372564
rect 522356 372524 535460 372552
rect 522356 372512 522362 372524
rect 535454 372512 535460 372524
rect 535512 372512 535518 372564
rect 484302 369792 484308 369844
rect 484360 369832 484366 369844
rect 535454 369832 535460 369844
rect 484360 369804 535460 369832
rect 484360 369792 484366 369804
rect 535454 369792 535460 369804
rect 535512 369792 535518 369844
rect 520918 367072 520924 367124
rect 520976 367112 520982 367124
rect 535454 367112 535460 367124
rect 520976 367084 535460 367112
rect 520976 367072 520982 367084
rect 535454 367072 535460 367084
rect 535512 367072 535518 367124
rect 515398 365712 515404 365764
rect 515456 365752 515462 365764
rect 535454 365752 535460 365764
rect 515456 365724 535460 365752
rect 515456 365712 515462 365724
rect 535454 365712 535460 365724
rect 535512 365712 535518 365764
rect 522298 361564 522304 361616
rect 522356 361604 522362 361616
rect 535454 361604 535460 361616
rect 522356 361576 535460 361604
rect 522356 361564 522362 361576
rect 535454 361564 535460 361576
rect 535512 361564 535518 361616
rect 470234 358487 470854 358493
rect 470234 358435 470262 358487
rect 470314 358435 470326 358487
rect 470378 358435 470390 358487
rect 470442 358435 470454 358487
rect 470506 358435 470518 358487
rect 470570 358435 470582 358487
rect 470634 358435 470646 358487
rect 470698 358435 470710 358487
rect 470762 358435 470774 358487
rect 470826 358435 470854 358487
rect 470234 358423 470854 358435
rect 470234 358371 470262 358423
rect 470314 358371 470326 358423
rect 470378 358371 470390 358423
rect 470442 358371 470454 358423
rect 470506 358371 470518 358423
rect 470570 358371 470582 358423
rect 470634 358371 470646 358423
rect 470698 358371 470710 358423
rect 470762 358371 470774 358423
rect 470826 358371 470854 358423
rect 470234 358359 470854 358371
rect 470234 358307 470262 358359
rect 470314 358307 470326 358359
rect 470378 358307 470390 358359
rect 470442 358307 470454 358359
rect 470506 358307 470518 358359
rect 470570 358307 470582 358359
rect 470634 358307 470646 358359
rect 470698 358307 470710 358359
rect 470762 358307 470774 358359
rect 470826 358307 470854 358359
rect 470234 358295 470854 358307
rect 470234 358243 470262 358295
rect 470314 358243 470326 358295
rect 470378 358243 470390 358295
rect 470442 358243 470454 358295
rect 470506 358243 470518 358295
rect 470570 358243 470582 358295
rect 470634 358243 470646 358295
rect 470698 358243 470710 358295
rect 470762 358243 470774 358295
rect 470826 358243 470854 358295
rect 470234 358231 470854 358243
rect 470234 358179 470262 358231
rect 470314 358179 470326 358231
rect 470378 358179 470390 358231
rect 470442 358179 470454 358231
rect 470506 358179 470518 358231
rect 470570 358179 470582 358231
rect 470634 358179 470646 358231
rect 470698 358179 470710 358231
rect 470762 358179 470774 358231
rect 470826 358179 470854 358231
rect 470234 358173 470854 358179
rect 471698 357552 471704 357604
rect 471756 357592 471762 357604
rect 473648 357592 473676 357664
rect 475102 357620 475108 357672
rect 475160 357620 475166 357672
rect 478874 357631 478880 357683
rect 478932 357631 478938 357683
rect 481818 357631 481824 357683
rect 481876 357631 481882 357683
rect 484946 357631 484952 357683
rect 485004 357631 485010 357683
rect 471756 357564 473676 357592
rect 471756 357552 471762 357564
rect 468994 357401 469614 357407
rect 468994 357349 469022 357401
rect 469074 357349 469086 357401
rect 469138 357349 469150 357401
rect 469202 357349 469214 357401
rect 469266 357349 469278 357401
rect 469330 357349 469342 357401
rect 469394 357349 469406 357401
rect 469458 357349 469470 357401
rect 469522 357349 469534 357401
rect 469586 357349 469614 357401
rect 468994 357337 469614 357349
rect 468994 357285 469022 357337
rect 469074 357285 469086 357337
rect 469138 357285 469150 357337
rect 469202 357285 469214 357337
rect 469266 357285 469278 357337
rect 469330 357285 469342 357337
rect 469394 357285 469406 357337
rect 469458 357285 469470 357337
rect 469522 357285 469534 357337
rect 469586 357285 469614 357337
rect 468994 357273 469614 357285
rect 468994 357221 469022 357273
rect 469074 357221 469086 357273
rect 469138 357221 469150 357273
rect 469202 357221 469214 357273
rect 469266 357221 469278 357273
rect 469330 357221 469342 357273
rect 469394 357221 469406 357273
rect 469458 357221 469470 357273
rect 469522 357221 469534 357273
rect 469586 357221 469614 357273
rect 468994 357209 469614 357221
rect 468994 357157 469022 357209
rect 469074 357157 469086 357209
rect 469138 357157 469150 357209
rect 469202 357157 469214 357209
rect 469266 357157 469278 357209
rect 469330 357157 469342 357209
rect 469394 357157 469406 357209
rect 469458 357157 469470 357209
rect 469522 357157 469534 357209
rect 469586 357157 469614 357209
rect 468994 357145 469614 357157
rect 468994 357093 469022 357145
rect 469074 357093 469086 357145
rect 469138 357093 469150 357145
rect 469202 357093 469214 357145
rect 469266 357093 469278 357145
rect 469330 357093 469342 357145
rect 469394 357093 469406 357145
rect 469458 357093 469470 357145
rect 469522 357093 469534 357145
rect 469586 357093 469614 357145
rect 468994 357087 469614 357093
rect 477034 356804 477040 356856
rect 477092 356853 477098 356856
rect 480162 356853 480168 356856
rect 477092 356847 477137 356853
rect 477125 356813 477137 356847
rect 477092 356807 477137 356813
rect 480131 356847 480168 356853
rect 480131 356813 480143 356847
rect 480131 356807 480168 356813
rect 477092 356804 477098 356807
rect 480162 356804 480168 356807
rect 480220 356804 480226 356856
rect 483198 356435 483204 356487
rect 483256 356435 483262 356487
rect 486234 356435 486240 356487
rect 486292 356435 486298 356487
rect 489288 356436 489316 356461
rect 492122 356436 492128 356448
rect 489288 356408 492128 356436
rect 492122 356396 492128 356408
rect 492180 356396 492186 356448
rect 470234 356314 470854 356320
rect 470234 356262 470262 356314
rect 470314 356262 470326 356314
rect 470378 356262 470390 356314
rect 470442 356262 470454 356314
rect 470506 356262 470518 356314
rect 470570 356262 470582 356314
rect 470634 356262 470646 356314
rect 470698 356262 470710 356314
rect 470762 356262 470774 356314
rect 470826 356262 470854 356314
rect 470234 356250 470854 356262
rect 470234 356198 470262 356250
rect 470314 356198 470326 356250
rect 470378 356198 470390 356250
rect 470442 356198 470454 356250
rect 470506 356198 470518 356250
rect 470570 356198 470582 356250
rect 470634 356198 470646 356250
rect 470698 356198 470710 356250
rect 470762 356198 470774 356250
rect 470826 356198 470854 356250
rect 470234 356186 470854 356198
rect 470234 356134 470262 356186
rect 470314 356134 470326 356186
rect 470378 356134 470390 356186
rect 470442 356134 470454 356186
rect 470506 356134 470518 356186
rect 470570 356134 470582 356186
rect 470634 356134 470646 356186
rect 470698 356134 470710 356186
rect 470762 356134 470774 356186
rect 470826 356134 470854 356186
rect 470234 356122 470854 356134
rect 470234 356070 470262 356122
rect 470314 356070 470326 356122
rect 470378 356070 470390 356122
rect 470442 356070 470454 356122
rect 470506 356070 470518 356122
rect 470570 356070 470582 356122
rect 470634 356070 470646 356122
rect 470698 356070 470710 356122
rect 470762 356070 470774 356122
rect 470826 356070 470854 356122
rect 470234 356058 470854 356070
rect 470234 356006 470262 356058
rect 470314 356006 470326 356058
rect 470378 356006 470390 356058
rect 470442 356006 470454 356058
rect 470506 356006 470518 356058
rect 470570 356006 470582 356058
rect 470634 356006 470646 356058
rect 470698 356006 470710 356058
rect 470762 356006 470774 356058
rect 470826 356006 470854 356058
rect 470234 356000 470854 356006
rect 480162 354628 480168 354680
rect 480220 354668 480226 354680
rect 516778 354668 516784 354680
rect 480220 354640 516784 354668
rect 480220 354628 480226 354640
rect 516778 354628 516784 354640
rect 516836 354628 516842 354680
rect 483198 354560 483204 354612
rect 483256 354600 483262 354612
rect 520918 354600 520924 354612
rect 483256 354572 520924 354600
rect 483256 354560 483262 354572
rect 520918 354560 520924 354572
rect 520976 354560 520982 354612
rect 477126 354492 477132 354544
rect 477184 354532 477190 354544
rect 496078 354532 496084 354544
rect 477184 354504 496084 354532
rect 477184 354492 477190 354504
rect 496078 354492 496084 354504
rect 496136 354492 496142 354544
rect 486234 353608 486240 353660
rect 486292 353648 486298 353660
rect 486292 353620 489914 353648
rect 486292 353608 486298 353620
rect 489886 353308 489914 353620
rect 525058 353308 525064 353320
rect 489886 353280 525064 353308
rect 525058 353268 525064 353280
rect 525116 353268 525122 353320
rect 470234 342486 470854 342492
rect 470234 342434 470262 342486
rect 470314 342434 470326 342486
rect 470378 342434 470390 342486
rect 470442 342434 470454 342486
rect 470506 342434 470518 342486
rect 470570 342434 470582 342486
rect 470634 342434 470646 342486
rect 470698 342434 470710 342486
rect 470762 342434 470774 342486
rect 470826 342434 470854 342486
rect 470234 342422 470854 342434
rect 470234 342370 470262 342422
rect 470314 342370 470326 342422
rect 470378 342370 470390 342422
rect 470442 342370 470454 342422
rect 470506 342370 470518 342422
rect 470570 342370 470582 342422
rect 470634 342370 470646 342422
rect 470698 342370 470710 342422
rect 470762 342370 470774 342422
rect 470826 342370 470854 342422
rect 470234 342358 470854 342370
rect 470234 342306 470262 342358
rect 470314 342306 470326 342358
rect 470378 342306 470390 342358
rect 470442 342306 470454 342358
rect 470506 342306 470518 342358
rect 470570 342306 470582 342358
rect 470634 342306 470646 342358
rect 470698 342306 470710 342358
rect 470762 342306 470774 342358
rect 470826 342306 470854 342358
rect 470234 342294 470854 342306
rect 470234 342242 470262 342294
rect 470314 342242 470326 342294
rect 470378 342242 470390 342294
rect 470442 342242 470454 342294
rect 470506 342242 470518 342294
rect 470570 342242 470582 342294
rect 470634 342242 470646 342294
rect 470698 342242 470710 342294
rect 470762 342242 470774 342294
rect 470826 342242 470854 342294
rect 470234 342230 470854 342242
rect 470234 342178 470262 342230
rect 470314 342178 470326 342230
rect 470378 342178 470390 342230
rect 470442 342178 470454 342230
rect 470506 342178 470518 342230
rect 470570 342178 470582 342230
rect 470634 342178 470646 342230
rect 470698 342178 470710 342230
rect 470762 342178 470774 342230
rect 470826 342178 470854 342230
rect 470234 342172 470854 342178
rect 471698 341776 471704 341828
rect 471756 341776 471762 341828
rect 471238 341708 471244 341760
rect 471296 341748 471302 341760
rect 471716 341748 471744 341776
rect 471296 341720 471744 341748
rect 471296 341708 471302 341720
rect 471716 341663 471744 341720
rect 468994 341399 469614 341405
rect 468994 341347 469022 341399
rect 469074 341347 469086 341399
rect 469138 341347 469150 341399
rect 469202 341347 469214 341399
rect 469266 341347 469278 341399
rect 469330 341347 469342 341399
rect 469394 341347 469406 341399
rect 469458 341347 469470 341399
rect 469522 341347 469534 341399
rect 469586 341347 469614 341399
rect 468994 341335 469614 341347
rect 468994 341283 469022 341335
rect 469074 341283 469086 341335
rect 469138 341283 469150 341335
rect 469202 341283 469214 341335
rect 469266 341283 469278 341335
rect 469330 341283 469342 341335
rect 469394 341283 469406 341335
rect 469458 341283 469470 341335
rect 469522 341283 469534 341335
rect 469586 341283 469614 341335
rect 468994 341271 469614 341283
rect 468994 341219 469022 341271
rect 469074 341219 469086 341271
rect 469138 341219 469150 341271
rect 469202 341219 469214 341271
rect 469266 341219 469278 341271
rect 469330 341219 469342 341271
rect 469394 341219 469406 341271
rect 469458 341219 469470 341271
rect 469522 341219 469534 341271
rect 469586 341219 469614 341271
rect 468994 341207 469614 341219
rect 468994 341155 469022 341207
rect 469074 341155 469086 341207
rect 469138 341155 469150 341207
rect 469202 341155 469214 341207
rect 469266 341155 469278 341207
rect 469330 341155 469342 341207
rect 469394 341155 469406 341207
rect 469458 341155 469470 341207
rect 469522 341155 469534 341207
rect 469586 341155 469614 341207
rect 468994 341143 469614 341155
rect 468994 341091 469022 341143
rect 469074 341091 469086 341143
rect 469138 341091 469150 341143
rect 469202 341091 469214 341143
rect 469266 341091 469278 341143
rect 469330 341091 469342 341143
rect 469394 341091 469406 341143
rect 469458 341091 469470 341143
rect 469522 341091 469534 341143
rect 469586 341091 469614 341143
rect 468994 341085 469614 341091
rect 482094 340873 482100 340876
rect 482063 340867 482100 340873
rect 474642 340803 474648 340855
rect 474700 340803 474706 340855
rect 482063 340833 482075 340867
rect 482063 340827 482100 340833
rect 482094 340824 482100 340827
rect 482152 340824 482158 340876
rect 485590 340478 485596 340490
rect 485438 340450 485596 340478
rect 485590 340438 485596 340450
rect 485648 340438 485654 340490
rect 475470 340397 475476 340400
rect 475430 340391 475476 340397
rect 475430 340357 475442 340391
rect 475430 340351 475476 340357
rect 475470 340348 475476 340351
rect 475528 340348 475534 340400
rect 478782 340397 478788 340400
rect 478747 340391 478788 340397
rect 478747 340357 478759 340391
rect 478747 340351 478788 340357
rect 478782 340348 478788 340351
rect 478840 340348 478846 340400
rect 488736 340388 488764 340464
rect 492214 340388 492220 340400
rect 488736 340360 492220 340388
rect 492214 340348 492220 340360
rect 492272 340348 492278 340400
rect 470234 340314 470854 340320
rect 470234 340262 470262 340314
rect 470314 340262 470326 340314
rect 470378 340262 470390 340314
rect 470442 340262 470454 340314
rect 470506 340262 470518 340314
rect 470570 340262 470582 340314
rect 470634 340262 470646 340314
rect 470698 340262 470710 340314
rect 470762 340262 470774 340314
rect 470826 340262 470854 340314
rect 470234 340250 470854 340262
rect 470234 340198 470262 340250
rect 470314 340198 470326 340250
rect 470378 340198 470390 340250
rect 470442 340198 470454 340250
rect 470506 340198 470518 340250
rect 470570 340198 470582 340250
rect 470634 340198 470646 340250
rect 470698 340198 470710 340250
rect 470762 340198 470774 340250
rect 470826 340198 470854 340250
rect 470234 340186 470854 340198
rect 470234 340134 470262 340186
rect 470314 340134 470326 340186
rect 470378 340134 470390 340186
rect 470442 340134 470454 340186
rect 470506 340134 470518 340186
rect 470570 340134 470582 340186
rect 470634 340134 470646 340186
rect 470698 340134 470710 340186
rect 470762 340134 470774 340186
rect 470826 340134 470854 340186
rect 470234 340122 470854 340134
rect 470234 340070 470262 340122
rect 470314 340070 470326 340122
rect 470378 340070 470390 340122
rect 470442 340070 470454 340122
rect 470506 340070 470518 340122
rect 470570 340070 470582 340122
rect 470634 340070 470646 340122
rect 470698 340070 470710 340122
rect 470762 340070 470774 340122
rect 470826 340070 470854 340122
rect 470234 340058 470854 340070
rect 470234 340006 470262 340058
rect 470314 340006 470326 340058
rect 470378 340006 470390 340058
rect 470442 340006 470454 340058
rect 470506 340006 470518 340058
rect 470570 340006 470582 340058
rect 470634 340006 470646 340058
rect 470698 340006 470710 340058
rect 470762 340006 470774 340058
rect 470826 340006 470854 340058
rect 470234 340000 470854 340006
rect 475470 339396 475476 339448
rect 475528 339396 475534 339448
rect 478782 339396 478788 339448
rect 478840 339436 478846 339448
rect 536374 339436 536380 339448
rect 478840 339408 536380 339436
rect 478840 339396 478846 339408
rect 536374 339396 536380 339408
rect 536432 339396 536438 339448
rect 475488 339300 475516 339396
rect 482094 339328 482100 339380
rect 482152 339368 482158 339380
rect 515398 339368 515404 339380
rect 482152 339340 515404 339368
rect 482152 339328 482158 339340
rect 515398 339328 515404 339340
rect 515456 339328 515462 339380
rect 497458 339300 497464 339312
rect 475488 339272 497464 339300
rect 497458 339260 497464 339272
rect 497516 339260 497522 339312
rect 523678 338036 523684 338088
rect 523736 338076 523742 338088
rect 535454 338076 535460 338088
rect 523736 338048 535460 338076
rect 523736 338036 523742 338048
rect 535454 338036 535460 338048
rect 535512 338036 535518 338088
rect 525058 332528 525064 332580
rect 525116 332568 525122 332580
rect 535454 332568 535460 332580
rect 525116 332540 535460 332568
rect 525116 332528 525122 332540
rect 535454 332528 535460 332540
rect 535512 332528 535518 332580
rect 485682 331168 485688 331220
rect 485740 331208 485746 331220
rect 535454 331208 535460 331220
rect 485740 331180 535460 331208
rect 485740 331168 485746 331180
rect 535454 331168 535460 331180
rect 535512 331168 535518 331220
rect 523678 325660 523684 325712
rect 523736 325700 523742 325712
rect 535454 325700 535460 325712
rect 523736 325672 535460 325700
rect 523736 325660 523742 325672
rect 535454 325660 535460 325672
rect 535512 325660 535518 325712
rect 470234 322486 470854 322492
rect 470234 322434 470262 322486
rect 470314 322434 470326 322486
rect 470378 322434 470390 322486
rect 470442 322434 470454 322486
rect 470506 322434 470518 322486
rect 470570 322434 470582 322486
rect 470634 322434 470646 322486
rect 470698 322434 470710 322486
rect 470762 322434 470774 322486
rect 470826 322434 470854 322486
rect 470234 322422 470854 322434
rect 470234 322370 470262 322422
rect 470314 322370 470326 322422
rect 470378 322370 470390 322422
rect 470442 322370 470454 322422
rect 470506 322370 470518 322422
rect 470570 322370 470582 322422
rect 470634 322370 470646 322422
rect 470698 322370 470710 322422
rect 470762 322370 470774 322422
rect 470826 322370 470854 322422
rect 470234 322358 470854 322370
rect 470234 322306 470262 322358
rect 470314 322306 470326 322358
rect 470378 322306 470390 322358
rect 470442 322306 470454 322358
rect 470506 322306 470518 322358
rect 470570 322306 470582 322358
rect 470634 322306 470646 322358
rect 470698 322306 470710 322358
rect 470762 322306 470774 322358
rect 470826 322306 470854 322358
rect 470234 322294 470854 322306
rect 470234 322242 470262 322294
rect 470314 322242 470326 322294
rect 470378 322242 470390 322294
rect 470442 322242 470454 322294
rect 470506 322242 470518 322294
rect 470570 322242 470582 322294
rect 470634 322242 470646 322294
rect 470698 322242 470710 322294
rect 470762 322242 470774 322294
rect 470826 322242 470854 322294
rect 470234 322230 470854 322242
rect 470234 322178 470262 322230
rect 470314 322178 470326 322230
rect 470378 322178 470390 322230
rect 470442 322178 470454 322230
rect 470506 322178 470518 322230
rect 470570 322178 470582 322230
rect 470634 322178 470646 322230
rect 470698 322178 470710 322230
rect 470762 322178 470774 322230
rect 470826 322178 470854 322230
rect 470234 322172 470854 322178
rect 471238 321580 471244 321632
rect 471296 321620 471302 321632
rect 471624 321620 471652 321663
rect 471296 321592 471652 321620
rect 471296 321580 471302 321592
rect 468994 321399 469614 321405
rect 468994 321347 469022 321399
rect 469074 321347 469086 321399
rect 469138 321347 469150 321399
rect 469202 321347 469214 321399
rect 469266 321347 469278 321399
rect 469330 321347 469342 321399
rect 469394 321347 469406 321399
rect 469458 321347 469470 321399
rect 469522 321347 469534 321399
rect 469586 321347 469614 321399
rect 468994 321335 469614 321347
rect 468994 321283 469022 321335
rect 469074 321283 469086 321335
rect 469138 321283 469150 321335
rect 469202 321283 469214 321335
rect 469266 321283 469278 321335
rect 469330 321283 469342 321335
rect 469394 321283 469406 321335
rect 469458 321283 469470 321335
rect 469522 321283 469534 321335
rect 469586 321283 469614 321335
rect 468994 321271 469614 321283
rect 468994 321219 469022 321271
rect 469074 321219 469086 321271
rect 469138 321219 469150 321271
rect 469202 321219 469214 321271
rect 469266 321219 469278 321271
rect 469330 321219 469342 321271
rect 469394 321219 469406 321271
rect 469458 321219 469470 321271
rect 469522 321219 469534 321271
rect 469586 321219 469614 321271
rect 468994 321207 469614 321219
rect 468994 321155 469022 321207
rect 469074 321155 469086 321207
rect 469138 321155 469150 321207
rect 469202 321155 469214 321207
rect 469266 321155 469278 321207
rect 469330 321155 469342 321207
rect 469394 321155 469406 321207
rect 469458 321155 469470 321207
rect 469522 321155 469534 321207
rect 469586 321155 469614 321207
rect 468994 321143 469614 321155
rect 468994 321091 469022 321143
rect 469074 321091 469086 321143
rect 469138 321091 469150 321143
rect 469202 321091 469214 321143
rect 469266 321091 469278 321143
rect 469330 321091 469342 321143
rect 469394 321091 469406 321143
rect 469458 321091 469470 321143
rect 469522 321091 469534 321143
rect 469586 321091 469614 321143
rect 468994 321085 469614 321091
rect 475470 320435 475476 320487
rect 475528 320435 475534 320487
rect 482370 320424 482376 320476
rect 482428 320424 482434 320476
rect 478927 320399 478985 320405
rect 478927 320365 478939 320399
rect 478973 320396 478985 320399
rect 479058 320396 479064 320408
rect 478973 320368 479064 320396
rect 478973 320365 478985 320368
rect 478927 320359 478985 320365
rect 479058 320356 479064 320368
rect 479116 320356 479122 320408
rect 485815 320399 485873 320405
rect 485815 320365 485827 320399
rect 485861 320396 485873 320399
rect 485958 320396 485964 320408
rect 485861 320368 485964 320396
rect 485861 320365 485873 320368
rect 485815 320359 485873 320365
rect 485958 320356 485964 320368
rect 486016 320356 486022 320408
rect 489288 320396 489316 320461
rect 492306 320396 492312 320408
rect 489288 320368 492312 320396
rect 492306 320356 492312 320368
rect 492364 320356 492370 320408
rect 470234 320314 470854 320320
rect 470234 320262 470262 320314
rect 470314 320262 470326 320314
rect 470378 320262 470390 320314
rect 470442 320262 470454 320314
rect 470506 320262 470518 320314
rect 470570 320262 470582 320314
rect 470634 320262 470646 320314
rect 470698 320262 470710 320314
rect 470762 320262 470774 320314
rect 470826 320262 470854 320314
rect 470234 320250 470854 320262
rect 470234 320198 470262 320250
rect 470314 320198 470326 320250
rect 470378 320198 470390 320250
rect 470442 320198 470454 320250
rect 470506 320198 470518 320250
rect 470570 320198 470582 320250
rect 470634 320198 470646 320250
rect 470698 320198 470710 320250
rect 470762 320198 470774 320250
rect 470826 320198 470854 320250
rect 470234 320186 470854 320198
rect 470234 320134 470262 320186
rect 470314 320134 470326 320186
rect 470378 320134 470390 320186
rect 470442 320134 470454 320186
rect 470506 320134 470518 320186
rect 470570 320134 470582 320186
rect 470634 320134 470646 320186
rect 470698 320134 470710 320186
rect 470762 320134 470774 320186
rect 470826 320134 470854 320186
rect 470234 320122 470854 320134
rect 470234 320070 470262 320122
rect 470314 320070 470326 320122
rect 470378 320070 470390 320122
rect 470442 320070 470454 320122
rect 470506 320070 470518 320122
rect 470570 320070 470582 320122
rect 470634 320070 470646 320122
rect 470698 320070 470710 320122
rect 470762 320070 470774 320122
rect 470826 320070 470854 320122
rect 470234 320058 470854 320070
rect 470234 320006 470262 320058
rect 470314 320006 470326 320058
rect 470378 320006 470390 320058
rect 470442 320006 470454 320058
rect 470506 320006 470518 320058
rect 470570 320006 470582 320058
rect 470634 320006 470646 320058
rect 470698 320006 470710 320058
rect 470762 320006 470774 320058
rect 470826 320006 470854 320058
rect 470234 320000 470854 320006
rect 475470 318724 475476 318776
rect 475528 318724 475534 318776
rect 479058 318724 479064 318776
rect 479116 318764 479122 318776
rect 536282 318764 536288 318776
rect 479116 318736 536288 318764
rect 479116 318724 479122 318736
rect 536282 318724 536288 318736
rect 536340 318724 536346 318776
rect 475488 318560 475516 318724
rect 482370 318656 482376 318708
rect 482428 318696 482434 318708
rect 536558 318696 536564 318708
rect 482428 318668 536564 318696
rect 482428 318656 482434 318668
rect 536558 318656 536564 318668
rect 536616 318656 536622 318708
rect 485958 318588 485964 318640
rect 486016 318628 486022 318640
rect 536006 318628 536012 318640
rect 486016 318600 536012 318628
rect 486016 318588 486022 318600
rect 536006 318588 536012 318600
rect 536064 318588 536070 318640
rect 498838 318560 498844 318572
rect 475488 318532 498844 318560
rect 498838 318520 498844 318532
rect 498896 318520 498902 318572
rect 470234 307086 470854 307092
rect 470234 307034 470262 307086
rect 470314 307034 470326 307086
rect 470378 307034 470390 307086
rect 470442 307034 470454 307086
rect 470506 307034 470518 307086
rect 470570 307034 470582 307086
rect 470634 307034 470646 307086
rect 470698 307034 470710 307086
rect 470762 307034 470774 307086
rect 470826 307034 470854 307086
rect 470234 307022 470854 307034
rect 470234 306970 470262 307022
rect 470314 306970 470326 307022
rect 470378 306970 470390 307022
rect 470442 306970 470454 307022
rect 470506 306970 470518 307022
rect 470570 306970 470582 307022
rect 470634 306970 470646 307022
rect 470698 306970 470710 307022
rect 470762 306970 470774 307022
rect 470826 306970 470854 307022
rect 470234 306958 470854 306970
rect 470234 306906 470262 306958
rect 470314 306906 470326 306958
rect 470378 306906 470390 306958
rect 470442 306906 470454 306958
rect 470506 306906 470518 306958
rect 470570 306906 470582 306958
rect 470634 306906 470646 306958
rect 470698 306906 470710 306958
rect 470762 306906 470774 306958
rect 470826 306906 470854 306958
rect 470234 306894 470854 306906
rect 470234 306842 470262 306894
rect 470314 306842 470326 306894
rect 470378 306842 470390 306894
rect 470442 306842 470454 306894
rect 470506 306842 470518 306894
rect 470570 306842 470582 306894
rect 470634 306842 470646 306894
rect 470698 306842 470710 306894
rect 470762 306842 470774 306894
rect 470826 306842 470854 306894
rect 470234 306830 470854 306842
rect 470234 306778 470262 306830
rect 470314 306778 470326 306830
rect 470378 306778 470390 306830
rect 470442 306778 470454 306830
rect 470506 306778 470518 306830
rect 470570 306778 470582 306830
rect 470634 306778 470646 306830
rect 470698 306778 470710 306830
rect 470762 306778 470774 306830
rect 470826 306778 470854 306830
rect 470234 306772 470854 306778
rect 471238 306280 471244 306332
rect 471296 306320 471302 306332
rect 471296 306292 471652 306320
rect 471296 306280 471302 306292
rect 471624 306264 471652 306292
rect 473722 306232 473728 306284
rect 473780 306232 473786 306284
rect 468994 306001 469614 306007
rect 468994 305949 469022 306001
rect 469074 305949 469086 306001
rect 469138 305949 469150 306001
rect 469202 305949 469214 306001
rect 469266 305949 469278 306001
rect 469330 305949 469342 306001
rect 469394 305949 469406 306001
rect 469458 305949 469470 306001
rect 469522 305949 469534 306001
rect 469586 305949 469614 306001
rect 468994 305937 469614 305949
rect 468994 305885 469022 305937
rect 469074 305885 469086 305937
rect 469138 305885 469150 305937
rect 469202 305885 469214 305937
rect 469266 305885 469278 305937
rect 469330 305885 469342 305937
rect 469394 305885 469406 305937
rect 469458 305885 469470 305937
rect 469522 305885 469534 305937
rect 469586 305885 469614 305937
rect 468994 305873 469614 305885
rect 468994 305821 469022 305873
rect 469074 305821 469086 305873
rect 469138 305821 469150 305873
rect 469202 305821 469214 305873
rect 469266 305821 469278 305873
rect 469330 305821 469342 305873
rect 469394 305821 469406 305873
rect 469458 305821 469470 305873
rect 469522 305821 469534 305873
rect 469586 305821 469614 305873
rect 468994 305809 469614 305821
rect 468994 305757 469022 305809
rect 469074 305757 469086 305809
rect 469138 305757 469150 305809
rect 469202 305757 469214 305809
rect 469266 305757 469278 305809
rect 469330 305757 469342 305809
rect 469394 305757 469406 305809
rect 469458 305757 469470 305809
rect 469522 305757 469534 305809
rect 469586 305757 469614 305809
rect 468994 305745 469614 305757
rect 468994 305693 469022 305745
rect 469074 305693 469086 305745
rect 469138 305693 469150 305745
rect 469202 305693 469214 305745
rect 469266 305693 469278 305745
rect 469330 305693 469342 305745
rect 469394 305693 469406 305745
rect 469458 305693 469470 305745
rect 469522 305693 469534 305745
rect 469586 305693 469614 305745
rect 468994 305687 469614 305693
rect 478598 305445 478604 305448
rect 478568 305439 478604 305445
rect 478568 305405 478580 305439
rect 478568 305399 478604 305405
rect 478598 305396 478604 305399
rect 478656 305396 478662 305448
rect 485130 305445 485136 305448
rect 485098 305439 485136 305445
rect 485098 305405 485110 305439
rect 485098 305399 485136 305405
rect 485130 305396 485136 305399
rect 485188 305396 485194 305448
rect 475286 305036 475292 305088
rect 475344 305036 475350 305088
rect 481818 305036 481824 305088
rect 481876 305036 481882 305088
rect 488382 305048 488672 305076
rect 488644 305028 488672 305048
rect 490558 305028 490564 305040
rect 488644 305000 490564 305028
rect 490558 304988 490564 305000
rect 490616 304988 490622 305040
rect 470234 304914 470854 304920
rect 470234 304862 470262 304914
rect 470314 304862 470326 304914
rect 470378 304862 470390 304914
rect 470442 304862 470454 304914
rect 470506 304862 470518 304914
rect 470570 304862 470582 304914
rect 470634 304862 470646 304914
rect 470698 304862 470710 304914
rect 470762 304862 470774 304914
rect 470826 304862 470854 304914
rect 470234 304850 470854 304862
rect 470234 304798 470262 304850
rect 470314 304798 470326 304850
rect 470378 304798 470390 304850
rect 470442 304798 470454 304850
rect 470506 304798 470518 304850
rect 470570 304798 470582 304850
rect 470634 304798 470646 304850
rect 470698 304798 470710 304850
rect 470762 304798 470774 304850
rect 470826 304798 470854 304850
rect 470234 304786 470854 304798
rect 470234 304734 470262 304786
rect 470314 304734 470326 304786
rect 470378 304734 470390 304786
rect 470442 304734 470454 304786
rect 470506 304734 470518 304786
rect 470570 304734 470582 304786
rect 470634 304734 470646 304786
rect 470698 304734 470710 304786
rect 470762 304734 470774 304786
rect 470826 304734 470854 304786
rect 470234 304722 470854 304734
rect 470234 304670 470262 304722
rect 470314 304670 470326 304722
rect 470378 304670 470390 304722
rect 470442 304670 470454 304722
rect 470506 304670 470518 304722
rect 470570 304670 470582 304722
rect 470634 304670 470646 304722
rect 470698 304670 470710 304722
rect 470762 304670 470774 304722
rect 470826 304670 470854 304722
rect 470234 304658 470854 304670
rect 470234 304606 470262 304658
rect 470314 304606 470326 304658
rect 470378 304606 470390 304658
rect 470442 304606 470454 304658
rect 470506 304606 470518 304658
rect 470570 304606 470582 304658
rect 470634 304606 470646 304658
rect 470698 304606 470710 304658
rect 470762 304606 470774 304658
rect 470826 304606 470854 304658
rect 470234 304600 470854 304606
rect 485056 303640 485268 303668
rect 475286 303560 475292 303612
rect 475344 303560 475350 303612
rect 478598 303560 478604 303612
rect 478656 303600 478662 303612
rect 478656 303572 480254 303600
rect 478656 303560 478662 303572
rect 475304 303396 475332 303560
rect 480226 303464 480254 303572
rect 481818 303560 481824 303612
rect 481876 303600 481882 303612
rect 485056 303600 485084 303640
rect 481876 303572 485084 303600
rect 481876 303560 481882 303572
rect 485130 303560 485136 303612
rect 485188 303560 485194 303612
rect 485240 303600 485268 303640
rect 536466 303600 536472 303612
rect 485240 303572 536472 303600
rect 536466 303560 536472 303572
rect 536524 303560 536530 303612
rect 485148 303532 485176 303560
rect 536650 303532 536656 303544
rect 485148 303504 536656 303532
rect 536650 303492 536656 303504
rect 536708 303492 536714 303544
rect 518158 303464 518164 303476
rect 480226 303436 518164 303464
rect 518158 303424 518164 303436
rect 518216 303424 518222 303476
rect 500218 303396 500224 303408
rect 475304 303368 500224 303396
rect 500218 303356 500224 303368
rect 500276 303356 500282 303408
rect 491938 300772 491944 300824
rect 491996 300812 492002 300824
rect 535454 300812 535460 300824
rect 491996 300784 535460 300812
rect 491996 300772 492002 300784
rect 535454 300772 535460 300784
rect 535512 300772 535518 300824
rect 492030 299412 492036 299464
rect 492088 299452 492094 299464
rect 535454 299452 535460 299464
rect 492088 299424 535460 299452
rect 492088 299412 492094 299424
rect 535454 299412 535460 299424
rect 535512 299412 535518 299464
rect 490742 298052 490748 298104
rect 490800 298092 490806 298104
rect 535454 298092 535460 298104
rect 490800 298064 535460 298092
rect 490800 298052 490806 298064
rect 535454 298052 535460 298064
rect 535512 298052 535518 298104
rect 492122 296624 492128 296676
rect 492180 296664 492186 296676
rect 535546 296664 535552 296676
rect 492180 296636 535552 296664
rect 492180 296624 492186 296636
rect 535546 296624 535552 296636
rect 535604 296624 535610 296676
rect 493318 296556 493324 296608
rect 493376 296596 493382 296608
rect 535454 296596 535460 296608
rect 493376 296568 535460 296596
rect 493376 296556 493382 296568
rect 535454 296556 535460 296568
rect 535512 296556 535518 296608
rect 492214 295264 492220 295316
rect 492272 295304 492278 295316
rect 535454 295304 535460 295316
rect 492272 295276 535460 295304
rect 492272 295264 492278 295276
rect 535454 295264 535460 295276
rect 535512 295264 535518 295316
rect 492306 293904 492312 293956
rect 492364 293944 492370 293956
rect 535546 293944 535552 293956
rect 492364 293916 535552 293944
rect 492364 293904 492370 293916
rect 535546 293904 535552 293916
rect 535604 293904 535610 293956
rect 490558 292476 490564 292528
rect 490616 292516 490622 292528
rect 535454 292516 535460 292528
rect 490616 292488 535460 292516
rect 490616 292476 490622 292488
rect 535454 292476 535460 292488
rect 535512 292476 535518 292528
rect 492950 289824 492956 289876
rect 493008 289864 493014 289876
rect 535454 289864 535460 289876
rect 493008 289836 535460 289864
rect 493008 289824 493014 289836
rect 535454 289824 535460 289836
rect 535512 289824 535518 289876
rect 491938 288396 491944 288448
rect 491996 288436 492002 288448
rect 535454 288436 535460 288448
rect 491996 288408 535460 288436
rect 491996 288396 492002 288408
rect 535454 288396 535460 288408
rect 535512 288396 535518 288448
rect 470234 287487 470854 287493
rect 470234 287435 470262 287487
rect 470314 287435 470326 287487
rect 470378 287435 470390 287487
rect 470442 287435 470454 287487
rect 470506 287435 470518 287487
rect 470570 287435 470582 287487
rect 470634 287435 470646 287487
rect 470698 287435 470710 287487
rect 470762 287435 470774 287487
rect 470826 287435 470854 287487
rect 470234 287423 470854 287435
rect 470234 287371 470262 287423
rect 470314 287371 470326 287423
rect 470378 287371 470390 287423
rect 470442 287371 470454 287423
rect 470506 287371 470518 287423
rect 470570 287371 470582 287423
rect 470634 287371 470646 287423
rect 470698 287371 470710 287423
rect 470762 287371 470774 287423
rect 470826 287371 470854 287423
rect 470234 287359 470854 287371
rect 470234 287307 470262 287359
rect 470314 287307 470326 287359
rect 470378 287307 470390 287359
rect 470442 287307 470454 287359
rect 470506 287307 470518 287359
rect 470570 287307 470582 287359
rect 470634 287307 470646 287359
rect 470698 287307 470710 287359
rect 470762 287307 470774 287359
rect 470826 287307 470854 287359
rect 470234 287295 470854 287307
rect 470234 287243 470262 287295
rect 470314 287243 470326 287295
rect 470378 287243 470390 287295
rect 470442 287243 470454 287295
rect 470506 287243 470518 287295
rect 470570 287243 470582 287295
rect 470634 287243 470646 287295
rect 470698 287243 470710 287295
rect 470762 287243 470774 287295
rect 470826 287243 470854 287295
rect 470234 287231 470854 287243
rect 470234 287179 470262 287231
rect 470314 287179 470326 287231
rect 470378 287179 470390 287231
rect 470442 287179 470454 287231
rect 470506 287179 470518 287231
rect 470570 287179 470582 287231
rect 470634 287179 470646 287231
rect 470698 287179 470710 287231
rect 470762 287179 470774 287231
rect 470826 287179 470854 287231
rect 470234 287173 470854 287179
rect 488632 286680 488684 286686
rect 471238 286628 471244 286680
rect 471296 286668 471302 286680
rect 471296 286640 471652 286668
rect 471296 286628 471302 286640
rect 471624 286532 471652 286640
rect 488632 286622 488684 286628
rect 471698 286532 471704 286544
rect 471624 286504 471704 286532
rect 471698 286492 471704 286504
rect 471756 286492 471762 286544
rect 468994 286402 469614 286408
rect 468994 286350 469022 286402
rect 469074 286350 469086 286402
rect 469138 286350 469150 286402
rect 469202 286350 469214 286402
rect 469266 286350 469278 286402
rect 469330 286350 469342 286402
rect 469394 286350 469406 286402
rect 469458 286350 469470 286402
rect 469522 286350 469534 286402
rect 469586 286350 469614 286402
rect 468994 286338 469614 286350
rect 468994 286286 469022 286338
rect 469074 286286 469086 286338
rect 469138 286286 469150 286338
rect 469202 286286 469214 286338
rect 469266 286286 469278 286338
rect 469330 286286 469342 286338
rect 469394 286286 469406 286338
rect 469458 286286 469470 286338
rect 469522 286286 469534 286338
rect 469586 286286 469614 286338
rect 468994 286274 469614 286286
rect 468994 286222 469022 286274
rect 469074 286222 469086 286274
rect 469138 286222 469150 286274
rect 469202 286222 469214 286274
rect 469266 286222 469278 286274
rect 469330 286222 469342 286274
rect 469394 286222 469406 286274
rect 469458 286222 469470 286274
rect 469522 286222 469534 286274
rect 469586 286222 469614 286274
rect 468994 286210 469614 286222
rect 468994 286158 469022 286210
rect 469074 286158 469086 286210
rect 469138 286158 469150 286210
rect 469202 286158 469214 286210
rect 469266 286158 469278 286210
rect 469330 286158 469342 286210
rect 469394 286158 469406 286210
rect 469458 286158 469470 286210
rect 469522 286158 469534 286210
rect 469586 286158 469614 286210
rect 468994 286146 469614 286158
rect 468994 286094 469022 286146
rect 469074 286094 469086 286146
rect 469138 286094 469150 286146
rect 469202 286094 469214 286146
rect 469266 286094 469278 286146
rect 469330 286094 469342 286146
rect 469394 286094 469406 286146
rect 469458 286094 469470 286146
rect 469522 286094 469534 286146
rect 469586 286094 469614 286146
rect 468994 286088 469614 286094
rect 490598 285991 490656 285997
rect 490598 285957 490610 285991
rect 490644 285988 490656 285991
rect 490644 285960 490880 285988
rect 490644 285957 490656 285960
rect 490598 285951 490656 285957
rect 479426 285812 479432 285864
rect 479484 285861 479490 285864
rect 479484 285855 479520 285861
rect 479508 285821 479520 285855
rect 479484 285815 479520 285821
rect 479484 285812 479490 285815
rect 490852 285648 490880 285960
rect 492950 285648 492956 285660
rect 490852 285620 492956 285648
rect 492950 285608 492956 285620
rect 493008 285608 493014 285660
rect 475746 285436 475752 285488
rect 475804 285436 475810 285488
rect 483198 285436 483204 285488
rect 483256 285436 483262 285488
rect 486878 285436 486884 285488
rect 486936 285436 486942 285488
rect 470234 285314 470854 285320
rect 470234 285262 470262 285314
rect 470314 285262 470326 285314
rect 470378 285262 470390 285314
rect 470442 285262 470454 285314
rect 470506 285262 470518 285314
rect 470570 285262 470582 285314
rect 470634 285262 470646 285314
rect 470698 285262 470710 285314
rect 470762 285262 470774 285314
rect 470826 285262 470854 285314
rect 470234 285250 470854 285262
rect 470234 285198 470262 285250
rect 470314 285198 470326 285250
rect 470378 285198 470390 285250
rect 470442 285198 470454 285250
rect 470506 285198 470518 285250
rect 470570 285198 470582 285250
rect 470634 285198 470646 285250
rect 470698 285198 470710 285250
rect 470762 285198 470774 285250
rect 470826 285198 470854 285250
rect 470234 285186 470854 285198
rect 470234 285134 470262 285186
rect 470314 285134 470326 285186
rect 470378 285134 470390 285186
rect 470442 285134 470454 285186
rect 470506 285134 470518 285186
rect 470570 285134 470582 285186
rect 470634 285134 470646 285186
rect 470698 285134 470710 285186
rect 470762 285134 470774 285186
rect 470826 285134 470854 285186
rect 470234 285122 470854 285134
rect 470234 285070 470262 285122
rect 470314 285070 470326 285122
rect 470378 285070 470390 285122
rect 470442 285070 470454 285122
rect 470506 285070 470518 285122
rect 470570 285070 470582 285122
rect 470634 285070 470646 285122
rect 470698 285070 470710 285122
rect 470762 285070 470774 285122
rect 470826 285070 470854 285122
rect 470234 285058 470854 285070
rect 470234 285006 470262 285058
rect 470314 285006 470326 285058
rect 470378 285006 470390 285058
rect 470442 285006 470454 285058
rect 470506 285006 470518 285058
rect 470570 285006 470582 285058
rect 470634 285006 470646 285058
rect 470698 285006 470710 285058
rect 470762 285006 470774 285058
rect 470826 285006 470854 285058
rect 470234 285000 470854 285006
rect 475746 284248 475752 284300
rect 475804 284248 475810 284300
rect 479426 284248 479432 284300
rect 479484 284288 479490 284300
rect 536098 284288 536104 284300
rect 479484 284260 536104 284288
rect 479484 284248 479490 284260
rect 536098 284248 536104 284260
rect 536156 284248 536162 284300
rect 475764 284084 475792 284248
rect 483198 284180 483204 284232
rect 483256 284180 483262 284232
rect 522298 284220 522304 284232
rect 485746 284192 522304 284220
rect 483216 284152 483244 284180
rect 485746 284152 485774 284192
rect 522298 284180 522304 284192
rect 522356 284180 522362 284232
rect 483216 284124 485774 284152
rect 486878 284112 486884 284164
rect 486936 284152 486942 284164
rect 523678 284152 523684 284164
rect 486936 284124 523684 284152
rect 486936 284112 486942 284124
rect 523678 284112 523684 284124
rect 523736 284112 523742 284164
rect 501598 284084 501604 284096
rect 475764 284056 501604 284084
rect 501598 284044 501604 284056
rect 501656 284044 501662 284096
rect 471698 270444 471704 270496
rect 471756 270484 471762 270496
rect 473722 270484 473728 270496
rect 471756 270456 473728 270484
rect 471756 270444 471762 270456
rect 473722 270444 473728 270456
rect 473780 270444 473786 270496
rect 470234 267487 470854 267493
rect 470234 267435 470262 267487
rect 470314 267435 470326 267487
rect 470378 267435 470390 267487
rect 470442 267435 470454 267487
rect 470506 267435 470518 267487
rect 470570 267435 470582 267487
rect 470634 267435 470646 267487
rect 470698 267435 470710 267487
rect 470762 267435 470774 267487
rect 470826 267435 470854 267487
rect 470234 267423 470854 267435
rect 470234 267371 470262 267423
rect 470314 267371 470326 267423
rect 470378 267371 470390 267423
rect 470442 267371 470454 267423
rect 470506 267371 470518 267423
rect 470570 267371 470582 267423
rect 470634 267371 470646 267423
rect 470698 267371 470710 267423
rect 470762 267371 470774 267423
rect 470826 267371 470854 267423
rect 470234 267359 470854 267371
rect 470234 267307 470262 267359
rect 470314 267307 470326 267359
rect 470378 267307 470390 267359
rect 470442 267307 470454 267359
rect 470506 267307 470518 267359
rect 470570 267307 470582 267359
rect 470634 267307 470646 267359
rect 470698 267307 470710 267359
rect 470762 267307 470774 267359
rect 470826 267307 470854 267359
rect 470234 267295 470854 267307
rect 470234 267243 470262 267295
rect 470314 267243 470326 267295
rect 470378 267243 470390 267295
rect 470442 267243 470454 267295
rect 470506 267243 470518 267295
rect 470570 267243 470582 267295
rect 470634 267243 470646 267295
rect 470698 267243 470710 267295
rect 470762 267243 470774 267295
rect 470826 267243 470854 267295
rect 470234 267231 470854 267243
rect 470234 267179 470262 267231
rect 470314 267179 470326 267231
rect 470378 267179 470390 267231
rect 470442 267179 470454 267231
rect 470506 267179 470518 267231
rect 470570 267179 470582 267231
rect 470634 267179 470646 267231
rect 470698 267179 470710 267231
rect 470762 267179 470774 267231
rect 470826 267179 470854 267231
rect 470234 267173 470854 267179
rect 473648 266540 473676 266664
rect 473722 266540 473728 266552
rect 473648 266512 473728 266540
rect 473722 266500 473728 266512
rect 473780 266500 473786 266552
rect 468994 266401 469614 266407
rect 468994 266349 469022 266401
rect 469074 266349 469086 266401
rect 469138 266349 469150 266401
rect 469202 266349 469214 266401
rect 469266 266349 469278 266401
rect 469330 266349 469342 266401
rect 469394 266349 469406 266401
rect 469458 266349 469470 266401
rect 469522 266349 469534 266401
rect 469586 266349 469614 266401
rect 468994 266337 469614 266349
rect 468994 266285 469022 266337
rect 469074 266285 469086 266337
rect 469138 266285 469150 266337
rect 469202 266285 469214 266337
rect 469266 266285 469278 266337
rect 469330 266285 469342 266337
rect 469394 266285 469406 266337
rect 469458 266285 469470 266337
rect 469522 266285 469534 266337
rect 469586 266285 469614 266337
rect 468994 266273 469614 266285
rect 468994 266221 469022 266273
rect 469074 266221 469086 266273
rect 469138 266221 469150 266273
rect 469202 266221 469214 266273
rect 469266 266221 469278 266273
rect 469330 266221 469342 266273
rect 469394 266221 469406 266273
rect 469458 266221 469470 266273
rect 469522 266221 469534 266273
rect 469586 266221 469614 266273
rect 468994 266209 469614 266221
rect 468994 266157 469022 266209
rect 469074 266157 469086 266209
rect 469138 266157 469150 266209
rect 469202 266157 469214 266209
rect 469266 266157 469278 266209
rect 469330 266157 469342 266209
rect 469394 266157 469406 266209
rect 469458 266157 469470 266209
rect 469522 266157 469534 266209
rect 469586 266157 469614 266209
rect 468994 266145 469614 266157
rect 468994 266093 469022 266145
rect 469074 266093 469086 266145
rect 469138 266093 469150 266145
rect 469202 266093 469214 266145
rect 469266 266093 469278 266145
rect 469330 266093 469342 266145
rect 469394 266093 469406 266145
rect 469458 266093 469470 266145
rect 469522 266093 469534 266145
rect 469586 266093 469614 266145
rect 468994 266087 469614 266093
rect 491938 265996 491944 266008
rect 489288 265968 491944 265996
rect 477126 265869 477132 265872
rect 477089 265863 477132 265869
rect 477089 265829 477101 265863
rect 477089 265823 477132 265829
rect 477126 265820 477132 265823
rect 477184 265820 477190 265872
rect 489288 265731 489316 265968
rect 491938 265956 491944 265968
rect 491996 265956 492002 266008
rect 480162 265435 480168 265487
rect 480220 265435 480226 265487
rect 483198 265435 483204 265487
rect 483256 265435 483262 265487
rect 486234 265435 486240 265487
rect 486292 265435 486298 265487
rect 470234 265314 470854 265320
rect 470234 265262 470262 265314
rect 470314 265262 470326 265314
rect 470378 265262 470390 265314
rect 470442 265262 470454 265314
rect 470506 265262 470518 265314
rect 470570 265262 470582 265314
rect 470634 265262 470646 265314
rect 470698 265262 470710 265314
rect 470762 265262 470774 265314
rect 470826 265262 470854 265314
rect 470234 265250 470854 265262
rect 470234 265198 470262 265250
rect 470314 265198 470326 265250
rect 470378 265198 470390 265250
rect 470442 265198 470454 265250
rect 470506 265198 470518 265250
rect 470570 265198 470582 265250
rect 470634 265198 470646 265250
rect 470698 265198 470710 265250
rect 470762 265198 470774 265250
rect 470826 265198 470854 265250
rect 470234 265186 470854 265198
rect 470234 265134 470262 265186
rect 470314 265134 470326 265186
rect 470378 265134 470390 265186
rect 470442 265134 470454 265186
rect 470506 265134 470518 265186
rect 470570 265134 470582 265186
rect 470634 265134 470646 265186
rect 470698 265134 470710 265186
rect 470762 265134 470774 265186
rect 470826 265134 470854 265186
rect 470234 265122 470854 265134
rect 470234 265070 470262 265122
rect 470314 265070 470326 265122
rect 470378 265070 470390 265122
rect 470442 265070 470454 265122
rect 470506 265070 470518 265122
rect 470570 265070 470582 265122
rect 470634 265070 470646 265122
rect 470698 265070 470710 265122
rect 470762 265070 470774 265122
rect 470826 265070 470854 265122
rect 470234 265058 470854 265070
rect 470234 265006 470262 265058
rect 470314 265006 470326 265058
rect 470378 265006 470390 265058
rect 470442 265006 470454 265058
rect 470506 265006 470518 265058
rect 470570 265006 470582 265058
rect 470634 265006 470646 265058
rect 470698 265006 470710 265058
rect 470762 265006 470774 265058
rect 470826 265006 470854 265058
rect 470234 265000 470854 265006
rect 494716 263588 494928 263616
rect 477126 263508 477132 263560
rect 477184 263508 477190 263560
rect 480162 263508 480168 263560
rect 480220 263548 480226 263560
rect 480220 263508 480254 263548
rect 483198 263508 483204 263560
rect 483256 263508 483262 263560
rect 486234 263508 486240 263560
rect 486292 263548 486298 263560
rect 494716 263548 494744 263588
rect 486292 263520 494744 263548
rect 494900 263548 494928 263588
rect 494900 263520 495020 263548
rect 486292 263508 486298 263520
rect 477144 263344 477172 263508
rect 480226 263412 480254 263508
rect 483216 263480 483244 263508
rect 494790 263480 494796 263492
rect 483216 263452 494796 263480
rect 494790 263440 494796 263452
rect 494848 263440 494854 263492
rect 494992 263480 495020 263520
rect 495066 263508 495072 263560
rect 495124 263548 495130 263560
rect 535914 263548 535920 263560
rect 495124 263520 535920 263548
rect 495124 263508 495130 263520
rect 535914 263508 535920 263520
rect 535972 263508 535978 263560
rect 536374 263480 536380 263492
rect 494992 263452 536380 263480
rect 536374 263440 536380 263452
rect 536432 263440 536438 263492
rect 519538 263412 519544 263424
rect 480226 263384 519544 263412
rect 519538 263372 519544 263384
rect 519596 263372 519602 263424
rect 502978 263344 502984 263356
rect 477144 263316 502984 263344
rect 502978 263304 502984 263316
rect 503036 263304 503042 263356
rect 473722 206932 473728 206984
rect 473780 206972 473786 206984
rect 580166 206972 580172 206984
rect 473780 206944 580172 206972
rect 473780 206932 473786 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
<< via1 >>
rect 470262 451433 470314 451485
rect 470326 451433 470378 451485
rect 470390 451433 470442 451485
rect 470454 451433 470506 451485
rect 470518 451433 470570 451485
rect 470582 451433 470634 451485
rect 470646 451433 470698 451485
rect 470710 451433 470762 451485
rect 470774 451433 470826 451485
rect 470262 451369 470314 451421
rect 470326 451369 470378 451421
rect 470390 451369 470442 451421
rect 470454 451369 470506 451421
rect 470518 451369 470570 451421
rect 470582 451369 470634 451421
rect 470646 451369 470698 451421
rect 470710 451369 470762 451421
rect 470774 451369 470826 451421
rect 470262 451305 470314 451357
rect 470326 451305 470378 451357
rect 470390 451305 470442 451357
rect 470454 451305 470506 451357
rect 470518 451305 470570 451357
rect 470582 451305 470634 451357
rect 470646 451305 470698 451357
rect 470710 451305 470762 451357
rect 470774 451305 470826 451357
rect 470262 451241 470314 451293
rect 470326 451241 470378 451293
rect 470390 451241 470442 451293
rect 470454 451241 470506 451293
rect 470518 451241 470570 451293
rect 470582 451241 470634 451293
rect 470646 451241 470698 451293
rect 470710 451241 470762 451293
rect 470774 451241 470826 451293
rect 470262 451177 470314 451229
rect 470326 451177 470378 451229
rect 470390 451177 470442 451229
rect 470454 451177 470506 451229
rect 470518 451177 470570 451229
rect 470582 451177 470634 451229
rect 470646 451177 470698 451229
rect 470710 451177 470762 451229
rect 470774 451177 470826 451229
rect 471336 450644 471388 450696
rect 469022 450347 469074 450399
rect 469086 450347 469138 450399
rect 469150 450347 469202 450399
rect 469214 450347 469266 450399
rect 469278 450347 469330 450399
rect 469342 450347 469394 450399
rect 469406 450347 469458 450399
rect 469470 450347 469522 450399
rect 469534 450347 469586 450399
rect 469022 450283 469074 450335
rect 469086 450283 469138 450335
rect 469150 450283 469202 450335
rect 469214 450283 469266 450335
rect 469278 450283 469330 450335
rect 469342 450283 469394 450335
rect 469406 450283 469458 450335
rect 469470 450283 469522 450335
rect 469534 450283 469586 450335
rect 469022 450219 469074 450271
rect 469086 450219 469138 450271
rect 469150 450219 469202 450271
rect 469214 450219 469266 450271
rect 469278 450219 469330 450271
rect 469342 450219 469394 450271
rect 469406 450219 469458 450271
rect 469470 450219 469522 450271
rect 469534 450219 469586 450271
rect 469022 450155 469074 450207
rect 469086 450155 469138 450207
rect 469150 450155 469202 450207
rect 469214 450155 469266 450207
rect 469278 450155 469330 450207
rect 469342 450155 469394 450207
rect 469406 450155 469458 450207
rect 469470 450155 469522 450207
rect 469534 450155 469586 450207
rect 469022 450091 469074 450143
rect 469086 450091 469138 450143
rect 469150 450091 469202 450143
rect 469214 450091 469266 450143
rect 469278 450091 469330 450143
rect 469342 450091 469394 450143
rect 469406 450091 469458 450143
rect 469470 450091 469522 450143
rect 469534 450091 469586 450143
rect 475384 449436 475436 449488
rect 478696 449436 478748 449488
rect 482008 449436 482060 449488
rect 485320 449436 485372 449488
rect 491944 449352 491996 449404
rect 470262 449262 470314 449314
rect 470326 449262 470378 449314
rect 470390 449262 470442 449314
rect 470454 449262 470506 449314
rect 470518 449262 470570 449314
rect 470582 449262 470634 449314
rect 470646 449262 470698 449314
rect 470710 449262 470762 449314
rect 470774 449262 470826 449314
rect 470262 449198 470314 449250
rect 470326 449198 470378 449250
rect 470390 449198 470442 449250
rect 470454 449198 470506 449250
rect 470518 449198 470570 449250
rect 470582 449198 470634 449250
rect 470646 449198 470698 449250
rect 470710 449198 470762 449250
rect 470774 449198 470826 449250
rect 470262 449134 470314 449186
rect 470326 449134 470378 449186
rect 470390 449134 470442 449186
rect 470454 449134 470506 449186
rect 470518 449134 470570 449186
rect 470582 449134 470634 449186
rect 470646 449134 470698 449186
rect 470710 449134 470762 449186
rect 470774 449134 470826 449186
rect 470262 449070 470314 449122
rect 470326 449070 470378 449122
rect 470390 449070 470442 449122
rect 470454 449070 470506 449122
rect 470518 449070 470570 449122
rect 470582 449070 470634 449122
rect 470646 449070 470698 449122
rect 470710 449070 470762 449122
rect 470774 449070 470826 449122
rect 470262 449006 470314 449058
rect 470326 449006 470378 449058
rect 470390 449006 470442 449058
rect 470454 449006 470506 449058
rect 470518 449006 470570 449058
rect 470582 449006 470634 449058
rect 470646 449006 470698 449058
rect 470710 449006 470762 449058
rect 470774 449006 470826 449058
rect 478696 446224 478748 446276
rect 515404 445884 515456 445936
rect 482008 445816 482060 445868
rect 485320 445816 485372 445868
rect 523684 445816 523736 445868
rect 520924 445748 520976 445800
rect 475384 445680 475436 445732
rect 535460 445680 535512 445732
rect 490564 442960 490616 443012
rect 535460 442960 535512 443012
rect 493324 441600 493376 441652
rect 535460 441600 535512 441652
rect 494704 440240 494756 440292
rect 535460 440240 535512 440292
rect 496084 438880 496136 438932
rect 535460 438880 535512 438932
rect 497464 437452 497516 437504
rect 535460 437452 535512 437504
rect 498844 436092 498896 436144
rect 535460 436092 535512 436144
rect 500224 434732 500276 434784
rect 535460 434732 535512 434784
rect 501604 433304 501656 433356
rect 535460 433304 535512 433356
rect 470262 433034 470314 433086
rect 470326 433034 470378 433086
rect 470390 433034 470442 433086
rect 470454 433034 470506 433086
rect 470518 433034 470570 433086
rect 470582 433034 470634 433086
rect 470646 433034 470698 433086
rect 470710 433034 470762 433086
rect 470774 433034 470826 433086
rect 470262 432970 470314 433022
rect 470326 432970 470378 433022
rect 470390 432970 470442 433022
rect 470454 432970 470506 433022
rect 470518 432970 470570 433022
rect 470582 432970 470634 433022
rect 470646 432970 470698 433022
rect 470710 432970 470762 433022
rect 470774 432970 470826 433022
rect 470262 432906 470314 432958
rect 470326 432906 470378 432958
rect 470390 432906 470442 432958
rect 470454 432906 470506 432958
rect 470518 432906 470570 432958
rect 470582 432906 470634 432958
rect 470646 432906 470698 432958
rect 470710 432906 470762 432958
rect 470774 432906 470826 432958
rect 470262 432842 470314 432894
rect 470326 432842 470378 432894
rect 470390 432842 470442 432894
rect 470454 432842 470506 432894
rect 470518 432842 470570 432894
rect 470582 432842 470634 432894
rect 470646 432842 470698 432894
rect 470710 432842 470762 432894
rect 470774 432842 470826 432894
rect 470262 432778 470314 432830
rect 470326 432778 470378 432830
rect 470390 432778 470442 432830
rect 470454 432778 470506 432830
rect 470518 432778 470570 432830
rect 470582 432778 470634 432830
rect 470646 432778 470698 432830
rect 470710 432778 470762 432830
rect 470774 432778 470826 432830
rect 471612 432238 471664 432290
rect 469022 431947 469074 431999
rect 469086 431947 469138 431999
rect 469150 431947 469202 431999
rect 469214 431947 469266 431999
rect 469278 431947 469330 431999
rect 469342 431947 469394 431999
rect 469406 431947 469458 431999
rect 469470 431947 469522 431999
rect 469534 431947 469586 431999
rect 502984 431944 503036 431996
rect 535460 431944 535512 431996
rect 469022 431883 469074 431935
rect 469086 431883 469138 431935
rect 469150 431883 469202 431935
rect 469214 431883 469266 431935
rect 469278 431883 469330 431935
rect 469342 431883 469394 431935
rect 469406 431883 469458 431935
rect 469470 431883 469522 431935
rect 469534 431883 469586 431935
rect 469022 431819 469074 431871
rect 469086 431819 469138 431871
rect 469150 431819 469202 431871
rect 469214 431819 469266 431871
rect 469278 431819 469330 431871
rect 469342 431819 469394 431871
rect 469406 431819 469458 431871
rect 469470 431819 469522 431871
rect 469534 431819 469586 431871
rect 469022 431755 469074 431807
rect 469086 431755 469138 431807
rect 469150 431755 469202 431807
rect 469214 431755 469266 431807
rect 469278 431755 469330 431807
rect 469342 431755 469394 431807
rect 469406 431755 469458 431807
rect 469470 431755 469522 431807
rect 469534 431755 469586 431807
rect 469022 431691 469074 431743
rect 469086 431691 469138 431743
rect 469150 431691 469202 431743
rect 469214 431691 469266 431743
rect 469278 431691 469330 431743
rect 469342 431691 469394 431743
rect 469406 431691 469458 431743
rect 469470 431691 469522 431743
rect 469534 431691 469586 431743
rect 478972 431443 479024 431452
rect 478972 431409 478977 431443
rect 478977 431409 479024 431443
rect 478972 431400 479024 431409
rect 485780 431443 485832 431452
rect 485780 431409 485831 431443
rect 485831 431409 485832 431443
rect 485780 431400 485832 431409
rect 475476 431035 475528 431087
rect 482376 431035 482428 431087
rect 492036 430992 492088 431044
rect 470262 430862 470314 430914
rect 470326 430862 470378 430914
rect 470390 430862 470442 430914
rect 470454 430862 470506 430914
rect 470518 430862 470570 430914
rect 470582 430862 470634 430914
rect 470646 430862 470698 430914
rect 470710 430862 470762 430914
rect 470774 430862 470826 430914
rect 470262 430798 470314 430850
rect 470326 430798 470378 430850
rect 470390 430798 470442 430850
rect 470454 430798 470506 430850
rect 470518 430798 470570 430850
rect 470582 430798 470634 430850
rect 470646 430798 470698 430850
rect 470710 430798 470762 430850
rect 470774 430798 470826 430850
rect 470262 430734 470314 430786
rect 470326 430734 470378 430786
rect 470390 430734 470442 430786
rect 470454 430734 470506 430786
rect 470518 430734 470570 430786
rect 470582 430734 470634 430786
rect 470646 430734 470698 430786
rect 470710 430734 470762 430786
rect 470774 430734 470826 430786
rect 470262 430670 470314 430722
rect 470326 430670 470378 430722
rect 470390 430670 470442 430722
rect 470454 430670 470506 430722
rect 470518 430670 470570 430722
rect 470582 430670 470634 430722
rect 470646 430670 470698 430722
rect 470710 430670 470762 430722
rect 470774 430670 470826 430722
rect 470262 430606 470314 430658
rect 470326 430606 470378 430658
rect 470390 430606 470442 430658
rect 470454 430606 470506 430658
rect 470518 430606 470570 430658
rect 470582 430606 470634 430658
rect 470646 430606 470698 430658
rect 470710 430606 470762 430658
rect 470774 430606 470826 430658
rect 475476 429088 475528 429140
rect 490564 429088 490616 429140
rect 482376 427796 482428 427848
rect 522304 427796 522356 427848
rect 470262 412034 470314 412086
rect 470326 412034 470378 412086
rect 470390 412034 470442 412086
rect 470454 412034 470506 412086
rect 470518 412034 470570 412086
rect 470582 412034 470634 412086
rect 470646 412034 470698 412086
rect 470710 412034 470762 412086
rect 470774 412034 470826 412086
rect 470262 411970 470314 412022
rect 470326 411970 470378 412022
rect 470390 411970 470442 412022
rect 470454 411970 470506 412022
rect 470518 411970 470570 412022
rect 470582 411970 470634 412022
rect 470646 411970 470698 412022
rect 470710 411970 470762 412022
rect 470774 411970 470826 412022
rect 470262 411906 470314 411958
rect 470326 411906 470378 411958
rect 470390 411906 470442 411958
rect 470454 411906 470506 411958
rect 470518 411906 470570 411958
rect 470582 411906 470634 411958
rect 470646 411906 470698 411958
rect 470710 411906 470762 411958
rect 470774 411906 470826 411958
rect 470262 411842 470314 411894
rect 470326 411842 470378 411894
rect 470390 411842 470442 411894
rect 470454 411842 470506 411894
rect 470518 411842 470570 411894
rect 470582 411842 470634 411894
rect 470646 411842 470698 411894
rect 470710 411842 470762 411894
rect 470774 411842 470826 411894
rect 470262 411778 470314 411830
rect 470326 411778 470378 411830
rect 470390 411778 470442 411830
rect 470454 411778 470506 411830
rect 470518 411778 470570 411830
rect 470582 411778 470634 411830
rect 470646 411778 470698 411830
rect 470710 411778 470762 411830
rect 470774 411778 470826 411830
rect 471244 411204 471296 411256
rect 473728 411232 473780 411284
rect 469022 410948 469074 411000
rect 469086 410948 469138 411000
rect 469150 410948 469202 411000
rect 469214 410948 469266 411000
rect 469278 410948 469330 411000
rect 469342 410948 469394 411000
rect 469406 410948 469458 411000
rect 469470 410948 469522 411000
rect 469534 410948 469586 411000
rect 469022 410884 469074 410936
rect 469086 410884 469138 410936
rect 469150 410884 469202 410936
rect 469214 410884 469266 410936
rect 469278 410884 469330 410936
rect 469342 410884 469394 410936
rect 469406 410884 469458 410936
rect 469470 410884 469522 410936
rect 469534 410884 469586 410936
rect 469022 410820 469074 410872
rect 469086 410820 469138 410872
rect 469150 410820 469202 410872
rect 469214 410820 469266 410872
rect 469278 410820 469330 410872
rect 469342 410820 469394 410872
rect 469406 410820 469458 410872
rect 469470 410820 469522 410872
rect 469534 410820 469586 410872
rect 469022 410756 469074 410808
rect 469086 410756 469138 410808
rect 469150 410756 469202 410808
rect 469214 410756 469266 410808
rect 469278 410756 469330 410808
rect 469342 410756 469394 410808
rect 469406 410756 469458 410808
rect 469470 410756 469522 410808
rect 469534 410756 469586 410808
rect 469022 410692 469074 410744
rect 469086 410692 469138 410744
rect 469150 410692 469202 410744
rect 469214 410692 469266 410744
rect 469278 410692 469330 410744
rect 469342 410692 469394 410744
rect 469406 410692 469458 410744
rect 469470 410692 469522 410744
rect 469534 410692 469586 410744
rect 478420 410388 478472 410440
rect 478604 410431 478656 410440
rect 478604 410397 478615 410431
rect 478615 410397 478656 410431
rect 478604 410388 478656 410397
rect 485136 410431 485188 410440
rect 485136 410397 485145 410431
rect 485145 410397 485188 410431
rect 485136 410388 485188 410397
rect 475292 410036 475344 410088
rect 481824 410036 481876 410088
rect 490748 409980 490800 410032
rect 470262 409862 470314 409914
rect 470326 409862 470378 409914
rect 470390 409862 470442 409914
rect 470454 409862 470506 409914
rect 470518 409862 470570 409914
rect 470582 409862 470634 409914
rect 470646 409862 470698 409914
rect 470710 409862 470762 409914
rect 470774 409862 470826 409914
rect 470262 409798 470314 409850
rect 470326 409798 470378 409850
rect 470390 409798 470442 409850
rect 470454 409798 470506 409850
rect 470518 409798 470570 409850
rect 470582 409798 470634 409850
rect 470646 409798 470698 409850
rect 470710 409798 470762 409850
rect 470774 409798 470826 409850
rect 470262 409734 470314 409786
rect 470326 409734 470378 409786
rect 470390 409734 470442 409786
rect 470454 409734 470506 409786
rect 470518 409734 470570 409786
rect 470582 409734 470634 409786
rect 470646 409734 470698 409786
rect 470710 409734 470762 409786
rect 470774 409734 470826 409786
rect 515404 409776 515456 409828
rect 535460 409776 535512 409828
rect 470262 409670 470314 409722
rect 470326 409670 470378 409722
rect 470390 409670 470442 409722
rect 470454 409670 470506 409722
rect 470518 409670 470570 409722
rect 470582 409670 470634 409722
rect 470646 409670 470698 409722
rect 470710 409670 470762 409722
rect 470774 409670 470826 409722
rect 470262 409606 470314 409658
rect 470326 409606 470378 409658
rect 470390 409606 470442 409658
rect 470454 409606 470506 409658
rect 470518 409606 470570 409658
rect 470582 409606 470634 409658
rect 470646 409606 470698 409658
rect 470710 409606 470762 409658
rect 470774 409606 470826 409658
rect 475292 408416 475344 408468
rect 493324 408416 493376 408468
rect 478604 407056 478656 407108
rect 535460 407056 535512 407108
rect 515404 404336 515456 404388
rect 535460 404336 535512 404388
rect 516784 402976 516836 403028
rect 535460 402976 535512 403028
rect 518164 398828 518216 398880
rect 535460 398828 535512 398880
rect 519544 396040 519596 396092
rect 535460 396040 535512 396092
rect 470262 391035 470314 391087
rect 470326 391035 470378 391087
rect 470390 391035 470442 391087
rect 470454 391035 470506 391087
rect 470518 391035 470570 391087
rect 470582 391035 470634 391087
rect 470646 391035 470698 391087
rect 470710 391035 470762 391087
rect 470774 391035 470826 391087
rect 470262 390971 470314 391023
rect 470326 390971 470378 391023
rect 470390 390971 470442 391023
rect 470454 390971 470506 391023
rect 470518 390971 470570 391023
rect 470582 390971 470634 391023
rect 470646 390971 470698 391023
rect 470710 390971 470762 391023
rect 470774 390971 470826 391023
rect 470262 390907 470314 390959
rect 470326 390907 470378 390959
rect 470390 390907 470442 390959
rect 470454 390907 470506 390959
rect 470518 390907 470570 390959
rect 470582 390907 470634 390959
rect 470646 390907 470698 390959
rect 470710 390907 470762 390959
rect 470774 390907 470826 390959
rect 470262 390843 470314 390895
rect 470326 390843 470378 390895
rect 470390 390843 470442 390895
rect 470454 390843 470506 390895
rect 470518 390843 470570 390895
rect 470582 390843 470634 390895
rect 470646 390843 470698 390895
rect 470710 390843 470762 390895
rect 470774 390843 470826 390895
rect 470262 390779 470314 390831
rect 470326 390779 470378 390831
rect 470390 390779 470442 390831
rect 470454 390779 470506 390831
rect 470518 390779 470570 390831
rect 470582 390779 470634 390831
rect 470646 390779 470698 390831
rect 470710 390779 470762 390831
rect 470774 390779 470826 390831
rect 471244 390260 471296 390312
rect 471704 390056 471756 390108
rect 469022 389952 469074 390004
rect 469086 389952 469138 390004
rect 469150 389952 469202 390004
rect 469214 389952 469266 390004
rect 469278 389952 469330 390004
rect 469342 389952 469394 390004
rect 469406 389952 469458 390004
rect 469470 389952 469522 390004
rect 469534 389952 469586 390004
rect 469022 389888 469074 389940
rect 469086 389888 469138 389940
rect 469150 389888 469202 389940
rect 469214 389888 469266 389940
rect 469278 389888 469330 389940
rect 469342 389888 469394 389940
rect 469406 389888 469458 389940
rect 469470 389888 469522 389940
rect 469534 389888 469586 389940
rect 469022 389824 469074 389876
rect 469086 389824 469138 389876
rect 469150 389824 469202 389876
rect 469214 389824 469266 389876
rect 469278 389824 469330 389876
rect 469342 389824 469394 389876
rect 469406 389824 469458 389876
rect 469470 389824 469522 389876
rect 469534 389824 469586 389876
rect 469022 389760 469074 389812
rect 469086 389760 469138 389812
rect 469150 389760 469202 389812
rect 469214 389760 469266 389812
rect 469278 389760 469330 389812
rect 469342 389760 469394 389812
rect 469406 389760 469458 389812
rect 469470 389760 469522 389812
rect 469534 389760 469586 389812
rect 469022 389696 469074 389748
rect 469086 389696 469138 389748
rect 469150 389696 469202 389748
rect 469214 389696 469266 389748
rect 469278 389696 469330 389748
rect 469342 389696 469394 389748
rect 469406 389696 469458 389748
rect 469470 389696 469522 389748
rect 469534 389696 469586 389748
rect 479432 389487 479484 389496
rect 479432 389453 479474 389487
rect 479474 389453 479484 389487
rect 479432 389444 479484 389453
rect 493324 389444 493376 389496
rect 475752 389036 475804 389088
rect 483204 389036 483256 389088
rect 486884 389036 486936 389088
rect 470262 388862 470314 388914
rect 470326 388862 470378 388914
rect 470390 388862 470442 388914
rect 470454 388862 470506 388914
rect 470518 388862 470570 388914
rect 470582 388862 470634 388914
rect 470646 388862 470698 388914
rect 470710 388862 470762 388914
rect 470774 388862 470826 388914
rect 470262 388798 470314 388850
rect 470326 388798 470378 388850
rect 470390 388798 470442 388850
rect 470454 388798 470506 388850
rect 470518 388798 470570 388850
rect 470582 388798 470634 388850
rect 470646 388798 470698 388850
rect 470710 388798 470762 388850
rect 470774 388798 470826 388850
rect 470262 388734 470314 388786
rect 470326 388734 470378 388786
rect 470390 388734 470442 388786
rect 470454 388734 470506 388786
rect 470518 388734 470570 388786
rect 470582 388734 470634 388786
rect 470646 388734 470698 388786
rect 470710 388734 470762 388786
rect 470774 388734 470826 388786
rect 470262 388670 470314 388722
rect 470326 388670 470378 388722
rect 470390 388670 470442 388722
rect 470454 388670 470506 388722
rect 470518 388670 470570 388722
rect 470582 388670 470634 388722
rect 470646 388670 470698 388722
rect 470710 388670 470762 388722
rect 470774 388670 470826 388722
rect 470262 388606 470314 388658
rect 470326 388606 470378 388658
rect 470390 388606 470442 388658
rect 470454 388606 470506 388658
rect 470518 388606 470570 388658
rect 470582 388606 470634 388658
rect 470646 388606 470698 388658
rect 470710 388606 470762 388658
rect 470774 388606 470826 388658
rect 475752 387744 475804 387796
rect 479432 387744 479484 387796
rect 515404 387744 515456 387796
rect 494704 387676 494756 387728
rect 483204 386384 483256 386436
rect 484308 386384 484360 386436
rect 520924 373940 520976 373992
rect 535460 373940 535512 373992
rect 536196 373396 536248 373448
rect 522304 372512 522356 372564
rect 535460 372512 535512 372564
rect 484308 369792 484360 369844
rect 535460 369792 535512 369844
rect 520924 367072 520976 367124
rect 535460 367072 535512 367124
rect 515404 365712 515456 365764
rect 535460 365712 535512 365764
rect 522304 361564 522356 361616
rect 535460 361564 535512 361616
rect 470262 358435 470314 358487
rect 470326 358435 470378 358487
rect 470390 358435 470442 358487
rect 470454 358435 470506 358487
rect 470518 358435 470570 358487
rect 470582 358435 470634 358487
rect 470646 358435 470698 358487
rect 470710 358435 470762 358487
rect 470774 358435 470826 358487
rect 470262 358371 470314 358423
rect 470326 358371 470378 358423
rect 470390 358371 470442 358423
rect 470454 358371 470506 358423
rect 470518 358371 470570 358423
rect 470582 358371 470634 358423
rect 470646 358371 470698 358423
rect 470710 358371 470762 358423
rect 470774 358371 470826 358423
rect 470262 358307 470314 358359
rect 470326 358307 470378 358359
rect 470390 358307 470442 358359
rect 470454 358307 470506 358359
rect 470518 358307 470570 358359
rect 470582 358307 470634 358359
rect 470646 358307 470698 358359
rect 470710 358307 470762 358359
rect 470774 358307 470826 358359
rect 470262 358243 470314 358295
rect 470326 358243 470378 358295
rect 470390 358243 470442 358295
rect 470454 358243 470506 358295
rect 470518 358243 470570 358295
rect 470582 358243 470634 358295
rect 470646 358243 470698 358295
rect 470710 358243 470762 358295
rect 470774 358243 470826 358295
rect 470262 358179 470314 358231
rect 470326 358179 470378 358231
rect 470390 358179 470442 358231
rect 470454 358179 470506 358231
rect 470518 358179 470570 358231
rect 470582 358179 470634 358231
rect 470646 358179 470698 358231
rect 470710 358179 470762 358231
rect 470774 358179 470826 358231
rect 471704 357552 471756 357604
rect 475108 357620 475160 357672
rect 478880 357631 478932 357683
rect 481824 357631 481876 357683
rect 484952 357631 485004 357683
rect 469022 357349 469074 357401
rect 469086 357349 469138 357401
rect 469150 357349 469202 357401
rect 469214 357349 469266 357401
rect 469278 357349 469330 357401
rect 469342 357349 469394 357401
rect 469406 357349 469458 357401
rect 469470 357349 469522 357401
rect 469534 357349 469586 357401
rect 469022 357285 469074 357337
rect 469086 357285 469138 357337
rect 469150 357285 469202 357337
rect 469214 357285 469266 357337
rect 469278 357285 469330 357337
rect 469342 357285 469394 357337
rect 469406 357285 469458 357337
rect 469470 357285 469522 357337
rect 469534 357285 469586 357337
rect 469022 357221 469074 357273
rect 469086 357221 469138 357273
rect 469150 357221 469202 357273
rect 469214 357221 469266 357273
rect 469278 357221 469330 357273
rect 469342 357221 469394 357273
rect 469406 357221 469458 357273
rect 469470 357221 469522 357273
rect 469534 357221 469586 357273
rect 469022 357157 469074 357209
rect 469086 357157 469138 357209
rect 469150 357157 469202 357209
rect 469214 357157 469266 357209
rect 469278 357157 469330 357209
rect 469342 357157 469394 357209
rect 469406 357157 469458 357209
rect 469470 357157 469522 357209
rect 469534 357157 469586 357209
rect 469022 357093 469074 357145
rect 469086 357093 469138 357145
rect 469150 357093 469202 357145
rect 469214 357093 469266 357145
rect 469278 357093 469330 357145
rect 469342 357093 469394 357145
rect 469406 357093 469458 357145
rect 469470 357093 469522 357145
rect 469534 357093 469586 357145
rect 477040 356847 477092 356856
rect 477040 356813 477091 356847
rect 477091 356813 477092 356847
rect 477040 356804 477092 356813
rect 480168 356847 480220 356856
rect 480168 356813 480177 356847
rect 480177 356813 480220 356847
rect 480168 356804 480220 356813
rect 483204 356435 483256 356487
rect 486240 356435 486292 356487
rect 492128 356396 492180 356448
rect 470262 356262 470314 356314
rect 470326 356262 470378 356314
rect 470390 356262 470442 356314
rect 470454 356262 470506 356314
rect 470518 356262 470570 356314
rect 470582 356262 470634 356314
rect 470646 356262 470698 356314
rect 470710 356262 470762 356314
rect 470774 356262 470826 356314
rect 470262 356198 470314 356250
rect 470326 356198 470378 356250
rect 470390 356198 470442 356250
rect 470454 356198 470506 356250
rect 470518 356198 470570 356250
rect 470582 356198 470634 356250
rect 470646 356198 470698 356250
rect 470710 356198 470762 356250
rect 470774 356198 470826 356250
rect 470262 356134 470314 356186
rect 470326 356134 470378 356186
rect 470390 356134 470442 356186
rect 470454 356134 470506 356186
rect 470518 356134 470570 356186
rect 470582 356134 470634 356186
rect 470646 356134 470698 356186
rect 470710 356134 470762 356186
rect 470774 356134 470826 356186
rect 470262 356070 470314 356122
rect 470326 356070 470378 356122
rect 470390 356070 470442 356122
rect 470454 356070 470506 356122
rect 470518 356070 470570 356122
rect 470582 356070 470634 356122
rect 470646 356070 470698 356122
rect 470710 356070 470762 356122
rect 470774 356070 470826 356122
rect 470262 356006 470314 356058
rect 470326 356006 470378 356058
rect 470390 356006 470442 356058
rect 470454 356006 470506 356058
rect 470518 356006 470570 356058
rect 470582 356006 470634 356058
rect 470646 356006 470698 356058
rect 470710 356006 470762 356058
rect 470774 356006 470826 356058
rect 480168 354628 480220 354680
rect 516784 354628 516836 354680
rect 483204 354560 483256 354612
rect 520924 354560 520976 354612
rect 477132 354492 477184 354544
rect 496084 354492 496136 354544
rect 486240 353608 486292 353660
rect 525064 353268 525116 353320
rect 470262 342434 470314 342486
rect 470326 342434 470378 342486
rect 470390 342434 470442 342486
rect 470454 342434 470506 342486
rect 470518 342434 470570 342486
rect 470582 342434 470634 342486
rect 470646 342434 470698 342486
rect 470710 342434 470762 342486
rect 470774 342434 470826 342486
rect 470262 342370 470314 342422
rect 470326 342370 470378 342422
rect 470390 342370 470442 342422
rect 470454 342370 470506 342422
rect 470518 342370 470570 342422
rect 470582 342370 470634 342422
rect 470646 342370 470698 342422
rect 470710 342370 470762 342422
rect 470774 342370 470826 342422
rect 470262 342306 470314 342358
rect 470326 342306 470378 342358
rect 470390 342306 470442 342358
rect 470454 342306 470506 342358
rect 470518 342306 470570 342358
rect 470582 342306 470634 342358
rect 470646 342306 470698 342358
rect 470710 342306 470762 342358
rect 470774 342306 470826 342358
rect 470262 342242 470314 342294
rect 470326 342242 470378 342294
rect 470390 342242 470442 342294
rect 470454 342242 470506 342294
rect 470518 342242 470570 342294
rect 470582 342242 470634 342294
rect 470646 342242 470698 342294
rect 470710 342242 470762 342294
rect 470774 342242 470826 342294
rect 470262 342178 470314 342230
rect 470326 342178 470378 342230
rect 470390 342178 470442 342230
rect 470454 342178 470506 342230
rect 470518 342178 470570 342230
rect 470582 342178 470634 342230
rect 470646 342178 470698 342230
rect 470710 342178 470762 342230
rect 470774 342178 470826 342230
rect 471704 341776 471756 341828
rect 471244 341708 471296 341760
rect 469022 341347 469074 341399
rect 469086 341347 469138 341399
rect 469150 341347 469202 341399
rect 469214 341347 469266 341399
rect 469278 341347 469330 341399
rect 469342 341347 469394 341399
rect 469406 341347 469458 341399
rect 469470 341347 469522 341399
rect 469534 341347 469586 341399
rect 469022 341283 469074 341335
rect 469086 341283 469138 341335
rect 469150 341283 469202 341335
rect 469214 341283 469266 341335
rect 469278 341283 469330 341335
rect 469342 341283 469394 341335
rect 469406 341283 469458 341335
rect 469470 341283 469522 341335
rect 469534 341283 469586 341335
rect 469022 341219 469074 341271
rect 469086 341219 469138 341271
rect 469150 341219 469202 341271
rect 469214 341219 469266 341271
rect 469278 341219 469330 341271
rect 469342 341219 469394 341271
rect 469406 341219 469458 341271
rect 469470 341219 469522 341271
rect 469534 341219 469586 341271
rect 469022 341155 469074 341207
rect 469086 341155 469138 341207
rect 469150 341155 469202 341207
rect 469214 341155 469266 341207
rect 469278 341155 469330 341207
rect 469342 341155 469394 341207
rect 469406 341155 469458 341207
rect 469470 341155 469522 341207
rect 469534 341155 469586 341207
rect 469022 341091 469074 341143
rect 469086 341091 469138 341143
rect 469150 341091 469202 341143
rect 469214 341091 469266 341143
rect 469278 341091 469330 341143
rect 469342 341091 469394 341143
rect 469406 341091 469458 341143
rect 469470 341091 469522 341143
rect 469534 341091 469586 341143
rect 482100 340867 482152 340876
rect 474648 340803 474700 340855
rect 482100 340833 482109 340867
rect 482109 340833 482152 340867
rect 482100 340824 482152 340833
rect 485596 340438 485648 340490
rect 475476 340348 475528 340400
rect 478788 340391 478840 340400
rect 478788 340357 478793 340391
rect 478793 340357 478840 340391
rect 478788 340348 478840 340357
rect 492220 340348 492272 340400
rect 470262 340262 470314 340314
rect 470326 340262 470378 340314
rect 470390 340262 470442 340314
rect 470454 340262 470506 340314
rect 470518 340262 470570 340314
rect 470582 340262 470634 340314
rect 470646 340262 470698 340314
rect 470710 340262 470762 340314
rect 470774 340262 470826 340314
rect 470262 340198 470314 340250
rect 470326 340198 470378 340250
rect 470390 340198 470442 340250
rect 470454 340198 470506 340250
rect 470518 340198 470570 340250
rect 470582 340198 470634 340250
rect 470646 340198 470698 340250
rect 470710 340198 470762 340250
rect 470774 340198 470826 340250
rect 470262 340134 470314 340186
rect 470326 340134 470378 340186
rect 470390 340134 470442 340186
rect 470454 340134 470506 340186
rect 470518 340134 470570 340186
rect 470582 340134 470634 340186
rect 470646 340134 470698 340186
rect 470710 340134 470762 340186
rect 470774 340134 470826 340186
rect 470262 340070 470314 340122
rect 470326 340070 470378 340122
rect 470390 340070 470442 340122
rect 470454 340070 470506 340122
rect 470518 340070 470570 340122
rect 470582 340070 470634 340122
rect 470646 340070 470698 340122
rect 470710 340070 470762 340122
rect 470774 340070 470826 340122
rect 470262 340006 470314 340058
rect 470326 340006 470378 340058
rect 470390 340006 470442 340058
rect 470454 340006 470506 340058
rect 470518 340006 470570 340058
rect 470582 340006 470634 340058
rect 470646 340006 470698 340058
rect 470710 340006 470762 340058
rect 470774 340006 470826 340058
rect 475476 339396 475528 339448
rect 478788 339396 478840 339448
rect 536380 339396 536432 339448
rect 482100 339328 482152 339380
rect 515404 339328 515456 339380
rect 497464 339260 497516 339312
rect 523684 338036 523736 338088
rect 535460 338036 535512 338088
rect 525064 332528 525116 332580
rect 535460 332528 535512 332580
rect 485688 331168 485740 331220
rect 535460 331168 535512 331220
rect 523684 325660 523736 325712
rect 535460 325660 535512 325712
rect 470262 322434 470314 322486
rect 470326 322434 470378 322486
rect 470390 322434 470442 322486
rect 470454 322434 470506 322486
rect 470518 322434 470570 322486
rect 470582 322434 470634 322486
rect 470646 322434 470698 322486
rect 470710 322434 470762 322486
rect 470774 322434 470826 322486
rect 470262 322370 470314 322422
rect 470326 322370 470378 322422
rect 470390 322370 470442 322422
rect 470454 322370 470506 322422
rect 470518 322370 470570 322422
rect 470582 322370 470634 322422
rect 470646 322370 470698 322422
rect 470710 322370 470762 322422
rect 470774 322370 470826 322422
rect 470262 322306 470314 322358
rect 470326 322306 470378 322358
rect 470390 322306 470442 322358
rect 470454 322306 470506 322358
rect 470518 322306 470570 322358
rect 470582 322306 470634 322358
rect 470646 322306 470698 322358
rect 470710 322306 470762 322358
rect 470774 322306 470826 322358
rect 470262 322242 470314 322294
rect 470326 322242 470378 322294
rect 470390 322242 470442 322294
rect 470454 322242 470506 322294
rect 470518 322242 470570 322294
rect 470582 322242 470634 322294
rect 470646 322242 470698 322294
rect 470710 322242 470762 322294
rect 470774 322242 470826 322294
rect 470262 322178 470314 322230
rect 470326 322178 470378 322230
rect 470390 322178 470442 322230
rect 470454 322178 470506 322230
rect 470518 322178 470570 322230
rect 470582 322178 470634 322230
rect 470646 322178 470698 322230
rect 470710 322178 470762 322230
rect 470774 322178 470826 322230
rect 471244 321580 471296 321632
rect 469022 321347 469074 321399
rect 469086 321347 469138 321399
rect 469150 321347 469202 321399
rect 469214 321347 469266 321399
rect 469278 321347 469330 321399
rect 469342 321347 469394 321399
rect 469406 321347 469458 321399
rect 469470 321347 469522 321399
rect 469534 321347 469586 321399
rect 469022 321283 469074 321335
rect 469086 321283 469138 321335
rect 469150 321283 469202 321335
rect 469214 321283 469266 321335
rect 469278 321283 469330 321335
rect 469342 321283 469394 321335
rect 469406 321283 469458 321335
rect 469470 321283 469522 321335
rect 469534 321283 469586 321335
rect 469022 321219 469074 321271
rect 469086 321219 469138 321271
rect 469150 321219 469202 321271
rect 469214 321219 469266 321271
rect 469278 321219 469330 321271
rect 469342 321219 469394 321271
rect 469406 321219 469458 321271
rect 469470 321219 469522 321271
rect 469534 321219 469586 321271
rect 469022 321155 469074 321207
rect 469086 321155 469138 321207
rect 469150 321155 469202 321207
rect 469214 321155 469266 321207
rect 469278 321155 469330 321207
rect 469342 321155 469394 321207
rect 469406 321155 469458 321207
rect 469470 321155 469522 321207
rect 469534 321155 469586 321207
rect 469022 321091 469074 321143
rect 469086 321091 469138 321143
rect 469150 321091 469202 321143
rect 469214 321091 469266 321143
rect 469278 321091 469330 321143
rect 469342 321091 469394 321143
rect 469406 321091 469458 321143
rect 469470 321091 469522 321143
rect 469534 321091 469586 321143
rect 475476 320435 475528 320487
rect 482376 320424 482428 320476
rect 479064 320356 479116 320408
rect 485964 320356 486016 320408
rect 492312 320356 492364 320408
rect 470262 320262 470314 320314
rect 470326 320262 470378 320314
rect 470390 320262 470442 320314
rect 470454 320262 470506 320314
rect 470518 320262 470570 320314
rect 470582 320262 470634 320314
rect 470646 320262 470698 320314
rect 470710 320262 470762 320314
rect 470774 320262 470826 320314
rect 470262 320198 470314 320250
rect 470326 320198 470378 320250
rect 470390 320198 470442 320250
rect 470454 320198 470506 320250
rect 470518 320198 470570 320250
rect 470582 320198 470634 320250
rect 470646 320198 470698 320250
rect 470710 320198 470762 320250
rect 470774 320198 470826 320250
rect 470262 320134 470314 320186
rect 470326 320134 470378 320186
rect 470390 320134 470442 320186
rect 470454 320134 470506 320186
rect 470518 320134 470570 320186
rect 470582 320134 470634 320186
rect 470646 320134 470698 320186
rect 470710 320134 470762 320186
rect 470774 320134 470826 320186
rect 470262 320070 470314 320122
rect 470326 320070 470378 320122
rect 470390 320070 470442 320122
rect 470454 320070 470506 320122
rect 470518 320070 470570 320122
rect 470582 320070 470634 320122
rect 470646 320070 470698 320122
rect 470710 320070 470762 320122
rect 470774 320070 470826 320122
rect 470262 320006 470314 320058
rect 470326 320006 470378 320058
rect 470390 320006 470442 320058
rect 470454 320006 470506 320058
rect 470518 320006 470570 320058
rect 470582 320006 470634 320058
rect 470646 320006 470698 320058
rect 470710 320006 470762 320058
rect 470774 320006 470826 320058
rect 475476 318724 475528 318776
rect 479064 318724 479116 318776
rect 536288 318724 536340 318776
rect 482376 318656 482428 318708
rect 536564 318656 536616 318708
rect 485964 318588 486016 318640
rect 536012 318588 536064 318640
rect 498844 318520 498896 318572
rect 470262 307034 470314 307086
rect 470326 307034 470378 307086
rect 470390 307034 470442 307086
rect 470454 307034 470506 307086
rect 470518 307034 470570 307086
rect 470582 307034 470634 307086
rect 470646 307034 470698 307086
rect 470710 307034 470762 307086
rect 470774 307034 470826 307086
rect 470262 306970 470314 307022
rect 470326 306970 470378 307022
rect 470390 306970 470442 307022
rect 470454 306970 470506 307022
rect 470518 306970 470570 307022
rect 470582 306970 470634 307022
rect 470646 306970 470698 307022
rect 470710 306970 470762 307022
rect 470774 306970 470826 307022
rect 470262 306906 470314 306958
rect 470326 306906 470378 306958
rect 470390 306906 470442 306958
rect 470454 306906 470506 306958
rect 470518 306906 470570 306958
rect 470582 306906 470634 306958
rect 470646 306906 470698 306958
rect 470710 306906 470762 306958
rect 470774 306906 470826 306958
rect 470262 306842 470314 306894
rect 470326 306842 470378 306894
rect 470390 306842 470442 306894
rect 470454 306842 470506 306894
rect 470518 306842 470570 306894
rect 470582 306842 470634 306894
rect 470646 306842 470698 306894
rect 470710 306842 470762 306894
rect 470774 306842 470826 306894
rect 470262 306778 470314 306830
rect 470326 306778 470378 306830
rect 470390 306778 470442 306830
rect 470454 306778 470506 306830
rect 470518 306778 470570 306830
rect 470582 306778 470634 306830
rect 470646 306778 470698 306830
rect 470710 306778 470762 306830
rect 470774 306778 470826 306830
rect 471244 306280 471296 306332
rect 473728 306232 473780 306284
rect 469022 305949 469074 306001
rect 469086 305949 469138 306001
rect 469150 305949 469202 306001
rect 469214 305949 469266 306001
rect 469278 305949 469330 306001
rect 469342 305949 469394 306001
rect 469406 305949 469458 306001
rect 469470 305949 469522 306001
rect 469534 305949 469586 306001
rect 469022 305885 469074 305937
rect 469086 305885 469138 305937
rect 469150 305885 469202 305937
rect 469214 305885 469266 305937
rect 469278 305885 469330 305937
rect 469342 305885 469394 305937
rect 469406 305885 469458 305937
rect 469470 305885 469522 305937
rect 469534 305885 469586 305937
rect 469022 305821 469074 305873
rect 469086 305821 469138 305873
rect 469150 305821 469202 305873
rect 469214 305821 469266 305873
rect 469278 305821 469330 305873
rect 469342 305821 469394 305873
rect 469406 305821 469458 305873
rect 469470 305821 469522 305873
rect 469534 305821 469586 305873
rect 469022 305757 469074 305809
rect 469086 305757 469138 305809
rect 469150 305757 469202 305809
rect 469214 305757 469266 305809
rect 469278 305757 469330 305809
rect 469342 305757 469394 305809
rect 469406 305757 469458 305809
rect 469470 305757 469522 305809
rect 469534 305757 469586 305809
rect 469022 305693 469074 305745
rect 469086 305693 469138 305745
rect 469150 305693 469202 305745
rect 469214 305693 469266 305745
rect 469278 305693 469330 305745
rect 469342 305693 469394 305745
rect 469406 305693 469458 305745
rect 469470 305693 469522 305745
rect 469534 305693 469586 305745
rect 478604 305439 478656 305448
rect 478604 305405 478614 305439
rect 478614 305405 478656 305439
rect 478604 305396 478656 305405
rect 485136 305439 485188 305448
rect 485136 305405 485144 305439
rect 485144 305405 485188 305439
rect 485136 305396 485188 305405
rect 475292 305036 475344 305088
rect 481824 305036 481876 305088
rect 490564 304988 490616 305040
rect 470262 304862 470314 304914
rect 470326 304862 470378 304914
rect 470390 304862 470442 304914
rect 470454 304862 470506 304914
rect 470518 304862 470570 304914
rect 470582 304862 470634 304914
rect 470646 304862 470698 304914
rect 470710 304862 470762 304914
rect 470774 304862 470826 304914
rect 470262 304798 470314 304850
rect 470326 304798 470378 304850
rect 470390 304798 470442 304850
rect 470454 304798 470506 304850
rect 470518 304798 470570 304850
rect 470582 304798 470634 304850
rect 470646 304798 470698 304850
rect 470710 304798 470762 304850
rect 470774 304798 470826 304850
rect 470262 304734 470314 304786
rect 470326 304734 470378 304786
rect 470390 304734 470442 304786
rect 470454 304734 470506 304786
rect 470518 304734 470570 304786
rect 470582 304734 470634 304786
rect 470646 304734 470698 304786
rect 470710 304734 470762 304786
rect 470774 304734 470826 304786
rect 470262 304670 470314 304722
rect 470326 304670 470378 304722
rect 470390 304670 470442 304722
rect 470454 304670 470506 304722
rect 470518 304670 470570 304722
rect 470582 304670 470634 304722
rect 470646 304670 470698 304722
rect 470710 304670 470762 304722
rect 470774 304670 470826 304722
rect 470262 304606 470314 304658
rect 470326 304606 470378 304658
rect 470390 304606 470442 304658
rect 470454 304606 470506 304658
rect 470518 304606 470570 304658
rect 470582 304606 470634 304658
rect 470646 304606 470698 304658
rect 470710 304606 470762 304658
rect 470774 304606 470826 304658
rect 475292 303560 475344 303612
rect 478604 303560 478656 303612
rect 481824 303560 481876 303612
rect 485136 303560 485188 303612
rect 536472 303560 536524 303612
rect 536656 303492 536708 303544
rect 518164 303424 518216 303476
rect 500224 303356 500276 303408
rect 491944 300772 491996 300824
rect 535460 300772 535512 300824
rect 492036 299412 492088 299464
rect 535460 299412 535512 299464
rect 490748 298052 490800 298104
rect 535460 298052 535512 298104
rect 492128 296624 492180 296676
rect 535552 296624 535604 296676
rect 493324 296556 493376 296608
rect 535460 296556 535512 296608
rect 492220 295264 492272 295316
rect 535460 295264 535512 295316
rect 492312 293904 492364 293956
rect 535552 293904 535604 293956
rect 490564 292476 490616 292528
rect 535460 292476 535512 292528
rect 492956 289824 493008 289876
rect 535460 289824 535512 289876
rect 491944 288396 491996 288448
rect 535460 288396 535512 288448
rect 470262 287435 470314 287487
rect 470326 287435 470378 287487
rect 470390 287435 470442 287487
rect 470454 287435 470506 287487
rect 470518 287435 470570 287487
rect 470582 287435 470634 287487
rect 470646 287435 470698 287487
rect 470710 287435 470762 287487
rect 470774 287435 470826 287487
rect 470262 287371 470314 287423
rect 470326 287371 470378 287423
rect 470390 287371 470442 287423
rect 470454 287371 470506 287423
rect 470518 287371 470570 287423
rect 470582 287371 470634 287423
rect 470646 287371 470698 287423
rect 470710 287371 470762 287423
rect 470774 287371 470826 287423
rect 470262 287307 470314 287359
rect 470326 287307 470378 287359
rect 470390 287307 470442 287359
rect 470454 287307 470506 287359
rect 470518 287307 470570 287359
rect 470582 287307 470634 287359
rect 470646 287307 470698 287359
rect 470710 287307 470762 287359
rect 470774 287307 470826 287359
rect 470262 287243 470314 287295
rect 470326 287243 470378 287295
rect 470390 287243 470442 287295
rect 470454 287243 470506 287295
rect 470518 287243 470570 287295
rect 470582 287243 470634 287295
rect 470646 287243 470698 287295
rect 470710 287243 470762 287295
rect 470774 287243 470826 287295
rect 470262 287179 470314 287231
rect 470326 287179 470378 287231
rect 470390 287179 470442 287231
rect 470454 287179 470506 287231
rect 470518 287179 470570 287231
rect 470582 287179 470634 287231
rect 470646 287179 470698 287231
rect 470710 287179 470762 287231
rect 470774 287179 470826 287231
rect 471244 286628 471296 286680
rect 488632 286628 488684 286680
rect 471704 286492 471756 286544
rect 469022 286350 469074 286402
rect 469086 286350 469138 286402
rect 469150 286350 469202 286402
rect 469214 286350 469266 286402
rect 469278 286350 469330 286402
rect 469342 286350 469394 286402
rect 469406 286350 469458 286402
rect 469470 286350 469522 286402
rect 469534 286350 469586 286402
rect 469022 286286 469074 286338
rect 469086 286286 469138 286338
rect 469150 286286 469202 286338
rect 469214 286286 469266 286338
rect 469278 286286 469330 286338
rect 469342 286286 469394 286338
rect 469406 286286 469458 286338
rect 469470 286286 469522 286338
rect 469534 286286 469586 286338
rect 469022 286222 469074 286274
rect 469086 286222 469138 286274
rect 469150 286222 469202 286274
rect 469214 286222 469266 286274
rect 469278 286222 469330 286274
rect 469342 286222 469394 286274
rect 469406 286222 469458 286274
rect 469470 286222 469522 286274
rect 469534 286222 469586 286274
rect 469022 286158 469074 286210
rect 469086 286158 469138 286210
rect 469150 286158 469202 286210
rect 469214 286158 469266 286210
rect 469278 286158 469330 286210
rect 469342 286158 469394 286210
rect 469406 286158 469458 286210
rect 469470 286158 469522 286210
rect 469534 286158 469586 286210
rect 469022 286094 469074 286146
rect 469086 286094 469138 286146
rect 469150 286094 469202 286146
rect 469214 286094 469266 286146
rect 469278 286094 469330 286146
rect 469342 286094 469394 286146
rect 469406 286094 469458 286146
rect 469470 286094 469522 286146
rect 469534 286094 469586 286146
rect 479432 285855 479484 285864
rect 479432 285821 479474 285855
rect 479474 285821 479484 285855
rect 479432 285812 479484 285821
rect 492956 285608 493008 285660
rect 475752 285436 475804 285488
rect 483204 285436 483256 285488
rect 486884 285436 486936 285488
rect 470262 285262 470314 285314
rect 470326 285262 470378 285314
rect 470390 285262 470442 285314
rect 470454 285262 470506 285314
rect 470518 285262 470570 285314
rect 470582 285262 470634 285314
rect 470646 285262 470698 285314
rect 470710 285262 470762 285314
rect 470774 285262 470826 285314
rect 470262 285198 470314 285250
rect 470326 285198 470378 285250
rect 470390 285198 470442 285250
rect 470454 285198 470506 285250
rect 470518 285198 470570 285250
rect 470582 285198 470634 285250
rect 470646 285198 470698 285250
rect 470710 285198 470762 285250
rect 470774 285198 470826 285250
rect 470262 285134 470314 285186
rect 470326 285134 470378 285186
rect 470390 285134 470442 285186
rect 470454 285134 470506 285186
rect 470518 285134 470570 285186
rect 470582 285134 470634 285186
rect 470646 285134 470698 285186
rect 470710 285134 470762 285186
rect 470774 285134 470826 285186
rect 470262 285070 470314 285122
rect 470326 285070 470378 285122
rect 470390 285070 470442 285122
rect 470454 285070 470506 285122
rect 470518 285070 470570 285122
rect 470582 285070 470634 285122
rect 470646 285070 470698 285122
rect 470710 285070 470762 285122
rect 470774 285070 470826 285122
rect 470262 285006 470314 285058
rect 470326 285006 470378 285058
rect 470390 285006 470442 285058
rect 470454 285006 470506 285058
rect 470518 285006 470570 285058
rect 470582 285006 470634 285058
rect 470646 285006 470698 285058
rect 470710 285006 470762 285058
rect 470774 285006 470826 285058
rect 475752 284248 475804 284300
rect 479432 284248 479484 284300
rect 536104 284248 536156 284300
rect 483204 284180 483256 284232
rect 522304 284180 522356 284232
rect 486884 284112 486936 284164
rect 523684 284112 523736 284164
rect 501604 284044 501656 284096
rect 471704 270444 471756 270496
rect 473728 270444 473780 270496
rect 470262 267435 470314 267487
rect 470326 267435 470378 267487
rect 470390 267435 470442 267487
rect 470454 267435 470506 267487
rect 470518 267435 470570 267487
rect 470582 267435 470634 267487
rect 470646 267435 470698 267487
rect 470710 267435 470762 267487
rect 470774 267435 470826 267487
rect 470262 267371 470314 267423
rect 470326 267371 470378 267423
rect 470390 267371 470442 267423
rect 470454 267371 470506 267423
rect 470518 267371 470570 267423
rect 470582 267371 470634 267423
rect 470646 267371 470698 267423
rect 470710 267371 470762 267423
rect 470774 267371 470826 267423
rect 470262 267307 470314 267359
rect 470326 267307 470378 267359
rect 470390 267307 470442 267359
rect 470454 267307 470506 267359
rect 470518 267307 470570 267359
rect 470582 267307 470634 267359
rect 470646 267307 470698 267359
rect 470710 267307 470762 267359
rect 470774 267307 470826 267359
rect 470262 267243 470314 267295
rect 470326 267243 470378 267295
rect 470390 267243 470442 267295
rect 470454 267243 470506 267295
rect 470518 267243 470570 267295
rect 470582 267243 470634 267295
rect 470646 267243 470698 267295
rect 470710 267243 470762 267295
rect 470774 267243 470826 267295
rect 470262 267179 470314 267231
rect 470326 267179 470378 267231
rect 470390 267179 470442 267231
rect 470454 267179 470506 267231
rect 470518 267179 470570 267231
rect 470582 267179 470634 267231
rect 470646 267179 470698 267231
rect 470710 267179 470762 267231
rect 470774 267179 470826 267231
rect 473728 266500 473780 266552
rect 469022 266349 469074 266401
rect 469086 266349 469138 266401
rect 469150 266349 469202 266401
rect 469214 266349 469266 266401
rect 469278 266349 469330 266401
rect 469342 266349 469394 266401
rect 469406 266349 469458 266401
rect 469470 266349 469522 266401
rect 469534 266349 469586 266401
rect 469022 266285 469074 266337
rect 469086 266285 469138 266337
rect 469150 266285 469202 266337
rect 469214 266285 469266 266337
rect 469278 266285 469330 266337
rect 469342 266285 469394 266337
rect 469406 266285 469458 266337
rect 469470 266285 469522 266337
rect 469534 266285 469586 266337
rect 469022 266221 469074 266273
rect 469086 266221 469138 266273
rect 469150 266221 469202 266273
rect 469214 266221 469266 266273
rect 469278 266221 469330 266273
rect 469342 266221 469394 266273
rect 469406 266221 469458 266273
rect 469470 266221 469522 266273
rect 469534 266221 469586 266273
rect 469022 266157 469074 266209
rect 469086 266157 469138 266209
rect 469150 266157 469202 266209
rect 469214 266157 469266 266209
rect 469278 266157 469330 266209
rect 469342 266157 469394 266209
rect 469406 266157 469458 266209
rect 469470 266157 469522 266209
rect 469534 266157 469586 266209
rect 469022 266093 469074 266145
rect 469086 266093 469138 266145
rect 469150 266093 469202 266145
rect 469214 266093 469266 266145
rect 469278 266093 469330 266145
rect 469342 266093 469394 266145
rect 469406 266093 469458 266145
rect 469470 266093 469522 266145
rect 469534 266093 469586 266145
rect 477132 265863 477184 265872
rect 477132 265829 477135 265863
rect 477135 265829 477184 265863
rect 477132 265820 477184 265829
rect 491944 265956 491996 266008
rect 480168 265435 480220 265487
rect 483204 265435 483256 265487
rect 486240 265435 486292 265487
rect 470262 265262 470314 265314
rect 470326 265262 470378 265314
rect 470390 265262 470442 265314
rect 470454 265262 470506 265314
rect 470518 265262 470570 265314
rect 470582 265262 470634 265314
rect 470646 265262 470698 265314
rect 470710 265262 470762 265314
rect 470774 265262 470826 265314
rect 470262 265198 470314 265250
rect 470326 265198 470378 265250
rect 470390 265198 470442 265250
rect 470454 265198 470506 265250
rect 470518 265198 470570 265250
rect 470582 265198 470634 265250
rect 470646 265198 470698 265250
rect 470710 265198 470762 265250
rect 470774 265198 470826 265250
rect 470262 265134 470314 265186
rect 470326 265134 470378 265186
rect 470390 265134 470442 265186
rect 470454 265134 470506 265186
rect 470518 265134 470570 265186
rect 470582 265134 470634 265186
rect 470646 265134 470698 265186
rect 470710 265134 470762 265186
rect 470774 265134 470826 265186
rect 470262 265070 470314 265122
rect 470326 265070 470378 265122
rect 470390 265070 470442 265122
rect 470454 265070 470506 265122
rect 470518 265070 470570 265122
rect 470582 265070 470634 265122
rect 470646 265070 470698 265122
rect 470710 265070 470762 265122
rect 470774 265070 470826 265122
rect 470262 265006 470314 265058
rect 470326 265006 470378 265058
rect 470390 265006 470442 265058
rect 470454 265006 470506 265058
rect 470518 265006 470570 265058
rect 470582 265006 470634 265058
rect 470646 265006 470698 265058
rect 470710 265006 470762 265058
rect 470774 265006 470826 265058
rect 477132 263508 477184 263560
rect 480168 263508 480220 263560
rect 483204 263508 483256 263560
rect 486240 263508 486292 263560
rect 494796 263440 494848 263492
rect 495072 263508 495124 263560
rect 535920 263508 535972 263560
rect 536380 263440 536432 263492
rect 519544 263372 519596 263424
rect 502984 263304 503036 263356
rect 473728 206932 473780 206984
rect 580172 206932 580224 206984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 470262 451485 470826 451491
rect 470314 451479 470326 451485
rect 470378 451479 470390 451485
rect 470442 451479 470454 451485
rect 470506 451479 470518 451485
rect 470570 451479 470582 451485
rect 470634 451479 470646 451485
rect 470698 451479 470710 451485
rect 470762 451479 470774 451485
rect 470506 451433 470516 451479
rect 470572 451433 470582 451479
rect 470262 451423 470276 451433
rect 470332 451423 470356 451433
rect 470412 451423 470436 451433
rect 470492 451423 470516 451433
rect 470572 451423 470596 451433
rect 470652 451423 470676 451433
rect 470732 451423 470756 451433
rect 470812 451423 470826 451433
rect 470262 451421 470826 451423
rect 470314 451399 470326 451421
rect 470378 451399 470390 451421
rect 470442 451399 470454 451421
rect 470506 451399 470518 451421
rect 470570 451399 470582 451421
rect 470634 451399 470646 451421
rect 470698 451399 470710 451421
rect 470762 451399 470774 451421
rect 470506 451369 470516 451399
rect 470572 451369 470582 451399
rect 470262 451357 470276 451369
rect 470332 451357 470356 451369
rect 470412 451357 470436 451369
rect 470492 451357 470516 451369
rect 470572 451357 470596 451369
rect 470652 451357 470676 451369
rect 470732 451357 470756 451369
rect 470812 451357 470826 451369
rect 470506 451343 470516 451357
rect 470572 451343 470582 451357
rect 470314 451319 470326 451343
rect 470378 451319 470390 451343
rect 470442 451319 470454 451343
rect 470506 451319 470518 451343
rect 470570 451319 470582 451343
rect 470634 451319 470646 451343
rect 470698 451319 470710 451343
rect 470762 451319 470774 451343
rect 470506 451305 470516 451319
rect 470572 451305 470582 451319
rect 470262 451293 470276 451305
rect 470332 451293 470356 451305
rect 470412 451293 470436 451305
rect 470492 451293 470516 451305
rect 470572 451293 470596 451305
rect 470652 451293 470676 451305
rect 470732 451293 470756 451305
rect 470812 451293 470826 451305
rect 470506 451263 470516 451293
rect 470572 451263 470582 451293
rect 470314 451241 470326 451263
rect 470378 451241 470390 451263
rect 470442 451241 470454 451263
rect 470506 451241 470518 451263
rect 470570 451241 470582 451263
rect 470634 451241 470646 451263
rect 470698 451241 470710 451263
rect 470762 451241 470774 451263
rect 470262 451239 470826 451241
rect 470262 451229 470276 451239
rect 470332 451229 470356 451239
rect 470412 451229 470436 451239
rect 470492 451229 470516 451239
rect 470572 451229 470596 451239
rect 470652 451229 470676 451239
rect 470732 451229 470756 451239
rect 470812 451229 470826 451239
rect 470506 451183 470516 451229
rect 470572 451183 470582 451229
rect 470314 451177 470326 451183
rect 470378 451177 470390 451183
rect 470442 451177 470454 451183
rect 470506 451177 470518 451183
rect 470570 451177 470582 451183
rect 470634 451177 470646 451183
rect 470698 451177 470710 451183
rect 470762 451177 470774 451183
rect 470262 451171 470826 451177
rect 471256 450758 471376 450786
rect 469022 450399 469586 450405
rect 469074 450393 469086 450399
rect 469138 450393 469150 450399
rect 469202 450393 469214 450399
rect 469266 450393 469278 450399
rect 469330 450393 469342 450399
rect 469394 450393 469406 450399
rect 469458 450393 469470 450399
rect 469522 450393 469534 450399
rect 469266 450347 469276 450393
rect 469332 450347 469342 450393
rect 469022 450337 469036 450347
rect 469092 450337 469116 450347
rect 469172 450337 469196 450347
rect 469252 450337 469276 450347
rect 469332 450337 469356 450347
rect 469412 450337 469436 450347
rect 469492 450337 469516 450347
rect 469572 450337 469586 450347
rect 469022 450335 469586 450337
rect 469074 450313 469086 450335
rect 469138 450313 469150 450335
rect 469202 450313 469214 450335
rect 469266 450313 469278 450335
rect 469330 450313 469342 450335
rect 469394 450313 469406 450335
rect 469458 450313 469470 450335
rect 469522 450313 469534 450335
rect 469266 450283 469276 450313
rect 469332 450283 469342 450313
rect 469022 450271 469036 450283
rect 469092 450271 469116 450283
rect 469172 450271 469196 450283
rect 469252 450271 469276 450283
rect 469332 450271 469356 450283
rect 469412 450271 469436 450283
rect 469492 450271 469516 450283
rect 469572 450271 469586 450283
rect 469266 450257 469276 450271
rect 469332 450257 469342 450271
rect 469074 450233 469086 450257
rect 469138 450233 469150 450257
rect 469202 450233 469214 450257
rect 469266 450233 469278 450257
rect 469330 450233 469342 450257
rect 469394 450233 469406 450257
rect 469458 450233 469470 450257
rect 469522 450233 469534 450257
rect 469266 450219 469276 450233
rect 469332 450219 469342 450233
rect 469022 450207 469036 450219
rect 469092 450207 469116 450219
rect 469172 450207 469196 450219
rect 469252 450207 469276 450219
rect 469332 450207 469356 450219
rect 469412 450207 469436 450219
rect 469492 450207 469516 450219
rect 469572 450207 469586 450219
rect 469266 450177 469276 450207
rect 469332 450177 469342 450207
rect 469074 450155 469086 450177
rect 469138 450155 469150 450177
rect 469202 450155 469214 450177
rect 469266 450155 469278 450177
rect 469330 450155 469342 450177
rect 469394 450155 469406 450177
rect 469458 450155 469470 450177
rect 469522 450155 469534 450177
rect 469022 450153 469586 450155
rect 469022 450143 469036 450153
rect 469092 450143 469116 450153
rect 469172 450143 469196 450153
rect 469252 450143 469276 450153
rect 469332 450143 469356 450153
rect 469412 450143 469436 450153
rect 469492 450143 469516 450153
rect 469572 450143 469586 450153
rect 469266 450097 469276 450143
rect 469332 450097 469342 450143
rect 469074 450091 469086 450097
rect 469138 450091 469150 450097
rect 469202 450091 469214 450097
rect 469266 450091 469278 450097
rect 469330 450091 469342 450097
rect 469394 450091 469406 450097
rect 469458 450091 469470 450097
rect 469522 450091 469534 450097
rect 469022 450085 469586 450091
rect 470262 449314 470826 449320
rect 470314 449308 470326 449314
rect 470378 449308 470390 449314
rect 470442 449308 470454 449314
rect 470506 449308 470518 449314
rect 470570 449308 470582 449314
rect 470634 449308 470646 449314
rect 470698 449308 470710 449314
rect 470762 449308 470774 449314
rect 470506 449262 470516 449308
rect 470572 449262 470582 449308
rect 470262 449252 470276 449262
rect 470332 449252 470356 449262
rect 470412 449252 470436 449262
rect 470492 449252 470516 449262
rect 470572 449252 470596 449262
rect 470652 449252 470676 449262
rect 470732 449252 470756 449262
rect 470812 449252 470826 449262
rect 470262 449250 470826 449252
rect 470314 449228 470326 449250
rect 470378 449228 470390 449250
rect 470442 449228 470454 449250
rect 470506 449228 470518 449250
rect 470570 449228 470582 449250
rect 470634 449228 470646 449250
rect 470698 449228 470710 449250
rect 470762 449228 470774 449250
rect 470506 449198 470516 449228
rect 470572 449198 470582 449228
rect 470262 449186 470276 449198
rect 470332 449186 470356 449198
rect 470412 449186 470436 449198
rect 470492 449186 470516 449198
rect 470572 449186 470596 449198
rect 470652 449186 470676 449198
rect 470732 449186 470756 449198
rect 470812 449186 470826 449198
rect 470506 449172 470516 449186
rect 470572 449172 470582 449186
rect 470314 449148 470326 449172
rect 470378 449148 470390 449172
rect 470442 449148 470454 449172
rect 470506 449148 470518 449172
rect 470570 449148 470582 449172
rect 470634 449148 470646 449172
rect 470698 449148 470710 449172
rect 470762 449148 470774 449172
rect 470506 449134 470516 449148
rect 470572 449134 470582 449148
rect 470262 449122 470276 449134
rect 470332 449122 470356 449134
rect 470412 449122 470436 449134
rect 470492 449122 470516 449134
rect 470572 449122 470596 449134
rect 470652 449122 470676 449134
rect 470732 449122 470756 449134
rect 470812 449122 470826 449134
rect 470506 449092 470516 449122
rect 470572 449092 470582 449122
rect 470314 449070 470326 449092
rect 470378 449070 470390 449092
rect 470442 449070 470454 449092
rect 470506 449070 470518 449092
rect 470570 449070 470582 449092
rect 470634 449070 470646 449092
rect 470698 449070 470710 449092
rect 470762 449070 470774 449092
rect 470262 449068 470826 449070
rect 470262 449058 470276 449068
rect 470332 449058 470356 449068
rect 470412 449058 470436 449068
rect 470492 449058 470516 449068
rect 470572 449058 470596 449068
rect 470652 449058 470676 449068
rect 470732 449058 470756 449068
rect 470812 449058 470826 449068
rect 470506 449012 470516 449058
rect 470572 449012 470582 449058
rect 470314 449006 470326 449012
rect 470378 449006 470390 449012
rect 470442 449006 470454 449012
rect 470506 449006 470518 449012
rect 470570 449006 470582 449012
rect 470634 449006 470646 449012
rect 470698 449006 470710 449012
rect 470762 449006 470774 449012
rect 470262 449000 470826 449006
rect 470262 433086 470826 433092
rect 470314 433080 470326 433086
rect 470378 433080 470390 433086
rect 470442 433080 470454 433086
rect 470506 433080 470518 433086
rect 470570 433080 470582 433086
rect 470634 433080 470646 433086
rect 470698 433080 470710 433086
rect 470762 433080 470774 433086
rect 470506 433034 470516 433080
rect 470572 433034 470582 433080
rect 470262 433024 470276 433034
rect 470332 433024 470356 433034
rect 470412 433024 470436 433034
rect 470492 433024 470516 433034
rect 470572 433024 470596 433034
rect 470652 433024 470676 433034
rect 470732 433024 470756 433034
rect 470812 433024 470826 433034
rect 470262 433022 470826 433024
rect 470314 433000 470326 433022
rect 470378 433000 470390 433022
rect 470442 433000 470454 433022
rect 470506 433000 470518 433022
rect 470570 433000 470582 433022
rect 470634 433000 470646 433022
rect 470698 433000 470710 433022
rect 470762 433000 470774 433022
rect 470506 432970 470516 433000
rect 470572 432970 470582 433000
rect 470262 432958 470276 432970
rect 470332 432958 470356 432970
rect 470412 432958 470436 432970
rect 470492 432958 470516 432970
rect 470572 432958 470596 432970
rect 470652 432958 470676 432970
rect 470732 432958 470756 432970
rect 470812 432958 470826 432970
rect 470506 432944 470516 432958
rect 470572 432944 470582 432958
rect 470314 432920 470326 432944
rect 470378 432920 470390 432944
rect 470442 432920 470454 432944
rect 470506 432920 470518 432944
rect 470570 432920 470582 432944
rect 470634 432920 470646 432944
rect 470698 432920 470710 432944
rect 470762 432920 470774 432944
rect 470506 432906 470516 432920
rect 470572 432906 470582 432920
rect 470262 432894 470276 432906
rect 470332 432894 470356 432906
rect 470412 432894 470436 432906
rect 470492 432894 470516 432906
rect 470572 432894 470596 432906
rect 470652 432894 470676 432906
rect 470732 432894 470756 432906
rect 470812 432894 470826 432906
rect 470506 432864 470516 432894
rect 470572 432864 470582 432894
rect 470314 432842 470326 432864
rect 470378 432842 470390 432864
rect 470442 432842 470454 432864
rect 470506 432842 470518 432864
rect 470570 432842 470582 432864
rect 470634 432842 470646 432864
rect 470698 432842 470710 432864
rect 470762 432842 470774 432864
rect 470262 432840 470826 432842
rect 470262 432830 470276 432840
rect 470332 432830 470356 432840
rect 470412 432830 470436 432840
rect 470492 432830 470516 432840
rect 470572 432830 470596 432840
rect 470652 432830 470676 432840
rect 470732 432830 470756 432840
rect 470812 432830 470826 432840
rect 470506 432784 470516 432830
rect 470572 432784 470582 432830
rect 470314 432778 470326 432784
rect 470378 432778 470390 432784
rect 470442 432778 470454 432784
rect 470506 432778 470518 432784
rect 470570 432778 470582 432784
rect 470634 432778 470646 432784
rect 470698 432778 470710 432784
rect 470762 432778 470774 432784
rect 470262 432772 470826 432778
rect 471256 432290 471284 450758
rect 471348 450702 471376 450758
rect 471336 450696 471388 450702
rect 471336 450638 471388 450644
rect 474108 450350 474554 450378
rect 474108 449721 474136 450350
rect 477843 450256 477899 450265
rect 477843 450191 477899 450200
rect 481160 450256 481216 450265
rect 481160 450191 481216 450200
rect 484477 450256 484533 450265
rect 484477 450191 484533 450200
rect 487793 450256 487849 450265
rect 487793 450191 487849 450200
rect 474094 449712 474150 449721
rect 474094 449647 474150 449656
rect 475384 449488 475436 449494
rect 475384 449430 475436 449436
rect 478696 449488 478748 449494
rect 478696 449430 478748 449436
rect 482008 449488 482060 449494
rect 482008 449430 482060 449436
rect 485320 449488 485372 449494
rect 485320 449430 485372 449436
rect 475396 445738 475424 449430
rect 478708 446282 478736 449430
rect 478696 446276 478748 446282
rect 478696 446218 478748 446224
rect 482020 445874 482048 449430
rect 485332 445874 485360 449430
rect 491944 449404 491996 449410
rect 491944 449346 491996 449352
rect 482008 445868 482060 445874
rect 482008 445810 482060 445816
rect 485320 445868 485372 445874
rect 485320 445810 485372 445816
rect 475384 445732 475436 445738
rect 475384 445674 475436 445680
rect 490564 443012 490616 443018
rect 490564 442954 490616 442960
rect 483570 432304 483626 432313
rect 471612 432290 471664 432296
rect 471256 432262 471612 432290
rect 469022 431999 469586 432005
rect 469074 431993 469086 431999
rect 469138 431993 469150 431999
rect 469202 431993 469214 431999
rect 469266 431993 469278 431999
rect 469330 431993 469342 431999
rect 469394 431993 469406 431999
rect 469458 431993 469470 431999
rect 469522 431993 469534 431999
rect 469266 431947 469276 431993
rect 469332 431947 469342 431993
rect 469022 431937 469036 431947
rect 469092 431937 469116 431947
rect 469172 431937 469196 431947
rect 469252 431937 469276 431947
rect 469332 431937 469356 431947
rect 469412 431937 469436 431947
rect 469492 431937 469516 431947
rect 469572 431937 469586 431947
rect 469022 431935 469586 431937
rect 469074 431913 469086 431935
rect 469138 431913 469150 431935
rect 469202 431913 469214 431935
rect 469266 431913 469278 431935
rect 469330 431913 469342 431935
rect 469394 431913 469406 431935
rect 469458 431913 469470 431935
rect 469522 431913 469534 431935
rect 469266 431883 469276 431913
rect 469332 431883 469342 431913
rect 469022 431871 469036 431883
rect 469092 431871 469116 431883
rect 469172 431871 469196 431883
rect 469252 431871 469276 431883
rect 469332 431871 469356 431883
rect 469412 431871 469436 431883
rect 469492 431871 469516 431883
rect 469572 431871 469586 431883
rect 469266 431857 469276 431871
rect 469332 431857 469342 431871
rect 469074 431833 469086 431857
rect 469138 431833 469150 431857
rect 469202 431833 469214 431857
rect 469266 431833 469278 431857
rect 469330 431833 469342 431857
rect 469394 431833 469406 431857
rect 469458 431833 469470 431857
rect 469522 431833 469534 431857
rect 469266 431819 469276 431833
rect 469332 431819 469342 431833
rect 469022 431807 469036 431819
rect 469092 431807 469116 431819
rect 469172 431807 469196 431819
rect 469252 431807 469276 431819
rect 469332 431807 469356 431819
rect 469412 431807 469436 431819
rect 469492 431807 469516 431819
rect 469572 431807 469586 431819
rect 469266 431777 469276 431807
rect 469332 431777 469342 431807
rect 469074 431755 469086 431777
rect 469138 431755 469150 431777
rect 469202 431755 469214 431777
rect 469266 431755 469278 431777
rect 469330 431755 469342 431777
rect 469394 431755 469406 431777
rect 469458 431755 469470 431777
rect 469522 431755 469534 431777
rect 469022 431753 469586 431755
rect 469022 431743 469036 431753
rect 469092 431743 469116 431753
rect 469172 431743 469196 431753
rect 469252 431743 469276 431753
rect 469332 431743 469356 431753
rect 469412 431743 469436 431753
rect 469492 431743 469516 431753
rect 469572 431743 469586 431753
rect 469266 431697 469276 431743
rect 469332 431697 469342 431743
rect 469074 431691 469086 431697
rect 469138 431691 469150 431697
rect 469202 431691 469214 431697
rect 469266 431691 469278 431697
rect 469330 431691 469342 431697
rect 469394 431691 469406 431697
rect 469458 431691 469470 431697
rect 469522 431691 469534 431697
rect 469022 431685 469586 431691
rect 470262 430914 470826 430920
rect 470314 430908 470326 430914
rect 470378 430908 470390 430914
rect 470442 430908 470454 430914
rect 470506 430908 470518 430914
rect 470570 430908 470582 430914
rect 470634 430908 470646 430914
rect 470698 430908 470710 430914
rect 470762 430908 470774 430914
rect 470506 430862 470516 430908
rect 470572 430862 470582 430908
rect 470262 430852 470276 430862
rect 470332 430852 470356 430862
rect 470412 430852 470436 430862
rect 470492 430852 470516 430862
rect 470572 430852 470596 430862
rect 470652 430852 470676 430862
rect 470732 430852 470756 430862
rect 470812 430852 470826 430862
rect 470262 430850 470826 430852
rect 470314 430828 470326 430850
rect 470378 430828 470390 430850
rect 470442 430828 470454 430850
rect 470506 430828 470518 430850
rect 470570 430828 470582 430850
rect 470634 430828 470646 430850
rect 470698 430828 470710 430850
rect 470762 430828 470774 430850
rect 470506 430798 470516 430828
rect 470572 430798 470582 430828
rect 470262 430786 470276 430798
rect 470332 430786 470356 430798
rect 470412 430786 470436 430798
rect 470492 430786 470516 430798
rect 470572 430786 470596 430798
rect 470652 430786 470676 430798
rect 470732 430786 470756 430798
rect 470812 430786 470826 430798
rect 470506 430772 470516 430786
rect 470572 430772 470582 430786
rect 470314 430748 470326 430772
rect 470378 430748 470390 430772
rect 470442 430748 470454 430772
rect 470506 430748 470518 430772
rect 470570 430748 470582 430772
rect 470634 430748 470646 430772
rect 470698 430748 470710 430772
rect 470762 430748 470774 430772
rect 470506 430734 470516 430748
rect 470572 430734 470582 430748
rect 470262 430722 470276 430734
rect 470332 430722 470356 430734
rect 470412 430722 470436 430734
rect 470492 430722 470516 430734
rect 470572 430722 470596 430734
rect 470652 430722 470676 430734
rect 470732 430722 470756 430734
rect 470812 430722 470826 430734
rect 470506 430692 470516 430722
rect 470572 430692 470582 430722
rect 470314 430670 470326 430692
rect 470378 430670 470390 430692
rect 470442 430670 470454 430692
rect 470506 430670 470518 430692
rect 470570 430670 470582 430692
rect 470634 430670 470646 430692
rect 470698 430670 470710 430692
rect 470762 430670 470774 430692
rect 470262 430668 470826 430670
rect 470262 430658 470276 430668
rect 470332 430658 470356 430668
rect 470412 430658 470436 430668
rect 470492 430658 470516 430668
rect 470572 430658 470596 430668
rect 470652 430658 470676 430668
rect 470732 430658 470756 430668
rect 470812 430658 470826 430668
rect 470506 430612 470516 430658
rect 470572 430612 470582 430658
rect 470314 430606 470326 430612
rect 470378 430606 470390 430612
rect 470442 430606 470454 430612
rect 470506 430606 470518 430612
rect 470570 430606 470582 430612
rect 470634 430606 470646 430612
rect 470698 430606 470710 430612
rect 470762 430606 470774 430612
rect 470262 430600 470826 430606
rect 470262 412086 470826 412092
rect 470314 412080 470326 412086
rect 470378 412080 470390 412086
rect 470442 412080 470454 412086
rect 470506 412080 470518 412086
rect 470570 412080 470582 412086
rect 470634 412080 470646 412086
rect 470698 412080 470710 412086
rect 470762 412080 470774 412086
rect 470506 412034 470516 412080
rect 470572 412034 470582 412080
rect 470262 412024 470276 412034
rect 470332 412024 470356 412034
rect 470412 412024 470436 412034
rect 470492 412024 470516 412034
rect 470572 412024 470596 412034
rect 470652 412024 470676 412034
rect 470732 412024 470756 412034
rect 470812 412024 470826 412034
rect 470262 412022 470826 412024
rect 470314 412000 470326 412022
rect 470378 412000 470390 412022
rect 470442 412000 470454 412022
rect 470506 412000 470518 412022
rect 470570 412000 470582 412022
rect 470634 412000 470646 412022
rect 470698 412000 470710 412022
rect 470762 412000 470774 412022
rect 470506 411970 470516 412000
rect 470572 411970 470582 412000
rect 470262 411958 470276 411970
rect 470332 411958 470356 411970
rect 470412 411958 470436 411970
rect 470492 411958 470516 411970
rect 470572 411958 470596 411970
rect 470652 411958 470676 411970
rect 470732 411958 470756 411970
rect 470812 411958 470826 411970
rect 470506 411944 470516 411958
rect 470572 411944 470582 411958
rect 470314 411920 470326 411944
rect 470378 411920 470390 411944
rect 470442 411920 470454 411944
rect 470506 411920 470518 411944
rect 470570 411920 470582 411944
rect 470634 411920 470646 411944
rect 470698 411920 470710 411944
rect 470762 411920 470774 411944
rect 470506 411906 470516 411920
rect 470572 411906 470582 411920
rect 470262 411894 470276 411906
rect 470332 411894 470356 411906
rect 470412 411894 470436 411906
rect 470492 411894 470516 411906
rect 470572 411894 470596 411906
rect 470652 411894 470676 411906
rect 470732 411894 470756 411906
rect 470812 411894 470826 411906
rect 470506 411864 470516 411894
rect 470572 411864 470582 411894
rect 470314 411842 470326 411864
rect 470378 411842 470390 411864
rect 470442 411842 470454 411864
rect 470506 411842 470518 411864
rect 470570 411842 470582 411864
rect 470634 411842 470646 411864
rect 470698 411842 470710 411864
rect 470762 411842 470774 411864
rect 470262 411840 470826 411842
rect 470262 411830 470276 411840
rect 470332 411830 470356 411840
rect 470412 411830 470436 411840
rect 470492 411830 470516 411840
rect 470572 411830 470596 411840
rect 470652 411830 470676 411840
rect 470732 411830 470756 411840
rect 470812 411830 470826 411840
rect 470506 411784 470516 411830
rect 470572 411784 470582 411830
rect 470314 411778 470326 411784
rect 470378 411778 470390 411784
rect 470442 411778 470454 411784
rect 470506 411778 470518 411784
rect 470570 411778 470582 411784
rect 470634 411778 470646 411784
rect 470698 411778 470710 411784
rect 470762 411778 470774 411784
rect 470262 411772 470826 411778
rect 471256 411262 471284 432262
rect 483143 432262 483570 432290
rect 483570 432239 483626 432248
rect 471612 432232 471664 432238
rect 481270 432168 481326 432177
rect 481326 432126 481573 432154
rect 481270 432103 481326 432112
rect 474292 431990 474685 432018
rect 488092 431990 488461 432018
rect 474292 431905 474320 431990
rect 488092 431905 488120 431990
rect 474278 431896 474334 431905
rect 474278 431831 474334 431840
rect 488078 431896 488134 431905
rect 488078 431831 488134 431840
rect 478102 431624 478158 431633
rect 478102 431559 478158 431568
rect 478972 431452 479024 431458
rect 478972 431394 479024 431400
rect 485780 431452 485832 431458
rect 485780 431394 485832 431400
rect 475476 431087 475528 431093
rect 475476 431029 475528 431035
rect 475488 429146 475516 431029
rect 475476 429140 475528 429146
rect 475476 429082 475528 429088
rect 478984 427961 479012 431394
rect 482376 431087 482428 431093
rect 482376 431029 482428 431035
rect 478970 427952 479026 427961
rect 478970 427887 479026 427896
rect 482388 427854 482416 431029
rect 485792 427961 485820 431394
rect 490576 429146 490604 442954
rect 490564 429140 490616 429146
rect 490564 429082 490616 429088
rect 485778 427952 485834 427961
rect 485778 427887 485834 427896
rect 482376 427848 482428 427854
rect 482376 427790 482428 427796
rect 473728 411284 473780 411290
rect 471244 411256 471296 411262
rect 473728 411226 473780 411232
rect 471244 411198 471296 411204
rect 469022 411000 469586 411006
rect 469074 410994 469086 411000
rect 469138 410994 469150 411000
rect 469202 410994 469214 411000
rect 469266 410994 469278 411000
rect 469330 410994 469342 411000
rect 469394 410994 469406 411000
rect 469458 410994 469470 411000
rect 469522 410994 469534 411000
rect 469266 410948 469276 410994
rect 469332 410948 469342 410994
rect 469022 410938 469036 410948
rect 469092 410938 469116 410948
rect 469172 410938 469196 410948
rect 469252 410938 469276 410948
rect 469332 410938 469356 410948
rect 469412 410938 469436 410948
rect 469492 410938 469516 410948
rect 469572 410938 469586 410948
rect 469022 410936 469586 410938
rect 469074 410914 469086 410936
rect 469138 410914 469150 410936
rect 469202 410914 469214 410936
rect 469266 410914 469278 410936
rect 469330 410914 469342 410936
rect 469394 410914 469406 410936
rect 469458 410914 469470 410936
rect 469522 410914 469534 410936
rect 469266 410884 469276 410914
rect 469332 410884 469342 410914
rect 469022 410872 469036 410884
rect 469092 410872 469116 410884
rect 469172 410872 469196 410884
rect 469252 410872 469276 410884
rect 469332 410872 469356 410884
rect 469412 410872 469436 410884
rect 469492 410872 469516 410884
rect 469572 410872 469586 410884
rect 469266 410858 469276 410872
rect 469332 410858 469342 410872
rect 469074 410834 469086 410858
rect 469138 410834 469150 410858
rect 469202 410834 469214 410858
rect 469266 410834 469278 410858
rect 469330 410834 469342 410858
rect 469394 410834 469406 410858
rect 469458 410834 469470 410858
rect 469522 410834 469534 410858
rect 469266 410820 469276 410834
rect 469332 410820 469342 410834
rect 469022 410808 469036 410820
rect 469092 410808 469116 410820
rect 469172 410808 469196 410820
rect 469252 410808 469276 410820
rect 469332 410808 469356 410820
rect 469412 410808 469436 410820
rect 469492 410808 469516 410820
rect 469572 410808 469586 410820
rect 469266 410778 469276 410808
rect 469332 410778 469342 410808
rect 469074 410756 469086 410778
rect 469138 410756 469150 410778
rect 469202 410756 469214 410778
rect 469266 410756 469278 410778
rect 469330 410756 469342 410778
rect 469394 410756 469406 410778
rect 469458 410756 469470 410778
rect 469522 410756 469534 410778
rect 469022 410754 469586 410756
rect 469022 410744 469036 410754
rect 469092 410744 469116 410754
rect 469172 410744 469196 410754
rect 469252 410744 469276 410754
rect 469332 410744 469356 410754
rect 469412 410744 469436 410754
rect 469492 410744 469516 410754
rect 469572 410744 469586 410754
rect 469266 410698 469276 410744
rect 469332 410698 469342 410744
rect 469074 410692 469086 410698
rect 469138 410692 469150 410698
rect 469202 410692 469214 410698
rect 469266 410692 469278 410698
rect 469330 410692 469342 410698
rect 469394 410692 469406 410698
rect 469458 410692 469470 410698
rect 469522 410692 469534 410698
rect 469022 410686 469586 410692
rect 470262 409914 470826 409920
rect 470314 409908 470326 409914
rect 470378 409908 470390 409914
rect 470442 409908 470454 409914
rect 470506 409908 470518 409914
rect 470570 409908 470582 409914
rect 470634 409908 470646 409914
rect 470698 409908 470710 409914
rect 470762 409908 470774 409914
rect 470506 409862 470516 409908
rect 470572 409862 470582 409908
rect 470262 409852 470276 409862
rect 470332 409852 470356 409862
rect 470412 409852 470436 409862
rect 470492 409852 470516 409862
rect 470572 409852 470596 409862
rect 470652 409852 470676 409862
rect 470732 409852 470756 409862
rect 470812 409852 470826 409862
rect 470262 409850 470826 409852
rect 470314 409828 470326 409850
rect 470378 409828 470390 409850
rect 470442 409828 470454 409850
rect 470506 409828 470518 409850
rect 470570 409828 470582 409850
rect 470634 409828 470646 409850
rect 470698 409828 470710 409850
rect 470762 409828 470774 409850
rect 470506 409798 470516 409828
rect 470572 409798 470582 409828
rect 470262 409786 470276 409798
rect 470332 409786 470356 409798
rect 470412 409786 470436 409798
rect 470492 409786 470516 409798
rect 470572 409786 470596 409798
rect 470652 409786 470676 409798
rect 470732 409786 470756 409798
rect 470812 409786 470826 409798
rect 470506 409772 470516 409786
rect 470572 409772 470582 409786
rect 470314 409748 470326 409772
rect 470378 409748 470390 409772
rect 470442 409748 470454 409772
rect 470506 409748 470518 409772
rect 470570 409748 470582 409772
rect 470634 409748 470646 409772
rect 470698 409748 470710 409772
rect 470762 409748 470774 409772
rect 470506 409734 470516 409748
rect 470572 409734 470582 409748
rect 470262 409722 470276 409734
rect 470332 409722 470356 409734
rect 470412 409722 470436 409734
rect 470492 409722 470516 409734
rect 470572 409722 470596 409734
rect 470652 409722 470676 409734
rect 470732 409722 470756 409734
rect 470812 409722 470826 409734
rect 470506 409692 470516 409722
rect 470572 409692 470582 409722
rect 470314 409670 470326 409692
rect 470378 409670 470390 409692
rect 470442 409670 470454 409692
rect 470506 409670 470518 409692
rect 470570 409670 470582 409692
rect 470634 409670 470646 409692
rect 470698 409670 470710 409692
rect 470762 409670 470774 409692
rect 470262 409668 470826 409670
rect 470262 409658 470276 409668
rect 470332 409658 470356 409668
rect 470412 409658 470436 409668
rect 470492 409658 470516 409668
rect 470572 409658 470596 409668
rect 470652 409658 470676 409668
rect 470732 409658 470756 409668
rect 470812 409658 470826 409668
rect 470506 409612 470516 409658
rect 470572 409612 470582 409658
rect 470314 409606 470326 409612
rect 470378 409606 470390 409612
rect 470442 409606 470454 409612
rect 470506 409606 470518 409612
rect 470570 409606 470582 409612
rect 470634 409606 470646 409612
rect 470698 409606 470710 409612
rect 470762 409606 470774 409612
rect 470262 409600 470826 409606
rect 470262 391087 470826 391093
rect 470314 391081 470326 391087
rect 470378 391081 470390 391087
rect 470442 391081 470454 391087
rect 470506 391081 470518 391087
rect 470570 391081 470582 391087
rect 470634 391081 470646 391087
rect 470698 391081 470710 391087
rect 470762 391081 470774 391087
rect 470506 391035 470516 391081
rect 470572 391035 470582 391081
rect 470262 391025 470276 391035
rect 470332 391025 470356 391035
rect 470412 391025 470436 391035
rect 470492 391025 470516 391035
rect 470572 391025 470596 391035
rect 470652 391025 470676 391035
rect 470732 391025 470756 391035
rect 470812 391025 470826 391035
rect 470262 391023 470826 391025
rect 470314 391001 470326 391023
rect 470378 391001 470390 391023
rect 470442 391001 470454 391023
rect 470506 391001 470518 391023
rect 470570 391001 470582 391023
rect 470634 391001 470646 391023
rect 470698 391001 470710 391023
rect 470762 391001 470774 391023
rect 470506 390971 470516 391001
rect 470572 390971 470582 391001
rect 470262 390959 470276 390971
rect 470332 390959 470356 390971
rect 470412 390959 470436 390971
rect 470492 390959 470516 390971
rect 470572 390959 470596 390971
rect 470652 390959 470676 390971
rect 470732 390959 470756 390971
rect 470812 390959 470826 390971
rect 470506 390945 470516 390959
rect 470572 390945 470582 390959
rect 470314 390921 470326 390945
rect 470378 390921 470390 390945
rect 470442 390921 470454 390945
rect 470506 390921 470518 390945
rect 470570 390921 470582 390945
rect 470634 390921 470646 390945
rect 470698 390921 470710 390945
rect 470762 390921 470774 390945
rect 470506 390907 470516 390921
rect 470572 390907 470582 390921
rect 470262 390895 470276 390907
rect 470332 390895 470356 390907
rect 470412 390895 470436 390907
rect 470492 390895 470516 390907
rect 470572 390895 470596 390907
rect 470652 390895 470676 390907
rect 470732 390895 470756 390907
rect 470812 390895 470826 390907
rect 470506 390865 470516 390895
rect 470572 390865 470582 390895
rect 470314 390843 470326 390865
rect 470378 390843 470390 390865
rect 470442 390843 470454 390865
rect 470506 390843 470518 390865
rect 470570 390843 470582 390865
rect 470634 390843 470646 390865
rect 470698 390843 470710 390865
rect 470762 390843 470774 390865
rect 470262 390841 470826 390843
rect 470262 390831 470276 390841
rect 470332 390831 470356 390841
rect 470412 390831 470436 390841
rect 470492 390831 470516 390841
rect 470572 390831 470596 390841
rect 470652 390831 470676 390841
rect 470732 390831 470756 390841
rect 470812 390831 470826 390841
rect 470506 390785 470516 390831
rect 470572 390785 470582 390831
rect 470314 390779 470326 390785
rect 470378 390779 470390 390785
rect 470442 390779 470454 390785
rect 470506 390779 470518 390785
rect 470570 390779 470582 390785
rect 470634 390779 470646 390785
rect 470698 390779 470710 390785
rect 470762 390779 470774 390785
rect 470262 390773 470826 390779
rect 471256 390318 471284 411198
rect 473740 410961 473768 411226
rect 473726 410952 473782 410961
rect 473726 410887 473782 410896
rect 478420 410440 478472 410446
rect 478420 410382 478472 410388
rect 478604 410440 478656 410446
rect 478604 410382 478656 410388
rect 478432 410145 478460 410382
rect 478418 410136 478474 410145
rect 475292 410088 475344 410094
rect 478418 410071 478474 410080
rect 475292 410030 475344 410036
rect 475304 408474 475332 410030
rect 475292 408468 475344 408474
rect 475292 408410 475344 408416
rect 478616 407114 478644 410382
rect 481019 410258 481047 410516
rect 484136 410502 484298 410530
rect 484136 410417 484164 410502
rect 485136 410440 485188 410446
rect 484122 410408 484178 410417
rect 485136 410382 485188 410388
rect 484122 410343 484178 410352
rect 481019 410230 481128 410258
rect 481100 410122 481128 410230
rect 481362 410136 481418 410145
rect 481100 410094 481362 410122
rect 481362 410071 481418 410080
rect 481824 410088 481876 410094
rect 481824 410030 481876 410036
rect 481836 407153 481864 410030
rect 485148 407153 485176 410382
rect 487549 410258 487577 410516
rect 487549 410230 487660 410258
rect 487632 410122 487660 410230
rect 487802 410136 487858 410145
rect 487632 410094 487802 410122
rect 487802 410071 487858 410080
rect 490748 410032 490800 410038
rect 490748 409974 490800 409980
rect 481822 407144 481878 407153
rect 478604 407108 478656 407114
rect 481822 407079 481878 407088
rect 485134 407144 485190 407153
rect 485134 407079 485190 407088
rect 478604 407050 478656 407056
rect 471244 390312 471296 390318
rect 471244 390254 471296 390260
rect 488552 390238 488658 390266
rect 488552 390153 488580 390238
rect 488538 390144 488594 390153
rect 471704 390108 471756 390114
rect 488538 390079 488594 390088
rect 471704 390050 471756 390056
rect 469022 390004 469586 390010
rect 469074 389998 469086 390004
rect 469138 389998 469150 390004
rect 469202 389998 469214 390004
rect 469266 389998 469278 390004
rect 469330 389998 469342 390004
rect 469394 389998 469406 390004
rect 469458 389998 469470 390004
rect 469522 389998 469534 390004
rect 469266 389952 469276 389998
rect 469332 389952 469342 389998
rect 469022 389942 469036 389952
rect 469092 389942 469116 389952
rect 469172 389942 469196 389952
rect 469252 389942 469276 389952
rect 469332 389942 469356 389952
rect 469412 389942 469436 389952
rect 469492 389942 469516 389952
rect 469572 389942 469586 389952
rect 469022 389940 469586 389942
rect 469074 389918 469086 389940
rect 469138 389918 469150 389940
rect 469202 389918 469214 389940
rect 469266 389918 469278 389940
rect 469330 389918 469342 389940
rect 469394 389918 469406 389940
rect 469458 389918 469470 389940
rect 469522 389918 469534 389940
rect 469266 389888 469276 389918
rect 469332 389888 469342 389918
rect 469022 389876 469036 389888
rect 469092 389876 469116 389888
rect 469172 389876 469196 389888
rect 469252 389876 469276 389888
rect 469332 389876 469356 389888
rect 469412 389876 469436 389888
rect 469492 389876 469516 389888
rect 469572 389876 469586 389888
rect 469266 389862 469276 389876
rect 469332 389862 469342 389876
rect 469074 389838 469086 389862
rect 469138 389838 469150 389862
rect 469202 389838 469214 389862
rect 469266 389838 469278 389862
rect 469330 389838 469342 389862
rect 469394 389838 469406 389862
rect 469458 389838 469470 389862
rect 469522 389838 469534 389862
rect 469266 389824 469276 389838
rect 469332 389824 469342 389838
rect 469022 389812 469036 389824
rect 469092 389812 469116 389824
rect 469172 389812 469196 389824
rect 469252 389812 469276 389824
rect 469332 389812 469356 389824
rect 469412 389812 469436 389824
rect 469492 389812 469516 389824
rect 469572 389812 469586 389824
rect 469266 389782 469276 389812
rect 469332 389782 469342 389812
rect 469074 389760 469086 389782
rect 469138 389760 469150 389782
rect 469202 389760 469214 389782
rect 469266 389760 469278 389782
rect 469330 389760 469342 389782
rect 469394 389760 469406 389782
rect 469458 389760 469470 389782
rect 469522 389760 469534 389782
rect 469022 389758 469586 389760
rect 469022 389748 469036 389758
rect 469092 389748 469116 389758
rect 469172 389748 469196 389758
rect 469252 389748 469276 389758
rect 469332 389748 469356 389758
rect 469412 389748 469436 389758
rect 469492 389748 469516 389758
rect 469572 389748 469586 389758
rect 469266 389702 469276 389748
rect 469332 389702 469342 389748
rect 469074 389696 469086 389702
rect 469138 389696 469150 389702
rect 469202 389696 469214 389702
rect 469266 389696 469278 389702
rect 469330 389696 469342 389702
rect 469394 389696 469406 389702
rect 469458 389696 469470 389702
rect 469522 389696 469534 389702
rect 469022 389690 469586 389696
rect 470262 388914 470826 388920
rect 470314 388908 470326 388914
rect 470378 388908 470390 388914
rect 470442 388908 470454 388914
rect 470506 388908 470518 388914
rect 470570 388908 470582 388914
rect 470634 388908 470646 388914
rect 470698 388908 470710 388914
rect 470762 388908 470774 388914
rect 470506 388862 470516 388908
rect 470572 388862 470582 388908
rect 470262 388852 470276 388862
rect 470332 388852 470356 388862
rect 470412 388852 470436 388862
rect 470492 388852 470516 388862
rect 470572 388852 470596 388862
rect 470652 388852 470676 388862
rect 470732 388852 470756 388862
rect 470812 388852 470826 388862
rect 470262 388850 470826 388852
rect 470314 388828 470326 388850
rect 470378 388828 470390 388850
rect 470442 388828 470454 388850
rect 470506 388828 470518 388850
rect 470570 388828 470582 388850
rect 470634 388828 470646 388850
rect 470698 388828 470710 388850
rect 470762 388828 470774 388850
rect 470506 388798 470516 388828
rect 470572 388798 470582 388828
rect 470262 388786 470276 388798
rect 470332 388786 470356 388798
rect 470412 388786 470436 388798
rect 470492 388786 470516 388798
rect 470572 388786 470596 388798
rect 470652 388786 470676 388798
rect 470732 388786 470756 388798
rect 470812 388786 470826 388798
rect 470506 388772 470516 388786
rect 470572 388772 470582 388786
rect 470314 388748 470326 388772
rect 470378 388748 470390 388772
rect 470442 388748 470454 388772
rect 470506 388748 470518 388772
rect 470570 388748 470582 388772
rect 470634 388748 470646 388772
rect 470698 388748 470710 388772
rect 470762 388748 470774 388772
rect 470506 388734 470516 388748
rect 470572 388734 470582 388748
rect 470262 388722 470276 388734
rect 470332 388722 470356 388734
rect 470412 388722 470436 388734
rect 470492 388722 470516 388734
rect 470572 388722 470596 388734
rect 470652 388722 470676 388734
rect 470732 388722 470756 388734
rect 470812 388722 470826 388734
rect 470506 388692 470516 388722
rect 470572 388692 470582 388722
rect 470314 388670 470326 388692
rect 470378 388670 470390 388692
rect 470442 388670 470454 388692
rect 470506 388670 470518 388692
rect 470570 388670 470582 388692
rect 470634 388670 470646 388692
rect 470698 388670 470710 388692
rect 470762 388670 470774 388692
rect 470262 388668 470826 388670
rect 470262 388658 470276 388668
rect 470332 388658 470356 388668
rect 470412 388658 470436 388668
rect 470492 388658 470516 388668
rect 470572 388658 470596 388668
rect 470652 388658 470676 388668
rect 470732 388658 470756 388668
rect 470812 388658 470826 388668
rect 470506 388612 470516 388658
rect 470572 388612 470582 388658
rect 470314 388606 470326 388612
rect 470378 388606 470390 388612
rect 470442 388606 470454 388612
rect 470506 388606 470518 388612
rect 470570 388606 470582 388612
rect 470634 388606 470646 388612
rect 470698 388606 470710 388612
rect 470762 388606 470774 388612
rect 470262 388600 470826 388606
rect 470262 358487 470826 358493
rect 470314 358481 470326 358487
rect 470378 358481 470390 358487
rect 470442 358481 470454 358487
rect 470506 358481 470518 358487
rect 470570 358481 470582 358487
rect 470634 358481 470646 358487
rect 470698 358481 470710 358487
rect 470762 358481 470774 358487
rect 470506 358435 470516 358481
rect 470572 358435 470582 358481
rect 470262 358425 470276 358435
rect 470332 358425 470356 358435
rect 470412 358425 470436 358435
rect 470492 358425 470516 358435
rect 470572 358425 470596 358435
rect 470652 358425 470676 358435
rect 470732 358425 470756 358435
rect 470812 358425 470826 358435
rect 470262 358423 470826 358425
rect 470314 358401 470326 358423
rect 470378 358401 470390 358423
rect 470442 358401 470454 358423
rect 470506 358401 470518 358423
rect 470570 358401 470582 358423
rect 470634 358401 470646 358423
rect 470698 358401 470710 358423
rect 470762 358401 470774 358423
rect 470506 358371 470516 358401
rect 470572 358371 470582 358401
rect 470262 358359 470276 358371
rect 470332 358359 470356 358371
rect 470412 358359 470436 358371
rect 470492 358359 470516 358371
rect 470572 358359 470596 358371
rect 470652 358359 470676 358371
rect 470732 358359 470756 358371
rect 470812 358359 470826 358371
rect 470506 358345 470516 358359
rect 470572 358345 470582 358359
rect 470314 358321 470326 358345
rect 470378 358321 470390 358345
rect 470442 358321 470454 358345
rect 470506 358321 470518 358345
rect 470570 358321 470582 358345
rect 470634 358321 470646 358345
rect 470698 358321 470710 358345
rect 470762 358321 470774 358345
rect 470506 358307 470516 358321
rect 470572 358307 470582 358321
rect 470262 358295 470276 358307
rect 470332 358295 470356 358307
rect 470412 358295 470436 358307
rect 470492 358295 470516 358307
rect 470572 358295 470596 358307
rect 470652 358295 470676 358307
rect 470732 358295 470756 358307
rect 470812 358295 470826 358307
rect 470506 358265 470516 358295
rect 470572 358265 470582 358295
rect 470314 358243 470326 358265
rect 470378 358243 470390 358265
rect 470442 358243 470454 358265
rect 470506 358243 470518 358265
rect 470570 358243 470582 358265
rect 470634 358243 470646 358265
rect 470698 358243 470710 358265
rect 470762 358243 470774 358265
rect 470262 358241 470826 358243
rect 470262 358231 470276 358241
rect 470332 358231 470356 358241
rect 470412 358231 470436 358241
rect 470492 358231 470516 358241
rect 470572 358231 470596 358241
rect 470652 358231 470676 358241
rect 470732 358231 470756 358241
rect 470812 358231 470826 358241
rect 470506 358185 470516 358231
rect 470572 358185 470582 358231
rect 470314 358179 470326 358185
rect 470378 358179 470390 358185
rect 470442 358179 470454 358185
rect 470506 358179 470518 358185
rect 470570 358179 470582 358185
rect 470634 358179 470646 358185
rect 470698 358179 470710 358185
rect 470762 358179 470774 358185
rect 470262 358173 470826 358179
rect 471716 357610 471744 390050
rect 479432 389496 479484 389502
rect 479432 389438 479484 389444
rect 482098 389464 482154 389473
rect 474936 389337 474964 389436
rect 478648 389337 478676 389436
rect 474922 389328 474978 389337
rect 474922 389263 474978 389272
rect 478634 389328 478690 389337
rect 478634 389263 478690 389272
rect 475752 389088 475804 389094
rect 475752 389030 475804 389036
rect 475764 387802 475792 389030
rect 479444 387802 479472 389438
rect 482154 389422 482374 389450
rect 482098 389399 482154 389408
rect 483204 389088 483256 389094
rect 483204 389030 483256 389036
rect 486884 389088 486936 389094
rect 486884 389030 486936 389036
rect 475752 387796 475804 387802
rect 475752 387738 475804 387744
rect 479432 387796 479484 387802
rect 479432 387738 479484 387744
rect 483216 386442 483244 389030
rect 486896 386481 486924 389030
rect 486882 386472 486938 386481
rect 483204 386436 483256 386442
rect 483204 386378 483256 386384
rect 484308 386436 484360 386442
rect 486882 386407 486938 386416
rect 484308 386378 484360 386384
rect 484320 369850 484348 386378
rect 484308 369844 484360 369850
rect 484308 369786 484360 369792
rect 478878 358048 478934 358057
rect 478878 357983 478934 357992
rect 481822 358048 481878 358057
rect 481822 357983 481878 357992
rect 484950 358048 485006 358057
rect 484950 357983 485006 357992
rect 488354 358048 488410 358057
rect 488354 357983 488410 357992
rect 478892 357689 478920 357983
rect 481836 357689 481864 357983
rect 484964 357689 484992 357983
rect 478880 357683 478932 357689
rect 475108 357672 475160 357678
rect 478880 357625 478932 357631
rect 481824 357683 481876 357689
rect 481824 357625 481876 357631
rect 484952 357683 485004 357689
rect 484952 357625 485004 357631
rect 475108 357614 475160 357620
rect 471704 357604 471756 357610
rect 471704 357546 471756 357552
rect 469022 357401 469586 357407
rect 469074 357395 469086 357401
rect 469138 357395 469150 357401
rect 469202 357395 469214 357401
rect 469266 357395 469278 357401
rect 469330 357395 469342 357401
rect 469394 357395 469406 357401
rect 469458 357395 469470 357401
rect 469522 357395 469534 357401
rect 469266 357349 469276 357395
rect 469332 357349 469342 357395
rect 469022 357339 469036 357349
rect 469092 357339 469116 357349
rect 469172 357339 469196 357349
rect 469252 357339 469276 357349
rect 469332 357339 469356 357349
rect 469412 357339 469436 357349
rect 469492 357339 469516 357349
rect 469572 357339 469586 357349
rect 469022 357337 469586 357339
rect 469074 357315 469086 357337
rect 469138 357315 469150 357337
rect 469202 357315 469214 357337
rect 469266 357315 469278 357337
rect 469330 357315 469342 357337
rect 469394 357315 469406 357337
rect 469458 357315 469470 357337
rect 469522 357315 469534 357337
rect 469266 357285 469276 357315
rect 469332 357285 469342 357315
rect 469022 357273 469036 357285
rect 469092 357273 469116 357285
rect 469172 357273 469196 357285
rect 469252 357273 469276 357285
rect 469332 357273 469356 357285
rect 469412 357273 469436 357285
rect 469492 357273 469516 357285
rect 469572 357273 469586 357285
rect 469266 357259 469276 357273
rect 469332 357259 469342 357273
rect 469074 357235 469086 357259
rect 469138 357235 469150 357259
rect 469202 357235 469214 357259
rect 469266 357235 469278 357259
rect 469330 357235 469342 357259
rect 469394 357235 469406 357259
rect 469458 357235 469470 357259
rect 469522 357235 469534 357259
rect 469266 357221 469276 357235
rect 469332 357221 469342 357235
rect 469022 357209 469036 357221
rect 469092 357209 469116 357221
rect 469172 357209 469196 357221
rect 469252 357209 469276 357221
rect 469332 357209 469356 357221
rect 469412 357209 469436 357221
rect 469492 357209 469516 357221
rect 469572 357209 469586 357221
rect 469266 357179 469276 357209
rect 469332 357179 469342 357209
rect 469074 357157 469086 357179
rect 469138 357157 469150 357179
rect 469202 357157 469214 357179
rect 469266 357157 469278 357179
rect 469330 357157 469342 357179
rect 469394 357157 469406 357179
rect 469458 357157 469470 357179
rect 469522 357157 469534 357179
rect 469022 357155 469586 357157
rect 469022 357145 469036 357155
rect 469092 357145 469116 357155
rect 469172 357145 469196 357155
rect 469252 357145 469276 357155
rect 469332 357145 469356 357155
rect 469412 357145 469436 357155
rect 469492 357145 469516 357155
rect 469572 357145 469586 357155
rect 469266 357099 469276 357145
rect 469332 357099 469342 357145
rect 469074 357093 469086 357099
rect 469138 357093 469150 357099
rect 469202 357093 469214 357099
rect 469266 357093 469278 357099
rect 469330 357093 469342 357099
rect 469394 357093 469406 357099
rect 469458 357093 469470 357099
rect 469522 357093 469534 357099
rect 469022 357087 469586 357093
rect 470262 356314 470826 356320
rect 470314 356308 470326 356314
rect 470378 356308 470390 356314
rect 470442 356308 470454 356314
rect 470506 356308 470518 356314
rect 470570 356308 470582 356314
rect 470634 356308 470646 356314
rect 470698 356308 470710 356314
rect 470762 356308 470774 356314
rect 470506 356262 470516 356308
rect 470572 356262 470582 356308
rect 470262 356252 470276 356262
rect 470332 356252 470356 356262
rect 470412 356252 470436 356262
rect 470492 356252 470516 356262
rect 470572 356252 470596 356262
rect 470652 356252 470676 356262
rect 470732 356252 470756 356262
rect 470812 356252 470826 356262
rect 470262 356250 470826 356252
rect 470314 356228 470326 356250
rect 470378 356228 470390 356250
rect 470442 356228 470454 356250
rect 470506 356228 470518 356250
rect 470570 356228 470582 356250
rect 470634 356228 470646 356250
rect 470698 356228 470710 356250
rect 470762 356228 470774 356250
rect 470506 356198 470516 356228
rect 470572 356198 470582 356228
rect 470262 356186 470276 356198
rect 470332 356186 470356 356198
rect 470412 356186 470436 356198
rect 470492 356186 470516 356198
rect 470572 356186 470596 356198
rect 470652 356186 470676 356198
rect 470732 356186 470756 356198
rect 470812 356186 470826 356198
rect 470506 356172 470516 356186
rect 470572 356172 470582 356186
rect 470314 356148 470326 356172
rect 470378 356148 470390 356172
rect 470442 356148 470454 356172
rect 470506 356148 470518 356172
rect 470570 356148 470582 356172
rect 470634 356148 470646 356172
rect 470698 356148 470710 356172
rect 470762 356148 470774 356172
rect 470506 356134 470516 356148
rect 470572 356134 470582 356148
rect 470262 356122 470276 356134
rect 470332 356122 470356 356134
rect 470412 356122 470436 356134
rect 470492 356122 470516 356134
rect 470572 356122 470596 356134
rect 470652 356122 470676 356134
rect 470732 356122 470756 356134
rect 470812 356122 470826 356134
rect 470506 356092 470516 356122
rect 470572 356092 470582 356122
rect 470314 356070 470326 356092
rect 470378 356070 470390 356092
rect 470442 356070 470454 356092
rect 470506 356070 470518 356092
rect 470570 356070 470582 356092
rect 470634 356070 470646 356092
rect 470698 356070 470710 356092
rect 470762 356070 470774 356092
rect 470262 356068 470826 356070
rect 470262 356058 470276 356068
rect 470332 356058 470356 356068
rect 470412 356058 470436 356068
rect 470492 356058 470516 356068
rect 470572 356058 470596 356068
rect 470652 356058 470676 356068
rect 470732 356058 470756 356068
rect 470812 356058 470826 356068
rect 470506 356012 470516 356058
rect 470572 356012 470582 356058
rect 470314 356006 470326 356012
rect 470378 356006 470390 356012
rect 470442 356006 470454 356012
rect 470506 356006 470518 356012
rect 470570 356006 470582 356012
rect 470634 356006 470646 356012
rect 470698 356006 470710 356012
rect 470762 356006 470774 356012
rect 470262 356000 470826 356006
rect 471716 354674 471744 357546
rect 475014 357504 475070 357513
rect 475120 357490 475148 357614
rect 475070 357462 475148 357490
rect 488368 357490 488396 357983
rect 488368 357462 488487 357490
rect 475014 357439 475070 357448
rect 477040 356856 477092 356862
rect 477040 356798 477092 356804
rect 480168 356856 480220 356862
rect 480168 356798 480220 356804
rect 477052 354674 477080 356798
rect 480180 354686 480208 356798
rect 483204 356487 483256 356493
rect 483204 356429 483256 356435
rect 486240 356487 486292 356493
rect 486240 356429 486292 356435
rect 480168 354680 480220 354686
rect 471716 354646 471928 354674
rect 477052 354646 477172 354674
rect 471900 345014 471928 354646
rect 477144 354550 477172 354646
rect 480168 354622 480220 354628
rect 483216 354618 483244 356429
rect 483204 354612 483256 354618
rect 483204 354554 483256 354560
rect 477132 354544 477184 354550
rect 477132 354486 477184 354492
rect 486252 353666 486280 356429
rect 486240 353660 486292 353666
rect 486240 353602 486292 353608
rect 471716 344986 471928 345014
rect 470262 342486 470826 342492
rect 470314 342480 470326 342486
rect 470378 342480 470390 342486
rect 470442 342480 470454 342486
rect 470506 342480 470518 342486
rect 470570 342480 470582 342486
rect 470634 342480 470646 342486
rect 470698 342480 470710 342486
rect 470762 342480 470774 342486
rect 470506 342434 470516 342480
rect 470572 342434 470582 342480
rect 470262 342424 470276 342434
rect 470332 342424 470356 342434
rect 470412 342424 470436 342434
rect 470492 342424 470516 342434
rect 470572 342424 470596 342434
rect 470652 342424 470676 342434
rect 470732 342424 470756 342434
rect 470812 342424 470826 342434
rect 470262 342422 470826 342424
rect 470314 342400 470326 342422
rect 470378 342400 470390 342422
rect 470442 342400 470454 342422
rect 470506 342400 470518 342422
rect 470570 342400 470582 342422
rect 470634 342400 470646 342422
rect 470698 342400 470710 342422
rect 470762 342400 470774 342422
rect 470506 342370 470516 342400
rect 470572 342370 470582 342400
rect 470262 342358 470276 342370
rect 470332 342358 470356 342370
rect 470412 342358 470436 342370
rect 470492 342358 470516 342370
rect 470572 342358 470596 342370
rect 470652 342358 470676 342370
rect 470732 342358 470756 342370
rect 470812 342358 470826 342370
rect 470506 342344 470516 342358
rect 470572 342344 470582 342358
rect 470314 342320 470326 342344
rect 470378 342320 470390 342344
rect 470442 342320 470454 342344
rect 470506 342320 470518 342344
rect 470570 342320 470582 342344
rect 470634 342320 470646 342344
rect 470698 342320 470710 342344
rect 470762 342320 470774 342344
rect 470506 342306 470516 342320
rect 470572 342306 470582 342320
rect 470262 342294 470276 342306
rect 470332 342294 470356 342306
rect 470412 342294 470436 342306
rect 470492 342294 470516 342306
rect 470572 342294 470596 342306
rect 470652 342294 470676 342306
rect 470732 342294 470756 342306
rect 470812 342294 470826 342306
rect 470506 342264 470516 342294
rect 470572 342264 470582 342294
rect 470314 342242 470326 342264
rect 470378 342242 470390 342264
rect 470442 342242 470454 342264
rect 470506 342242 470518 342264
rect 470570 342242 470582 342264
rect 470634 342242 470646 342264
rect 470698 342242 470710 342264
rect 470762 342242 470774 342264
rect 470262 342240 470826 342242
rect 470262 342230 470276 342240
rect 470332 342230 470356 342240
rect 470412 342230 470436 342240
rect 470492 342230 470516 342240
rect 470572 342230 470596 342240
rect 470652 342230 470676 342240
rect 470732 342230 470756 342240
rect 470812 342230 470826 342240
rect 470506 342184 470516 342230
rect 470572 342184 470582 342230
rect 470314 342178 470326 342184
rect 470378 342178 470390 342184
rect 470442 342178 470454 342184
rect 470506 342178 470518 342184
rect 470570 342178 470582 342184
rect 470634 342178 470646 342184
rect 470698 342178 470710 342184
rect 470762 342178 470774 342184
rect 470262 342172 470826 342178
rect 471716 341834 471744 344986
rect 471704 341828 471756 341834
rect 471704 341770 471756 341776
rect 471244 341760 471296 341766
rect 471244 341702 471296 341708
rect 469022 341399 469586 341405
rect 469074 341393 469086 341399
rect 469138 341393 469150 341399
rect 469202 341393 469214 341399
rect 469266 341393 469278 341399
rect 469330 341393 469342 341399
rect 469394 341393 469406 341399
rect 469458 341393 469470 341399
rect 469522 341393 469534 341399
rect 469266 341347 469276 341393
rect 469332 341347 469342 341393
rect 469022 341337 469036 341347
rect 469092 341337 469116 341347
rect 469172 341337 469196 341347
rect 469252 341337 469276 341347
rect 469332 341337 469356 341347
rect 469412 341337 469436 341347
rect 469492 341337 469516 341347
rect 469572 341337 469586 341347
rect 469022 341335 469586 341337
rect 469074 341313 469086 341335
rect 469138 341313 469150 341335
rect 469202 341313 469214 341335
rect 469266 341313 469278 341335
rect 469330 341313 469342 341335
rect 469394 341313 469406 341335
rect 469458 341313 469470 341335
rect 469522 341313 469534 341335
rect 469266 341283 469276 341313
rect 469332 341283 469342 341313
rect 469022 341271 469036 341283
rect 469092 341271 469116 341283
rect 469172 341271 469196 341283
rect 469252 341271 469276 341283
rect 469332 341271 469356 341283
rect 469412 341271 469436 341283
rect 469492 341271 469516 341283
rect 469572 341271 469586 341283
rect 469266 341257 469276 341271
rect 469332 341257 469342 341271
rect 469074 341233 469086 341257
rect 469138 341233 469150 341257
rect 469202 341233 469214 341257
rect 469266 341233 469278 341257
rect 469330 341233 469342 341257
rect 469394 341233 469406 341257
rect 469458 341233 469470 341257
rect 469522 341233 469534 341257
rect 469266 341219 469276 341233
rect 469332 341219 469342 341233
rect 469022 341207 469036 341219
rect 469092 341207 469116 341219
rect 469172 341207 469196 341219
rect 469252 341207 469276 341219
rect 469332 341207 469356 341219
rect 469412 341207 469436 341219
rect 469492 341207 469516 341219
rect 469572 341207 469586 341219
rect 469266 341177 469276 341207
rect 469332 341177 469342 341207
rect 469074 341155 469086 341177
rect 469138 341155 469150 341177
rect 469202 341155 469214 341177
rect 469266 341155 469278 341177
rect 469330 341155 469342 341177
rect 469394 341155 469406 341177
rect 469458 341155 469470 341177
rect 469522 341155 469534 341177
rect 469022 341153 469586 341155
rect 469022 341143 469036 341153
rect 469092 341143 469116 341153
rect 469172 341143 469196 341153
rect 469252 341143 469276 341153
rect 469332 341143 469356 341153
rect 469412 341143 469436 341153
rect 469492 341143 469516 341153
rect 469572 341143 469586 341153
rect 469266 341097 469276 341143
rect 469332 341097 469342 341143
rect 469074 341091 469086 341097
rect 469138 341091 469150 341097
rect 469202 341091 469214 341097
rect 469266 341091 469278 341097
rect 469330 341091 469342 341097
rect 469394 341091 469406 341097
rect 469458 341091 469470 341097
rect 469522 341091 469534 341097
rect 469022 341085 469586 341091
rect 470262 340314 470826 340320
rect 470314 340308 470326 340314
rect 470378 340308 470390 340314
rect 470442 340308 470454 340314
rect 470506 340308 470518 340314
rect 470570 340308 470582 340314
rect 470634 340308 470646 340314
rect 470698 340308 470710 340314
rect 470762 340308 470774 340314
rect 470506 340262 470516 340308
rect 470572 340262 470582 340308
rect 470262 340252 470276 340262
rect 470332 340252 470356 340262
rect 470412 340252 470436 340262
rect 470492 340252 470516 340262
rect 470572 340252 470596 340262
rect 470652 340252 470676 340262
rect 470732 340252 470756 340262
rect 470812 340252 470826 340262
rect 470262 340250 470826 340252
rect 470314 340228 470326 340250
rect 470378 340228 470390 340250
rect 470442 340228 470454 340250
rect 470506 340228 470518 340250
rect 470570 340228 470582 340250
rect 470634 340228 470646 340250
rect 470698 340228 470710 340250
rect 470762 340228 470774 340250
rect 470506 340198 470516 340228
rect 470572 340198 470582 340228
rect 470262 340186 470276 340198
rect 470332 340186 470356 340198
rect 470412 340186 470436 340198
rect 470492 340186 470516 340198
rect 470572 340186 470596 340198
rect 470652 340186 470676 340198
rect 470732 340186 470756 340198
rect 470812 340186 470826 340198
rect 470506 340172 470516 340186
rect 470572 340172 470582 340186
rect 470314 340148 470326 340172
rect 470378 340148 470390 340172
rect 470442 340148 470454 340172
rect 470506 340148 470518 340172
rect 470570 340148 470582 340172
rect 470634 340148 470646 340172
rect 470698 340148 470710 340172
rect 470762 340148 470774 340172
rect 470506 340134 470516 340148
rect 470572 340134 470582 340148
rect 470262 340122 470276 340134
rect 470332 340122 470356 340134
rect 470412 340122 470436 340134
rect 470492 340122 470516 340134
rect 470572 340122 470596 340134
rect 470652 340122 470676 340134
rect 470732 340122 470756 340134
rect 470812 340122 470826 340134
rect 470506 340092 470516 340122
rect 470572 340092 470582 340122
rect 470314 340070 470326 340092
rect 470378 340070 470390 340092
rect 470442 340070 470454 340092
rect 470506 340070 470518 340092
rect 470570 340070 470582 340092
rect 470634 340070 470646 340092
rect 470698 340070 470710 340092
rect 470762 340070 470774 340092
rect 470262 340068 470826 340070
rect 470262 340058 470276 340068
rect 470332 340058 470356 340068
rect 470412 340058 470436 340068
rect 470492 340058 470516 340068
rect 470572 340058 470596 340068
rect 470652 340058 470676 340068
rect 470732 340058 470756 340068
rect 470812 340058 470826 340068
rect 470506 340012 470516 340058
rect 470572 340012 470582 340058
rect 470314 340006 470326 340012
rect 470378 340006 470390 340012
rect 470442 340006 470454 340012
rect 470506 340006 470518 340012
rect 470570 340006 470582 340012
rect 470634 340006 470646 340012
rect 470698 340006 470710 340012
rect 470762 340006 470774 340012
rect 470262 340000 470826 340006
rect 470262 322486 470826 322492
rect 470314 322480 470326 322486
rect 470378 322480 470390 322486
rect 470442 322480 470454 322486
rect 470506 322480 470518 322486
rect 470570 322480 470582 322486
rect 470634 322480 470646 322486
rect 470698 322480 470710 322486
rect 470762 322480 470774 322486
rect 470506 322434 470516 322480
rect 470572 322434 470582 322480
rect 470262 322424 470276 322434
rect 470332 322424 470356 322434
rect 470412 322424 470436 322434
rect 470492 322424 470516 322434
rect 470572 322424 470596 322434
rect 470652 322424 470676 322434
rect 470732 322424 470756 322434
rect 470812 322424 470826 322434
rect 470262 322422 470826 322424
rect 470314 322400 470326 322422
rect 470378 322400 470390 322422
rect 470442 322400 470454 322422
rect 470506 322400 470518 322422
rect 470570 322400 470582 322422
rect 470634 322400 470646 322422
rect 470698 322400 470710 322422
rect 470762 322400 470774 322422
rect 470506 322370 470516 322400
rect 470572 322370 470582 322400
rect 470262 322358 470276 322370
rect 470332 322358 470356 322370
rect 470412 322358 470436 322370
rect 470492 322358 470516 322370
rect 470572 322358 470596 322370
rect 470652 322358 470676 322370
rect 470732 322358 470756 322370
rect 470812 322358 470826 322370
rect 470506 322344 470516 322358
rect 470572 322344 470582 322358
rect 470314 322320 470326 322344
rect 470378 322320 470390 322344
rect 470442 322320 470454 322344
rect 470506 322320 470518 322344
rect 470570 322320 470582 322344
rect 470634 322320 470646 322344
rect 470698 322320 470710 322344
rect 470762 322320 470774 322344
rect 470506 322306 470516 322320
rect 470572 322306 470582 322320
rect 470262 322294 470276 322306
rect 470332 322294 470356 322306
rect 470412 322294 470436 322306
rect 470492 322294 470516 322306
rect 470572 322294 470596 322306
rect 470652 322294 470676 322306
rect 470732 322294 470756 322306
rect 470812 322294 470826 322306
rect 470506 322264 470516 322294
rect 470572 322264 470582 322294
rect 470314 322242 470326 322264
rect 470378 322242 470390 322264
rect 470442 322242 470454 322264
rect 470506 322242 470518 322264
rect 470570 322242 470582 322264
rect 470634 322242 470646 322264
rect 470698 322242 470710 322264
rect 470762 322242 470774 322264
rect 470262 322240 470826 322242
rect 470262 322230 470276 322240
rect 470332 322230 470356 322240
rect 470412 322230 470436 322240
rect 470492 322230 470516 322240
rect 470572 322230 470596 322240
rect 470652 322230 470676 322240
rect 470732 322230 470756 322240
rect 470812 322230 470826 322240
rect 470506 322184 470516 322230
rect 470572 322184 470582 322230
rect 470314 322178 470326 322184
rect 470378 322178 470390 322184
rect 470442 322178 470454 322184
rect 470506 322178 470518 322184
rect 470570 322178 470582 322184
rect 470634 322178 470646 322184
rect 470698 322178 470710 322184
rect 470762 322178 470774 322184
rect 470262 322172 470826 322178
rect 471256 321638 471284 341702
rect 484504 341414 484577 341442
rect 484504 341306 484532 341414
rect 484412 341278 484532 341306
rect 484412 341057 484440 341278
rect 484398 341048 484454 341057
rect 477906 340992 477915 341048
rect 477971 340992 477980 341048
rect 481223 340992 481232 341048
rect 481288 340992 481297 341048
rect 487885 340992 487894 341048
rect 487950 340992 487959 341048
rect 484398 340983 484454 340992
rect 482100 340876 482152 340882
rect 474648 340855 474700 340861
rect 482100 340818 482152 340824
rect 474648 340797 474700 340803
rect 474554 340504 474610 340513
rect 474660 340490 474688 340797
rect 474610 340462 474688 340490
rect 474554 340439 474610 340448
rect 475476 340400 475528 340406
rect 475476 340342 475528 340348
rect 478788 340400 478840 340406
rect 478788 340342 478840 340348
rect 475488 339454 475516 340342
rect 478800 339454 478828 340342
rect 475476 339448 475528 339454
rect 475476 339390 475528 339396
rect 478788 339448 478840 339454
rect 478788 339390 478840 339396
rect 482112 339386 482140 340818
rect 485596 340490 485648 340496
rect 485596 340432 485648 340438
rect 482100 339380 482152 339386
rect 482100 339322 482152 339328
rect 485608 335354 485636 340432
rect 485608 335326 485728 335354
rect 485700 331226 485728 335326
rect 485688 331220 485740 331226
rect 485688 331162 485740 331168
rect 471244 321632 471296 321638
rect 471244 321574 471296 321580
rect 469022 321399 469586 321405
rect 469074 321393 469086 321399
rect 469138 321393 469150 321399
rect 469202 321393 469214 321399
rect 469266 321393 469278 321399
rect 469330 321393 469342 321399
rect 469394 321393 469406 321399
rect 469458 321393 469470 321399
rect 469522 321393 469534 321399
rect 469266 321347 469276 321393
rect 469332 321347 469342 321393
rect 469022 321337 469036 321347
rect 469092 321337 469116 321347
rect 469172 321337 469196 321347
rect 469252 321337 469276 321347
rect 469332 321337 469356 321347
rect 469412 321337 469436 321347
rect 469492 321337 469516 321347
rect 469572 321337 469586 321347
rect 469022 321335 469586 321337
rect 469074 321313 469086 321335
rect 469138 321313 469150 321335
rect 469202 321313 469214 321335
rect 469266 321313 469278 321335
rect 469330 321313 469342 321335
rect 469394 321313 469406 321335
rect 469458 321313 469470 321335
rect 469522 321313 469534 321335
rect 469266 321283 469276 321313
rect 469332 321283 469342 321313
rect 469022 321271 469036 321283
rect 469092 321271 469116 321283
rect 469172 321271 469196 321283
rect 469252 321271 469276 321283
rect 469332 321271 469356 321283
rect 469412 321271 469436 321283
rect 469492 321271 469516 321283
rect 469572 321271 469586 321283
rect 469266 321257 469276 321271
rect 469332 321257 469342 321271
rect 469074 321233 469086 321257
rect 469138 321233 469150 321257
rect 469202 321233 469214 321257
rect 469266 321233 469278 321257
rect 469330 321233 469342 321257
rect 469394 321233 469406 321257
rect 469458 321233 469470 321257
rect 469522 321233 469534 321257
rect 469266 321219 469276 321233
rect 469332 321219 469342 321233
rect 469022 321207 469036 321219
rect 469092 321207 469116 321219
rect 469172 321207 469196 321219
rect 469252 321207 469276 321219
rect 469332 321207 469356 321219
rect 469412 321207 469436 321219
rect 469492 321207 469516 321219
rect 469572 321207 469586 321219
rect 469266 321177 469276 321207
rect 469332 321177 469342 321207
rect 469074 321155 469086 321177
rect 469138 321155 469150 321177
rect 469202 321155 469214 321177
rect 469266 321155 469278 321177
rect 469330 321155 469342 321177
rect 469394 321155 469406 321177
rect 469458 321155 469470 321177
rect 469522 321155 469534 321177
rect 469022 321153 469586 321155
rect 469022 321143 469036 321153
rect 469092 321143 469116 321153
rect 469172 321143 469196 321153
rect 469252 321143 469276 321153
rect 469332 321143 469356 321153
rect 469412 321143 469436 321153
rect 469492 321143 469516 321153
rect 469572 321143 469586 321153
rect 469266 321097 469276 321143
rect 469332 321097 469342 321143
rect 469074 321091 469086 321097
rect 469138 321091 469150 321097
rect 469202 321091 469214 321097
rect 469266 321091 469278 321097
rect 469330 321091 469342 321097
rect 469394 321091 469406 321097
rect 469458 321091 469470 321097
rect 469522 321091 469534 321097
rect 469022 321085 469586 321091
rect 470262 320314 470826 320320
rect 470314 320308 470326 320314
rect 470378 320308 470390 320314
rect 470442 320308 470454 320314
rect 470506 320308 470518 320314
rect 470570 320308 470582 320314
rect 470634 320308 470646 320314
rect 470698 320308 470710 320314
rect 470762 320308 470774 320314
rect 470506 320262 470516 320308
rect 470572 320262 470582 320308
rect 470262 320252 470276 320262
rect 470332 320252 470356 320262
rect 470412 320252 470436 320262
rect 470492 320252 470516 320262
rect 470572 320252 470596 320262
rect 470652 320252 470676 320262
rect 470732 320252 470756 320262
rect 470812 320252 470826 320262
rect 470262 320250 470826 320252
rect 470314 320228 470326 320250
rect 470378 320228 470390 320250
rect 470442 320228 470454 320250
rect 470506 320228 470518 320250
rect 470570 320228 470582 320250
rect 470634 320228 470646 320250
rect 470698 320228 470710 320250
rect 470762 320228 470774 320250
rect 470506 320198 470516 320228
rect 470572 320198 470582 320228
rect 470262 320186 470276 320198
rect 470332 320186 470356 320198
rect 470412 320186 470436 320198
rect 470492 320186 470516 320198
rect 470572 320186 470596 320198
rect 470652 320186 470676 320198
rect 470732 320186 470756 320198
rect 470812 320186 470826 320198
rect 470506 320172 470516 320186
rect 470572 320172 470582 320186
rect 470314 320148 470326 320172
rect 470378 320148 470390 320172
rect 470442 320148 470454 320172
rect 470506 320148 470518 320172
rect 470570 320148 470582 320172
rect 470634 320148 470646 320172
rect 470698 320148 470710 320172
rect 470762 320148 470774 320172
rect 470506 320134 470516 320148
rect 470572 320134 470582 320148
rect 470262 320122 470276 320134
rect 470332 320122 470356 320134
rect 470412 320122 470436 320134
rect 470492 320122 470516 320134
rect 470572 320122 470596 320134
rect 470652 320122 470676 320134
rect 470732 320122 470756 320134
rect 470812 320122 470826 320134
rect 470506 320092 470516 320122
rect 470572 320092 470582 320122
rect 470314 320070 470326 320092
rect 470378 320070 470390 320092
rect 470442 320070 470454 320092
rect 470506 320070 470518 320092
rect 470570 320070 470582 320092
rect 470634 320070 470646 320092
rect 470698 320070 470710 320092
rect 470762 320070 470774 320092
rect 470262 320068 470826 320070
rect 470262 320058 470276 320068
rect 470332 320058 470356 320068
rect 470412 320058 470436 320068
rect 470492 320058 470516 320068
rect 470572 320058 470596 320068
rect 470652 320058 470676 320068
rect 470732 320058 470756 320068
rect 470812 320058 470826 320068
rect 470506 320012 470516 320058
rect 470572 320012 470582 320058
rect 470314 320006 470326 320012
rect 470378 320006 470390 320012
rect 470442 320006 470454 320012
rect 470506 320006 470518 320012
rect 470570 320006 470582 320012
rect 470634 320006 470646 320012
rect 470698 320006 470710 320012
rect 470762 320006 470774 320012
rect 470262 320000 470826 320006
rect 470262 307086 470826 307092
rect 470314 307080 470326 307086
rect 470378 307080 470390 307086
rect 470442 307080 470454 307086
rect 470506 307080 470518 307086
rect 470570 307080 470582 307086
rect 470634 307080 470646 307086
rect 470698 307080 470710 307086
rect 470762 307080 470774 307086
rect 470506 307034 470516 307080
rect 470572 307034 470582 307080
rect 470262 307024 470276 307034
rect 470332 307024 470356 307034
rect 470412 307024 470436 307034
rect 470492 307024 470516 307034
rect 470572 307024 470596 307034
rect 470652 307024 470676 307034
rect 470732 307024 470756 307034
rect 470812 307024 470826 307034
rect 470262 307022 470826 307024
rect 470314 307000 470326 307022
rect 470378 307000 470390 307022
rect 470442 307000 470454 307022
rect 470506 307000 470518 307022
rect 470570 307000 470582 307022
rect 470634 307000 470646 307022
rect 470698 307000 470710 307022
rect 470762 307000 470774 307022
rect 470506 306970 470516 307000
rect 470572 306970 470582 307000
rect 470262 306958 470276 306970
rect 470332 306958 470356 306970
rect 470412 306958 470436 306970
rect 470492 306958 470516 306970
rect 470572 306958 470596 306970
rect 470652 306958 470676 306970
rect 470732 306958 470756 306970
rect 470812 306958 470826 306970
rect 470506 306944 470516 306958
rect 470572 306944 470582 306958
rect 470314 306920 470326 306944
rect 470378 306920 470390 306944
rect 470442 306920 470454 306944
rect 470506 306920 470518 306944
rect 470570 306920 470582 306944
rect 470634 306920 470646 306944
rect 470698 306920 470710 306944
rect 470762 306920 470774 306944
rect 470506 306906 470516 306920
rect 470572 306906 470582 306920
rect 470262 306894 470276 306906
rect 470332 306894 470356 306906
rect 470412 306894 470436 306906
rect 470492 306894 470516 306906
rect 470572 306894 470596 306906
rect 470652 306894 470676 306906
rect 470732 306894 470756 306906
rect 470812 306894 470826 306906
rect 470506 306864 470516 306894
rect 470572 306864 470582 306894
rect 470314 306842 470326 306864
rect 470378 306842 470390 306864
rect 470442 306842 470454 306864
rect 470506 306842 470518 306864
rect 470570 306842 470582 306864
rect 470634 306842 470646 306864
rect 470698 306842 470710 306864
rect 470762 306842 470774 306864
rect 470262 306840 470826 306842
rect 470262 306830 470276 306840
rect 470332 306830 470356 306840
rect 470412 306830 470436 306840
rect 470492 306830 470516 306840
rect 470572 306830 470596 306840
rect 470652 306830 470676 306840
rect 470732 306830 470756 306840
rect 470812 306830 470826 306840
rect 470506 306784 470516 306830
rect 470572 306784 470582 306830
rect 470314 306778 470326 306784
rect 470378 306778 470390 306784
rect 470442 306778 470454 306784
rect 470506 306778 470518 306784
rect 470570 306778 470582 306784
rect 470634 306778 470646 306784
rect 470698 306778 470710 306784
rect 470762 306778 470774 306784
rect 470262 306772 470826 306778
rect 471256 306338 471284 321574
rect 474278 321328 474334 321337
rect 484582 321328 484638 321337
rect 474334 321286 474680 321314
rect 474278 321263 474334 321272
rect 484638 321286 485012 321314
rect 484582 321263 484638 321272
rect 488170 321056 488226 321065
rect 478125 321014 478184 321042
rect 478156 320929 478184 321014
rect 481560 320929 481588 321042
rect 488226 321014 488456 321042
rect 488170 320991 488226 321000
rect 478142 320920 478198 320929
rect 478142 320855 478198 320864
rect 481546 320920 481602 320929
rect 481546 320855 481602 320864
rect 475476 320487 475528 320493
rect 475476 320429 475528 320435
rect 482376 320476 482428 320482
rect 475488 318782 475516 320429
rect 482376 320418 482428 320424
rect 479064 320408 479116 320414
rect 479064 320350 479116 320356
rect 479076 318782 479104 320350
rect 475476 318776 475528 318782
rect 475476 318718 475528 318724
rect 479064 318776 479116 318782
rect 479064 318718 479116 318724
rect 482388 318714 482416 320418
rect 485964 320408 486016 320414
rect 485964 320350 486016 320356
rect 482376 318708 482428 318714
rect 482376 318650 482428 318656
rect 485976 318646 486004 320350
rect 485964 318640 486016 318646
rect 485964 318582 486016 318588
rect 471244 306332 471296 306338
rect 471244 306274 471296 306280
rect 473728 306284 473780 306290
rect 469022 306001 469586 306007
rect 469074 305995 469086 306001
rect 469138 305995 469150 306001
rect 469202 305995 469214 306001
rect 469266 305995 469278 306001
rect 469330 305995 469342 306001
rect 469394 305995 469406 306001
rect 469458 305995 469470 306001
rect 469522 305995 469534 306001
rect 469266 305949 469276 305995
rect 469332 305949 469342 305995
rect 469022 305939 469036 305949
rect 469092 305939 469116 305949
rect 469172 305939 469196 305949
rect 469252 305939 469276 305949
rect 469332 305939 469356 305949
rect 469412 305939 469436 305949
rect 469492 305939 469516 305949
rect 469572 305939 469586 305949
rect 469022 305937 469586 305939
rect 469074 305915 469086 305937
rect 469138 305915 469150 305937
rect 469202 305915 469214 305937
rect 469266 305915 469278 305937
rect 469330 305915 469342 305937
rect 469394 305915 469406 305937
rect 469458 305915 469470 305937
rect 469522 305915 469534 305937
rect 469266 305885 469276 305915
rect 469332 305885 469342 305915
rect 469022 305873 469036 305885
rect 469092 305873 469116 305885
rect 469172 305873 469196 305885
rect 469252 305873 469276 305885
rect 469332 305873 469356 305885
rect 469412 305873 469436 305885
rect 469492 305873 469516 305885
rect 469572 305873 469586 305885
rect 469266 305859 469276 305873
rect 469332 305859 469342 305873
rect 469074 305835 469086 305859
rect 469138 305835 469150 305859
rect 469202 305835 469214 305859
rect 469266 305835 469278 305859
rect 469330 305835 469342 305859
rect 469394 305835 469406 305859
rect 469458 305835 469470 305859
rect 469522 305835 469534 305859
rect 469266 305821 469276 305835
rect 469332 305821 469342 305835
rect 469022 305809 469036 305821
rect 469092 305809 469116 305821
rect 469172 305809 469196 305821
rect 469252 305809 469276 305821
rect 469332 305809 469356 305821
rect 469412 305809 469436 305821
rect 469492 305809 469516 305821
rect 469572 305809 469586 305821
rect 469266 305779 469276 305809
rect 469332 305779 469342 305809
rect 469074 305757 469086 305779
rect 469138 305757 469150 305779
rect 469202 305757 469214 305779
rect 469266 305757 469278 305779
rect 469330 305757 469342 305779
rect 469394 305757 469406 305779
rect 469458 305757 469470 305779
rect 469522 305757 469534 305779
rect 469022 305755 469586 305757
rect 469022 305745 469036 305755
rect 469092 305745 469116 305755
rect 469172 305745 469196 305755
rect 469252 305745 469276 305755
rect 469332 305745 469356 305755
rect 469412 305745 469436 305755
rect 469492 305745 469516 305755
rect 469572 305745 469586 305755
rect 469266 305699 469276 305745
rect 469332 305699 469342 305745
rect 469074 305693 469086 305699
rect 469138 305693 469150 305699
rect 469202 305693 469214 305699
rect 469266 305693 469278 305699
rect 469330 305693 469342 305699
rect 469394 305693 469406 305699
rect 469458 305693 469470 305699
rect 469522 305693 469534 305699
rect 469022 305687 469586 305693
rect 470262 304914 470826 304920
rect 470314 304908 470326 304914
rect 470378 304908 470390 304914
rect 470442 304908 470454 304914
rect 470506 304908 470518 304914
rect 470570 304908 470582 304914
rect 470634 304908 470646 304914
rect 470698 304908 470710 304914
rect 470762 304908 470774 304914
rect 470506 304862 470516 304908
rect 470572 304862 470582 304908
rect 470262 304852 470276 304862
rect 470332 304852 470356 304862
rect 470412 304852 470436 304862
rect 470492 304852 470516 304862
rect 470572 304852 470596 304862
rect 470652 304852 470676 304862
rect 470732 304852 470756 304862
rect 470812 304852 470826 304862
rect 470262 304850 470826 304852
rect 470314 304828 470326 304850
rect 470378 304828 470390 304850
rect 470442 304828 470454 304850
rect 470506 304828 470518 304850
rect 470570 304828 470582 304850
rect 470634 304828 470646 304850
rect 470698 304828 470710 304850
rect 470762 304828 470774 304850
rect 470506 304798 470516 304828
rect 470572 304798 470582 304828
rect 470262 304786 470276 304798
rect 470332 304786 470356 304798
rect 470412 304786 470436 304798
rect 470492 304786 470516 304798
rect 470572 304786 470596 304798
rect 470652 304786 470676 304798
rect 470732 304786 470756 304798
rect 470812 304786 470826 304798
rect 470506 304772 470516 304786
rect 470572 304772 470582 304786
rect 470314 304748 470326 304772
rect 470378 304748 470390 304772
rect 470442 304748 470454 304772
rect 470506 304748 470518 304772
rect 470570 304748 470582 304772
rect 470634 304748 470646 304772
rect 470698 304748 470710 304772
rect 470762 304748 470774 304772
rect 470506 304734 470516 304748
rect 470572 304734 470582 304748
rect 470262 304722 470276 304734
rect 470332 304722 470356 304734
rect 470412 304722 470436 304734
rect 470492 304722 470516 304734
rect 470572 304722 470596 304734
rect 470652 304722 470676 304734
rect 470732 304722 470756 304734
rect 470812 304722 470826 304734
rect 470506 304692 470516 304722
rect 470572 304692 470582 304722
rect 470314 304670 470326 304692
rect 470378 304670 470390 304692
rect 470442 304670 470454 304692
rect 470506 304670 470518 304692
rect 470570 304670 470582 304692
rect 470634 304670 470646 304692
rect 470698 304670 470710 304692
rect 470762 304670 470774 304692
rect 470262 304668 470826 304670
rect 470262 304658 470276 304668
rect 470332 304658 470356 304668
rect 470412 304658 470436 304668
rect 470492 304658 470516 304668
rect 470572 304658 470596 304668
rect 470652 304658 470676 304668
rect 470732 304658 470756 304668
rect 470812 304658 470826 304668
rect 470506 304612 470516 304658
rect 470572 304612 470582 304658
rect 470314 304606 470326 304612
rect 470378 304606 470390 304612
rect 470442 304606 470454 304612
rect 470506 304606 470518 304612
rect 470570 304606 470582 304612
rect 470634 304606 470646 304612
rect 470698 304606 470710 304612
rect 470762 304606 470774 304612
rect 470262 304600 470826 304606
rect 470262 287487 470826 287493
rect 470314 287481 470326 287487
rect 470378 287481 470390 287487
rect 470442 287481 470454 287487
rect 470506 287481 470518 287487
rect 470570 287481 470582 287487
rect 470634 287481 470646 287487
rect 470698 287481 470710 287487
rect 470762 287481 470774 287487
rect 470506 287435 470516 287481
rect 470572 287435 470582 287481
rect 470262 287425 470276 287435
rect 470332 287425 470356 287435
rect 470412 287425 470436 287435
rect 470492 287425 470516 287435
rect 470572 287425 470596 287435
rect 470652 287425 470676 287435
rect 470732 287425 470756 287435
rect 470812 287425 470826 287435
rect 470262 287423 470826 287425
rect 470314 287401 470326 287423
rect 470378 287401 470390 287423
rect 470442 287401 470454 287423
rect 470506 287401 470518 287423
rect 470570 287401 470582 287423
rect 470634 287401 470646 287423
rect 470698 287401 470710 287423
rect 470762 287401 470774 287423
rect 470506 287371 470516 287401
rect 470572 287371 470582 287401
rect 470262 287359 470276 287371
rect 470332 287359 470356 287371
rect 470412 287359 470436 287371
rect 470492 287359 470516 287371
rect 470572 287359 470596 287371
rect 470652 287359 470676 287371
rect 470732 287359 470756 287371
rect 470812 287359 470826 287371
rect 470506 287345 470516 287359
rect 470572 287345 470582 287359
rect 470314 287321 470326 287345
rect 470378 287321 470390 287345
rect 470442 287321 470454 287345
rect 470506 287321 470518 287345
rect 470570 287321 470582 287345
rect 470634 287321 470646 287345
rect 470698 287321 470710 287345
rect 470762 287321 470774 287345
rect 470506 287307 470516 287321
rect 470572 287307 470582 287321
rect 470262 287295 470276 287307
rect 470332 287295 470356 287307
rect 470412 287295 470436 287307
rect 470492 287295 470516 287307
rect 470572 287295 470596 287307
rect 470652 287295 470676 287307
rect 470732 287295 470756 287307
rect 470812 287295 470826 287307
rect 470506 287265 470516 287295
rect 470572 287265 470582 287295
rect 470314 287243 470326 287265
rect 470378 287243 470390 287265
rect 470442 287243 470454 287265
rect 470506 287243 470518 287265
rect 470570 287243 470582 287265
rect 470634 287243 470646 287265
rect 470698 287243 470710 287265
rect 470762 287243 470774 287265
rect 470262 287241 470826 287243
rect 470262 287231 470276 287241
rect 470332 287231 470356 287241
rect 470412 287231 470436 287241
rect 470492 287231 470516 287241
rect 470572 287231 470596 287241
rect 470652 287231 470676 287241
rect 470732 287231 470756 287241
rect 470812 287231 470826 287241
rect 470506 287185 470516 287231
rect 470572 287185 470582 287231
rect 470314 287179 470326 287185
rect 470378 287179 470390 287185
rect 470442 287179 470454 287185
rect 470506 287179 470518 287185
rect 470570 287179 470582 287185
rect 470634 287179 470646 287185
rect 470698 287179 470710 287185
rect 470762 287179 470774 287185
rect 470262 287173 470826 287179
rect 471256 286686 471284 306274
rect 473728 306226 473780 306232
rect 473740 305969 473768 306226
rect 487525 306176 487534 306232
rect 487590 306176 487599 306232
rect 481004 306096 481060 306105
rect 481004 306031 481060 306040
rect 473726 305960 473782 305969
rect 473726 305895 473782 305904
rect 477739 305688 477795 305697
rect 477739 305623 477795 305632
rect 484122 305552 484178 305561
rect 484178 305510 484297 305538
rect 484122 305487 484178 305496
rect 478604 305448 478656 305454
rect 478604 305390 478656 305396
rect 485136 305448 485188 305454
rect 485136 305390 485188 305396
rect 475292 305088 475344 305094
rect 475292 305030 475344 305036
rect 475304 303618 475332 305030
rect 478616 303618 478644 305390
rect 481824 305088 481876 305094
rect 481824 305030 481876 305036
rect 481836 303618 481864 305030
rect 485148 303618 485176 305390
rect 490564 305040 490616 305046
rect 490564 304982 490616 304988
rect 475292 303612 475344 303618
rect 475292 303554 475344 303560
rect 478604 303612 478656 303618
rect 478604 303554 478656 303560
rect 481824 303612 481876 303618
rect 481824 303554 481876 303560
rect 485136 303612 485188 303618
rect 485136 303554 485188 303560
rect 490576 292534 490604 304982
rect 490760 298110 490788 409974
rect 491956 300830 491984 449346
rect 515404 445936 515456 445942
rect 515404 445878 515456 445884
rect 493324 441652 493376 441658
rect 493324 441594 493376 441600
rect 492036 431044 492088 431050
rect 492036 430986 492088 430992
rect 491944 300824 491996 300830
rect 491944 300766 491996 300772
rect 492048 299470 492076 430986
rect 493336 408474 493364 441594
rect 494704 440292 494756 440298
rect 494704 440234 494756 440240
rect 493324 408468 493376 408474
rect 493324 408410 493376 408416
rect 493324 389496 493376 389502
rect 493324 389438 493376 389444
rect 492128 356448 492180 356454
rect 492128 356390 492180 356396
rect 492036 299464 492088 299470
rect 492036 299406 492088 299412
rect 490748 298104 490800 298110
rect 490748 298046 490800 298052
rect 492140 296682 492168 356390
rect 492220 340400 492272 340406
rect 492220 340342 492272 340348
rect 492128 296676 492180 296682
rect 492128 296618 492180 296624
rect 492232 295322 492260 340342
rect 492312 320408 492364 320414
rect 492312 320350 492364 320356
rect 492220 295316 492272 295322
rect 492220 295258 492272 295264
rect 492324 293962 492352 320350
rect 493336 296614 493364 389438
rect 494716 387734 494744 440234
rect 496084 438932 496136 438938
rect 496084 438874 496136 438880
rect 494704 387728 494756 387734
rect 494704 387670 494756 387676
rect 496096 354550 496124 438874
rect 497464 437504 497516 437510
rect 497464 437446 497516 437452
rect 496084 354544 496136 354550
rect 496084 354486 496136 354492
rect 497476 339318 497504 437446
rect 498844 436144 498896 436150
rect 498844 436086 498896 436092
rect 497464 339312 497516 339318
rect 497464 339254 497516 339260
rect 498856 318578 498884 436086
rect 500224 434784 500276 434790
rect 500224 434726 500276 434732
rect 498844 318572 498896 318578
rect 498844 318514 498896 318520
rect 500236 303414 500264 434726
rect 501604 433356 501656 433362
rect 501604 433298 501656 433304
rect 500224 303408 500276 303414
rect 500224 303350 500276 303356
rect 493324 296608 493376 296614
rect 493324 296550 493376 296556
rect 492312 293956 492364 293962
rect 492312 293898 492364 293904
rect 490564 292528 490616 292534
rect 490564 292470 490616 292476
rect 492956 289876 493008 289882
rect 492956 289818 493008 289824
rect 491944 288448 491996 288454
rect 491944 288390 491996 288396
rect 478633 286920 478689 286929
rect 478633 286855 478689 286864
rect 471244 286680 471296 286686
rect 471244 286622 471296 286628
rect 474912 286592 474921 286648
rect 474977 286592 474986 286648
rect 478647 286620 478675 286855
rect 488632 286680 488684 286686
rect 488630 286648 488632 286657
rect 488684 286648 488686 286657
rect 488630 286583 488686 286592
rect 471704 286544 471756 286550
rect 471704 286486 471756 286492
rect 469022 286402 469586 286408
rect 469074 286396 469086 286402
rect 469138 286396 469150 286402
rect 469202 286396 469214 286402
rect 469266 286396 469278 286402
rect 469330 286396 469342 286402
rect 469394 286396 469406 286402
rect 469458 286396 469470 286402
rect 469522 286396 469534 286402
rect 469266 286350 469276 286396
rect 469332 286350 469342 286396
rect 469022 286340 469036 286350
rect 469092 286340 469116 286350
rect 469172 286340 469196 286350
rect 469252 286340 469276 286350
rect 469332 286340 469356 286350
rect 469412 286340 469436 286350
rect 469492 286340 469516 286350
rect 469572 286340 469586 286350
rect 469022 286338 469586 286340
rect 469074 286316 469086 286338
rect 469138 286316 469150 286338
rect 469202 286316 469214 286338
rect 469266 286316 469278 286338
rect 469330 286316 469342 286338
rect 469394 286316 469406 286338
rect 469458 286316 469470 286338
rect 469522 286316 469534 286338
rect 469266 286286 469276 286316
rect 469332 286286 469342 286316
rect 469022 286274 469036 286286
rect 469092 286274 469116 286286
rect 469172 286274 469196 286286
rect 469252 286274 469276 286286
rect 469332 286274 469356 286286
rect 469412 286274 469436 286286
rect 469492 286274 469516 286286
rect 469572 286274 469586 286286
rect 469266 286260 469276 286274
rect 469332 286260 469342 286274
rect 469074 286236 469086 286260
rect 469138 286236 469150 286260
rect 469202 286236 469214 286260
rect 469266 286236 469278 286260
rect 469330 286236 469342 286260
rect 469394 286236 469406 286260
rect 469458 286236 469470 286260
rect 469522 286236 469534 286260
rect 469266 286222 469276 286236
rect 469332 286222 469342 286236
rect 469022 286210 469036 286222
rect 469092 286210 469116 286222
rect 469172 286210 469196 286222
rect 469252 286210 469276 286222
rect 469332 286210 469356 286222
rect 469412 286210 469436 286222
rect 469492 286210 469516 286222
rect 469572 286210 469586 286222
rect 469266 286180 469276 286210
rect 469332 286180 469342 286210
rect 469074 286158 469086 286180
rect 469138 286158 469150 286180
rect 469202 286158 469214 286180
rect 469266 286158 469278 286180
rect 469330 286158 469342 286180
rect 469394 286158 469406 286180
rect 469458 286158 469470 286180
rect 469522 286158 469534 286180
rect 469022 286156 469586 286158
rect 469022 286146 469036 286156
rect 469092 286146 469116 286156
rect 469172 286146 469196 286156
rect 469252 286146 469276 286156
rect 469332 286146 469356 286156
rect 469412 286146 469436 286156
rect 469492 286146 469516 286156
rect 469572 286146 469586 286156
rect 469266 286100 469276 286146
rect 469332 286100 469342 286146
rect 469074 286094 469086 286100
rect 469138 286094 469150 286100
rect 469202 286094 469214 286100
rect 469266 286094 469278 286100
rect 469330 286094 469342 286100
rect 469394 286094 469406 286100
rect 469458 286094 469470 286100
rect 469522 286094 469534 286100
rect 469022 286088 469586 286094
rect 470262 285314 470826 285320
rect 470314 285308 470326 285314
rect 470378 285308 470390 285314
rect 470442 285308 470454 285314
rect 470506 285308 470518 285314
rect 470570 285308 470582 285314
rect 470634 285308 470646 285314
rect 470698 285308 470710 285314
rect 470762 285308 470774 285314
rect 470506 285262 470516 285308
rect 470572 285262 470582 285308
rect 470262 285252 470276 285262
rect 470332 285252 470356 285262
rect 470412 285252 470436 285262
rect 470492 285252 470516 285262
rect 470572 285252 470596 285262
rect 470652 285252 470676 285262
rect 470732 285252 470756 285262
rect 470812 285252 470826 285262
rect 470262 285250 470826 285252
rect 470314 285228 470326 285250
rect 470378 285228 470390 285250
rect 470442 285228 470454 285250
rect 470506 285228 470518 285250
rect 470570 285228 470582 285250
rect 470634 285228 470646 285250
rect 470698 285228 470710 285250
rect 470762 285228 470774 285250
rect 470506 285198 470516 285228
rect 470572 285198 470582 285228
rect 470262 285186 470276 285198
rect 470332 285186 470356 285198
rect 470412 285186 470436 285198
rect 470492 285186 470516 285198
rect 470572 285186 470596 285198
rect 470652 285186 470676 285198
rect 470732 285186 470756 285198
rect 470812 285186 470826 285198
rect 470506 285172 470516 285186
rect 470572 285172 470582 285186
rect 470314 285148 470326 285172
rect 470378 285148 470390 285172
rect 470442 285148 470454 285172
rect 470506 285148 470518 285172
rect 470570 285148 470582 285172
rect 470634 285148 470646 285172
rect 470698 285148 470710 285172
rect 470762 285148 470774 285172
rect 470506 285134 470516 285148
rect 470572 285134 470582 285148
rect 470262 285122 470276 285134
rect 470332 285122 470356 285134
rect 470412 285122 470436 285134
rect 470492 285122 470516 285134
rect 470572 285122 470596 285134
rect 470652 285122 470676 285134
rect 470732 285122 470756 285134
rect 470812 285122 470826 285134
rect 470506 285092 470516 285122
rect 470572 285092 470582 285122
rect 470314 285070 470326 285092
rect 470378 285070 470390 285092
rect 470442 285070 470454 285092
rect 470506 285070 470518 285092
rect 470570 285070 470582 285092
rect 470634 285070 470646 285092
rect 470698 285070 470710 285092
rect 470762 285070 470774 285092
rect 470262 285068 470826 285070
rect 470262 285058 470276 285068
rect 470332 285058 470356 285068
rect 470412 285058 470436 285068
rect 470492 285058 470516 285068
rect 470572 285058 470596 285068
rect 470652 285058 470676 285068
rect 470732 285058 470756 285068
rect 470812 285058 470826 285068
rect 470506 285012 470516 285058
rect 470572 285012 470582 285058
rect 470314 285006 470326 285012
rect 470378 285006 470390 285012
rect 470442 285006 470454 285012
rect 470506 285006 470518 285012
rect 470570 285006 470582 285012
rect 470634 285006 470646 285012
rect 470698 285006 470710 285012
rect 470762 285006 470774 285012
rect 470262 285000 470826 285006
rect 471716 270502 471744 286486
rect 479432 285864 479484 285870
rect 485870 285832 485926 285841
rect 479432 285806 479484 285812
rect 475752 285488 475804 285494
rect 475752 285430 475804 285436
rect 475764 284306 475792 285430
rect 479444 284306 479472 285806
rect 482336 285776 482345 285832
rect 482401 285776 482410 285832
rect 485926 285790 486085 285818
rect 485870 285767 485926 285776
rect 483204 285488 483256 285494
rect 483204 285430 483256 285436
rect 486884 285488 486936 285494
rect 486884 285430 486936 285436
rect 475752 284300 475804 284306
rect 475752 284242 475804 284248
rect 479432 284300 479484 284306
rect 479432 284242 479484 284248
rect 483216 284238 483244 285430
rect 483204 284232 483256 284238
rect 483204 284174 483256 284180
rect 486896 284170 486924 285430
rect 486884 284164 486936 284170
rect 486884 284106 486936 284112
rect 471704 270496 471756 270502
rect 471704 270438 471756 270444
rect 473728 270496 473780 270502
rect 473728 270438 473780 270444
rect 470262 267487 470826 267493
rect 470314 267481 470326 267487
rect 470378 267481 470390 267487
rect 470442 267481 470454 267487
rect 470506 267481 470518 267487
rect 470570 267481 470582 267487
rect 470634 267481 470646 267487
rect 470698 267481 470710 267487
rect 470762 267481 470774 267487
rect 470506 267435 470516 267481
rect 470572 267435 470582 267481
rect 470262 267425 470276 267435
rect 470332 267425 470356 267435
rect 470412 267425 470436 267435
rect 470492 267425 470516 267435
rect 470572 267425 470596 267435
rect 470652 267425 470676 267435
rect 470732 267425 470756 267435
rect 470812 267425 470826 267435
rect 470262 267423 470826 267425
rect 470314 267401 470326 267423
rect 470378 267401 470390 267423
rect 470442 267401 470454 267423
rect 470506 267401 470518 267423
rect 470570 267401 470582 267423
rect 470634 267401 470646 267423
rect 470698 267401 470710 267423
rect 470762 267401 470774 267423
rect 470506 267371 470516 267401
rect 470572 267371 470582 267401
rect 470262 267359 470276 267371
rect 470332 267359 470356 267371
rect 470412 267359 470436 267371
rect 470492 267359 470516 267371
rect 470572 267359 470596 267371
rect 470652 267359 470676 267371
rect 470732 267359 470756 267371
rect 470812 267359 470826 267371
rect 470506 267345 470516 267359
rect 470572 267345 470582 267359
rect 470314 267321 470326 267345
rect 470378 267321 470390 267345
rect 470442 267321 470454 267345
rect 470506 267321 470518 267345
rect 470570 267321 470582 267345
rect 470634 267321 470646 267345
rect 470698 267321 470710 267345
rect 470762 267321 470774 267345
rect 470506 267307 470516 267321
rect 470572 267307 470582 267321
rect 470262 267295 470276 267307
rect 470332 267295 470356 267307
rect 470412 267295 470436 267307
rect 470492 267295 470516 267307
rect 470572 267295 470596 267307
rect 470652 267295 470676 267307
rect 470732 267295 470756 267307
rect 470812 267295 470826 267307
rect 470506 267265 470516 267295
rect 470572 267265 470582 267295
rect 470314 267243 470326 267265
rect 470378 267243 470390 267265
rect 470442 267243 470454 267265
rect 470506 267243 470518 267265
rect 470570 267243 470582 267265
rect 470634 267243 470646 267265
rect 470698 267243 470710 267265
rect 470762 267243 470774 267265
rect 470262 267241 470826 267243
rect 470262 267231 470276 267241
rect 470332 267231 470356 267241
rect 470412 267231 470436 267241
rect 470492 267231 470516 267241
rect 470572 267231 470596 267241
rect 470652 267231 470676 267241
rect 470732 267231 470756 267241
rect 470812 267231 470826 267241
rect 470506 267185 470516 267231
rect 470572 267185 470582 267231
rect 470314 267179 470326 267185
rect 470378 267179 470390 267185
rect 470442 267179 470454 267185
rect 470506 267179 470518 267185
rect 470570 267179 470582 267185
rect 470634 267179 470646 267185
rect 470698 267179 470710 267185
rect 470762 267179 470774 267185
rect 470262 267173 470826 267179
rect 473740 266558 473768 270438
rect 473728 266552 473780 266558
rect 473728 266494 473780 266500
rect 469022 266401 469586 266407
rect 469074 266395 469086 266401
rect 469138 266395 469150 266401
rect 469202 266395 469214 266401
rect 469266 266395 469278 266401
rect 469330 266395 469342 266401
rect 469394 266395 469406 266401
rect 469458 266395 469470 266401
rect 469522 266395 469534 266401
rect 469266 266349 469276 266395
rect 469332 266349 469342 266395
rect 469022 266339 469036 266349
rect 469092 266339 469116 266349
rect 469172 266339 469196 266349
rect 469252 266339 469276 266349
rect 469332 266339 469356 266349
rect 469412 266339 469436 266349
rect 469492 266339 469516 266349
rect 469572 266339 469586 266349
rect 469022 266337 469586 266339
rect 469074 266315 469086 266337
rect 469138 266315 469150 266337
rect 469202 266315 469214 266337
rect 469266 266315 469278 266337
rect 469330 266315 469342 266337
rect 469394 266315 469406 266337
rect 469458 266315 469470 266337
rect 469522 266315 469534 266337
rect 469266 266285 469276 266315
rect 469332 266285 469342 266315
rect 469022 266273 469036 266285
rect 469092 266273 469116 266285
rect 469172 266273 469196 266285
rect 469252 266273 469276 266285
rect 469332 266273 469356 266285
rect 469412 266273 469436 266285
rect 469492 266273 469516 266285
rect 469572 266273 469586 266285
rect 469266 266259 469276 266273
rect 469332 266259 469342 266273
rect 469074 266235 469086 266259
rect 469138 266235 469150 266259
rect 469202 266235 469214 266259
rect 469266 266235 469278 266259
rect 469330 266235 469342 266259
rect 469394 266235 469406 266259
rect 469458 266235 469470 266259
rect 469522 266235 469534 266259
rect 469266 266221 469276 266235
rect 469332 266221 469342 266235
rect 469022 266209 469036 266221
rect 469092 266209 469116 266221
rect 469172 266209 469196 266221
rect 469252 266209 469276 266221
rect 469332 266209 469356 266221
rect 469412 266209 469436 266221
rect 469492 266209 469516 266221
rect 469572 266209 469586 266221
rect 469266 266179 469276 266209
rect 469332 266179 469342 266209
rect 469074 266157 469086 266179
rect 469138 266157 469150 266179
rect 469202 266157 469214 266179
rect 469266 266157 469278 266179
rect 469330 266157 469342 266179
rect 469394 266157 469406 266179
rect 469458 266157 469470 266179
rect 469522 266157 469534 266179
rect 469022 266155 469586 266157
rect 469022 266145 469036 266155
rect 469092 266145 469116 266155
rect 469172 266145 469196 266155
rect 469252 266145 469276 266155
rect 469332 266145 469356 266155
rect 469412 266145 469436 266155
rect 469492 266145 469516 266155
rect 469572 266145 469586 266155
rect 469266 266099 469276 266145
rect 469332 266099 469342 266145
rect 469074 266093 469086 266099
rect 469138 266093 469150 266099
rect 469202 266093 469214 266099
rect 469266 266093 469278 266099
rect 469330 266093 469342 266099
rect 469394 266093 469406 266099
rect 469458 266093 469470 266099
rect 469522 266093 469534 266099
rect 469022 266087 469586 266093
rect 470262 265314 470826 265320
rect 470314 265308 470326 265314
rect 470378 265308 470390 265314
rect 470442 265308 470454 265314
rect 470506 265308 470518 265314
rect 470570 265308 470582 265314
rect 470634 265308 470646 265314
rect 470698 265308 470710 265314
rect 470762 265308 470774 265314
rect 470506 265262 470516 265308
rect 470572 265262 470582 265308
rect 470262 265252 470276 265262
rect 470332 265252 470356 265262
rect 470412 265252 470436 265262
rect 470492 265252 470516 265262
rect 470572 265252 470596 265262
rect 470652 265252 470676 265262
rect 470732 265252 470756 265262
rect 470812 265252 470826 265262
rect 470262 265250 470826 265252
rect 470314 265228 470326 265250
rect 470378 265228 470390 265250
rect 470442 265228 470454 265250
rect 470506 265228 470518 265250
rect 470570 265228 470582 265250
rect 470634 265228 470646 265250
rect 470698 265228 470710 265250
rect 470762 265228 470774 265250
rect 470506 265198 470516 265228
rect 470572 265198 470582 265228
rect 470262 265186 470276 265198
rect 470332 265186 470356 265198
rect 470412 265186 470436 265198
rect 470492 265186 470516 265198
rect 470572 265186 470596 265198
rect 470652 265186 470676 265198
rect 470732 265186 470756 265198
rect 470812 265186 470826 265198
rect 470506 265172 470516 265186
rect 470572 265172 470582 265186
rect 470314 265148 470326 265172
rect 470378 265148 470390 265172
rect 470442 265148 470454 265172
rect 470506 265148 470518 265172
rect 470570 265148 470582 265172
rect 470634 265148 470646 265172
rect 470698 265148 470710 265172
rect 470762 265148 470774 265172
rect 470506 265134 470516 265148
rect 470572 265134 470582 265148
rect 470262 265122 470276 265134
rect 470332 265122 470356 265134
rect 470412 265122 470436 265134
rect 470492 265122 470516 265134
rect 470572 265122 470596 265134
rect 470652 265122 470676 265134
rect 470732 265122 470756 265134
rect 470812 265122 470826 265134
rect 470506 265092 470516 265122
rect 470572 265092 470582 265122
rect 470314 265070 470326 265092
rect 470378 265070 470390 265092
rect 470442 265070 470454 265092
rect 470506 265070 470518 265092
rect 470570 265070 470582 265092
rect 470634 265070 470646 265092
rect 470698 265070 470710 265092
rect 470762 265070 470774 265092
rect 470262 265068 470826 265070
rect 470262 265058 470276 265068
rect 470332 265058 470356 265068
rect 470412 265058 470436 265068
rect 470492 265058 470516 265068
rect 470572 265058 470596 265068
rect 470652 265058 470676 265068
rect 470732 265058 470756 265068
rect 470812 265058 470826 265068
rect 470506 265012 470516 265058
rect 470572 265012 470582 265058
rect 470314 265006 470326 265012
rect 470378 265006 470390 265012
rect 470442 265006 470454 265012
rect 470506 265006 470518 265012
rect 470570 265006 470582 265012
rect 470634 265006 470646 265012
rect 470698 265006 470710 265012
rect 470762 265006 470774 265012
rect 470262 265000 470826 265006
rect 473740 206990 473768 266494
rect 491956 266014 491984 288390
rect 492968 285666 492996 289818
rect 492956 285660 493008 285666
rect 492956 285602 493008 285608
rect 501616 284102 501644 433298
rect 502984 431996 503036 432002
rect 502984 431938 503036 431944
rect 501604 284096 501656 284102
rect 501604 284038 501656 284044
rect 491944 266008 491996 266014
rect 479062 265976 479118 265985
rect 479118 265948 479341 265962
rect 491944 265950 491996 265956
rect 479118 265934 479355 265948
rect 479062 265911 479118 265920
rect 477132 265872 477184 265878
rect 477132 265814 477184 265820
rect 476275 265690 476303 265812
rect 476275 265662 476344 265690
rect 476316 265010 476344 265662
rect 476486 265024 476542 265033
rect 476316 264982 476486 265010
rect 476486 264959 476542 264968
rect 477144 263566 477172 265814
rect 479327 265690 479355 265934
rect 482379 265690 482407 265812
rect 485431 265690 485459 265812
rect 479327 265662 479380 265690
rect 482379 265662 482416 265690
rect 485431 265662 485728 265690
rect 479352 265010 479380 265662
rect 480168 265487 480220 265493
rect 480168 265429 480220 265435
rect 479522 265024 479578 265033
rect 479352 264982 479522 265010
rect 479522 264959 479578 264968
rect 480180 263566 480208 265429
rect 482388 265010 482416 265662
rect 483204 265487 483256 265493
rect 483204 265429 483256 265435
rect 482834 265024 482890 265033
rect 482388 264982 482834 265010
rect 482834 264959 482890 264968
rect 483216 263566 483244 265429
rect 485700 265033 485728 265662
rect 488483 265554 488511 265812
rect 488722 265568 488778 265577
rect 488483 265526 488722 265554
rect 488722 265503 488778 265512
rect 486240 265487 486292 265493
rect 486240 265429 486292 265435
rect 485686 265024 485742 265033
rect 485686 264959 485742 264968
rect 486252 263566 486280 265429
rect 477132 263560 477184 263566
rect 477132 263502 477184 263508
rect 480168 263560 480220 263566
rect 480168 263502 480220 263508
rect 483204 263560 483256 263566
rect 483204 263502 483256 263508
rect 486240 263560 486292 263566
rect 495072 263560 495124 263566
rect 486240 263502 486292 263508
rect 494808 263508 495072 263514
rect 494808 263502 495124 263508
rect 494808 263498 495112 263502
rect 494796 263492 495112 263498
rect 494848 263486 495112 263492
rect 494796 263434 494848 263440
rect 502996 263362 503024 431938
rect 515416 409834 515444 445878
rect 523684 445868 523736 445874
rect 523684 445810 523736 445816
rect 520924 445800 520976 445806
rect 520924 445742 520976 445748
rect 515404 409828 515456 409834
rect 515404 409770 515456 409776
rect 515404 404388 515456 404394
rect 515404 404330 515456 404336
rect 515416 387802 515444 404330
rect 516784 403028 516836 403034
rect 516784 402970 516836 402976
rect 515404 387796 515456 387802
rect 515404 387738 515456 387744
rect 515404 365764 515456 365770
rect 515404 365706 515456 365712
rect 515416 339386 515444 365706
rect 516796 354686 516824 402970
rect 518164 398880 518216 398886
rect 518164 398822 518216 398828
rect 516784 354680 516836 354686
rect 516784 354622 516836 354628
rect 515404 339380 515456 339386
rect 515404 339322 515456 339328
rect 518176 303482 518204 398822
rect 519544 396092 519596 396098
rect 519544 396034 519596 396040
rect 518164 303476 518216 303482
rect 518164 303418 518216 303424
rect 519556 263430 519584 396034
rect 520936 373998 520964 445742
rect 522304 427848 522356 427854
rect 522304 427790 522356 427796
rect 520924 373992 520976 373998
rect 520924 373934 520976 373940
rect 522316 372570 522344 427790
rect 522304 372564 522356 372570
rect 522304 372506 522356 372512
rect 520924 367124 520976 367130
rect 520924 367066 520976 367072
rect 520936 354618 520964 367066
rect 522304 361616 522356 361622
rect 522304 361558 522356 361564
rect 520924 354612 520976 354618
rect 520924 354554 520976 354560
rect 522316 284238 522344 361558
rect 523696 338094 523724 445810
rect 535460 445732 535512 445738
rect 535460 445674 535512 445680
rect 535472 444825 535500 445674
rect 538692 445182 539258 445210
rect 546710 445182 547368 445210
rect 535458 444816 535514 444825
rect 535458 444751 535514 444760
rect 535458 443456 535514 443465
rect 535458 443391 535514 443400
rect 535472 443018 535500 443391
rect 535460 443012 535512 443018
rect 535460 442954 535512 442960
rect 535458 442096 535514 442105
rect 535458 442031 535514 442040
rect 535472 441658 535500 442031
rect 535460 441652 535512 441658
rect 535460 441594 535512 441600
rect 535458 440736 535514 440745
rect 535458 440671 535514 440680
rect 535472 440298 535500 440671
rect 535460 440292 535512 440298
rect 535460 440234 535512 440240
rect 535458 439376 535514 439385
rect 535458 439311 535514 439320
rect 535472 438938 535500 439311
rect 535460 438932 535512 438938
rect 535460 438874 535512 438880
rect 535458 438016 535514 438025
rect 535458 437951 535514 437960
rect 535472 437510 535500 437951
rect 535460 437504 535512 437510
rect 535460 437446 535512 437452
rect 535458 436656 535514 436665
rect 535458 436591 535514 436600
rect 535472 436150 535500 436591
rect 535460 436144 535512 436150
rect 535460 436086 535512 436092
rect 535458 435296 535514 435305
rect 535458 435231 535514 435240
rect 535472 434790 535500 435231
rect 535460 434784 535512 434790
rect 535460 434726 535512 434732
rect 535458 433936 535514 433945
rect 535458 433871 535514 433880
rect 535472 433362 535500 433871
rect 535460 433356 535512 433362
rect 535460 433298 535512 433304
rect 535458 432576 535514 432585
rect 535458 432511 535514 432520
rect 535472 432002 535500 432511
rect 535460 431996 535512 432002
rect 535460 431938 535512 431944
rect 536746 424416 536802 424425
rect 536746 424351 536802 424360
rect 535460 409828 535512 409834
rect 535460 409770 535512 409776
rect 535472 409329 535500 409770
rect 535458 409320 535514 409329
rect 535458 409255 535514 409264
rect 535460 407108 535512 407114
rect 535460 407050 535512 407056
rect 535472 406609 535500 407050
rect 535458 406600 535514 406609
rect 535458 406535 535514 406544
rect 535458 404560 535514 404569
rect 535458 404495 535514 404504
rect 535472 404394 535500 404495
rect 535460 404388 535512 404394
rect 535460 404330 535512 404336
rect 535458 403200 535514 403209
rect 535458 403135 535514 403144
rect 535472 403034 535500 403135
rect 535460 403028 535512 403034
rect 535460 402970 535512 402976
rect 536378 401704 536434 401713
rect 536378 401639 536434 401648
rect 536286 400344 536342 400353
rect 536286 400279 536342 400288
rect 535458 399120 535514 399129
rect 535458 399055 535514 399064
rect 535472 398886 535500 399055
rect 535460 398880 535512 398886
rect 535460 398822 535512 398828
rect 536102 397488 536158 397497
rect 536102 397423 536158 397432
rect 535458 396400 535514 396409
rect 535458 396335 535514 396344
rect 535472 396098 535500 396335
rect 535460 396092 535512 396098
rect 535460 396034 535512 396040
rect 535460 373992 535512 373998
rect 535460 373934 535512 373940
rect 535472 372881 535500 373934
rect 535458 372872 535514 372881
rect 535458 372807 535514 372816
rect 535460 372564 535512 372570
rect 535460 372506 535512 372512
rect 535472 371521 535500 372506
rect 535458 371512 535514 371521
rect 535458 371447 535514 371456
rect 535460 369844 535512 369850
rect 535460 369786 535512 369792
rect 535472 368801 535500 369786
rect 535458 368792 535514 368801
rect 535458 368727 535514 368736
rect 535458 367432 535514 367441
rect 535458 367367 535514 367376
rect 535472 367130 535500 367367
rect 535460 367124 535512 367130
rect 535460 367066 535512 367072
rect 535458 366072 535514 366081
rect 535458 366007 535514 366016
rect 535472 365770 535500 366007
rect 535460 365764 535512 365770
rect 535460 365706 535512 365712
rect 535458 361992 535514 362001
rect 535458 361927 535514 361936
rect 535472 361622 535500 361927
rect 535460 361616 535512 361622
rect 535460 361558 535512 361564
rect 535918 360632 535974 360641
rect 535918 360567 535974 360576
rect 525064 353320 525116 353326
rect 525064 353262 525116 353268
rect 523684 338088 523736 338094
rect 523684 338030 523736 338036
rect 525076 332586 525104 353262
rect 535460 338088 535512 338094
rect 535460 338030 535512 338036
rect 535472 336841 535500 338030
rect 535458 336832 535514 336841
rect 535458 336767 535514 336776
rect 525064 332580 525116 332586
rect 525064 332522 525116 332528
rect 535460 332580 535512 332586
rect 535460 332522 535512 332528
rect 535472 331401 535500 332522
rect 535458 331392 535514 331401
rect 535458 331327 535514 331336
rect 535460 331220 535512 331226
rect 535460 331162 535512 331168
rect 535472 330041 535500 331162
rect 535458 330032 535514 330041
rect 535458 329967 535514 329976
rect 535458 325952 535514 325961
rect 535458 325887 535514 325896
rect 535472 325718 535500 325887
rect 523684 325712 523736 325718
rect 523684 325654 523736 325660
rect 535460 325712 535512 325718
rect 535460 325654 535512 325660
rect 522304 284232 522356 284238
rect 522304 284174 522356 284180
rect 523696 284170 523724 325654
rect 535460 300824 535512 300830
rect 535458 300792 535460 300801
rect 535512 300792 535514 300801
rect 535458 300727 535514 300736
rect 535460 299464 535512 299470
rect 535458 299432 535460 299441
rect 535512 299432 535514 299441
rect 535458 299367 535514 299376
rect 535460 298104 535512 298110
rect 535458 298072 535460 298081
rect 535512 298072 535514 298081
rect 535458 298007 535514 298016
rect 535458 296712 535514 296721
rect 535458 296647 535514 296656
rect 535552 296676 535604 296682
rect 535472 296614 535500 296647
rect 535552 296618 535604 296624
rect 535460 296608 535512 296614
rect 535460 296550 535512 296556
rect 535564 295361 535592 296618
rect 535550 295352 535606 295361
rect 535460 295316 535512 295322
rect 535550 295287 535606 295296
rect 535460 295258 535512 295264
rect 535472 294001 535500 295258
rect 535458 293992 535514 294001
rect 535458 293927 535514 293936
rect 535552 293956 535604 293962
rect 535552 293898 535604 293904
rect 535564 292641 535592 293898
rect 535550 292632 535606 292641
rect 535550 292567 535606 292576
rect 535460 292528 535512 292534
rect 535460 292470 535512 292476
rect 535472 291281 535500 292470
rect 535458 291272 535514 291281
rect 535458 291207 535514 291216
rect 535458 289912 535514 289921
rect 535458 289847 535460 289856
rect 535512 289847 535514 289856
rect 535460 289818 535512 289824
rect 535458 288552 535514 288561
rect 535458 288487 535514 288496
rect 535472 288454 535500 288487
rect 535460 288448 535512 288454
rect 535460 288390 535512 288396
rect 523684 284164 523736 284170
rect 523684 284106 523736 284112
rect 535932 263566 535960 360567
rect 536010 328672 536066 328681
rect 536010 328607 536066 328616
rect 536024 318646 536052 328607
rect 536012 318640 536064 318646
rect 536012 318582 536064 318588
rect 536116 284306 536144 397423
rect 536194 388376 536250 388385
rect 536194 388311 536250 388320
rect 536208 373454 536236 388311
rect 536196 373448 536248 373454
rect 536196 373390 536248 373396
rect 536208 359281 536236 373390
rect 536194 359272 536250 359281
rect 536194 359207 536250 359216
rect 536300 318782 536328 400279
rect 536392 339454 536420 401639
rect 536760 396001 536788 424351
rect 538692 422294 538720 445182
rect 541714 445088 541770 445097
rect 541714 445023 541770 445032
rect 544198 445088 544254 445097
rect 544198 445023 544254 445032
rect 538692 422266 538904 422294
rect 538876 409170 538904 422266
rect 547340 412634 547368 445182
rect 547064 412606 547368 412634
rect 547064 409714 547092 412606
rect 546710 409686 547368 409714
rect 541714 409320 541770 409329
rect 544290 409320 544346 409329
rect 544226 409278 544290 409306
rect 541714 409255 541770 409264
rect 544290 409255 544346 409264
rect 538784 409142 539258 409170
rect 536746 395992 536802 396001
rect 536746 395927 536802 395936
rect 538784 393314 538812 409142
rect 547340 404977 547368 409686
rect 547326 404968 547382 404977
rect 547326 404903 547382 404912
rect 538692 393286 538812 393314
rect 538692 383654 538720 393286
rect 538692 383626 538812 383654
rect 538784 373266 538812 383626
rect 547340 373994 547368 404903
rect 547064 373966 547368 373994
rect 544474 373416 544530 373425
rect 544226 373374 544474 373402
rect 544474 373351 544530 373360
rect 547064 373266 547092 373966
rect 538784 373238 539258 373266
rect 546710 373238 547092 373266
rect 536562 364712 536618 364721
rect 536562 364647 536618 364656
rect 536470 363352 536526 363361
rect 536470 363287 536526 363296
rect 536380 339448 536432 339454
rect 536380 339390 536432 339396
rect 536378 324592 536434 324601
rect 536378 324527 536434 324536
rect 536288 318776 536340 318782
rect 536288 318718 536340 318724
rect 536104 284300 536156 284306
rect 536104 284242 536156 284248
rect 535920 263560 535972 263566
rect 535920 263502 535972 263508
rect 536392 263498 536420 324527
rect 536484 303618 536512 363287
rect 536576 318714 536604 364647
rect 538784 354674 538812 373238
rect 541714 373144 541770 373153
rect 541714 373079 541770 373088
rect 547064 364334 547092 373238
rect 547064 364306 547368 364334
rect 538692 354646 538812 354674
rect 536746 352472 536802 352481
rect 536746 352407 536802 352416
rect 536654 327312 536710 327321
rect 536654 327247 536710 327256
rect 536564 318708 536616 318714
rect 536564 318650 536616 318656
rect 536472 303612 536524 303618
rect 536472 303554 536524 303560
rect 536668 303550 536696 327247
rect 536760 323241 536788 352407
rect 538692 345014 538720 354646
rect 547340 345014 547368 364306
rect 538692 344986 538904 345014
rect 538876 337770 538904 344986
rect 547064 344986 547368 345014
rect 541714 339552 541770 339561
rect 541714 339487 541770 339496
rect 544198 339552 544254 339561
rect 544198 339487 544254 339496
rect 538784 337742 539258 337770
rect 541728 337756 541756 339487
rect 544212 337756 544240 339487
rect 547064 337770 547092 344986
rect 546710 337742 547092 337770
rect 536746 323232 536802 323241
rect 536746 323167 536802 323176
rect 536746 316432 536802 316441
rect 536746 316367 536802 316376
rect 536656 303544 536708 303550
rect 536656 303486 536708 303492
rect 536760 287201 536788 316367
rect 538784 316034 538812 337742
rect 547064 335354 547092 337742
rect 547064 335326 547460 335354
rect 538784 316006 538904 316034
rect 538876 301730 538904 316006
rect 547432 306374 547460 335326
rect 547064 306346 547460 306374
rect 544198 303784 544254 303793
rect 544198 303719 544254 303728
rect 541714 303648 541770 303657
rect 541714 303583 541770 303592
rect 538692 301702 539258 301730
rect 541728 301716 541756 303583
rect 544212 301716 544240 303719
rect 547064 301730 547092 306346
rect 547326 303648 547382 303657
rect 547326 303583 547382 303592
rect 546710 301702 547092 301730
rect 536746 287192 536802 287201
rect 536746 287127 536802 287136
rect 536380 263492 536432 263498
rect 536380 263434 536432 263440
rect 519544 263424 519596 263430
rect 519544 263366 519596 263372
rect 502984 263356 503036 263362
rect 502984 263298 503036 263304
rect 538692 245585 538720 301702
rect 547340 300121 547368 303583
rect 547326 300112 547382 300121
rect 547326 300047 547382 300056
rect 580170 300112 580226 300121
rect 580170 300047 580226 300056
rect 580184 298761 580212 300047
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 538678 245576 538734 245585
rect 538678 245511 538734 245520
rect 473728 206984 473780 206990
rect 473728 206926 473780 206932
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 470276 451433 470314 451479
rect 470314 451433 470326 451479
rect 470326 451433 470332 451479
rect 470356 451433 470378 451479
rect 470378 451433 470390 451479
rect 470390 451433 470412 451479
rect 470436 451433 470442 451479
rect 470442 451433 470454 451479
rect 470454 451433 470492 451479
rect 470516 451433 470518 451479
rect 470518 451433 470570 451479
rect 470570 451433 470572 451479
rect 470596 451433 470634 451479
rect 470634 451433 470646 451479
rect 470646 451433 470652 451479
rect 470676 451433 470698 451479
rect 470698 451433 470710 451479
rect 470710 451433 470732 451479
rect 470756 451433 470762 451479
rect 470762 451433 470774 451479
rect 470774 451433 470812 451479
rect 470276 451423 470332 451433
rect 470356 451423 470412 451433
rect 470436 451423 470492 451433
rect 470516 451423 470572 451433
rect 470596 451423 470652 451433
rect 470676 451423 470732 451433
rect 470756 451423 470812 451433
rect 470276 451369 470314 451399
rect 470314 451369 470326 451399
rect 470326 451369 470332 451399
rect 470356 451369 470378 451399
rect 470378 451369 470390 451399
rect 470390 451369 470412 451399
rect 470436 451369 470442 451399
rect 470442 451369 470454 451399
rect 470454 451369 470492 451399
rect 470516 451369 470518 451399
rect 470518 451369 470570 451399
rect 470570 451369 470572 451399
rect 470596 451369 470634 451399
rect 470634 451369 470646 451399
rect 470646 451369 470652 451399
rect 470676 451369 470698 451399
rect 470698 451369 470710 451399
rect 470710 451369 470732 451399
rect 470756 451369 470762 451399
rect 470762 451369 470774 451399
rect 470774 451369 470812 451399
rect 470276 451357 470332 451369
rect 470356 451357 470412 451369
rect 470436 451357 470492 451369
rect 470516 451357 470572 451369
rect 470596 451357 470652 451369
rect 470676 451357 470732 451369
rect 470756 451357 470812 451369
rect 470276 451343 470314 451357
rect 470314 451343 470326 451357
rect 470326 451343 470332 451357
rect 470356 451343 470378 451357
rect 470378 451343 470390 451357
rect 470390 451343 470412 451357
rect 470436 451343 470442 451357
rect 470442 451343 470454 451357
rect 470454 451343 470492 451357
rect 470516 451343 470518 451357
rect 470518 451343 470570 451357
rect 470570 451343 470572 451357
rect 470596 451343 470634 451357
rect 470634 451343 470646 451357
rect 470646 451343 470652 451357
rect 470676 451343 470698 451357
rect 470698 451343 470710 451357
rect 470710 451343 470732 451357
rect 470756 451343 470762 451357
rect 470762 451343 470774 451357
rect 470774 451343 470812 451357
rect 470276 451305 470314 451319
rect 470314 451305 470326 451319
rect 470326 451305 470332 451319
rect 470356 451305 470378 451319
rect 470378 451305 470390 451319
rect 470390 451305 470412 451319
rect 470436 451305 470442 451319
rect 470442 451305 470454 451319
rect 470454 451305 470492 451319
rect 470516 451305 470518 451319
rect 470518 451305 470570 451319
rect 470570 451305 470572 451319
rect 470596 451305 470634 451319
rect 470634 451305 470646 451319
rect 470646 451305 470652 451319
rect 470676 451305 470698 451319
rect 470698 451305 470710 451319
rect 470710 451305 470732 451319
rect 470756 451305 470762 451319
rect 470762 451305 470774 451319
rect 470774 451305 470812 451319
rect 470276 451293 470332 451305
rect 470356 451293 470412 451305
rect 470436 451293 470492 451305
rect 470516 451293 470572 451305
rect 470596 451293 470652 451305
rect 470676 451293 470732 451305
rect 470756 451293 470812 451305
rect 470276 451263 470314 451293
rect 470314 451263 470326 451293
rect 470326 451263 470332 451293
rect 470356 451263 470378 451293
rect 470378 451263 470390 451293
rect 470390 451263 470412 451293
rect 470436 451263 470442 451293
rect 470442 451263 470454 451293
rect 470454 451263 470492 451293
rect 470516 451263 470518 451293
rect 470518 451263 470570 451293
rect 470570 451263 470572 451293
rect 470596 451263 470634 451293
rect 470634 451263 470646 451293
rect 470646 451263 470652 451293
rect 470676 451263 470698 451293
rect 470698 451263 470710 451293
rect 470710 451263 470732 451293
rect 470756 451263 470762 451293
rect 470762 451263 470774 451293
rect 470774 451263 470812 451293
rect 470276 451229 470332 451239
rect 470356 451229 470412 451239
rect 470436 451229 470492 451239
rect 470516 451229 470572 451239
rect 470596 451229 470652 451239
rect 470676 451229 470732 451239
rect 470756 451229 470812 451239
rect 470276 451183 470314 451229
rect 470314 451183 470326 451229
rect 470326 451183 470332 451229
rect 470356 451183 470378 451229
rect 470378 451183 470390 451229
rect 470390 451183 470412 451229
rect 470436 451183 470442 451229
rect 470442 451183 470454 451229
rect 470454 451183 470492 451229
rect 470516 451183 470518 451229
rect 470518 451183 470570 451229
rect 470570 451183 470572 451229
rect 470596 451183 470634 451229
rect 470634 451183 470646 451229
rect 470646 451183 470652 451229
rect 470676 451183 470698 451229
rect 470698 451183 470710 451229
rect 470710 451183 470732 451229
rect 470756 451183 470762 451229
rect 470762 451183 470774 451229
rect 470774 451183 470812 451229
rect 469036 450347 469074 450393
rect 469074 450347 469086 450393
rect 469086 450347 469092 450393
rect 469116 450347 469138 450393
rect 469138 450347 469150 450393
rect 469150 450347 469172 450393
rect 469196 450347 469202 450393
rect 469202 450347 469214 450393
rect 469214 450347 469252 450393
rect 469276 450347 469278 450393
rect 469278 450347 469330 450393
rect 469330 450347 469332 450393
rect 469356 450347 469394 450393
rect 469394 450347 469406 450393
rect 469406 450347 469412 450393
rect 469436 450347 469458 450393
rect 469458 450347 469470 450393
rect 469470 450347 469492 450393
rect 469516 450347 469522 450393
rect 469522 450347 469534 450393
rect 469534 450347 469572 450393
rect 469036 450337 469092 450347
rect 469116 450337 469172 450347
rect 469196 450337 469252 450347
rect 469276 450337 469332 450347
rect 469356 450337 469412 450347
rect 469436 450337 469492 450347
rect 469516 450337 469572 450347
rect 469036 450283 469074 450313
rect 469074 450283 469086 450313
rect 469086 450283 469092 450313
rect 469116 450283 469138 450313
rect 469138 450283 469150 450313
rect 469150 450283 469172 450313
rect 469196 450283 469202 450313
rect 469202 450283 469214 450313
rect 469214 450283 469252 450313
rect 469276 450283 469278 450313
rect 469278 450283 469330 450313
rect 469330 450283 469332 450313
rect 469356 450283 469394 450313
rect 469394 450283 469406 450313
rect 469406 450283 469412 450313
rect 469436 450283 469458 450313
rect 469458 450283 469470 450313
rect 469470 450283 469492 450313
rect 469516 450283 469522 450313
rect 469522 450283 469534 450313
rect 469534 450283 469572 450313
rect 469036 450271 469092 450283
rect 469116 450271 469172 450283
rect 469196 450271 469252 450283
rect 469276 450271 469332 450283
rect 469356 450271 469412 450283
rect 469436 450271 469492 450283
rect 469516 450271 469572 450283
rect 469036 450257 469074 450271
rect 469074 450257 469086 450271
rect 469086 450257 469092 450271
rect 469116 450257 469138 450271
rect 469138 450257 469150 450271
rect 469150 450257 469172 450271
rect 469196 450257 469202 450271
rect 469202 450257 469214 450271
rect 469214 450257 469252 450271
rect 469276 450257 469278 450271
rect 469278 450257 469330 450271
rect 469330 450257 469332 450271
rect 469356 450257 469394 450271
rect 469394 450257 469406 450271
rect 469406 450257 469412 450271
rect 469436 450257 469458 450271
rect 469458 450257 469470 450271
rect 469470 450257 469492 450271
rect 469516 450257 469522 450271
rect 469522 450257 469534 450271
rect 469534 450257 469572 450271
rect 469036 450219 469074 450233
rect 469074 450219 469086 450233
rect 469086 450219 469092 450233
rect 469116 450219 469138 450233
rect 469138 450219 469150 450233
rect 469150 450219 469172 450233
rect 469196 450219 469202 450233
rect 469202 450219 469214 450233
rect 469214 450219 469252 450233
rect 469276 450219 469278 450233
rect 469278 450219 469330 450233
rect 469330 450219 469332 450233
rect 469356 450219 469394 450233
rect 469394 450219 469406 450233
rect 469406 450219 469412 450233
rect 469436 450219 469458 450233
rect 469458 450219 469470 450233
rect 469470 450219 469492 450233
rect 469516 450219 469522 450233
rect 469522 450219 469534 450233
rect 469534 450219 469572 450233
rect 469036 450207 469092 450219
rect 469116 450207 469172 450219
rect 469196 450207 469252 450219
rect 469276 450207 469332 450219
rect 469356 450207 469412 450219
rect 469436 450207 469492 450219
rect 469516 450207 469572 450219
rect 469036 450177 469074 450207
rect 469074 450177 469086 450207
rect 469086 450177 469092 450207
rect 469116 450177 469138 450207
rect 469138 450177 469150 450207
rect 469150 450177 469172 450207
rect 469196 450177 469202 450207
rect 469202 450177 469214 450207
rect 469214 450177 469252 450207
rect 469276 450177 469278 450207
rect 469278 450177 469330 450207
rect 469330 450177 469332 450207
rect 469356 450177 469394 450207
rect 469394 450177 469406 450207
rect 469406 450177 469412 450207
rect 469436 450177 469458 450207
rect 469458 450177 469470 450207
rect 469470 450177 469492 450207
rect 469516 450177 469522 450207
rect 469522 450177 469534 450207
rect 469534 450177 469572 450207
rect 469036 450143 469092 450153
rect 469116 450143 469172 450153
rect 469196 450143 469252 450153
rect 469276 450143 469332 450153
rect 469356 450143 469412 450153
rect 469436 450143 469492 450153
rect 469516 450143 469572 450153
rect 469036 450097 469074 450143
rect 469074 450097 469086 450143
rect 469086 450097 469092 450143
rect 469116 450097 469138 450143
rect 469138 450097 469150 450143
rect 469150 450097 469172 450143
rect 469196 450097 469202 450143
rect 469202 450097 469214 450143
rect 469214 450097 469252 450143
rect 469276 450097 469278 450143
rect 469278 450097 469330 450143
rect 469330 450097 469332 450143
rect 469356 450097 469394 450143
rect 469394 450097 469406 450143
rect 469406 450097 469412 450143
rect 469436 450097 469458 450143
rect 469458 450097 469470 450143
rect 469470 450097 469492 450143
rect 469516 450097 469522 450143
rect 469522 450097 469534 450143
rect 469534 450097 469572 450143
rect 470276 449262 470314 449308
rect 470314 449262 470326 449308
rect 470326 449262 470332 449308
rect 470356 449262 470378 449308
rect 470378 449262 470390 449308
rect 470390 449262 470412 449308
rect 470436 449262 470442 449308
rect 470442 449262 470454 449308
rect 470454 449262 470492 449308
rect 470516 449262 470518 449308
rect 470518 449262 470570 449308
rect 470570 449262 470572 449308
rect 470596 449262 470634 449308
rect 470634 449262 470646 449308
rect 470646 449262 470652 449308
rect 470676 449262 470698 449308
rect 470698 449262 470710 449308
rect 470710 449262 470732 449308
rect 470756 449262 470762 449308
rect 470762 449262 470774 449308
rect 470774 449262 470812 449308
rect 470276 449252 470332 449262
rect 470356 449252 470412 449262
rect 470436 449252 470492 449262
rect 470516 449252 470572 449262
rect 470596 449252 470652 449262
rect 470676 449252 470732 449262
rect 470756 449252 470812 449262
rect 470276 449198 470314 449228
rect 470314 449198 470326 449228
rect 470326 449198 470332 449228
rect 470356 449198 470378 449228
rect 470378 449198 470390 449228
rect 470390 449198 470412 449228
rect 470436 449198 470442 449228
rect 470442 449198 470454 449228
rect 470454 449198 470492 449228
rect 470516 449198 470518 449228
rect 470518 449198 470570 449228
rect 470570 449198 470572 449228
rect 470596 449198 470634 449228
rect 470634 449198 470646 449228
rect 470646 449198 470652 449228
rect 470676 449198 470698 449228
rect 470698 449198 470710 449228
rect 470710 449198 470732 449228
rect 470756 449198 470762 449228
rect 470762 449198 470774 449228
rect 470774 449198 470812 449228
rect 470276 449186 470332 449198
rect 470356 449186 470412 449198
rect 470436 449186 470492 449198
rect 470516 449186 470572 449198
rect 470596 449186 470652 449198
rect 470676 449186 470732 449198
rect 470756 449186 470812 449198
rect 470276 449172 470314 449186
rect 470314 449172 470326 449186
rect 470326 449172 470332 449186
rect 470356 449172 470378 449186
rect 470378 449172 470390 449186
rect 470390 449172 470412 449186
rect 470436 449172 470442 449186
rect 470442 449172 470454 449186
rect 470454 449172 470492 449186
rect 470516 449172 470518 449186
rect 470518 449172 470570 449186
rect 470570 449172 470572 449186
rect 470596 449172 470634 449186
rect 470634 449172 470646 449186
rect 470646 449172 470652 449186
rect 470676 449172 470698 449186
rect 470698 449172 470710 449186
rect 470710 449172 470732 449186
rect 470756 449172 470762 449186
rect 470762 449172 470774 449186
rect 470774 449172 470812 449186
rect 470276 449134 470314 449148
rect 470314 449134 470326 449148
rect 470326 449134 470332 449148
rect 470356 449134 470378 449148
rect 470378 449134 470390 449148
rect 470390 449134 470412 449148
rect 470436 449134 470442 449148
rect 470442 449134 470454 449148
rect 470454 449134 470492 449148
rect 470516 449134 470518 449148
rect 470518 449134 470570 449148
rect 470570 449134 470572 449148
rect 470596 449134 470634 449148
rect 470634 449134 470646 449148
rect 470646 449134 470652 449148
rect 470676 449134 470698 449148
rect 470698 449134 470710 449148
rect 470710 449134 470732 449148
rect 470756 449134 470762 449148
rect 470762 449134 470774 449148
rect 470774 449134 470812 449148
rect 470276 449122 470332 449134
rect 470356 449122 470412 449134
rect 470436 449122 470492 449134
rect 470516 449122 470572 449134
rect 470596 449122 470652 449134
rect 470676 449122 470732 449134
rect 470756 449122 470812 449134
rect 470276 449092 470314 449122
rect 470314 449092 470326 449122
rect 470326 449092 470332 449122
rect 470356 449092 470378 449122
rect 470378 449092 470390 449122
rect 470390 449092 470412 449122
rect 470436 449092 470442 449122
rect 470442 449092 470454 449122
rect 470454 449092 470492 449122
rect 470516 449092 470518 449122
rect 470518 449092 470570 449122
rect 470570 449092 470572 449122
rect 470596 449092 470634 449122
rect 470634 449092 470646 449122
rect 470646 449092 470652 449122
rect 470676 449092 470698 449122
rect 470698 449092 470710 449122
rect 470710 449092 470732 449122
rect 470756 449092 470762 449122
rect 470762 449092 470774 449122
rect 470774 449092 470812 449122
rect 470276 449058 470332 449068
rect 470356 449058 470412 449068
rect 470436 449058 470492 449068
rect 470516 449058 470572 449068
rect 470596 449058 470652 449068
rect 470676 449058 470732 449068
rect 470756 449058 470812 449068
rect 470276 449012 470314 449058
rect 470314 449012 470326 449058
rect 470326 449012 470332 449058
rect 470356 449012 470378 449058
rect 470378 449012 470390 449058
rect 470390 449012 470412 449058
rect 470436 449012 470442 449058
rect 470442 449012 470454 449058
rect 470454 449012 470492 449058
rect 470516 449012 470518 449058
rect 470518 449012 470570 449058
rect 470570 449012 470572 449058
rect 470596 449012 470634 449058
rect 470634 449012 470646 449058
rect 470646 449012 470652 449058
rect 470676 449012 470698 449058
rect 470698 449012 470710 449058
rect 470710 449012 470732 449058
rect 470756 449012 470762 449058
rect 470762 449012 470774 449058
rect 470774 449012 470812 449058
rect 470276 433034 470314 433080
rect 470314 433034 470326 433080
rect 470326 433034 470332 433080
rect 470356 433034 470378 433080
rect 470378 433034 470390 433080
rect 470390 433034 470412 433080
rect 470436 433034 470442 433080
rect 470442 433034 470454 433080
rect 470454 433034 470492 433080
rect 470516 433034 470518 433080
rect 470518 433034 470570 433080
rect 470570 433034 470572 433080
rect 470596 433034 470634 433080
rect 470634 433034 470646 433080
rect 470646 433034 470652 433080
rect 470676 433034 470698 433080
rect 470698 433034 470710 433080
rect 470710 433034 470732 433080
rect 470756 433034 470762 433080
rect 470762 433034 470774 433080
rect 470774 433034 470812 433080
rect 470276 433024 470332 433034
rect 470356 433024 470412 433034
rect 470436 433024 470492 433034
rect 470516 433024 470572 433034
rect 470596 433024 470652 433034
rect 470676 433024 470732 433034
rect 470756 433024 470812 433034
rect 470276 432970 470314 433000
rect 470314 432970 470326 433000
rect 470326 432970 470332 433000
rect 470356 432970 470378 433000
rect 470378 432970 470390 433000
rect 470390 432970 470412 433000
rect 470436 432970 470442 433000
rect 470442 432970 470454 433000
rect 470454 432970 470492 433000
rect 470516 432970 470518 433000
rect 470518 432970 470570 433000
rect 470570 432970 470572 433000
rect 470596 432970 470634 433000
rect 470634 432970 470646 433000
rect 470646 432970 470652 433000
rect 470676 432970 470698 433000
rect 470698 432970 470710 433000
rect 470710 432970 470732 433000
rect 470756 432970 470762 433000
rect 470762 432970 470774 433000
rect 470774 432970 470812 433000
rect 470276 432958 470332 432970
rect 470356 432958 470412 432970
rect 470436 432958 470492 432970
rect 470516 432958 470572 432970
rect 470596 432958 470652 432970
rect 470676 432958 470732 432970
rect 470756 432958 470812 432970
rect 470276 432944 470314 432958
rect 470314 432944 470326 432958
rect 470326 432944 470332 432958
rect 470356 432944 470378 432958
rect 470378 432944 470390 432958
rect 470390 432944 470412 432958
rect 470436 432944 470442 432958
rect 470442 432944 470454 432958
rect 470454 432944 470492 432958
rect 470516 432944 470518 432958
rect 470518 432944 470570 432958
rect 470570 432944 470572 432958
rect 470596 432944 470634 432958
rect 470634 432944 470646 432958
rect 470646 432944 470652 432958
rect 470676 432944 470698 432958
rect 470698 432944 470710 432958
rect 470710 432944 470732 432958
rect 470756 432944 470762 432958
rect 470762 432944 470774 432958
rect 470774 432944 470812 432958
rect 470276 432906 470314 432920
rect 470314 432906 470326 432920
rect 470326 432906 470332 432920
rect 470356 432906 470378 432920
rect 470378 432906 470390 432920
rect 470390 432906 470412 432920
rect 470436 432906 470442 432920
rect 470442 432906 470454 432920
rect 470454 432906 470492 432920
rect 470516 432906 470518 432920
rect 470518 432906 470570 432920
rect 470570 432906 470572 432920
rect 470596 432906 470634 432920
rect 470634 432906 470646 432920
rect 470646 432906 470652 432920
rect 470676 432906 470698 432920
rect 470698 432906 470710 432920
rect 470710 432906 470732 432920
rect 470756 432906 470762 432920
rect 470762 432906 470774 432920
rect 470774 432906 470812 432920
rect 470276 432894 470332 432906
rect 470356 432894 470412 432906
rect 470436 432894 470492 432906
rect 470516 432894 470572 432906
rect 470596 432894 470652 432906
rect 470676 432894 470732 432906
rect 470756 432894 470812 432906
rect 470276 432864 470314 432894
rect 470314 432864 470326 432894
rect 470326 432864 470332 432894
rect 470356 432864 470378 432894
rect 470378 432864 470390 432894
rect 470390 432864 470412 432894
rect 470436 432864 470442 432894
rect 470442 432864 470454 432894
rect 470454 432864 470492 432894
rect 470516 432864 470518 432894
rect 470518 432864 470570 432894
rect 470570 432864 470572 432894
rect 470596 432864 470634 432894
rect 470634 432864 470646 432894
rect 470646 432864 470652 432894
rect 470676 432864 470698 432894
rect 470698 432864 470710 432894
rect 470710 432864 470732 432894
rect 470756 432864 470762 432894
rect 470762 432864 470774 432894
rect 470774 432864 470812 432894
rect 470276 432830 470332 432840
rect 470356 432830 470412 432840
rect 470436 432830 470492 432840
rect 470516 432830 470572 432840
rect 470596 432830 470652 432840
rect 470676 432830 470732 432840
rect 470756 432830 470812 432840
rect 470276 432784 470314 432830
rect 470314 432784 470326 432830
rect 470326 432784 470332 432830
rect 470356 432784 470378 432830
rect 470378 432784 470390 432830
rect 470390 432784 470412 432830
rect 470436 432784 470442 432830
rect 470442 432784 470454 432830
rect 470454 432784 470492 432830
rect 470516 432784 470518 432830
rect 470518 432784 470570 432830
rect 470570 432784 470572 432830
rect 470596 432784 470634 432830
rect 470634 432784 470646 432830
rect 470646 432784 470652 432830
rect 470676 432784 470698 432830
rect 470698 432784 470710 432830
rect 470710 432784 470732 432830
rect 470756 432784 470762 432830
rect 470762 432784 470774 432830
rect 470774 432784 470812 432830
rect 477843 450200 477899 450256
rect 481160 450200 481216 450256
rect 484477 450200 484533 450256
rect 487793 450200 487849 450256
rect 474094 449656 474150 449712
rect 469036 431947 469074 431993
rect 469074 431947 469086 431993
rect 469086 431947 469092 431993
rect 469116 431947 469138 431993
rect 469138 431947 469150 431993
rect 469150 431947 469172 431993
rect 469196 431947 469202 431993
rect 469202 431947 469214 431993
rect 469214 431947 469252 431993
rect 469276 431947 469278 431993
rect 469278 431947 469330 431993
rect 469330 431947 469332 431993
rect 469356 431947 469394 431993
rect 469394 431947 469406 431993
rect 469406 431947 469412 431993
rect 469436 431947 469458 431993
rect 469458 431947 469470 431993
rect 469470 431947 469492 431993
rect 469516 431947 469522 431993
rect 469522 431947 469534 431993
rect 469534 431947 469572 431993
rect 469036 431937 469092 431947
rect 469116 431937 469172 431947
rect 469196 431937 469252 431947
rect 469276 431937 469332 431947
rect 469356 431937 469412 431947
rect 469436 431937 469492 431947
rect 469516 431937 469572 431947
rect 469036 431883 469074 431913
rect 469074 431883 469086 431913
rect 469086 431883 469092 431913
rect 469116 431883 469138 431913
rect 469138 431883 469150 431913
rect 469150 431883 469172 431913
rect 469196 431883 469202 431913
rect 469202 431883 469214 431913
rect 469214 431883 469252 431913
rect 469276 431883 469278 431913
rect 469278 431883 469330 431913
rect 469330 431883 469332 431913
rect 469356 431883 469394 431913
rect 469394 431883 469406 431913
rect 469406 431883 469412 431913
rect 469436 431883 469458 431913
rect 469458 431883 469470 431913
rect 469470 431883 469492 431913
rect 469516 431883 469522 431913
rect 469522 431883 469534 431913
rect 469534 431883 469572 431913
rect 469036 431871 469092 431883
rect 469116 431871 469172 431883
rect 469196 431871 469252 431883
rect 469276 431871 469332 431883
rect 469356 431871 469412 431883
rect 469436 431871 469492 431883
rect 469516 431871 469572 431883
rect 469036 431857 469074 431871
rect 469074 431857 469086 431871
rect 469086 431857 469092 431871
rect 469116 431857 469138 431871
rect 469138 431857 469150 431871
rect 469150 431857 469172 431871
rect 469196 431857 469202 431871
rect 469202 431857 469214 431871
rect 469214 431857 469252 431871
rect 469276 431857 469278 431871
rect 469278 431857 469330 431871
rect 469330 431857 469332 431871
rect 469356 431857 469394 431871
rect 469394 431857 469406 431871
rect 469406 431857 469412 431871
rect 469436 431857 469458 431871
rect 469458 431857 469470 431871
rect 469470 431857 469492 431871
rect 469516 431857 469522 431871
rect 469522 431857 469534 431871
rect 469534 431857 469572 431871
rect 469036 431819 469074 431833
rect 469074 431819 469086 431833
rect 469086 431819 469092 431833
rect 469116 431819 469138 431833
rect 469138 431819 469150 431833
rect 469150 431819 469172 431833
rect 469196 431819 469202 431833
rect 469202 431819 469214 431833
rect 469214 431819 469252 431833
rect 469276 431819 469278 431833
rect 469278 431819 469330 431833
rect 469330 431819 469332 431833
rect 469356 431819 469394 431833
rect 469394 431819 469406 431833
rect 469406 431819 469412 431833
rect 469436 431819 469458 431833
rect 469458 431819 469470 431833
rect 469470 431819 469492 431833
rect 469516 431819 469522 431833
rect 469522 431819 469534 431833
rect 469534 431819 469572 431833
rect 469036 431807 469092 431819
rect 469116 431807 469172 431819
rect 469196 431807 469252 431819
rect 469276 431807 469332 431819
rect 469356 431807 469412 431819
rect 469436 431807 469492 431819
rect 469516 431807 469572 431819
rect 469036 431777 469074 431807
rect 469074 431777 469086 431807
rect 469086 431777 469092 431807
rect 469116 431777 469138 431807
rect 469138 431777 469150 431807
rect 469150 431777 469172 431807
rect 469196 431777 469202 431807
rect 469202 431777 469214 431807
rect 469214 431777 469252 431807
rect 469276 431777 469278 431807
rect 469278 431777 469330 431807
rect 469330 431777 469332 431807
rect 469356 431777 469394 431807
rect 469394 431777 469406 431807
rect 469406 431777 469412 431807
rect 469436 431777 469458 431807
rect 469458 431777 469470 431807
rect 469470 431777 469492 431807
rect 469516 431777 469522 431807
rect 469522 431777 469534 431807
rect 469534 431777 469572 431807
rect 469036 431743 469092 431753
rect 469116 431743 469172 431753
rect 469196 431743 469252 431753
rect 469276 431743 469332 431753
rect 469356 431743 469412 431753
rect 469436 431743 469492 431753
rect 469516 431743 469572 431753
rect 469036 431697 469074 431743
rect 469074 431697 469086 431743
rect 469086 431697 469092 431743
rect 469116 431697 469138 431743
rect 469138 431697 469150 431743
rect 469150 431697 469172 431743
rect 469196 431697 469202 431743
rect 469202 431697 469214 431743
rect 469214 431697 469252 431743
rect 469276 431697 469278 431743
rect 469278 431697 469330 431743
rect 469330 431697 469332 431743
rect 469356 431697 469394 431743
rect 469394 431697 469406 431743
rect 469406 431697 469412 431743
rect 469436 431697 469458 431743
rect 469458 431697 469470 431743
rect 469470 431697 469492 431743
rect 469516 431697 469522 431743
rect 469522 431697 469534 431743
rect 469534 431697 469572 431743
rect 470276 430862 470314 430908
rect 470314 430862 470326 430908
rect 470326 430862 470332 430908
rect 470356 430862 470378 430908
rect 470378 430862 470390 430908
rect 470390 430862 470412 430908
rect 470436 430862 470442 430908
rect 470442 430862 470454 430908
rect 470454 430862 470492 430908
rect 470516 430862 470518 430908
rect 470518 430862 470570 430908
rect 470570 430862 470572 430908
rect 470596 430862 470634 430908
rect 470634 430862 470646 430908
rect 470646 430862 470652 430908
rect 470676 430862 470698 430908
rect 470698 430862 470710 430908
rect 470710 430862 470732 430908
rect 470756 430862 470762 430908
rect 470762 430862 470774 430908
rect 470774 430862 470812 430908
rect 470276 430852 470332 430862
rect 470356 430852 470412 430862
rect 470436 430852 470492 430862
rect 470516 430852 470572 430862
rect 470596 430852 470652 430862
rect 470676 430852 470732 430862
rect 470756 430852 470812 430862
rect 470276 430798 470314 430828
rect 470314 430798 470326 430828
rect 470326 430798 470332 430828
rect 470356 430798 470378 430828
rect 470378 430798 470390 430828
rect 470390 430798 470412 430828
rect 470436 430798 470442 430828
rect 470442 430798 470454 430828
rect 470454 430798 470492 430828
rect 470516 430798 470518 430828
rect 470518 430798 470570 430828
rect 470570 430798 470572 430828
rect 470596 430798 470634 430828
rect 470634 430798 470646 430828
rect 470646 430798 470652 430828
rect 470676 430798 470698 430828
rect 470698 430798 470710 430828
rect 470710 430798 470732 430828
rect 470756 430798 470762 430828
rect 470762 430798 470774 430828
rect 470774 430798 470812 430828
rect 470276 430786 470332 430798
rect 470356 430786 470412 430798
rect 470436 430786 470492 430798
rect 470516 430786 470572 430798
rect 470596 430786 470652 430798
rect 470676 430786 470732 430798
rect 470756 430786 470812 430798
rect 470276 430772 470314 430786
rect 470314 430772 470326 430786
rect 470326 430772 470332 430786
rect 470356 430772 470378 430786
rect 470378 430772 470390 430786
rect 470390 430772 470412 430786
rect 470436 430772 470442 430786
rect 470442 430772 470454 430786
rect 470454 430772 470492 430786
rect 470516 430772 470518 430786
rect 470518 430772 470570 430786
rect 470570 430772 470572 430786
rect 470596 430772 470634 430786
rect 470634 430772 470646 430786
rect 470646 430772 470652 430786
rect 470676 430772 470698 430786
rect 470698 430772 470710 430786
rect 470710 430772 470732 430786
rect 470756 430772 470762 430786
rect 470762 430772 470774 430786
rect 470774 430772 470812 430786
rect 470276 430734 470314 430748
rect 470314 430734 470326 430748
rect 470326 430734 470332 430748
rect 470356 430734 470378 430748
rect 470378 430734 470390 430748
rect 470390 430734 470412 430748
rect 470436 430734 470442 430748
rect 470442 430734 470454 430748
rect 470454 430734 470492 430748
rect 470516 430734 470518 430748
rect 470518 430734 470570 430748
rect 470570 430734 470572 430748
rect 470596 430734 470634 430748
rect 470634 430734 470646 430748
rect 470646 430734 470652 430748
rect 470676 430734 470698 430748
rect 470698 430734 470710 430748
rect 470710 430734 470732 430748
rect 470756 430734 470762 430748
rect 470762 430734 470774 430748
rect 470774 430734 470812 430748
rect 470276 430722 470332 430734
rect 470356 430722 470412 430734
rect 470436 430722 470492 430734
rect 470516 430722 470572 430734
rect 470596 430722 470652 430734
rect 470676 430722 470732 430734
rect 470756 430722 470812 430734
rect 470276 430692 470314 430722
rect 470314 430692 470326 430722
rect 470326 430692 470332 430722
rect 470356 430692 470378 430722
rect 470378 430692 470390 430722
rect 470390 430692 470412 430722
rect 470436 430692 470442 430722
rect 470442 430692 470454 430722
rect 470454 430692 470492 430722
rect 470516 430692 470518 430722
rect 470518 430692 470570 430722
rect 470570 430692 470572 430722
rect 470596 430692 470634 430722
rect 470634 430692 470646 430722
rect 470646 430692 470652 430722
rect 470676 430692 470698 430722
rect 470698 430692 470710 430722
rect 470710 430692 470732 430722
rect 470756 430692 470762 430722
rect 470762 430692 470774 430722
rect 470774 430692 470812 430722
rect 470276 430658 470332 430668
rect 470356 430658 470412 430668
rect 470436 430658 470492 430668
rect 470516 430658 470572 430668
rect 470596 430658 470652 430668
rect 470676 430658 470732 430668
rect 470756 430658 470812 430668
rect 470276 430612 470314 430658
rect 470314 430612 470326 430658
rect 470326 430612 470332 430658
rect 470356 430612 470378 430658
rect 470378 430612 470390 430658
rect 470390 430612 470412 430658
rect 470436 430612 470442 430658
rect 470442 430612 470454 430658
rect 470454 430612 470492 430658
rect 470516 430612 470518 430658
rect 470518 430612 470570 430658
rect 470570 430612 470572 430658
rect 470596 430612 470634 430658
rect 470634 430612 470646 430658
rect 470646 430612 470652 430658
rect 470676 430612 470698 430658
rect 470698 430612 470710 430658
rect 470710 430612 470732 430658
rect 470756 430612 470762 430658
rect 470762 430612 470774 430658
rect 470774 430612 470812 430658
rect 470276 412034 470314 412080
rect 470314 412034 470326 412080
rect 470326 412034 470332 412080
rect 470356 412034 470378 412080
rect 470378 412034 470390 412080
rect 470390 412034 470412 412080
rect 470436 412034 470442 412080
rect 470442 412034 470454 412080
rect 470454 412034 470492 412080
rect 470516 412034 470518 412080
rect 470518 412034 470570 412080
rect 470570 412034 470572 412080
rect 470596 412034 470634 412080
rect 470634 412034 470646 412080
rect 470646 412034 470652 412080
rect 470676 412034 470698 412080
rect 470698 412034 470710 412080
rect 470710 412034 470732 412080
rect 470756 412034 470762 412080
rect 470762 412034 470774 412080
rect 470774 412034 470812 412080
rect 470276 412024 470332 412034
rect 470356 412024 470412 412034
rect 470436 412024 470492 412034
rect 470516 412024 470572 412034
rect 470596 412024 470652 412034
rect 470676 412024 470732 412034
rect 470756 412024 470812 412034
rect 470276 411970 470314 412000
rect 470314 411970 470326 412000
rect 470326 411970 470332 412000
rect 470356 411970 470378 412000
rect 470378 411970 470390 412000
rect 470390 411970 470412 412000
rect 470436 411970 470442 412000
rect 470442 411970 470454 412000
rect 470454 411970 470492 412000
rect 470516 411970 470518 412000
rect 470518 411970 470570 412000
rect 470570 411970 470572 412000
rect 470596 411970 470634 412000
rect 470634 411970 470646 412000
rect 470646 411970 470652 412000
rect 470676 411970 470698 412000
rect 470698 411970 470710 412000
rect 470710 411970 470732 412000
rect 470756 411970 470762 412000
rect 470762 411970 470774 412000
rect 470774 411970 470812 412000
rect 470276 411958 470332 411970
rect 470356 411958 470412 411970
rect 470436 411958 470492 411970
rect 470516 411958 470572 411970
rect 470596 411958 470652 411970
rect 470676 411958 470732 411970
rect 470756 411958 470812 411970
rect 470276 411944 470314 411958
rect 470314 411944 470326 411958
rect 470326 411944 470332 411958
rect 470356 411944 470378 411958
rect 470378 411944 470390 411958
rect 470390 411944 470412 411958
rect 470436 411944 470442 411958
rect 470442 411944 470454 411958
rect 470454 411944 470492 411958
rect 470516 411944 470518 411958
rect 470518 411944 470570 411958
rect 470570 411944 470572 411958
rect 470596 411944 470634 411958
rect 470634 411944 470646 411958
rect 470646 411944 470652 411958
rect 470676 411944 470698 411958
rect 470698 411944 470710 411958
rect 470710 411944 470732 411958
rect 470756 411944 470762 411958
rect 470762 411944 470774 411958
rect 470774 411944 470812 411958
rect 470276 411906 470314 411920
rect 470314 411906 470326 411920
rect 470326 411906 470332 411920
rect 470356 411906 470378 411920
rect 470378 411906 470390 411920
rect 470390 411906 470412 411920
rect 470436 411906 470442 411920
rect 470442 411906 470454 411920
rect 470454 411906 470492 411920
rect 470516 411906 470518 411920
rect 470518 411906 470570 411920
rect 470570 411906 470572 411920
rect 470596 411906 470634 411920
rect 470634 411906 470646 411920
rect 470646 411906 470652 411920
rect 470676 411906 470698 411920
rect 470698 411906 470710 411920
rect 470710 411906 470732 411920
rect 470756 411906 470762 411920
rect 470762 411906 470774 411920
rect 470774 411906 470812 411920
rect 470276 411894 470332 411906
rect 470356 411894 470412 411906
rect 470436 411894 470492 411906
rect 470516 411894 470572 411906
rect 470596 411894 470652 411906
rect 470676 411894 470732 411906
rect 470756 411894 470812 411906
rect 470276 411864 470314 411894
rect 470314 411864 470326 411894
rect 470326 411864 470332 411894
rect 470356 411864 470378 411894
rect 470378 411864 470390 411894
rect 470390 411864 470412 411894
rect 470436 411864 470442 411894
rect 470442 411864 470454 411894
rect 470454 411864 470492 411894
rect 470516 411864 470518 411894
rect 470518 411864 470570 411894
rect 470570 411864 470572 411894
rect 470596 411864 470634 411894
rect 470634 411864 470646 411894
rect 470646 411864 470652 411894
rect 470676 411864 470698 411894
rect 470698 411864 470710 411894
rect 470710 411864 470732 411894
rect 470756 411864 470762 411894
rect 470762 411864 470774 411894
rect 470774 411864 470812 411894
rect 470276 411830 470332 411840
rect 470356 411830 470412 411840
rect 470436 411830 470492 411840
rect 470516 411830 470572 411840
rect 470596 411830 470652 411840
rect 470676 411830 470732 411840
rect 470756 411830 470812 411840
rect 470276 411784 470314 411830
rect 470314 411784 470326 411830
rect 470326 411784 470332 411830
rect 470356 411784 470378 411830
rect 470378 411784 470390 411830
rect 470390 411784 470412 411830
rect 470436 411784 470442 411830
rect 470442 411784 470454 411830
rect 470454 411784 470492 411830
rect 470516 411784 470518 411830
rect 470518 411784 470570 411830
rect 470570 411784 470572 411830
rect 470596 411784 470634 411830
rect 470634 411784 470646 411830
rect 470646 411784 470652 411830
rect 470676 411784 470698 411830
rect 470698 411784 470710 411830
rect 470710 411784 470732 411830
rect 470756 411784 470762 411830
rect 470762 411784 470774 411830
rect 470774 411784 470812 411830
rect 483570 432248 483626 432304
rect 481270 432112 481326 432168
rect 474278 431840 474334 431896
rect 488078 431840 488134 431896
rect 478102 431568 478158 431624
rect 478970 427896 479026 427952
rect 485778 427896 485834 427952
rect 469036 410948 469074 410994
rect 469074 410948 469086 410994
rect 469086 410948 469092 410994
rect 469116 410948 469138 410994
rect 469138 410948 469150 410994
rect 469150 410948 469172 410994
rect 469196 410948 469202 410994
rect 469202 410948 469214 410994
rect 469214 410948 469252 410994
rect 469276 410948 469278 410994
rect 469278 410948 469330 410994
rect 469330 410948 469332 410994
rect 469356 410948 469394 410994
rect 469394 410948 469406 410994
rect 469406 410948 469412 410994
rect 469436 410948 469458 410994
rect 469458 410948 469470 410994
rect 469470 410948 469492 410994
rect 469516 410948 469522 410994
rect 469522 410948 469534 410994
rect 469534 410948 469572 410994
rect 469036 410938 469092 410948
rect 469116 410938 469172 410948
rect 469196 410938 469252 410948
rect 469276 410938 469332 410948
rect 469356 410938 469412 410948
rect 469436 410938 469492 410948
rect 469516 410938 469572 410948
rect 469036 410884 469074 410914
rect 469074 410884 469086 410914
rect 469086 410884 469092 410914
rect 469116 410884 469138 410914
rect 469138 410884 469150 410914
rect 469150 410884 469172 410914
rect 469196 410884 469202 410914
rect 469202 410884 469214 410914
rect 469214 410884 469252 410914
rect 469276 410884 469278 410914
rect 469278 410884 469330 410914
rect 469330 410884 469332 410914
rect 469356 410884 469394 410914
rect 469394 410884 469406 410914
rect 469406 410884 469412 410914
rect 469436 410884 469458 410914
rect 469458 410884 469470 410914
rect 469470 410884 469492 410914
rect 469516 410884 469522 410914
rect 469522 410884 469534 410914
rect 469534 410884 469572 410914
rect 469036 410872 469092 410884
rect 469116 410872 469172 410884
rect 469196 410872 469252 410884
rect 469276 410872 469332 410884
rect 469356 410872 469412 410884
rect 469436 410872 469492 410884
rect 469516 410872 469572 410884
rect 469036 410858 469074 410872
rect 469074 410858 469086 410872
rect 469086 410858 469092 410872
rect 469116 410858 469138 410872
rect 469138 410858 469150 410872
rect 469150 410858 469172 410872
rect 469196 410858 469202 410872
rect 469202 410858 469214 410872
rect 469214 410858 469252 410872
rect 469276 410858 469278 410872
rect 469278 410858 469330 410872
rect 469330 410858 469332 410872
rect 469356 410858 469394 410872
rect 469394 410858 469406 410872
rect 469406 410858 469412 410872
rect 469436 410858 469458 410872
rect 469458 410858 469470 410872
rect 469470 410858 469492 410872
rect 469516 410858 469522 410872
rect 469522 410858 469534 410872
rect 469534 410858 469572 410872
rect 469036 410820 469074 410834
rect 469074 410820 469086 410834
rect 469086 410820 469092 410834
rect 469116 410820 469138 410834
rect 469138 410820 469150 410834
rect 469150 410820 469172 410834
rect 469196 410820 469202 410834
rect 469202 410820 469214 410834
rect 469214 410820 469252 410834
rect 469276 410820 469278 410834
rect 469278 410820 469330 410834
rect 469330 410820 469332 410834
rect 469356 410820 469394 410834
rect 469394 410820 469406 410834
rect 469406 410820 469412 410834
rect 469436 410820 469458 410834
rect 469458 410820 469470 410834
rect 469470 410820 469492 410834
rect 469516 410820 469522 410834
rect 469522 410820 469534 410834
rect 469534 410820 469572 410834
rect 469036 410808 469092 410820
rect 469116 410808 469172 410820
rect 469196 410808 469252 410820
rect 469276 410808 469332 410820
rect 469356 410808 469412 410820
rect 469436 410808 469492 410820
rect 469516 410808 469572 410820
rect 469036 410778 469074 410808
rect 469074 410778 469086 410808
rect 469086 410778 469092 410808
rect 469116 410778 469138 410808
rect 469138 410778 469150 410808
rect 469150 410778 469172 410808
rect 469196 410778 469202 410808
rect 469202 410778 469214 410808
rect 469214 410778 469252 410808
rect 469276 410778 469278 410808
rect 469278 410778 469330 410808
rect 469330 410778 469332 410808
rect 469356 410778 469394 410808
rect 469394 410778 469406 410808
rect 469406 410778 469412 410808
rect 469436 410778 469458 410808
rect 469458 410778 469470 410808
rect 469470 410778 469492 410808
rect 469516 410778 469522 410808
rect 469522 410778 469534 410808
rect 469534 410778 469572 410808
rect 469036 410744 469092 410754
rect 469116 410744 469172 410754
rect 469196 410744 469252 410754
rect 469276 410744 469332 410754
rect 469356 410744 469412 410754
rect 469436 410744 469492 410754
rect 469516 410744 469572 410754
rect 469036 410698 469074 410744
rect 469074 410698 469086 410744
rect 469086 410698 469092 410744
rect 469116 410698 469138 410744
rect 469138 410698 469150 410744
rect 469150 410698 469172 410744
rect 469196 410698 469202 410744
rect 469202 410698 469214 410744
rect 469214 410698 469252 410744
rect 469276 410698 469278 410744
rect 469278 410698 469330 410744
rect 469330 410698 469332 410744
rect 469356 410698 469394 410744
rect 469394 410698 469406 410744
rect 469406 410698 469412 410744
rect 469436 410698 469458 410744
rect 469458 410698 469470 410744
rect 469470 410698 469492 410744
rect 469516 410698 469522 410744
rect 469522 410698 469534 410744
rect 469534 410698 469572 410744
rect 470276 409862 470314 409908
rect 470314 409862 470326 409908
rect 470326 409862 470332 409908
rect 470356 409862 470378 409908
rect 470378 409862 470390 409908
rect 470390 409862 470412 409908
rect 470436 409862 470442 409908
rect 470442 409862 470454 409908
rect 470454 409862 470492 409908
rect 470516 409862 470518 409908
rect 470518 409862 470570 409908
rect 470570 409862 470572 409908
rect 470596 409862 470634 409908
rect 470634 409862 470646 409908
rect 470646 409862 470652 409908
rect 470676 409862 470698 409908
rect 470698 409862 470710 409908
rect 470710 409862 470732 409908
rect 470756 409862 470762 409908
rect 470762 409862 470774 409908
rect 470774 409862 470812 409908
rect 470276 409852 470332 409862
rect 470356 409852 470412 409862
rect 470436 409852 470492 409862
rect 470516 409852 470572 409862
rect 470596 409852 470652 409862
rect 470676 409852 470732 409862
rect 470756 409852 470812 409862
rect 470276 409798 470314 409828
rect 470314 409798 470326 409828
rect 470326 409798 470332 409828
rect 470356 409798 470378 409828
rect 470378 409798 470390 409828
rect 470390 409798 470412 409828
rect 470436 409798 470442 409828
rect 470442 409798 470454 409828
rect 470454 409798 470492 409828
rect 470516 409798 470518 409828
rect 470518 409798 470570 409828
rect 470570 409798 470572 409828
rect 470596 409798 470634 409828
rect 470634 409798 470646 409828
rect 470646 409798 470652 409828
rect 470676 409798 470698 409828
rect 470698 409798 470710 409828
rect 470710 409798 470732 409828
rect 470756 409798 470762 409828
rect 470762 409798 470774 409828
rect 470774 409798 470812 409828
rect 470276 409786 470332 409798
rect 470356 409786 470412 409798
rect 470436 409786 470492 409798
rect 470516 409786 470572 409798
rect 470596 409786 470652 409798
rect 470676 409786 470732 409798
rect 470756 409786 470812 409798
rect 470276 409772 470314 409786
rect 470314 409772 470326 409786
rect 470326 409772 470332 409786
rect 470356 409772 470378 409786
rect 470378 409772 470390 409786
rect 470390 409772 470412 409786
rect 470436 409772 470442 409786
rect 470442 409772 470454 409786
rect 470454 409772 470492 409786
rect 470516 409772 470518 409786
rect 470518 409772 470570 409786
rect 470570 409772 470572 409786
rect 470596 409772 470634 409786
rect 470634 409772 470646 409786
rect 470646 409772 470652 409786
rect 470676 409772 470698 409786
rect 470698 409772 470710 409786
rect 470710 409772 470732 409786
rect 470756 409772 470762 409786
rect 470762 409772 470774 409786
rect 470774 409772 470812 409786
rect 470276 409734 470314 409748
rect 470314 409734 470326 409748
rect 470326 409734 470332 409748
rect 470356 409734 470378 409748
rect 470378 409734 470390 409748
rect 470390 409734 470412 409748
rect 470436 409734 470442 409748
rect 470442 409734 470454 409748
rect 470454 409734 470492 409748
rect 470516 409734 470518 409748
rect 470518 409734 470570 409748
rect 470570 409734 470572 409748
rect 470596 409734 470634 409748
rect 470634 409734 470646 409748
rect 470646 409734 470652 409748
rect 470676 409734 470698 409748
rect 470698 409734 470710 409748
rect 470710 409734 470732 409748
rect 470756 409734 470762 409748
rect 470762 409734 470774 409748
rect 470774 409734 470812 409748
rect 470276 409722 470332 409734
rect 470356 409722 470412 409734
rect 470436 409722 470492 409734
rect 470516 409722 470572 409734
rect 470596 409722 470652 409734
rect 470676 409722 470732 409734
rect 470756 409722 470812 409734
rect 470276 409692 470314 409722
rect 470314 409692 470326 409722
rect 470326 409692 470332 409722
rect 470356 409692 470378 409722
rect 470378 409692 470390 409722
rect 470390 409692 470412 409722
rect 470436 409692 470442 409722
rect 470442 409692 470454 409722
rect 470454 409692 470492 409722
rect 470516 409692 470518 409722
rect 470518 409692 470570 409722
rect 470570 409692 470572 409722
rect 470596 409692 470634 409722
rect 470634 409692 470646 409722
rect 470646 409692 470652 409722
rect 470676 409692 470698 409722
rect 470698 409692 470710 409722
rect 470710 409692 470732 409722
rect 470756 409692 470762 409722
rect 470762 409692 470774 409722
rect 470774 409692 470812 409722
rect 470276 409658 470332 409668
rect 470356 409658 470412 409668
rect 470436 409658 470492 409668
rect 470516 409658 470572 409668
rect 470596 409658 470652 409668
rect 470676 409658 470732 409668
rect 470756 409658 470812 409668
rect 470276 409612 470314 409658
rect 470314 409612 470326 409658
rect 470326 409612 470332 409658
rect 470356 409612 470378 409658
rect 470378 409612 470390 409658
rect 470390 409612 470412 409658
rect 470436 409612 470442 409658
rect 470442 409612 470454 409658
rect 470454 409612 470492 409658
rect 470516 409612 470518 409658
rect 470518 409612 470570 409658
rect 470570 409612 470572 409658
rect 470596 409612 470634 409658
rect 470634 409612 470646 409658
rect 470646 409612 470652 409658
rect 470676 409612 470698 409658
rect 470698 409612 470710 409658
rect 470710 409612 470732 409658
rect 470756 409612 470762 409658
rect 470762 409612 470774 409658
rect 470774 409612 470812 409658
rect 470276 391035 470314 391081
rect 470314 391035 470326 391081
rect 470326 391035 470332 391081
rect 470356 391035 470378 391081
rect 470378 391035 470390 391081
rect 470390 391035 470412 391081
rect 470436 391035 470442 391081
rect 470442 391035 470454 391081
rect 470454 391035 470492 391081
rect 470516 391035 470518 391081
rect 470518 391035 470570 391081
rect 470570 391035 470572 391081
rect 470596 391035 470634 391081
rect 470634 391035 470646 391081
rect 470646 391035 470652 391081
rect 470676 391035 470698 391081
rect 470698 391035 470710 391081
rect 470710 391035 470732 391081
rect 470756 391035 470762 391081
rect 470762 391035 470774 391081
rect 470774 391035 470812 391081
rect 470276 391025 470332 391035
rect 470356 391025 470412 391035
rect 470436 391025 470492 391035
rect 470516 391025 470572 391035
rect 470596 391025 470652 391035
rect 470676 391025 470732 391035
rect 470756 391025 470812 391035
rect 470276 390971 470314 391001
rect 470314 390971 470326 391001
rect 470326 390971 470332 391001
rect 470356 390971 470378 391001
rect 470378 390971 470390 391001
rect 470390 390971 470412 391001
rect 470436 390971 470442 391001
rect 470442 390971 470454 391001
rect 470454 390971 470492 391001
rect 470516 390971 470518 391001
rect 470518 390971 470570 391001
rect 470570 390971 470572 391001
rect 470596 390971 470634 391001
rect 470634 390971 470646 391001
rect 470646 390971 470652 391001
rect 470676 390971 470698 391001
rect 470698 390971 470710 391001
rect 470710 390971 470732 391001
rect 470756 390971 470762 391001
rect 470762 390971 470774 391001
rect 470774 390971 470812 391001
rect 470276 390959 470332 390971
rect 470356 390959 470412 390971
rect 470436 390959 470492 390971
rect 470516 390959 470572 390971
rect 470596 390959 470652 390971
rect 470676 390959 470732 390971
rect 470756 390959 470812 390971
rect 470276 390945 470314 390959
rect 470314 390945 470326 390959
rect 470326 390945 470332 390959
rect 470356 390945 470378 390959
rect 470378 390945 470390 390959
rect 470390 390945 470412 390959
rect 470436 390945 470442 390959
rect 470442 390945 470454 390959
rect 470454 390945 470492 390959
rect 470516 390945 470518 390959
rect 470518 390945 470570 390959
rect 470570 390945 470572 390959
rect 470596 390945 470634 390959
rect 470634 390945 470646 390959
rect 470646 390945 470652 390959
rect 470676 390945 470698 390959
rect 470698 390945 470710 390959
rect 470710 390945 470732 390959
rect 470756 390945 470762 390959
rect 470762 390945 470774 390959
rect 470774 390945 470812 390959
rect 470276 390907 470314 390921
rect 470314 390907 470326 390921
rect 470326 390907 470332 390921
rect 470356 390907 470378 390921
rect 470378 390907 470390 390921
rect 470390 390907 470412 390921
rect 470436 390907 470442 390921
rect 470442 390907 470454 390921
rect 470454 390907 470492 390921
rect 470516 390907 470518 390921
rect 470518 390907 470570 390921
rect 470570 390907 470572 390921
rect 470596 390907 470634 390921
rect 470634 390907 470646 390921
rect 470646 390907 470652 390921
rect 470676 390907 470698 390921
rect 470698 390907 470710 390921
rect 470710 390907 470732 390921
rect 470756 390907 470762 390921
rect 470762 390907 470774 390921
rect 470774 390907 470812 390921
rect 470276 390895 470332 390907
rect 470356 390895 470412 390907
rect 470436 390895 470492 390907
rect 470516 390895 470572 390907
rect 470596 390895 470652 390907
rect 470676 390895 470732 390907
rect 470756 390895 470812 390907
rect 470276 390865 470314 390895
rect 470314 390865 470326 390895
rect 470326 390865 470332 390895
rect 470356 390865 470378 390895
rect 470378 390865 470390 390895
rect 470390 390865 470412 390895
rect 470436 390865 470442 390895
rect 470442 390865 470454 390895
rect 470454 390865 470492 390895
rect 470516 390865 470518 390895
rect 470518 390865 470570 390895
rect 470570 390865 470572 390895
rect 470596 390865 470634 390895
rect 470634 390865 470646 390895
rect 470646 390865 470652 390895
rect 470676 390865 470698 390895
rect 470698 390865 470710 390895
rect 470710 390865 470732 390895
rect 470756 390865 470762 390895
rect 470762 390865 470774 390895
rect 470774 390865 470812 390895
rect 470276 390831 470332 390841
rect 470356 390831 470412 390841
rect 470436 390831 470492 390841
rect 470516 390831 470572 390841
rect 470596 390831 470652 390841
rect 470676 390831 470732 390841
rect 470756 390831 470812 390841
rect 470276 390785 470314 390831
rect 470314 390785 470326 390831
rect 470326 390785 470332 390831
rect 470356 390785 470378 390831
rect 470378 390785 470390 390831
rect 470390 390785 470412 390831
rect 470436 390785 470442 390831
rect 470442 390785 470454 390831
rect 470454 390785 470492 390831
rect 470516 390785 470518 390831
rect 470518 390785 470570 390831
rect 470570 390785 470572 390831
rect 470596 390785 470634 390831
rect 470634 390785 470646 390831
rect 470646 390785 470652 390831
rect 470676 390785 470698 390831
rect 470698 390785 470710 390831
rect 470710 390785 470732 390831
rect 470756 390785 470762 390831
rect 470762 390785 470774 390831
rect 470774 390785 470812 390831
rect 473726 410896 473782 410952
rect 478418 410080 478474 410136
rect 484122 410352 484178 410408
rect 481362 410080 481418 410136
rect 487802 410080 487858 410136
rect 481822 407088 481878 407144
rect 485134 407088 485190 407144
rect 488538 390088 488594 390144
rect 469036 389952 469074 389998
rect 469074 389952 469086 389998
rect 469086 389952 469092 389998
rect 469116 389952 469138 389998
rect 469138 389952 469150 389998
rect 469150 389952 469172 389998
rect 469196 389952 469202 389998
rect 469202 389952 469214 389998
rect 469214 389952 469252 389998
rect 469276 389952 469278 389998
rect 469278 389952 469330 389998
rect 469330 389952 469332 389998
rect 469356 389952 469394 389998
rect 469394 389952 469406 389998
rect 469406 389952 469412 389998
rect 469436 389952 469458 389998
rect 469458 389952 469470 389998
rect 469470 389952 469492 389998
rect 469516 389952 469522 389998
rect 469522 389952 469534 389998
rect 469534 389952 469572 389998
rect 469036 389942 469092 389952
rect 469116 389942 469172 389952
rect 469196 389942 469252 389952
rect 469276 389942 469332 389952
rect 469356 389942 469412 389952
rect 469436 389942 469492 389952
rect 469516 389942 469572 389952
rect 469036 389888 469074 389918
rect 469074 389888 469086 389918
rect 469086 389888 469092 389918
rect 469116 389888 469138 389918
rect 469138 389888 469150 389918
rect 469150 389888 469172 389918
rect 469196 389888 469202 389918
rect 469202 389888 469214 389918
rect 469214 389888 469252 389918
rect 469276 389888 469278 389918
rect 469278 389888 469330 389918
rect 469330 389888 469332 389918
rect 469356 389888 469394 389918
rect 469394 389888 469406 389918
rect 469406 389888 469412 389918
rect 469436 389888 469458 389918
rect 469458 389888 469470 389918
rect 469470 389888 469492 389918
rect 469516 389888 469522 389918
rect 469522 389888 469534 389918
rect 469534 389888 469572 389918
rect 469036 389876 469092 389888
rect 469116 389876 469172 389888
rect 469196 389876 469252 389888
rect 469276 389876 469332 389888
rect 469356 389876 469412 389888
rect 469436 389876 469492 389888
rect 469516 389876 469572 389888
rect 469036 389862 469074 389876
rect 469074 389862 469086 389876
rect 469086 389862 469092 389876
rect 469116 389862 469138 389876
rect 469138 389862 469150 389876
rect 469150 389862 469172 389876
rect 469196 389862 469202 389876
rect 469202 389862 469214 389876
rect 469214 389862 469252 389876
rect 469276 389862 469278 389876
rect 469278 389862 469330 389876
rect 469330 389862 469332 389876
rect 469356 389862 469394 389876
rect 469394 389862 469406 389876
rect 469406 389862 469412 389876
rect 469436 389862 469458 389876
rect 469458 389862 469470 389876
rect 469470 389862 469492 389876
rect 469516 389862 469522 389876
rect 469522 389862 469534 389876
rect 469534 389862 469572 389876
rect 469036 389824 469074 389838
rect 469074 389824 469086 389838
rect 469086 389824 469092 389838
rect 469116 389824 469138 389838
rect 469138 389824 469150 389838
rect 469150 389824 469172 389838
rect 469196 389824 469202 389838
rect 469202 389824 469214 389838
rect 469214 389824 469252 389838
rect 469276 389824 469278 389838
rect 469278 389824 469330 389838
rect 469330 389824 469332 389838
rect 469356 389824 469394 389838
rect 469394 389824 469406 389838
rect 469406 389824 469412 389838
rect 469436 389824 469458 389838
rect 469458 389824 469470 389838
rect 469470 389824 469492 389838
rect 469516 389824 469522 389838
rect 469522 389824 469534 389838
rect 469534 389824 469572 389838
rect 469036 389812 469092 389824
rect 469116 389812 469172 389824
rect 469196 389812 469252 389824
rect 469276 389812 469332 389824
rect 469356 389812 469412 389824
rect 469436 389812 469492 389824
rect 469516 389812 469572 389824
rect 469036 389782 469074 389812
rect 469074 389782 469086 389812
rect 469086 389782 469092 389812
rect 469116 389782 469138 389812
rect 469138 389782 469150 389812
rect 469150 389782 469172 389812
rect 469196 389782 469202 389812
rect 469202 389782 469214 389812
rect 469214 389782 469252 389812
rect 469276 389782 469278 389812
rect 469278 389782 469330 389812
rect 469330 389782 469332 389812
rect 469356 389782 469394 389812
rect 469394 389782 469406 389812
rect 469406 389782 469412 389812
rect 469436 389782 469458 389812
rect 469458 389782 469470 389812
rect 469470 389782 469492 389812
rect 469516 389782 469522 389812
rect 469522 389782 469534 389812
rect 469534 389782 469572 389812
rect 469036 389748 469092 389758
rect 469116 389748 469172 389758
rect 469196 389748 469252 389758
rect 469276 389748 469332 389758
rect 469356 389748 469412 389758
rect 469436 389748 469492 389758
rect 469516 389748 469572 389758
rect 469036 389702 469074 389748
rect 469074 389702 469086 389748
rect 469086 389702 469092 389748
rect 469116 389702 469138 389748
rect 469138 389702 469150 389748
rect 469150 389702 469172 389748
rect 469196 389702 469202 389748
rect 469202 389702 469214 389748
rect 469214 389702 469252 389748
rect 469276 389702 469278 389748
rect 469278 389702 469330 389748
rect 469330 389702 469332 389748
rect 469356 389702 469394 389748
rect 469394 389702 469406 389748
rect 469406 389702 469412 389748
rect 469436 389702 469458 389748
rect 469458 389702 469470 389748
rect 469470 389702 469492 389748
rect 469516 389702 469522 389748
rect 469522 389702 469534 389748
rect 469534 389702 469572 389748
rect 470276 388862 470314 388908
rect 470314 388862 470326 388908
rect 470326 388862 470332 388908
rect 470356 388862 470378 388908
rect 470378 388862 470390 388908
rect 470390 388862 470412 388908
rect 470436 388862 470442 388908
rect 470442 388862 470454 388908
rect 470454 388862 470492 388908
rect 470516 388862 470518 388908
rect 470518 388862 470570 388908
rect 470570 388862 470572 388908
rect 470596 388862 470634 388908
rect 470634 388862 470646 388908
rect 470646 388862 470652 388908
rect 470676 388862 470698 388908
rect 470698 388862 470710 388908
rect 470710 388862 470732 388908
rect 470756 388862 470762 388908
rect 470762 388862 470774 388908
rect 470774 388862 470812 388908
rect 470276 388852 470332 388862
rect 470356 388852 470412 388862
rect 470436 388852 470492 388862
rect 470516 388852 470572 388862
rect 470596 388852 470652 388862
rect 470676 388852 470732 388862
rect 470756 388852 470812 388862
rect 470276 388798 470314 388828
rect 470314 388798 470326 388828
rect 470326 388798 470332 388828
rect 470356 388798 470378 388828
rect 470378 388798 470390 388828
rect 470390 388798 470412 388828
rect 470436 388798 470442 388828
rect 470442 388798 470454 388828
rect 470454 388798 470492 388828
rect 470516 388798 470518 388828
rect 470518 388798 470570 388828
rect 470570 388798 470572 388828
rect 470596 388798 470634 388828
rect 470634 388798 470646 388828
rect 470646 388798 470652 388828
rect 470676 388798 470698 388828
rect 470698 388798 470710 388828
rect 470710 388798 470732 388828
rect 470756 388798 470762 388828
rect 470762 388798 470774 388828
rect 470774 388798 470812 388828
rect 470276 388786 470332 388798
rect 470356 388786 470412 388798
rect 470436 388786 470492 388798
rect 470516 388786 470572 388798
rect 470596 388786 470652 388798
rect 470676 388786 470732 388798
rect 470756 388786 470812 388798
rect 470276 388772 470314 388786
rect 470314 388772 470326 388786
rect 470326 388772 470332 388786
rect 470356 388772 470378 388786
rect 470378 388772 470390 388786
rect 470390 388772 470412 388786
rect 470436 388772 470442 388786
rect 470442 388772 470454 388786
rect 470454 388772 470492 388786
rect 470516 388772 470518 388786
rect 470518 388772 470570 388786
rect 470570 388772 470572 388786
rect 470596 388772 470634 388786
rect 470634 388772 470646 388786
rect 470646 388772 470652 388786
rect 470676 388772 470698 388786
rect 470698 388772 470710 388786
rect 470710 388772 470732 388786
rect 470756 388772 470762 388786
rect 470762 388772 470774 388786
rect 470774 388772 470812 388786
rect 470276 388734 470314 388748
rect 470314 388734 470326 388748
rect 470326 388734 470332 388748
rect 470356 388734 470378 388748
rect 470378 388734 470390 388748
rect 470390 388734 470412 388748
rect 470436 388734 470442 388748
rect 470442 388734 470454 388748
rect 470454 388734 470492 388748
rect 470516 388734 470518 388748
rect 470518 388734 470570 388748
rect 470570 388734 470572 388748
rect 470596 388734 470634 388748
rect 470634 388734 470646 388748
rect 470646 388734 470652 388748
rect 470676 388734 470698 388748
rect 470698 388734 470710 388748
rect 470710 388734 470732 388748
rect 470756 388734 470762 388748
rect 470762 388734 470774 388748
rect 470774 388734 470812 388748
rect 470276 388722 470332 388734
rect 470356 388722 470412 388734
rect 470436 388722 470492 388734
rect 470516 388722 470572 388734
rect 470596 388722 470652 388734
rect 470676 388722 470732 388734
rect 470756 388722 470812 388734
rect 470276 388692 470314 388722
rect 470314 388692 470326 388722
rect 470326 388692 470332 388722
rect 470356 388692 470378 388722
rect 470378 388692 470390 388722
rect 470390 388692 470412 388722
rect 470436 388692 470442 388722
rect 470442 388692 470454 388722
rect 470454 388692 470492 388722
rect 470516 388692 470518 388722
rect 470518 388692 470570 388722
rect 470570 388692 470572 388722
rect 470596 388692 470634 388722
rect 470634 388692 470646 388722
rect 470646 388692 470652 388722
rect 470676 388692 470698 388722
rect 470698 388692 470710 388722
rect 470710 388692 470732 388722
rect 470756 388692 470762 388722
rect 470762 388692 470774 388722
rect 470774 388692 470812 388722
rect 470276 388658 470332 388668
rect 470356 388658 470412 388668
rect 470436 388658 470492 388668
rect 470516 388658 470572 388668
rect 470596 388658 470652 388668
rect 470676 388658 470732 388668
rect 470756 388658 470812 388668
rect 470276 388612 470314 388658
rect 470314 388612 470326 388658
rect 470326 388612 470332 388658
rect 470356 388612 470378 388658
rect 470378 388612 470390 388658
rect 470390 388612 470412 388658
rect 470436 388612 470442 388658
rect 470442 388612 470454 388658
rect 470454 388612 470492 388658
rect 470516 388612 470518 388658
rect 470518 388612 470570 388658
rect 470570 388612 470572 388658
rect 470596 388612 470634 388658
rect 470634 388612 470646 388658
rect 470646 388612 470652 388658
rect 470676 388612 470698 388658
rect 470698 388612 470710 388658
rect 470710 388612 470732 388658
rect 470756 388612 470762 388658
rect 470762 388612 470774 388658
rect 470774 388612 470812 388658
rect 470276 358435 470314 358481
rect 470314 358435 470326 358481
rect 470326 358435 470332 358481
rect 470356 358435 470378 358481
rect 470378 358435 470390 358481
rect 470390 358435 470412 358481
rect 470436 358435 470442 358481
rect 470442 358435 470454 358481
rect 470454 358435 470492 358481
rect 470516 358435 470518 358481
rect 470518 358435 470570 358481
rect 470570 358435 470572 358481
rect 470596 358435 470634 358481
rect 470634 358435 470646 358481
rect 470646 358435 470652 358481
rect 470676 358435 470698 358481
rect 470698 358435 470710 358481
rect 470710 358435 470732 358481
rect 470756 358435 470762 358481
rect 470762 358435 470774 358481
rect 470774 358435 470812 358481
rect 470276 358425 470332 358435
rect 470356 358425 470412 358435
rect 470436 358425 470492 358435
rect 470516 358425 470572 358435
rect 470596 358425 470652 358435
rect 470676 358425 470732 358435
rect 470756 358425 470812 358435
rect 470276 358371 470314 358401
rect 470314 358371 470326 358401
rect 470326 358371 470332 358401
rect 470356 358371 470378 358401
rect 470378 358371 470390 358401
rect 470390 358371 470412 358401
rect 470436 358371 470442 358401
rect 470442 358371 470454 358401
rect 470454 358371 470492 358401
rect 470516 358371 470518 358401
rect 470518 358371 470570 358401
rect 470570 358371 470572 358401
rect 470596 358371 470634 358401
rect 470634 358371 470646 358401
rect 470646 358371 470652 358401
rect 470676 358371 470698 358401
rect 470698 358371 470710 358401
rect 470710 358371 470732 358401
rect 470756 358371 470762 358401
rect 470762 358371 470774 358401
rect 470774 358371 470812 358401
rect 470276 358359 470332 358371
rect 470356 358359 470412 358371
rect 470436 358359 470492 358371
rect 470516 358359 470572 358371
rect 470596 358359 470652 358371
rect 470676 358359 470732 358371
rect 470756 358359 470812 358371
rect 470276 358345 470314 358359
rect 470314 358345 470326 358359
rect 470326 358345 470332 358359
rect 470356 358345 470378 358359
rect 470378 358345 470390 358359
rect 470390 358345 470412 358359
rect 470436 358345 470442 358359
rect 470442 358345 470454 358359
rect 470454 358345 470492 358359
rect 470516 358345 470518 358359
rect 470518 358345 470570 358359
rect 470570 358345 470572 358359
rect 470596 358345 470634 358359
rect 470634 358345 470646 358359
rect 470646 358345 470652 358359
rect 470676 358345 470698 358359
rect 470698 358345 470710 358359
rect 470710 358345 470732 358359
rect 470756 358345 470762 358359
rect 470762 358345 470774 358359
rect 470774 358345 470812 358359
rect 470276 358307 470314 358321
rect 470314 358307 470326 358321
rect 470326 358307 470332 358321
rect 470356 358307 470378 358321
rect 470378 358307 470390 358321
rect 470390 358307 470412 358321
rect 470436 358307 470442 358321
rect 470442 358307 470454 358321
rect 470454 358307 470492 358321
rect 470516 358307 470518 358321
rect 470518 358307 470570 358321
rect 470570 358307 470572 358321
rect 470596 358307 470634 358321
rect 470634 358307 470646 358321
rect 470646 358307 470652 358321
rect 470676 358307 470698 358321
rect 470698 358307 470710 358321
rect 470710 358307 470732 358321
rect 470756 358307 470762 358321
rect 470762 358307 470774 358321
rect 470774 358307 470812 358321
rect 470276 358295 470332 358307
rect 470356 358295 470412 358307
rect 470436 358295 470492 358307
rect 470516 358295 470572 358307
rect 470596 358295 470652 358307
rect 470676 358295 470732 358307
rect 470756 358295 470812 358307
rect 470276 358265 470314 358295
rect 470314 358265 470326 358295
rect 470326 358265 470332 358295
rect 470356 358265 470378 358295
rect 470378 358265 470390 358295
rect 470390 358265 470412 358295
rect 470436 358265 470442 358295
rect 470442 358265 470454 358295
rect 470454 358265 470492 358295
rect 470516 358265 470518 358295
rect 470518 358265 470570 358295
rect 470570 358265 470572 358295
rect 470596 358265 470634 358295
rect 470634 358265 470646 358295
rect 470646 358265 470652 358295
rect 470676 358265 470698 358295
rect 470698 358265 470710 358295
rect 470710 358265 470732 358295
rect 470756 358265 470762 358295
rect 470762 358265 470774 358295
rect 470774 358265 470812 358295
rect 470276 358231 470332 358241
rect 470356 358231 470412 358241
rect 470436 358231 470492 358241
rect 470516 358231 470572 358241
rect 470596 358231 470652 358241
rect 470676 358231 470732 358241
rect 470756 358231 470812 358241
rect 470276 358185 470314 358231
rect 470314 358185 470326 358231
rect 470326 358185 470332 358231
rect 470356 358185 470378 358231
rect 470378 358185 470390 358231
rect 470390 358185 470412 358231
rect 470436 358185 470442 358231
rect 470442 358185 470454 358231
rect 470454 358185 470492 358231
rect 470516 358185 470518 358231
rect 470518 358185 470570 358231
rect 470570 358185 470572 358231
rect 470596 358185 470634 358231
rect 470634 358185 470646 358231
rect 470646 358185 470652 358231
rect 470676 358185 470698 358231
rect 470698 358185 470710 358231
rect 470710 358185 470732 358231
rect 470756 358185 470762 358231
rect 470762 358185 470774 358231
rect 470774 358185 470812 358231
rect 474922 389272 474978 389328
rect 478634 389272 478690 389328
rect 482098 389408 482154 389464
rect 486882 386416 486938 386472
rect 478878 357992 478934 358048
rect 481822 357992 481878 358048
rect 484950 357992 485006 358048
rect 488354 357992 488410 358048
rect 469036 357349 469074 357395
rect 469074 357349 469086 357395
rect 469086 357349 469092 357395
rect 469116 357349 469138 357395
rect 469138 357349 469150 357395
rect 469150 357349 469172 357395
rect 469196 357349 469202 357395
rect 469202 357349 469214 357395
rect 469214 357349 469252 357395
rect 469276 357349 469278 357395
rect 469278 357349 469330 357395
rect 469330 357349 469332 357395
rect 469356 357349 469394 357395
rect 469394 357349 469406 357395
rect 469406 357349 469412 357395
rect 469436 357349 469458 357395
rect 469458 357349 469470 357395
rect 469470 357349 469492 357395
rect 469516 357349 469522 357395
rect 469522 357349 469534 357395
rect 469534 357349 469572 357395
rect 469036 357339 469092 357349
rect 469116 357339 469172 357349
rect 469196 357339 469252 357349
rect 469276 357339 469332 357349
rect 469356 357339 469412 357349
rect 469436 357339 469492 357349
rect 469516 357339 469572 357349
rect 469036 357285 469074 357315
rect 469074 357285 469086 357315
rect 469086 357285 469092 357315
rect 469116 357285 469138 357315
rect 469138 357285 469150 357315
rect 469150 357285 469172 357315
rect 469196 357285 469202 357315
rect 469202 357285 469214 357315
rect 469214 357285 469252 357315
rect 469276 357285 469278 357315
rect 469278 357285 469330 357315
rect 469330 357285 469332 357315
rect 469356 357285 469394 357315
rect 469394 357285 469406 357315
rect 469406 357285 469412 357315
rect 469436 357285 469458 357315
rect 469458 357285 469470 357315
rect 469470 357285 469492 357315
rect 469516 357285 469522 357315
rect 469522 357285 469534 357315
rect 469534 357285 469572 357315
rect 469036 357273 469092 357285
rect 469116 357273 469172 357285
rect 469196 357273 469252 357285
rect 469276 357273 469332 357285
rect 469356 357273 469412 357285
rect 469436 357273 469492 357285
rect 469516 357273 469572 357285
rect 469036 357259 469074 357273
rect 469074 357259 469086 357273
rect 469086 357259 469092 357273
rect 469116 357259 469138 357273
rect 469138 357259 469150 357273
rect 469150 357259 469172 357273
rect 469196 357259 469202 357273
rect 469202 357259 469214 357273
rect 469214 357259 469252 357273
rect 469276 357259 469278 357273
rect 469278 357259 469330 357273
rect 469330 357259 469332 357273
rect 469356 357259 469394 357273
rect 469394 357259 469406 357273
rect 469406 357259 469412 357273
rect 469436 357259 469458 357273
rect 469458 357259 469470 357273
rect 469470 357259 469492 357273
rect 469516 357259 469522 357273
rect 469522 357259 469534 357273
rect 469534 357259 469572 357273
rect 469036 357221 469074 357235
rect 469074 357221 469086 357235
rect 469086 357221 469092 357235
rect 469116 357221 469138 357235
rect 469138 357221 469150 357235
rect 469150 357221 469172 357235
rect 469196 357221 469202 357235
rect 469202 357221 469214 357235
rect 469214 357221 469252 357235
rect 469276 357221 469278 357235
rect 469278 357221 469330 357235
rect 469330 357221 469332 357235
rect 469356 357221 469394 357235
rect 469394 357221 469406 357235
rect 469406 357221 469412 357235
rect 469436 357221 469458 357235
rect 469458 357221 469470 357235
rect 469470 357221 469492 357235
rect 469516 357221 469522 357235
rect 469522 357221 469534 357235
rect 469534 357221 469572 357235
rect 469036 357209 469092 357221
rect 469116 357209 469172 357221
rect 469196 357209 469252 357221
rect 469276 357209 469332 357221
rect 469356 357209 469412 357221
rect 469436 357209 469492 357221
rect 469516 357209 469572 357221
rect 469036 357179 469074 357209
rect 469074 357179 469086 357209
rect 469086 357179 469092 357209
rect 469116 357179 469138 357209
rect 469138 357179 469150 357209
rect 469150 357179 469172 357209
rect 469196 357179 469202 357209
rect 469202 357179 469214 357209
rect 469214 357179 469252 357209
rect 469276 357179 469278 357209
rect 469278 357179 469330 357209
rect 469330 357179 469332 357209
rect 469356 357179 469394 357209
rect 469394 357179 469406 357209
rect 469406 357179 469412 357209
rect 469436 357179 469458 357209
rect 469458 357179 469470 357209
rect 469470 357179 469492 357209
rect 469516 357179 469522 357209
rect 469522 357179 469534 357209
rect 469534 357179 469572 357209
rect 469036 357145 469092 357155
rect 469116 357145 469172 357155
rect 469196 357145 469252 357155
rect 469276 357145 469332 357155
rect 469356 357145 469412 357155
rect 469436 357145 469492 357155
rect 469516 357145 469572 357155
rect 469036 357099 469074 357145
rect 469074 357099 469086 357145
rect 469086 357099 469092 357145
rect 469116 357099 469138 357145
rect 469138 357099 469150 357145
rect 469150 357099 469172 357145
rect 469196 357099 469202 357145
rect 469202 357099 469214 357145
rect 469214 357099 469252 357145
rect 469276 357099 469278 357145
rect 469278 357099 469330 357145
rect 469330 357099 469332 357145
rect 469356 357099 469394 357145
rect 469394 357099 469406 357145
rect 469406 357099 469412 357145
rect 469436 357099 469458 357145
rect 469458 357099 469470 357145
rect 469470 357099 469492 357145
rect 469516 357099 469522 357145
rect 469522 357099 469534 357145
rect 469534 357099 469572 357145
rect 470276 356262 470314 356308
rect 470314 356262 470326 356308
rect 470326 356262 470332 356308
rect 470356 356262 470378 356308
rect 470378 356262 470390 356308
rect 470390 356262 470412 356308
rect 470436 356262 470442 356308
rect 470442 356262 470454 356308
rect 470454 356262 470492 356308
rect 470516 356262 470518 356308
rect 470518 356262 470570 356308
rect 470570 356262 470572 356308
rect 470596 356262 470634 356308
rect 470634 356262 470646 356308
rect 470646 356262 470652 356308
rect 470676 356262 470698 356308
rect 470698 356262 470710 356308
rect 470710 356262 470732 356308
rect 470756 356262 470762 356308
rect 470762 356262 470774 356308
rect 470774 356262 470812 356308
rect 470276 356252 470332 356262
rect 470356 356252 470412 356262
rect 470436 356252 470492 356262
rect 470516 356252 470572 356262
rect 470596 356252 470652 356262
rect 470676 356252 470732 356262
rect 470756 356252 470812 356262
rect 470276 356198 470314 356228
rect 470314 356198 470326 356228
rect 470326 356198 470332 356228
rect 470356 356198 470378 356228
rect 470378 356198 470390 356228
rect 470390 356198 470412 356228
rect 470436 356198 470442 356228
rect 470442 356198 470454 356228
rect 470454 356198 470492 356228
rect 470516 356198 470518 356228
rect 470518 356198 470570 356228
rect 470570 356198 470572 356228
rect 470596 356198 470634 356228
rect 470634 356198 470646 356228
rect 470646 356198 470652 356228
rect 470676 356198 470698 356228
rect 470698 356198 470710 356228
rect 470710 356198 470732 356228
rect 470756 356198 470762 356228
rect 470762 356198 470774 356228
rect 470774 356198 470812 356228
rect 470276 356186 470332 356198
rect 470356 356186 470412 356198
rect 470436 356186 470492 356198
rect 470516 356186 470572 356198
rect 470596 356186 470652 356198
rect 470676 356186 470732 356198
rect 470756 356186 470812 356198
rect 470276 356172 470314 356186
rect 470314 356172 470326 356186
rect 470326 356172 470332 356186
rect 470356 356172 470378 356186
rect 470378 356172 470390 356186
rect 470390 356172 470412 356186
rect 470436 356172 470442 356186
rect 470442 356172 470454 356186
rect 470454 356172 470492 356186
rect 470516 356172 470518 356186
rect 470518 356172 470570 356186
rect 470570 356172 470572 356186
rect 470596 356172 470634 356186
rect 470634 356172 470646 356186
rect 470646 356172 470652 356186
rect 470676 356172 470698 356186
rect 470698 356172 470710 356186
rect 470710 356172 470732 356186
rect 470756 356172 470762 356186
rect 470762 356172 470774 356186
rect 470774 356172 470812 356186
rect 470276 356134 470314 356148
rect 470314 356134 470326 356148
rect 470326 356134 470332 356148
rect 470356 356134 470378 356148
rect 470378 356134 470390 356148
rect 470390 356134 470412 356148
rect 470436 356134 470442 356148
rect 470442 356134 470454 356148
rect 470454 356134 470492 356148
rect 470516 356134 470518 356148
rect 470518 356134 470570 356148
rect 470570 356134 470572 356148
rect 470596 356134 470634 356148
rect 470634 356134 470646 356148
rect 470646 356134 470652 356148
rect 470676 356134 470698 356148
rect 470698 356134 470710 356148
rect 470710 356134 470732 356148
rect 470756 356134 470762 356148
rect 470762 356134 470774 356148
rect 470774 356134 470812 356148
rect 470276 356122 470332 356134
rect 470356 356122 470412 356134
rect 470436 356122 470492 356134
rect 470516 356122 470572 356134
rect 470596 356122 470652 356134
rect 470676 356122 470732 356134
rect 470756 356122 470812 356134
rect 470276 356092 470314 356122
rect 470314 356092 470326 356122
rect 470326 356092 470332 356122
rect 470356 356092 470378 356122
rect 470378 356092 470390 356122
rect 470390 356092 470412 356122
rect 470436 356092 470442 356122
rect 470442 356092 470454 356122
rect 470454 356092 470492 356122
rect 470516 356092 470518 356122
rect 470518 356092 470570 356122
rect 470570 356092 470572 356122
rect 470596 356092 470634 356122
rect 470634 356092 470646 356122
rect 470646 356092 470652 356122
rect 470676 356092 470698 356122
rect 470698 356092 470710 356122
rect 470710 356092 470732 356122
rect 470756 356092 470762 356122
rect 470762 356092 470774 356122
rect 470774 356092 470812 356122
rect 470276 356058 470332 356068
rect 470356 356058 470412 356068
rect 470436 356058 470492 356068
rect 470516 356058 470572 356068
rect 470596 356058 470652 356068
rect 470676 356058 470732 356068
rect 470756 356058 470812 356068
rect 470276 356012 470314 356058
rect 470314 356012 470326 356058
rect 470326 356012 470332 356058
rect 470356 356012 470378 356058
rect 470378 356012 470390 356058
rect 470390 356012 470412 356058
rect 470436 356012 470442 356058
rect 470442 356012 470454 356058
rect 470454 356012 470492 356058
rect 470516 356012 470518 356058
rect 470518 356012 470570 356058
rect 470570 356012 470572 356058
rect 470596 356012 470634 356058
rect 470634 356012 470646 356058
rect 470646 356012 470652 356058
rect 470676 356012 470698 356058
rect 470698 356012 470710 356058
rect 470710 356012 470732 356058
rect 470756 356012 470762 356058
rect 470762 356012 470774 356058
rect 470774 356012 470812 356058
rect 475014 357448 475070 357504
rect 470276 342434 470314 342480
rect 470314 342434 470326 342480
rect 470326 342434 470332 342480
rect 470356 342434 470378 342480
rect 470378 342434 470390 342480
rect 470390 342434 470412 342480
rect 470436 342434 470442 342480
rect 470442 342434 470454 342480
rect 470454 342434 470492 342480
rect 470516 342434 470518 342480
rect 470518 342434 470570 342480
rect 470570 342434 470572 342480
rect 470596 342434 470634 342480
rect 470634 342434 470646 342480
rect 470646 342434 470652 342480
rect 470676 342434 470698 342480
rect 470698 342434 470710 342480
rect 470710 342434 470732 342480
rect 470756 342434 470762 342480
rect 470762 342434 470774 342480
rect 470774 342434 470812 342480
rect 470276 342424 470332 342434
rect 470356 342424 470412 342434
rect 470436 342424 470492 342434
rect 470516 342424 470572 342434
rect 470596 342424 470652 342434
rect 470676 342424 470732 342434
rect 470756 342424 470812 342434
rect 470276 342370 470314 342400
rect 470314 342370 470326 342400
rect 470326 342370 470332 342400
rect 470356 342370 470378 342400
rect 470378 342370 470390 342400
rect 470390 342370 470412 342400
rect 470436 342370 470442 342400
rect 470442 342370 470454 342400
rect 470454 342370 470492 342400
rect 470516 342370 470518 342400
rect 470518 342370 470570 342400
rect 470570 342370 470572 342400
rect 470596 342370 470634 342400
rect 470634 342370 470646 342400
rect 470646 342370 470652 342400
rect 470676 342370 470698 342400
rect 470698 342370 470710 342400
rect 470710 342370 470732 342400
rect 470756 342370 470762 342400
rect 470762 342370 470774 342400
rect 470774 342370 470812 342400
rect 470276 342358 470332 342370
rect 470356 342358 470412 342370
rect 470436 342358 470492 342370
rect 470516 342358 470572 342370
rect 470596 342358 470652 342370
rect 470676 342358 470732 342370
rect 470756 342358 470812 342370
rect 470276 342344 470314 342358
rect 470314 342344 470326 342358
rect 470326 342344 470332 342358
rect 470356 342344 470378 342358
rect 470378 342344 470390 342358
rect 470390 342344 470412 342358
rect 470436 342344 470442 342358
rect 470442 342344 470454 342358
rect 470454 342344 470492 342358
rect 470516 342344 470518 342358
rect 470518 342344 470570 342358
rect 470570 342344 470572 342358
rect 470596 342344 470634 342358
rect 470634 342344 470646 342358
rect 470646 342344 470652 342358
rect 470676 342344 470698 342358
rect 470698 342344 470710 342358
rect 470710 342344 470732 342358
rect 470756 342344 470762 342358
rect 470762 342344 470774 342358
rect 470774 342344 470812 342358
rect 470276 342306 470314 342320
rect 470314 342306 470326 342320
rect 470326 342306 470332 342320
rect 470356 342306 470378 342320
rect 470378 342306 470390 342320
rect 470390 342306 470412 342320
rect 470436 342306 470442 342320
rect 470442 342306 470454 342320
rect 470454 342306 470492 342320
rect 470516 342306 470518 342320
rect 470518 342306 470570 342320
rect 470570 342306 470572 342320
rect 470596 342306 470634 342320
rect 470634 342306 470646 342320
rect 470646 342306 470652 342320
rect 470676 342306 470698 342320
rect 470698 342306 470710 342320
rect 470710 342306 470732 342320
rect 470756 342306 470762 342320
rect 470762 342306 470774 342320
rect 470774 342306 470812 342320
rect 470276 342294 470332 342306
rect 470356 342294 470412 342306
rect 470436 342294 470492 342306
rect 470516 342294 470572 342306
rect 470596 342294 470652 342306
rect 470676 342294 470732 342306
rect 470756 342294 470812 342306
rect 470276 342264 470314 342294
rect 470314 342264 470326 342294
rect 470326 342264 470332 342294
rect 470356 342264 470378 342294
rect 470378 342264 470390 342294
rect 470390 342264 470412 342294
rect 470436 342264 470442 342294
rect 470442 342264 470454 342294
rect 470454 342264 470492 342294
rect 470516 342264 470518 342294
rect 470518 342264 470570 342294
rect 470570 342264 470572 342294
rect 470596 342264 470634 342294
rect 470634 342264 470646 342294
rect 470646 342264 470652 342294
rect 470676 342264 470698 342294
rect 470698 342264 470710 342294
rect 470710 342264 470732 342294
rect 470756 342264 470762 342294
rect 470762 342264 470774 342294
rect 470774 342264 470812 342294
rect 470276 342230 470332 342240
rect 470356 342230 470412 342240
rect 470436 342230 470492 342240
rect 470516 342230 470572 342240
rect 470596 342230 470652 342240
rect 470676 342230 470732 342240
rect 470756 342230 470812 342240
rect 470276 342184 470314 342230
rect 470314 342184 470326 342230
rect 470326 342184 470332 342230
rect 470356 342184 470378 342230
rect 470378 342184 470390 342230
rect 470390 342184 470412 342230
rect 470436 342184 470442 342230
rect 470442 342184 470454 342230
rect 470454 342184 470492 342230
rect 470516 342184 470518 342230
rect 470518 342184 470570 342230
rect 470570 342184 470572 342230
rect 470596 342184 470634 342230
rect 470634 342184 470646 342230
rect 470646 342184 470652 342230
rect 470676 342184 470698 342230
rect 470698 342184 470710 342230
rect 470710 342184 470732 342230
rect 470756 342184 470762 342230
rect 470762 342184 470774 342230
rect 470774 342184 470812 342230
rect 469036 341347 469074 341393
rect 469074 341347 469086 341393
rect 469086 341347 469092 341393
rect 469116 341347 469138 341393
rect 469138 341347 469150 341393
rect 469150 341347 469172 341393
rect 469196 341347 469202 341393
rect 469202 341347 469214 341393
rect 469214 341347 469252 341393
rect 469276 341347 469278 341393
rect 469278 341347 469330 341393
rect 469330 341347 469332 341393
rect 469356 341347 469394 341393
rect 469394 341347 469406 341393
rect 469406 341347 469412 341393
rect 469436 341347 469458 341393
rect 469458 341347 469470 341393
rect 469470 341347 469492 341393
rect 469516 341347 469522 341393
rect 469522 341347 469534 341393
rect 469534 341347 469572 341393
rect 469036 341337 469092 341347
rect 469116 341337 469172 341347
rect 469196 341337 469252 341347
rect 469276 341337 469332 341347
rect 469356 341337 469412 341347
rect 469436 341337 469492 341347
rect 469516 341337 469572 341347
rect 469036 341283 469074 341313
rect 469074 341283 469086 341313
rect 469086 341283 469092 341313
rect 469116 341283 469138 341313
rect 469138 341283 469150 341313
rect 469150 341283 469172 341313
rect 469196 341283 469202 341313
rect 469202 341283 469214 341313
rect 469214 341283 469252 341313
rect 469276 341283 469278 341313
rect 469278 341283 469330 341313
rect 469330 341283 469332 341313
rect 469356 341283 469394 341313
rect 469394 341283 469406 341313
rect 469406 341283 469412 341313
rect 469436 341283 469458 341313
rect 469458 341283 469470 341313
rect 469470 341283 469492 341313
rect 469516 341283 469522 341313
rect 469522 341283 469534 341313
rect 469534 341283 469572 341313
rect 469036 341271 469092 341283
rect 469116 341271 469172 341283
rect 469196 341271 469252 341283
rect 469276 341271 469332 341283
rect 469356 341271 469412 341283
rect 469436 341271 469492 341283
rect 469516 341271 469572 341283
rect 469036 341257 469074 341271
rect 469074 341257 469086 341271
rect 469086 341257 469092 341271
rect 469116 341257 469138 341271
rect 469138 341257 469150 341271
rect 469150 341257 469172 341271
rect 469196 341257 469202 341271
rect 469202 341257 469214 341271
rect 469214 341257 469252 341271
rect 469276 341257 469278 341271
rect 469278 341257 469330 341271
rect 469330 341257 469332 341271
rect 469356 341257 469394 341271
rect 469394 341257 469406 341271
rect 469406 341257 469412 341271
rect 469436 341257 469458 341271
rect 469458 341257 469470 341271
rect 469470 341257 469492 341271
rect 469516 341257 469522 341271
rect 469522 341257 469534 341271
rect 469534 341257 469572 341271
rect 469036 341219 469074 341233
rect 469074 341219 469086 341233
rect 469086 341219 469092 341233
rect 469116 341219 469138 341233
rect 469138 341219 469150 341233
rect 469150 341219 469172 341233
rect 469196 341219 469202 341233
rect 469202 341219 469214 341233
rect 469214 341219 469252 341233
rect 469276 341219 469278 341233
rect 469278 341219 469330 341233
rect 469330 341219 469332 341233
rect 469356 341219 469394 341233
rect 469394 341219 469406 341233
rect 469406 341219 469412 341233
rect 469436 341219 469458 341233
rect 469458 341219 469470 341233
rect 469470 341219 469492 341233
rect 469516 341219 469522 341233
rect 469522 341219 469534 341233
rect 469534 341219 469572 341233
rect 469036 341207 469092 341219
rect 469116 341207 469172 341219
rect 469196 341207 469252 341219
rect 469276 341207 469332 341219
rect 469356 341207 469412 341219
rect 469436 341207 469492 341219
rect 469516 341207 469572 341219
rect 469036 341177 469074 341207
rect 469074 341177 469086 341207
rect 469086 341177 469092 341207
rect 469116 341177 469138 341207
rect 469138 341177 469150 341207
rect 469150 341177 469172 341207
rect 469196 341177 469202 341207
rect 469202 341177 469214 341207
rect 469214 341177 469252 341207
rect 469276 341177 469278 341207
rect 469278 341177 469330 341207
rect 469330 341177 469332 341207
rect 469356 341177 469394 341207
rect 469394 341177 469406 341207
rect 469406 341177 469412 341207
rect 469436 341177 469458 341207
rect 469458 341177 469470 341207
rect 469470 341177 469492 341207
rect 469516 341177 469522 341207
rect 469522 341177 469534 341207
rect 469534 341177 469572 341207
rect 469036 341143 469092 341153
rect 469116 341143 469172 341153
rect 469196 341143 469252 341153
rect 469276 341143 469332 341153
rect 469356 341143 469412 341153
rect 469436 341143 469492 341153
rect 469516 341143 469572 341153
rect 469036 341097 469074 341143
rect 469074 341097 469086 341143
rect 469086 341097 469092 341143
rect 469116 341097 469138 341143
rect 469138 341097 469150 341143
rect 469150 341097 469172 341143
rect 469196 341097 469202 341143
rect 469202 341097 469214 341143
rect 469214 341097 469252 341143
rect 469276 341097 469278 341143
rect 469278 341097 469330 341143
rect 469330 341097 469332 341143
rect 469356 341097 469394 341143
rect 469394 341097 469406 341143
rect 469406 341097 469412 341143
rect 469436 341097 469458 341143
rect 469458 341097 469470 341143
rect 469470 341097 469492 341143
rect 469516 341097 469522 341143
rect 469522 341097 469534 341143
rect 469534 341097 469572 341143
rect 470276 340262 470314 340308
rect 470314 340262 470326 340308
rect 470326 340262 470332 340308
rect 470356 340262 470378 340308
rect 470378 340262 470390 340308
rect 470390 340262 470412 340308
rect 470436 340262 470442 340308
rect 470442 340262 470454 340308
rect 470454 340262 470492 340308
rect 470516 340262 470518 340308
rect 470518 340262 470570 340308
rect 470570 340262 470572 340308
rect 470596 340262 470634 340308
rect 470634 340262 470646 340308
rect 470646 340262 470652 340308
rect 470676 340262 470698 340308
rect 470698 340262 470710 340308
rect 470710 340262 470732 340308
rect 470756 340262 470762 340308
rect 470762 340262 470774 340308
rect 470774 340262 470812 340308
rect 470276 340252 470332 340262
rect 470356 340252 470412 340262
rect 470436 340252 470492 340262
rect 470516 340252 470572 340262
rect 470596 340252 470652 340262
rect 470676 340252 470732 340262
rect 470756 340252 470812 340262
rect 470276 340198 470314 340228
rect 470314 340198 470326 340228
rect 470326 340198 470332 340228
rect 470356 340198 470378 340228
rect 470378 340198 470390 340228
rect 470390 340198 470412 340228
rect 470436 340198 470442 340228
rect 470442 340198 470454 340228
rect 470454 340198 470492 340228
rect 470516 340198 470518 340228
rect 470518 340198 470570 340228
rect 470570 340198 470572 340228
rect 470596 340198 470634 340228
rect 470634 340198 470646 340228
rect 470646 340198 470652 340228
rect 470676 340198 470698 340228
rect 470698 340198 470710 340228
rect 470710 340198 470732 340228
rect 470756 340198 470762 340228
rect 470762 340198 470774 340228
rect 470774 340198 470812 340228
rect 470276 340186 470332 340198
rect 470356 340186 470412 340198
rect 470436 340186 470492 340198
rect 470516 340186 470572 340198
rect 470596 340186 470652 340198
rect 470676 340186 470732 340198
rect 470756 340186 470812 340198
rect 470276 340172 470314 340186
rect 470314 340172 470326 340186
rect 470326 340172 470332 340186
rect 470356 340172 470378 340186
rect 470378 340172 470390 340186
rect 470390 340172 470412 340186
rect 470436 340172 470442 340186
rect 470442 340172 470454 340186
rect 470454 340172 470492 340186
rect 470516 340172 470518 340186
rect 470518 340172 470570 340186
rect 470570 340172 470572 340186
rect 470596 340172 470634 340186
rect 470634 340172 470646 340186
rect 470646 340172 470652 340186
rect 470676 340172 470698 340186
rect 470698 340172 470710 340186
rect 470710 340172 470732 340186
rect 470756 340172 470762 340186
rect 470762 340172 470774 340186
rect 470774 340172 470812 340186
rect 470276 340134 470314 340148
rect 470314 340134 470326 340148
rect 470326 340134 470332 340148
rect 470356 340134 470378 340148
rect 470378 340134 470390 340148
rect 470390 340134 470412 340148
rect 470436 340134 470442 340148
rect 470442 340134 470454 340148
rect 470454 340134 470492 340148
rect 470516 340134 470518 340148
rect 470518 340134 470570 340148
rect 470570 340134 470572 340148
rect 470596 340134 470634 340148
rect 470634 340134 470646 340148
rect 470646 340134 470652 340148
rect 470676 340134 470698 340148
rect 470698 340134 470710 340148
rect 470710 340134 470732 340148
rect 470756 340134 470762 340148
rect 470762 340134 470774 340148
rect 470774 340134 470812 340148
rect 470276 340122 470332 340134
rect 470356 340122 470412 340134
rect 470436 340122 470492 340134
rect 470516 340122 470572 340134
rect 470596 340122 470652 340134
rect 470676 340122 470732 340134
rect 470756 340122 470812 340134
rect 470276 340092 470314 340122
rect 470314 340092 470326 340122
rect 470326 340092 470332 340122
rect 470356 340092 470378 340122
rect 470378 340092 470390 340122
rect 470390 340092 470412 340122
rect 470436 340092 470442 340122
rect 470442 340092 470454 340122
rect 470454 340092 470492 340122
rect 470516 340092 470518 340122
rect 470518 340092 470570 340122
rect 470570 340092 470572 340122
rect 470596 340092 470634 340122
rect 470634 340092 470646 340122
rect 470646 340092 470652 340122
rect 470676 340092 470698 340122
rect 470698 340092 470710 340122
rect 470710 340092 470732 340122
rect 470756 340092 470762 340122
rect 470762 340092 470774 340122
rect 470774 340092 470812 340122
rect 470276 340058 470332 340068
rect 470356 340058 470412 340068
rect 470436 340058 470492 340068
rect 470516 340058 470572 340068
rect 470596 340058 470652 340068
rect 470676 340058 470732 340068
rect 470756 340058 470812 340068
rect 470276 340012 470314 340058
rect 470314 340012 470326 340058
rect 470326 340012 470332 340058
rect 470356 340012 470378 340058
rect 470378 340012 470390 340058
rect 470390 340012 470412 340058
rect 470436 340012 470442 340058
rect 470442 340012 470454 340058
rect 470454 340012 470492 340058
rect 470516 340012 470518 340058
rect 470518 340012 470570 340058
rect 470570 340012 470572 340058
rect 470596 340012 470634 340058
rect 470634 340012 470646 340058
rect 470646 340012 470652 340058
rect 470676 340012 470698 340058
rect 470698 340012 470710 340058
rect 470710 340012 470732 340058
rect 470756 340012 470762 340058
rect 470762 340012 470774 340058
rect 470774 340012 470812 340058
rect 470276 322434 470314 322480
rect 470314 322434 470326 322480
rect 470326 322434 470332 322480
rect 470356 322434 470378 322480
rect 470378 322434 470390 322480
rect 470390 322434 470412 322480
rect 470436 322434 470442 322480
rect 470442 322434 470454 322480
rect 470454 322434 470492 322480
rect 470516 322434 470518 322480
rect 470518 322434 470570 322480
rect 470570 322434 470572 322480
rect 470596 322434 470634 322480
rect 470634 322434 470646 322480
rect 470646 322434 470652 322480
rect 470676 322434 470698 322480
rect 470698 322434 470710 322480
rect 470710 322434 470732 322480
rect 470756 322434 470762 322480
rect 470762 322434 470774 322480
rect 470774 322434 470812 322480
rect 470276 322424 470332 322434
rect 470356 322424 470412 322434
rect 470436 322424 470492 322434
rect 470516 322424 470572 322434
rect 470596 322424 470652 322434
rect 470676 322424 470732 322434
rect 470756 322424 470812 322434
rect 470276 322370 470314 322400
rect 470314 322370 470326 322400
rect 470326 322370 470332 322400
rect 470356 322370 470378 322400
rect 470378 322370 470390 322400
rect 470390 322370 470412 322400
rect 470436 322370 470442 322400
rect 470442 322370 470454 322400
rect 470454 322370 470492 322400
rect 470516 322370 470518 322400
rect 470518 322370 470570 322400
rect 470570 322370 470572 322400
rect 470596 322370 470634 322400
rect 470634 322370 470646 322400
rect 470646 322370 470652 322400
rect 470676 322370 470698 322400
rect 470698 322370 470710 322400
rect 470710 322370 470732 322400
rect 470756 322370 470762 322400
rect 470762 322370 470774 322400
rect 470774 322370 470812 322400
rect 470276 322358 470332 322370
rect 470356 322358 470412 322370
rect 470436 322358 470492 322370
rect 470516 322358 470572 322370
rect 470596 322358 470652 322370
rect 470676 322358 470732 322370
rect 470756 322358 470812 322370
rect 470276 322344 470314 322358
rect 470314 322344 470326 322358
rect 470326 322344 470332 322358
rect 470356 322344 470378 322358
rect 470378 322344 470390 322358
rect 470390 322344 470412 322358
rect 470436 322344 470442 322358
rect 470442 322344 470454 322358
rect 470454 322344 470492 322358
rect 470516 322344 470518 322358
rect 470518 322344 470570 322358
rect 470570 322344 470572 322358
rect 470596 322344 470634 322358
rect 470634 322344 470646 322358
rect 470646 322344 470652 322358
rect 470676 322344 470698 322358
rect 470698 322344 470710 322358
rect 470710 322344 470732 322358
rect 470756 322344 470762 322358
rect 470762 322344 470774 322358
rect 470774 322344 470812 322358
rect 470276 322306 470314 322320
rect 470314 322306 470326 322320
rect 470326 322306 470332 322320
rect 470356 322306 470378 322320
rect 470378 322306 470390 322320
rect 470390 322306 470412 322320
rect 470436 322306 470442 322320
rect 470442 322306 470454 322320
rect 470454 322306 470492 322320
rect 470516 322306 470518 322320
rect 470518 322306 470570 322320
rect 470570 322306 470572 322320
rect 470596 322306 470634 322320
rect 470634 322306 470646 322320
rect 470646 322306 470652 322320
rect 470676 322306 470698 322320
rect 470698 322306 470710 322320
rect 470710 322306 470732 322320
rect 470756 322306 470762 322320
rect 470762 322306 470774 322320
rect 470774 322306 470812 322320
rect 470276 322294 470332 322306
rect 470356 322294 470412 322306
rect 470436 322294 470492 322306
rect 470516 322294 470572 322306
rect 470596 322294 470652 322306
rect 470676 322294 470732 322306
rect 470756 322294 470812 322306
rect 470276 322264 470314 322294
rect 470314 322264 470326 322294
rect 470326 322264 470332 322294
rect 470356 322264 470378 322294
rect 470378 322264 470390 322294
rect 470390 322264 470412 322294
rect 470436 322264 470442 322294
rect 470442 322264 470454 322294
rect 470454 322264 470492 322294
rect 470516 322264 470518 322294
rect 470518 322264 470570 322294
rect 470570 322264 470572 322294
rect 470596 322264 470634 322294
rect 470634 322264 470646 322294
rect 470646 322264 470652 322294
rect 470676 322264 470698 322294
rect 470698 322264 470710 322294
rect 470710 322264 470732 322294
rect 470756 322264 470762 322294
rect 470762 322264 470774 322294
rect 470774 322264 470812 322294
rect 470276 322230 470332 322240
rect 470356 322230 470412 322240
rect 470436 322230 470492 322240
rect 470516 322230 470572 322240
rect 470596 322230 470652 322240
rect 470676 322230 470732 322240
rect 470756 322230 470812 322240
rect 470276 322184 470314 322230
rect 470314 322184 470326 322230
rect 470326 322184 470332 322230
rect 470356 322184 470378 322230
rect 470378 322184 470390 322230
rect 470390 322184 470412 322230
rect 470436 322184 470442 322230
rect 470442 322184 470454 322230
rect 470454 322184 470492 322230
rect 470516 322184 470518 322230
rect 470518 322184 470570 322230
rect 470570 322184 470572 322230
rect 470596 322184 470634 322230
rect 470634 322184 470646 322230
rect 470646 322184 470652 322230
rect 470676 322184 470698 322230
rect 470698 322184 470710 322230
rect 470710 322184 470732 322230
rect 470756 322184 470762 322230
rect 470762 322184 470774 322230
rect 470774 322184 470812 322230
rect 477915 340992 477971 341048
rect 481232 340992 481288 341048
rect 484398 340992 484454 341048
rect 487894 340992 487950 341048
rect 474554 340448 474610 340504
rect 469036 321347 469074 321393
rect 469074 321347 469086 321393
rect 469086 321347 469092 321393
rect 469116 321347 469138 321393
rect 469138 321347 469150 321393
rect 469150 321347 469172 321393
rect 469196 321347 469202 321393
rect 469202 321347 469214 321393
rect 469214 321347 469252 321393
rect 469276 321347 469278 321393
rect 469278 321347 469330 321393
rect 469330 321347 469332 321393
rect 469356 321347 469394 321393
rect 469394 321347 469406 321393
rect 469406 321347 469412 321393
rect 469436 321347 469458 321393
rect 469458 321347 469470 321393
rect 469470 321347 469492 321393
rect 469516 321347 469522 321393
rect 469522 321347 469534 321393
rect 469534 321347 469572 321393
rect 469036 321337 469092 321347
rect 469116 321337 469172 321347
rect 469196 321337 469252 321347
rect 469276 321337 469332 321347
rect 469356 321337 469412 321347
rect 469436 321337 469492 321347
rect 469516 321337 469572 321347
rect 469036 321283 469074 321313
rect 469074 321283 469086 321313
rect 469086 321283 469092 321313
rect 469116 321283 469138 321313
rect 469138 321283 469150 321313
rect 469150 321283 469172 321313
rect 469196 321283 469202 321313
rect 469202 321283 469214 321313
rect 469214 321283 469252 321313
rect 469276 321283 469278 321313
rect 469278 321283 469330 321313
rect 469330 321283 469332 321313
rect 469356 321283 469394 321313
rect 469394 321283 469406 321313
rect 469406 321283 469412 321313
rect 469436 321283 469458 321313
rect 469458 321283 469470 321313
rect 469470 321283 469492 321313
rect 469516 321283 469522 321313
rect 469522 321283 469534 321313
rect 469534 321283 469572 321313
rect 469036 321271 469092 321283
rect 469116 321271 469172 321283
rect 469196 321271 469252 321283
rect 469276 321271 469332 321283
rect 469356 321271 469412 321283
rect 469436 321271 469492 321283
rect 469516 321271 469572 321283
rect 469036 321257 469074 321271
rect 469074 321257 469086 321271
rect 469086 321257 469092 321271
rect 469116 321257 469138 321271
rect 469138 321257 469150 321271
rect 469150 321257 469172 321271
rect 469196 321257 469202 321271
rect 469202 321257 469214 321271
rect 469214 321257 469252 321271
rect 469276 321257 469278 321271
rect 469278 321257 469330 321271
rect 469330 321257 469332 321271
rect 469356 321257 469394 321271
rect 469394 321257 469406 321271
rect 469406 321257 469412 321271
rect 469436 321257 469458 321271
rect 469458 321257 469470 321271
rect 469470 321257 469492 321271
rect 469516 321257 469522 321271
rect 469522 321257 469534 321271
rect 469534 321257 469572 321271
rect 469036 321219 469074 321233
rect 469074 321219 469086 321233
rect 469086 321219 469092 321233
rect 469116 321219 469138 321233
rect 469138 321219 469150 321233
rect 469150 321219 469172 321233
rect 469196 321219 469202 321233
rect 469202 321219 469214 321233
rect 469214 321219 469252 321233
rect 469276 321219 469278 321233
rect 469278 321219 469330 321233
rect 469330 321219 469332 321233
rect 469356 321219 469394 321233
rect 469394 321219 469406 321233
rect 469406 321219 469412 321233
rect 469436 321219 469458 321233
rect 469458 321219 469470 321233
rect 469470 321219 469492 321233
rect 469516 321219 469522 321233
rect 469522 321219 469534 321233
rect 469534 321219 469572 321233
rect 469036 321207 469092 321219
rect 469116 321207 469172 321219
rect 469196 321207 469252 321219
rect 469276 321207 469332 321219
rect 469356 321207 469412 321219
rect 469436 321207 469492 321219
rect 469516 321207 469572 321219
rect 469036 321177 469074 321207
rect 469074 321177 469086 321207
rect 469086 321177 469092 321207
rect 469116 321177 469138 321207
rect 469138 321177 469150 321207
rect 469150 321177 469172 321207
rect 469196 321177 469202 321207
rect 469202 321177 469214 321207
rect 469214 321177 469252 321207
rect 469276 321177 469278 321207
rect 469278 321177 469330 321207
rect 469330 321177 469332 321207
rect 469356 321177 469394 321207
rect 469394 321177 469406 321207
rect 469406 321177 469412 321207
rect 469436 321177 469458 321207
rect 469458 321177 469470 321207
rect 469470 321177 469492 321207
rect 469516 321177 469522 321207
rect 469522 321177 469534 321207
rect 469534 321177 469572 321207
rect 469036 321143 469092 321153
rect 469116 321143 469172 321153
rect 469196 321143 469252 321153
rect 469276 321143 469332 321153
rect 469356 321143 469412 321153
rect 469436 321143 469492 321153
rect 469516 321143 469572 321153
rect 469036 321097 469074 321143
rect 469074 321097 469086 321143
rect 469086 321097 469092 321143
rect 469116 321097 469138 321143
rect 469138 321097 469150 321143
rect 469150 321097 469172 321143
rect 469196 321097 469202 321143
rect 469202 321097 469214 321143
rect 469214 321097 469252 321143
rect 469276 321097 469278 321143
rect 469278 321097 469330 321143
rect 469330 321097 469332 321143
rect 469356 321097 469394 321143
rect 469394 321097 469406 321143
rect 469406 321097 469412 321143
rect 469436 321097 469458 321143
rect 469458 321097 469470 321143
rect 469470 321097 469492 321143
rect 469516 321097 469522 321143
rect 469522 321097 469534 321143
rect 469534 321097 469572 321143
rect 470276 320262 470314 320308
rect 470314 320262 470326 320308
rect 470326 320262 470332 320308
rect 470356 320262 470378 320308
rect 470378 320262 470390 320308
rect 470390 320262 470412 320308
rect 470436 320262 470442 320308
rect 470442 320262 470454 320308
rect 470454 320262 470492 320308
rect 470516 320262 470518 320308
rect 470518 320262 470570 320308
rect 470570 320262 470572 320308
rect 470596 320262 470634 320308
rect 470634 320262 470646 320308
rect 470646 320262 470652 320308
rect 470676 320262 470698 320308
rect 470698 320262 470710 320308
rect 470710 320262 470732 320308
rect 470756 320262 470762 320308
rect 470762 320262 470774 320308
rect 470774 320262 470812 320308
rect 470276 320252 470332 320262
rect 470356 320252 470412 320262
rect 470436 320252 470492 320262
rect 470516 320252 470572 320262
rect 470596 320252 470652 320262
rect 470676 320252 470732 320262
rect 470756 320252 470812 320262
rect 470276 320198 470314 320228
rect 470314 320198 470326 320228
rect 470326 320198 470332 320228
rect 470356 320198 470378 320228
rect 470378 320198 470390 320228
rect 470390 320198 470412 320228
rect 470436 320198 470442 320228
rect 470442 320198 470454 320228
rect 470454 320198 470492 320228
rect 470516 320198 470518 320228
rect 470518 320198 470570 320228
rect 470570 320198 470572 320228
rect 470596 320198 470634 320228
rect 470634 320198 470646 320228
rect 470646 320198 470652 320228
rect 470676 320198 470698 320228
rect 470698 320198 470710 320228
rect 470710 320198 470732 320228
rect 470756 320198 470762 320228
rect 470762 320198 470774 320228
rect 470774 320198 470812 320228
rect 470276 320186 470332 320198
rect 470356 320186 470412 320198
rect 470436 320186 470492 320198
rect 470516 320186 470572 320198
rect 470596 320186 470652 320198
rect 470676 320186 470732 320198
rect 470756 320186 470812 320198
rect 470276 320172 470314 320186
rect 470314 320172 470326 320186
rect 470326 320172 470332 320186
rect 470356 320172 470378 320186
rect 470378 320172 470390 320186
rect 470390 320172 470412 320186
rect 470436 320172 470442 320186
rect 470442 320172 470454 320186
rect 470454 320172 470492 320186
rect 470516 320172 470518 320186
rect 470518 320172 470570 320186
rect 470570 320172 470572 320186
rect 470596 320172 470634 320186
rect 470634 320172 470646 320186
rect 470646 320172 470652 320186
rect 470676 320172 470698 320186
rect 470698 320172 470710 320186
rect 470710 320172 470732 320186
rect 470756 320172 470762 320186
rect 470762 320172 470774 320186
rect 470774 320172 470812 320186
rect 470276 320134 470314 320148
rect 470314 320134 470326 320148
rect 470326 320134 470332 320148
rect 470356 320134 470378 320148
rect 470378 320134 470390 320148
rect 470390 320134 470412 320148
rect 470436 320134 470442 320148
rect 470442 320134 470454 320148
rect 470454 320134 470492 320148
rect 470516 320134 470518 320148
rect 470518 320134 470570 320148
rect 470570 320134 470572 320148
rect 470596 320134 470634 320148
rect 470634 320134 470646 320148
rect 470646 320134 470652 320148
rect 470676 320134 470698 320148
rect 470698 320134 470710 320148
rect 470710 320134 470732 320148
rect 470756 320134 470762 320148
rect 470762 320134 470774 320148
rect 470774 320134 470812 320148
rect 470276 320122 470332 320134
rect 470356 320122 470412 320134
rect 470436 320122 470492 320134
rect 470516 320122 470572 320134
rect 470596 320122 470652 320134
rect 470676 320122 470732 320134
rect 470756 320122 470812 320134
rect 470276 320092 470314 320122
rect 470314 320092 470326 320122
rect 470326 320092 470332 320122
rect 470356 320092 470378 320122
rect 470378 320092 470390 320122
rect 470390 320092 470412 320122
rect 470436 320092 470442 320122
rect 470442 320092 470454 320122
rect 470454 320092 470492 320122
rect 470516 320092 470518 320122
rect 470518 320092 470570 320122
rect 470570 320092 470572 320122
rect 470596 320092 470634 320122
rect 470634 320092 470646 320122
rect 470646 320092 470652 320122
rect 470676 320092 470698 320122
rect 470698 320092 470710 320122
rect 470710 320092 470732 320122
rect 470756 320092 470762 320122
rect 470762 320092 470774 320122
rect 470774 320092 470812 320122
rect 470276 320058 470332 320068
rect 470356 320058 470412 320068
rect 470436 320058 470492 320068
rect 470516 320058 470572 320068
rect 470596 320058 470652 320068
rect 470676 320058 470732 320068
rect 470756 320058 470812 320068
rect 470276 320012 470314 320058
rect 470314 320012 470326 320058
rect 470326 320012 470332 320058
rect 470356 320012 470378 320058
rect 470378 320012 470390 320058
rect 470390 320012 470412 320058
rect 470436 320012 470442 320058
rect 470442 320012 470454 320058
rect 470454 320012 470492 320058
rect 470516 320012 470518 320058
rect 470518 320012 470570 320058
rect 470570 320012 470572 320058
rect 470596 320012 470634 320058
rect 470634 320012 470646 320058
rect 470646 320012 470652 320058
rect 470676 320012 470698 320058
rect 470698 320012 470710 320058
rect 470710 320012 470732 320058
rect 470756 320012 470762 320058
rect 470762 320012 470774 320058
rect 470774 320012 470812 320058
rect 470276 307034 470314 307080
rect 470314 307034 470326 307080
rect 470326 307034 470332 307080
rect 470356 307034 470378 307080
rect 470378 307034 470390 307080
rect 470390 307034 470412 307080
rect 470436 307034 470442 307080
rect 470442 307034 470454 307080
rect 470454 307034 470492 307080
rect 470516 307034 470518 307080
rect 470518 307034 470570 307080
rect 470570 307034 470572 307080
rect 470596 307034 470634 307080
rect 470634 307034 470646 307080
rect 470646 307034 470652 307080
rect 470676 307034 470698 307080
rect 470698 307034 470710 307080
rect 470710 307034 470732 307080
rect 470756 307034 470762 307080
rect 470762 307034 470774 307080
rect 470774 307034 470812 307080
rect 470276 307024 470332 307034
rect 470356 307024 470412 307034
rect 470436 307024 470492 307034
rect 470516 307024 470572 307034
rect 470596 307024 470652 307034
rect 470676 307024 470732 307034
rect 470756 307024 470812 307034
rect 470276 306970 470314 307000
rect 470314 306970 470326 307000
rect 470326 306970 470332 307000
rect 470356 306970 470378 307000
rect 470378 306970 470390 307000
rect 470390 306970 470412 307000
rect 470436 306970 470442 307000
rect 470442 306970 470454 307000
rect 470454 306970 470492 307000
rect 470516 306970 470518 307000
rect 470518 306970 470570 307000
rect 470570 306970 470572 307000
rect 470596 306970 470634 307000
rect 470634 306970 470646 307000
rect 470646 306970 470652 307000
rect 470676 306970 470698 307000
rect 470698 306970 470710 307000
rect 470710 306970 470732 307000
rect 470756 306970 470762 307000
rect 470762 306970 470774 307000
rect 470774 306970 470812 307000
rect 470276 306958 470332 306970
rect 470356 306958 470412 306970
rect 470436 306958 470492 306970
rect 470516 306958 470572 306970
rect 470596 306958 470652 306970
rect 470676 306958 470732 306970
rect 470756 306958 470812 306970
rect 470276 306944 470314 306958
rect 470314 306944 470326 306958
rect 470326 306944 470332 306958
rect 470356 306944 470378 306958
rect 470378 306944 470390 306958
rect 470390 306944 470412 306958
rect 470436 306944 470442 306958
rect 470442 306944 470454 306958
rect 470454 306944 470492 306958
rect 470516 306944 470518 306958
rect 470518 306944 470570 306958
rect 470570 306944 470572 306958
rect 470596 306944 470634 306958
rect 470634 306944 470646 306958
rect 470646 306944 470652 306958
rect 470676 306944 470698 306958
rect 470698 306944 470710 306958
rect 470710 306944 470732 306958
rect 470756 306944 470762 306958
rect 470762 306944 470774 306958
rect 470774 306944 470812 306958
rect 470276 306906 470314 306920
rect 470314 306906 470326 306920
rect 470326 306906 470332 306920
rect 470356 306906 470378 306920
rect 470378 306906 470390 306920
rect 470390 306906 470412 306920
rect 470436 306906 470442 306920
rect 470442 306906 470454 306920
rect 470454 306906 470492 306920
rect 470516 306906 470518 306920
rect 470518 306906 470570 306920
rect 470570 306906 470572 306920
rect 470596 306906 470634 306920
rect 470634 306906 470646 306920
rect 470646 306906 470652 306920
rect 470676 306906 470698 306920
rect 470698 306906 470710 306920
rect 470710 306906 470732 306920
rect 470756 306906 470762 306920
rect 470762 306906 470774 306920
rect 470774 306906 470812 306920
rect 470276 306894 470332 306906
rect 470356 306894 470412 306906
rect 470436 306894 470492 306906
rect 470516 306894 470572 306906
rect 470596 306894 470652 306906
rect 470676 306894 470732 306906
rect 470756 306894 470812 306906
rect 470276 306864 470314 306894
rect 470314 306864 470326 306894
rect 470326 306864 470332 306894
rect 470356 306864 470378 306894
rect 470378 306864 470390 306894
rect 470390 306864 470412 306894
rect 470436 306864 470442 306894
rect 470442 306864 470454 306894
rect 470454 306864 470492 306894
rect 470516 306864 470518 306894
rect 470518 306864 470570 306894
rect 470570 306864 470572 306894
rect 470596 306864 470634 306894
rect 470634 306864 470646 306894
rect 470646 306864 470652 306894
rect 470676 306864 470698 306894
rect 470698 306864 470710 306894
rect 470710 306864 470732 306894
rect 470756 306864 470762 306894
rect 470762 306864 470774 306894
rect 470774 306864 470812 306894
rect 470276 306830 470332 306840
rect 470356 306830 470412 306840
rect 470436 306830 470492 306840
rect 470516 306830 470572 306840
rect 470596 306830 470652 306840
rect 470676 306830 470732 306840
rect 470756 306830 470812 306840
rect 470276 306784 470314 306830
rect 470314 306784 470326 306830
rect 470326 306784 470332 306830
rect 470356 306784 470378 306830
rect 470378 306784 470390 306830
rect 470390 306784 470412 306830
rect 470436 306784 470442 306830
rect 470442 306784 470454 306830
rect 470454 306784 470492 306830
rect 470516 306784 470518 306830
rect 470518 306784 470570 306830
rect 470570 306784 470572 306830
rect 470596 306784 470634 306830
rect 470634 306784 470646 306830
rect 470646 306784 470652 306830
rect 470676 306784 470698 306830
rect 470698 306784 470710 306830
rect 470710 306784 470732 306830
rect 470756 306784 470762 306830
rect 470762 306784 470774 306830
rect 470774 306784 470812 306830
rect 474278 321272 474334 321328
rect 484582 321272 484638 321328
rect 488170 321000 488226 321056
rect 478142 320864 478198 320920
rect 481546 320864 481602 320920
rect 469036 305949 469074 305995
rect 469074 305949 469086 305995
rect 469086 305949 469092 305995
rect 469116 305949 469138 305995
rect 469138 305949 469150 305995
rect 469150 305949 469172 305995
rect 469196 305949 469202 305995
rect 469202 305949 469214 305995
rect 469214 305949 469252 305995
rect 469276 305949 469278 305995
rect 469278 305949 469330 305995
rect 469330 305949 469332 305995
rect 469356 305949 469394 305995
rect 469394 305949 469406 305995
rect 469406 305949 469412 305995
rect 469436 305949 469458 305995
rect 469458 305949 469470 305995
rect 469470 305949 469492 305995
rect 469516 305949 469522 305995
rect 469522 305949 469534 305995
rect 469534 305949 469572 305995
rect 469036 305939 469092 305949
rect 469116 305939 469172 305949
rect 469196 305939 469252 305949
rect 469276 305939 469332 305949
rect 469356 305939 469412 305949
rect 469436 305939 469492 305949
rect 469516 305939 469572 305949
rect 469036 305885 469074 305915
rect 469074 305885 469086 305915
rect 469086 305885 469092 305915
rect 469116 305885 469138 305915
rect 469138 305885 469150 305915
rect 469150 305885 469172 305915
rect 469196 305885 469202 305915
rect 469202 305885 469214 305915
rect 469214 305885 469252 305915
rect 469276 305885 469278 305915
rect 469278 305885 469330 305915
rect 469330 305885 469332 305915
rect 469356 305885 469394 305915
rect 469394 305885 469406 305915
rect 469406 305885 469412 305915
rect 469436 305885 469458 305915
rect 469458 305885 469470 305915
rect 469470 305885 469492 305915
rect 469516 305885 469522 305915
rect 469522 305885 469534 305915
rect 469534 305885 469572 305915
rect 469036 305873 469092 305885
rect 469116 305873 469172 305885
rect 469196 305873 469252 305885
rect 469276 305873 469332 305885
rect 469356 305873 469412 305885
rect 469436 305873 469492 305885
rect 469516 305873 469572 305885
rect 469036 305859 469074 305873
rect 469074 305859 469086 305873
rect 469086 305859 469092 305873
rect 469116 305859 469138 305873
rect 469138 305859 469150 305873
rect 469150 305859 469172 305873
rect 469196 305859 469202 305873
rect 469202 305859 469214 305873
rect 469214 305859 469252 305873
rect 469276 305859 469278 305873
rect 469278 305859 469330 305873
rect 469330 305859 469332 305873
rect 469356 305859 469394 305873
rect 469394 305859 469406 305873
rect 469406 305859 469412 305873
rect 469436 305859 469458 305873
rect 469458 305859 469470 305873
rect 469470 305859 469492 305873
rect 469516 305859 469522 305873
rect 469522 305859 469534 305873
rect 469534 305859 469572 305873
rect 469036 305821 469074 305835
rect 469074 305821 469086 305835
rect 469086 305821 469092 305835
rect 469116 305821 469138 305835
rect 469138 305821 469150 305835
rect 469150 305821 469172 305835
rect 469196 305821 469202 305835
rect 469202 305821 469214 305835
rect 469214 305821 469252 305835
rect 469276 305821 469278 305835
rect 469278 305821 469330 305835
rect 469330 305821 469332 305835
rect 469356 305821 469394 305835
rect 469394 305821 469406 305835
rect 469406 305821 469412 305835
rect 469436 305821 469458 305835
rect 469458 305821 469470 305835
rect 469470 305821 469492 305835
rect 469516 305821 469522 305835
rect 469522 305821 469534 305835
rect 469534 305821 469572 305835
rect 469036 305809 469092 305821
rect 469116 305809 469172 305821
rect 469196 305809 469252 305821
rect 469276 305809 469332 305821
rect 469356 305809 469412 305821
rect 469436 305809 469492 305821
rect 469516 305809 469572 305821
rect 469036 305779 469074 305809
rect 469074 305779 469086 305809
rect 469086 305779 469092 305809
rect 469116 305779 469138 305809
rect 469138 305779 469150 305809
rect 469150 305779 469172 305809
rect 469196 305779 469202 305809
rect 469202 305779 469214 305809
rect 469214 305779 469252 305809
rect 469276 305779 469278 305809
rect 469278 305779 469330 305809
rect 469330 305779 469332 305809
rect 469356 305779 469394 305809
rect 469394 305779 469406 305809
rect 469406 305779 469412 305809
rect 469436 305779 469458 305809
rect 469458 305779 469470 305809
rect 469470 305779 469492 305809
rect 469516 305779 469522 305809
rect 469522 305779 469534 305809
rect 469534 305779 469572 305809
rect 469036 305745 469092 305755
rect 469116 305745 469172 305755
rect 469196 305745 469252 305755
rect 469276 305745 469332 305755
rect 469356 305745 469412 305755
rect 469436 305745 469492 305755
rect 469516 305745 469572 305755
rect 469036 305699 469074 305745
rect 469074 305699 469086 305745
rect 469086 305699 469092 305745
rect 469116 305699 469138 305745
rect 469138 305699 469150 305745
rect 469150 305699 469172 305745
rect 469196 305699 469202 305745
rect 469202 305699 469214 305745
rect 469214 305699 469252 305745
rect 469276 305699 469278 305745
rect 469278 305699 469330 305745
rect 469330 305699 469332 305745
rect 469356 305699 469394 305745
rect 469394 305699 469406 305745
rect 469406 305699 469412 305745
rect 469436 305699 469458 305745
rect 469458 305699 469470 305745
rect 469470 305699 469492 305745
rect 469516 305699 469522 305745
rect 469522 305699 469534 305745
rect 469534 305699 469572 305745
rect 470276 304862 470314 304908
rect 470314 304862 470326 304908
rect 470326 304862 470332 304908
rect 470356 304862 470378 304908
rect 470378 304862 470390 304908
rect 470390 304862 470412 304908
rect 470436 304862 470442 304908
rect 470442 304862 470454 304908
rect 470454 304862 470492 304908
rect 470516 304862 470518 304908
rect 470518 304862 470570 304908
rect 470570 304862 470572 304908
rect 470596 304862 470634 304908
rect 470634 304862 470646 304908
rect 470646 304862 470652 304908
rect 470676 304862 470698 304908
rect 470698 304862 470710 304908
rect 470710 304862 470732 304908
rect 470756 304862 470762 304908
rect 470762 304862 470774 304908
rect 470774 304862 470812 304908
rect 470276 304852 470332 304862
rect 470356 304852 470412 304862
rect 470436 304852 470492 304862
rect 470516 304852 470572 304862
rect 470596 304852 470652 304862
rect 470676 304852 470732 304862
rect 470756 304852 470812 304862
rect 470276 304798 470314 304828
rect 470314 304798 470326 304828
rect 470326 304798 470332 304828
rect 470356 304798 470378 304828
rect 470378 304798 470390 304828
rect 470390 304798 470412 304828
rect 470436 304798 470442 304828
rect 470442 304798 470454 304828
rect 470454 304798 470492 304828
rect 470516 304798 470518 304828
rect 470518 304798 470570 304828
rect 470570 304798 470572 304828
rect 470596 304798 470634 304828
rect 470634 304798 470646 304828
rect 470646 304798 470652 304828
rect 470676 304798 470698 304828
rect 470698 304798 470710 304828
rect 470710 304798 470732 304828
rect 470756 304798 470762 304828
rect 470762 304798 470774 304828
rect 470774 304798 470812 304828
rect 470276 304786 470332 304798
rect 470356 304786 470412 304798
rect 470436 304786 470492 304798
rect 470516 304786 470572 304798
rect 470596 304786 470652 304798
rect 470676 304786 470732 304798
rect 470756 304786 470812 304798
rect 470276 304772 470314 304786
rect 470314 304772 470326 304786
rect 470326 304772 470332 304786
rect 470356 304772 470378 304786
rect 470378 304772 470390 304786
rect 470390 304772 470412 304786
rect 470436 304772 470442 304786
rect 470442 304772 470454 304786
rect 470454 304772 470492 304786
rect 470516 304772 470518 304786
rect 470518 304772 470570 304786
rect 470570 304772 470572 304786
rect 470596 304772 470634 304786
rect 470634 304772 470646 304786
rect 470646 304772 470652 304786
rect 470676 304772 470698 304786
rect 470698 304772 470710 304786
rect 470710 304772 470732 304786
rect 470756 304772 470762 304786
rect 470762 304772 470774 304786
rect 470774 304772 470812 304786
rect 470276 304734 470314 304748
rect 470314 304734 470326 304748
rect 470326 304734 470332 304748
rect 470356 304734 470378 304748
rect 470378 304734 470390 304748
rect 470390 304734 470412 304748
rect 470436 304734 470442 304748
rect 470442 304734 470454 304748
rect 470454 304734 470492 304748
rect 470516 304734 470518 304748
rect 470518 304734 470570 304748
rect 470570 304734 470572 304748
rect 470596 304734 470634 304748
rect 470634 304734 470646 304748
rect 470646 304734 470652 304748
rect 470676 304734 470698 304748
rect 470698 304734 470710 304748
rect 470710 304734 470732 304748
rect 470756 304734 470762 304748
rect 470762 304734 470774 304748
rect 470774 304734 470812 304748
rect 470276 304722 470332 304734
rect 470356 304722 470412 304734
rect 470436 304722 470492 304734
rect 470516 304722 470572 304734
rect 470596 304722 470652 304734
rect 470676 304722 470732 304734
rect 470756 304722 470812 304734
rect 470276 304692 470314 304722
rect 470314 304692 470326 304722
rect 470326 304692 470332 304722
rect 470356 304692 470378 304722
rect 470378 304692 470390 304722
rect 470390 304692 470412 304722
rect 470436 304692 470442 304722
rect 470442 304692 470454 304722
rect 470454 304692 470492 304722
rect 470516 304692 470518 304722
rect 470518 304692 470570 304722
rect 470570 304692 470572 304722
rect 470596 304692 470634 304722
rect 470634 304692 470646 304722
rect 470646 304692 470652 304722
rect 470676 304692 470698 304722
rect 470698 304692 470710 304722
rect 470710 304692 470732 304722
rect 470756 304692 470762 304722
rect 470762 304692 470774 304722
rect 470774 304692 470812 304722
rect 470276 304658 470332 304668
rect 470356 304658 470412 304668
rect 470436 304658 470492 304668
rect 470516 304658 470572 304668
rect 470596 304658 470652 304668
rect 470676 304658 470732 304668
rect 470756 304658 470812 304668
rect 470276 304612 470314 304658
rect 470314 304612 470326 304658
rect 470326 304612 470332 304658
rect 470356 304612 470378 304658
rect 470378 304612 470390 304658
rect 470390 304612 470412 304658
rect 470436 304612 470442 304658
rect 470442 304612 470454 304658
rect 470454 304612 470492 304658
rect 470516 304612 470518 304658
rect 470518 304612 470570 304658
rect 470570 304612 470572 304658
rect 470596 304612 470634 304658
rect 470634 304612 470646 304658
rect 470646 304612 470652 304658
rect 470676 304612 470698 304658
rect 470698 304612 470710 304658
rect 470710 304612 470732 304658
rect 470756 304612 470762 304658
rect 470762 304612 470774 304658
rect 470774 304612 470812 304658
rect 470276 287435 470314 287481
rect 470314 287435 470326 287481
rect 470326 287435 470332 287481
rect 470356 287435 470378 287481
rect 470378 287435 470390 287481
rect 470390 287435 470412 287481
rect 470436 287435 470442 287481
rect 470442 287435 470454 287481
rect 470454 287435 470492 287481
rect 470516 287435 470518 287481
rect 470518 287435 470570 287481
rect 470570 287435 470572 287481
rect 470596 287435 470634 287481
rect 470634 287435 470646 287481
rect 470646 287435 470652 287481
rect 470676 287435 470698 287481
rect 470698 287435 470710 287481
rect 470710 287435 470732 287481
rect 470756 287435 470762 287481
rect 470762 287435 470774 287481
rect 470774 287435 470812 287481
rect 470276 287425 470332 287435
rect 470356 287425 470412 287435
rect 470436 287425 470492 287435
rect 470516 287425 470572 287435
rect 470596 287425 470652 287435
rect 470676 287425 470732 287435
rect 470756 287425 470812 287435
rect 470276 287371 470314 287401
rect 470314 287371 470326 287401
rect 470326 287371 470332 287401
rect 470356 287371 470378 287401
rect 470378 287371 470390 287401
rect 470390 287371 470412 287401
rect 470436 287371 470442 287401
rect 470442 287371 470454 287401
rect 470454 287371 470492 287401
rect 470516 287371 470518 287401
rect 470518 287371 470570 287401
rect 470570 287371 470572 287401
rect 470596 287371 470634 287401
rect 470634 287371 470646 287401
rect 470646 287371 470652 287401
rect 470676 287371 470698 287401
rect 470698 287371 470710 287401
rect 470710 287371 470732 287401
rect 470756 287371 470762 287401
rect 470762 287371 470774 287401
rect 470774 287371 470812 287401
rect 470276 287359 470332 287371
rect 470356 287359 470412 287371
rect 470436 287359 470492 287371
rect 470516 287359 470572 287371
rect 470596 287359 470652 287371
rect 470676 287359 470732 287371
rect 470756 287359 470812 287371
rect 470276 287345 470314 287359
rect 470314 287345 470326 287359
rect 470326 287345 470332 287359
rect 470356 287345 470378 287359
rect 470378 287345 470390 287359
rect 470390 287345 470412 287359
rect 470436 287345 470442 287359
rect 470442 287345 470454 287359
rect 470454 287345 470492 287359
rect 470516 287345 470518 287359
rect 470518 287345 470570 287359
rect 470570 287345 470572 287359
rect 470596 287345 470634 287359
rect 470634 287345 470646 287359
rect 470646 287345 470652 287359
rect 470676 287345 470698 287359
rect 470698 287345 470710 287359
rect 470710 287345 470732 287359
rect 470756 287345 470762 287359
rect 470762 287345 470774 287359
rect 470774 287345 470812 287359
rect 470276 287307 470314 287321
rect 470314 287307 470326 287321
rect 470326 287307 470332 287321
rect 470356 287307 470378 287321
rect 470378 287307 470390 287321
rect 470390 287307 470412 287321
rect 470436 287307 470442 287321
rect 470442 287307 470454 287321
rect 470454 287307 470492 287321
rect 470516 287307 470518 287321
rect 470518 287307 470570 287321
rect 470570 287307 470572 287321
rect 470596 287307 470634 287321
rect 470634 287307 470646 287321
rect 470646 287307 470652 287321
rect 470676 287307 470698 287321
rect 470698 287307 470710 287321
rect 470710 287307 470732 287321
rect 470756 287307 470762 287321
rect 470762 287307 470774 287321
rect 470774 287307 470812 287321
rect 470276 287295 470332 287307
rect 470356 287295 470412 287307
rect 470436 287295 470492 287307
rect 470516 287295 470572 287307
rect 470596 287295 470652 287307
rect 470676 287295 470732 287307
rect 470756 287295 470812 287307
rect 470276 287265 470314 287295
rect 470314 287265 470326 287295
rect 470326 287265 470332 287295
rect 470356 287265 470378 287295
rect 470378 287265 470390 287295
rect 470390 287265 470412 287295
rect 470436 287265 470442 287295
rect 470442 287265 470454 287295
rect 470454 287265 470492 287295
rect 470516 287265 470518 287295
rect 470518 287265 470570 287295
rect 470570 287265 470572 287295
rect 470596 287265 470634 287295
rect 470634 287265 470646 287295
rect 470646 287265 470652 287295
rect 470676 287265 470698 287295
rect 470698 287265 470710 287295
rect 470710 287265 470732 287295
rect 470756 287265 470762 287295
rect 470762 287265 470774 287295
rect 470774 287265 470812 287295
rect 470276 287231 470332 287241
rect 470356 287231 470412 287241
rect 470436 287231 470492 287241
rect 470516 287231 470572 287241
rect 470596 287231 470652 287241
rect 470676 287231 470732 287241
rect 470756 287231 470812 287241
rect 470276 287185 470314 287231
rect 470314 287185 470326 287231
rect 470326 287185 470332 287231
rect 470356 287185 470378 287231
rect 470378 287185 470390 287231
rect 470390 287185 470412 287231
rect 470436 287185 470442 287231
rect 470442 287185 470454 287231
rect 470454 287185 470492 287231
rect 470516 287185 470518 287231
rect 470518 287185 470570 287231
rect 470570 287185 470572 287231
rect 470596 287185 470634 287231
rect 470634 287185 470646 287231
rect 470646 287185 470652 287231
rect 470676 287185 470698 287231
rect 470698 287185 470710 287231
rect 470710 287185 470732 287231
rect 470756 287185 470762 287231
rect 470762 287185 470774 287231
rect 470774 287185 470812 287231
rect 487534 306176 487590 306232
rect 481004 306040 481060 306096
rect 473726 305904 473782 305960
rect 477739 305632 477795 305688
rect 484122 305496 484178 305552
rect 478633 286864 478689 286920
rect 474921 286592 474977 286648
rect 488630 286628 488632 286648
rect 488632 286628 488684 286648
rect 488684 286628 488686 286648
rect 488630 286592 488686 286628
rect 469036 286350 469074 286396
rect 469074 286350 469086 286396
rect 469086 286350 469092 286396
rect 469116 286350 469138 286396
rect 469138 286350 469150 286396
rect 469150 286350 469172 286396
rect 469196 286350 469202 286396
rect 469202 286350 469214 286396
rect 469214 286350 469252 286396
rect 469276 286350 469278 286396
rect 469278 286350 469330 286396
rect 469330 286350 469332 286396
rect 469356 286350 469394 286396
rect 469394 286350 469406 286396
rect 469406 286350 469412 286396
rect 469436 286350 469458 286396
rect 469458 286350 469470 286396
rect 469470 286350 469492 286396
rect 469516 286350 469522 286396
rect 469522 286350 469534 286396
rect 469534 286350 469572 286396
rect 469036 286340 469092 286350
rect 469116 286340 469172 286350
rect 469196 286340 469252 286350
rect 469276 286340 469332 286350
rect 469356 286340 469412 286350
rect 469436 286340 469492 286350
rect 469516 286340 469572 286350
rect 469036 286286 469074 286316
rect 469074 286286 469086 286316
rect 469086 286286 469092 286316
rect 469116 286286 469138 286316
rect 469138 286286 469150 286316
rect 469150 286286 469172 286316
rect 469196 286286 469202 286316
rect 469202 286286 469214 286316
rect 469214 286286 469252 286316
rect 469276 286286 469278 286316
rect 469278 286286 469330 286316
rect 469330 286286 469332 286316
rect 469356 286286 469394 286316
rect 469394 286286 469406 286316
rect 469406 286286 469412 286316
rect 469436 286286 469458 286316
rect 469458 286286 469470 286316
rect 469470 286286 469492 286316
rect 469516 286286 469522 286316
rect 469522 286286 469534 286316
rect 469534 286286 469572 286316
rect 469036 286274 469092 286286
rect 469116 286274 469172 286286
rect 469196 286274 469252 286286
rect 469276 286274 469332 286286
rect 469356 286274 469412 286286
rect 469436 286274 469492 286286
rect 469516 286274 469572 286286
rect 469036 286260 469074 286274
rect 469074 286260 469086 286274
rect 469086 286260 469092 286274
rect 469116 286260 469138 286274
rect 469138 286260 469150 286274
rect 469150 286260 469172 286274
rect 469196 286260 469202 286274
rect 469202 286260 469214 286274
rect 469214 286260 469252 286274
rect 469276 286260 469278 286274
rect 469278 286260 469330 286274
rect 469330 286260 469332 286274
rect 469356 286260 469394 286274
rect 469394 286260 469406 286274
rect 469406 286260 469412 286274
rect 469436 286260 469458 286274
rect 469458 286260 469470 286274
rect 469470 286260 469492 286274
rect 469516 286260 469522 286274
rect 469522 286260 469534 286274
rect 469534 286260 469572 286274
rect 469036 286222 469074 286236
rect 469074 286222 469086 286236
rect 469086 286222 469092 286236
rect 469116 286222 469138 286236
rect 469138 286222 469150 286236
rect 469150 286222 469172 286236
rect 469196 286222 469202 286236
rect 469202 286222 469214 286236
rect 469214 286222 469252 286236
rect 469276 286222 469278 286236
rect 469278 286222 469330 286236
rect 469330 286222 469332 286236
rect 469356 286222 469394 286236
rect 469394 286222 469406 286236
rect 469406 286222 469412 286236
rect 469436 286222 469458 286236
rect 469458 286222 469470 286236
rect 469470 286222 469492 286236
rect 469516 286222 469522 286236
rect 469522 286222 469534 286236
rect 469534 286222 469572 286236
rect 469036 286210 469092 286222
rect 469116 286210 469172 286222
rect 469196 286210 469252 286222
rect 469276 286210 469332 286222
rect 469356 286210 469412 286222
rect 469436 286210 469492 286222
rect 469516 286210 469572 286222
rect 469036 286180 469074 286210
rect 469074 286180 469086 286210
rect 469086 286180 469092 286210
rect 469116 286180 469138 286210
rect 469138 286180 469150 286210
rect 469150 286180 469172 286210
rect 469196 286180 469202 286210
rect 469202 286180 469214 286210
rect 469214 286180 469252 286210
rect 469276 286180 469278 286210
rect 469278 286180 469330 286210
rect 469330 286180 469332 286210
rect 469356 286180 469394 286210
rect 469394 286180 469406 286210
rect 469406 286180 469412 286210
rect 469436 286180 469458 286210
rect 469458 286180 469470 286210
rect 469470 286180 469492 286210
rect 469516 286180 469522 286210
rect 469522 286180 469534 286210
rect 469534 286180 469572 286210
rect 469036 286146 469092 286156
rect 469116 286146 469172 286156
rect 469196 286146 469252 286156
rect 469276 286146 469332 286156
rect 469356 286146 469412 286156
rect 469436 286146 469492 286156
rect 469516 286146 469572 286156
rect 469036 286100 469074 286146
rect 469074 286100 469086 286146
rect 469086 286100 469092 286146
rect 469116 286100 469138 286146
rect 469138 286100 469150 286146
rect 469150 286100 469172 286146
rect 469196 286100 469202 286146
rect 469202 286100 469214 286146
rect 469214 286100 469252 286146
rect 469276 286100 469278 286146
rect 469278 286100 469330 286146
rect 469330 286100 469332 286146
rect 469356 286100 469394 286146
rect 469394 286100 469406 286146
rect 469406 286100 469412 286146
rect 469436 286100 469458 286146
rect 469458 286100 469470 286146
rect 469470 286100 469492 286146
rect 469516 286100 469522 286146
rect 469522 286100 469534 286146
rect 469534 286100 469572 286146
rect 470276 285262 470314 285308
rect 470314 285262 470326 285308
rect 470326 285262 470332 285308
rect 470356 285262 470378 285308
rect 470378 285262 470390 285308
rect 470390 285262 470412 285308
rect 470436 285262 470442 285308
rect 470442 285262 470454 285308
rect 470454 285262 470492 285308
rect 470516 285262 470518 285308
rect 470518 285262 470570 285308
rect 470570 285262 470572 285308
rect 470596 285262 470634 285308
rect 470634 285262 470646 285308
rect 470646 285262 470652 285308
rect 470676 285262 470698 285308
rect 470698 285262 470710 285308
rect 470710 285262 470732 285308
rect 470756 285262 470762 285308
rect 470762 285262 470774 285308
rect 470774 285262 470812 285308
rect 470276 285252 470332 285262
rect 470356 285252 470412 285262
rect 470436 285252 470492 285262
rect 470516 285252 470572 285262
rect 470596 285252 470652 285262
rect 470676 285252 470732 285262
rect 470756 285252 470812 285262
rect 470276 285198 470314 285228
rect 470314 285198 470326 285228
rect 470326 285198 470332 285228
rect 470356 285198 470378 285228
rect 470378 285198 470390 285228
rect 470390 285198 470412 285228
rect 470436 285198 470442 285228
rect 470442 285198 470454 285228
rect 470454 285198 470492 285228
rect 470516 285198 470518 285228
rect 470518 285198 470570 285228
rect 470570 285198 470572 285228
rect 470596 285198 470634 285228
rect 470634 285198 470646 285228
rect 470646 285198 470652 285228
rect 470676 285198 470698 285228
rect 470698 285198 470710 285228
rect 470710 285198 470732 285228
rect 470756 285198 470762 285228
rect 470762 285198 470774 285228
rect 470774 285198 470812 285228
rect 470276 285186 470332 285198
rect 470356 285186 470412 285198
rect 470436 285186 470492 285198
rect 470516 285186 470572 285198
rect 470596 285186 470652 285198
rect 470676 285186 470732 285198
rect 470756 285186 470812 285198
rect 470276 285172 470314 285186
rect 470314 285172 470326 285186
rect 470326 285172 470332 285186
rect 470356 285172 470378 285186
rect 470378 285172 470390 285186
rect 470390 285172 470412 285186
rect 470436 285172 470442 285186
rect 470442 285172 470454 285186
rect 470454 285172 470492 285186
rect 470516 285172 470518 285186
rect 470518 285172 470570 285186
rect 470570 285172 470572 285186
rect 470596 285172 470634 285186
rect 470634 285172 470646 285186
rect 470646 285172 470652 285186
rect 470676 285172 470698 285186
rect 470698 285172 470710 285186
rect 470710 285172 470732 285186
rect 470756 285172 470762 285186
rect 470762 285172 470774 285186
rect 470774 285172 470812 285186
rect 470276 285134 470314 285148
rect 470314 285134 470326 285148
rect 470326 285134 470332 285148
rect 470356 285134 470378 285148
rect 470378 285134 470390 285148
rect 470390 285134 470412 285148
rect 470436 285134 470442 285148
rect 470442 285134 470454 285148
rect 470454 285134 470492 285148
rect 470516 285134 470518 285148
rect 470518 285134 470570 285148
rect 470570 285134 470572 285148
rect 470596 285134 470634 285148
rect 470634 285134 470646 285148
rect 470646 285134 470652 285148
rect 470676 285134 470698 285148
rect 470698 285134 470710 285148
rect 470710 285134 470732 285148
rect 470756 285134 470762 285148
rect 470762 285134 470774 285148
rect 470774 285134 470812 285148
rect 470276 285122 470332 285134
rect 470356 285122 470412 285134
rect 470436 285122 470492 285134
rect 470516 285122 470572 285134
rect 470596 285122 470652 285134
rect 470676 285122 470732 285134
rect 470756 285122 470812 285134
rect 470276 285092 470314 285122
rect 470314 285092 470326 285122
rect 470326 285092 470332 285122
rect 470356 285092 470378 285122
rect 470378 285092 470390 285122
rect 470390 285092 470412 285122
rect 470436 285092 470442 285122
rect 470442 285092 470454 285122
rect 470454 285092 470492 285122
rect 470516 285092 470518 285122
rect 470518 285092 470570 285122
rect 470570 285092 470572 285122
rect 470596 285092 470634 285122
rect 470634 285092 470646 285122
rect 470646 285092 470652 285122
rect 470676 285092 470698 285122
rect 470698 285092 470710 285122
rect 470710 285092 470732 285122
rect 470756 285092 470762 285122
rect 470762 285092 470774 285122
rect 470774 285092 470812 285122
rect 470276 285058 470332 285068
rect 470356 285058 470412 285068
rect 470436 285058 470492 285068
rect 470516 285058 470572 285068
rect 470596 285058 470652 285068
rect 470676 285058 470732 285068
rect 470756 285058 470812 285068
rect 470276 285012 470314 285058
rect 470314 285012 470326 285058
rect 470326 285012 470332 285058
rect 470356 285012 470378 285058
rect 470378 285012 470390 285058
rect 470390 285012 470412 285058
rect 470436 285012 470442 285058
rect 470442 285012 470454 285058
rect 470454 285012 470492 285058
rect 470516 285012 470518 285058
rect 470518 285012 470570 285058
rect 470570 285012 470572 285058
rect 470596 285012 470634 285058
rect 470634 285012 470646 285058
rect 470646 285012 470652 285058
rect 470676 285012 470698 285058
rect 470698 285012 470710 285058
rect 470710 285012 470732 285058
rect 470756 285012 470762 285058
rect 470762 285012 470774 285058
rect 470774 285012 470812 285058
rect 482345 285776 482401 285832
rect 485870 285776 485926 285832
rect 470276 267435 470314 267481
rect 470314 267435 470326 267481
rect 470326 267435 470332 267481
rect 470356 267435 470378 267481
rect 470378 267435 470390 267481
rect 470390 267435 470412 267481
rect 470436 267435 470442 267481
rect 470442 267435 470454 267481
rect 470454 267435 470492 267481
rect 470516 267435 470518 267481
rect 470518 267435 470570 267481
rect 470570 267435 470572 267481
rect 470596 267435 470634 267481
rect 470634 267435 470646 267481
rect 470646 267435 470652 267481
rect 470676 267435 470698 267481
rect 470698 267435 470710 267481
rect 470710 267435 470732 267481
rect 470756 267435 470762 267481
rect 470762 267435 470774 267481
rect 470774 267435 470812 267481
rect 470276 267425 470332 267435
rect 470356 267425 470412 267435
rect 470436 267425 470492 267435
rect 470516 267425 470572 267435
rect 470596 267425 470652 267435
rect 470676 267425 470732 267435
rect 470756 267425 470812 267435
rect 470276 267371 470314 267401
rect 470314 267371 470326 267401
rect 470326 267371 470332 267401
rect 470356 267371 470378 267401
rect 470378 267371 470390 267401
rect 470390 267371 470412 267401
rect 470436 267371 470442 267401
rect 470442 267371 470454 267401
rect 470454 267371 470492 267401
rect 470516 267371 470518 267401
rect 470518 267371 470570 267401
rect 470570 267371 470572 267401
rect 470596 267371 470634 267401
rect 470634 267371 470646 267401
rect 470646 267371 470652 267401
rect 470676 267371 470698 267401
rect 470698 267371 470710 267401
rect 470710 267371 470732 267401
rect 470756 267371 470762 267401
rect 470762 267371 470774 267401
rect 470774 267371 470812 267401
rect 470276 267359 470332 267371
rect 470356 267359 470412 267371
rect 470436 267359 470492 267371
rect 470516 267359 470572 267371
rect 470596 267359 470652 267371
rect 470676 267359 470732 267371
rect 470756 267359 470812 267371
rect 470276 267345 470314 267359
rect 470314 267345 470326 267359
rect 470326 267345 470332 267359
rect 470356 267345 470378 267359
rect 470378 267345 470390 267359
rect 470390 267345 470412 267359
rect 470436 267345 470442 267359
rect 470442 267345 470454 267359
rect 470454 267345 470492 267359
rect 470516 267345 470518 267359
rect 470518 267345 470570 267359
rect 470570 267345 470572 267359
rect 470596 267345 470634 267359
rect 470634 267345 470646 267359
rect 470646 267345 470652 267359
rect 470676 267345 470698 267359
rect 470698 267345 470710 267359
rect 470710 267345 470732 267359
rect 470756 267345 470762 267359
rect 470762 267345 470774 267359
rect 470774 267345 470812 267359
rect 470276 267307 470314 267321
rect 470314 267307 470326 267321
rect 470326 267307 470332 267321
rect 470356 267307 470378 267321
rect 470378 267307 470390 267321
rect 470390 267307 470412 267321
rect 470436 267307 470442 267321
rect 470442 267307 470454 267321
rect 470454 267307 470492 267321
rect 470516 267307 470518 267321
rect 470518 267307 470570 267321
rect 470570 267307 470572 267321
rect 470596 267307 470634 267321
rect 470634 267307 470646 267321
rect 470646 267307 470652 267321
rect 470676 267307 470698 267321
rect 470698 267307 470710 267321
rect 470710 267307 470732 267321
rect 470756 267307 470762 267321
rect 470762 267307 470774 267321
rect 470774 267307 470812 267321
rect 470276 267295 470332 267307
rect 470356 267295 470412 267307
rect 470436 267295 470492 267307
rect 470516 267295 470572 267307
rect 470596 267295 470652 267307
rect 470676 267295 470732 267307
rect 470756 267295 470812 267307
rect 470276 267265 470314 267295
rect 470314 267265 470326 267295
rect 470326 267265 470332 267295
rect 470356 267265 470378 267295
rect 470378 267265 470390 267295
rect 470390 267265 470412 267295
rect 470436 267265 470442 267295
rect 470442 267265 470454 267295
rect 470454 267265 470492 267295
rect 470516 267265 470518 267295
rect 470518 267265 470570 267295
rect 470570 267265 470572 267295
rect 470596 267265 470634 267295
rect 470634 267265 470646 267295
rect 470646 267265 470652 267295
rect 470676 267265 470698 267295
rect 470698 267265 470710 267295
rect 470710 267265 470732 267295
rect 470756 267265 470762 267295
rect 470762 267265 470774 267295
rect 470774 267265 470812 267295
rect 470276 267231 470332 267241
rect 470356 267231 470412 267241
rect 470436 267231 470492 267241
rect 470516 267231 470572 267241
rect 470596 267231 470652 267241
rect 470676 267231 470732 267241
rect 470756 267231 470812 267241
rect 470276 267185 470314 267231
rect 470314 267185 470326 267231
rect 470326 267185 470332 267231
rect 470356 267185 470378 267231
rect 470378 267185 470390 267231
rect 470390 267185 470412 267231
rect 470436 267185 470442 267231
rect 470442 267185 470454 267231
rect 470454 267185 470492 267231
rect 470516 267185 470518 267231
rect 470518 267185 470570 267231
rect 470570 267185 470572 267231
rect 470596 267185 470634 267231
rect 470634 267185 470646 267231
rect 470646 267185 470652 267231
rect 470676 267185 470698 267231
rect 470698 267185 470710 267231
rect 470710 267185 470732 267231
rect 470756 267185 470762 267231
rect 470762 267185 470774 267231
rect 470774 267185 470812 267231
rect 469036 266349 469074 266395
rect 469074 266349 469086 266395
rect 469086 266349 469092 266395
rect 469116 266349 469138 266395
rect 469138 266349 469150 266395
rect 469150 266349 469172 266395
rect 469196 266349 469202 266395
rect 469202 266349 469214 266395
rect 469214 266349 469252 266395
rect 469276 266349 469278 266395
rect 469278 266349 469330 266395
rect 469330 266349 469332 266395
rect 469356 266349 469394 266395
rect 469394 266349 469406 266395
rect 469406 266349 469412 266395
rect 469436 266349 469458 266395
rect 469458 266349 469470 266395
rect 469470 266349 469492 266395
rect 469516 266349 469522 266395
rect 469522 266349 469534 266395
rect 469534 266349 469572 266395
rect 469036 266339 469092 266349
rect 469116 266339 469172 266349
rect 469196 266339 469252 266349
rect 469276 266339 469332 266349
rect 469356 266339 469412 266349
rect 469436 266339 469492 266349
rect 469516 266339 469572 266349
rect 469036 266285 469074 266315
rect 469074 266285 469086 266315
rect 469086 266285 469092 266315
rect 469116 266285 469138 266315
rect 469138 266285 469150 266315
rect 469150 266285 469172 266315
rect 469196 266285 469202 266315
rect 469202 266285 469214 266315
rect 469214 266285 469252 266315
rect 469276 266285 469278 266315
rect 469278 266285 469330 266315
rect 469330 266285 469332 266315
rect 469356 266285 469394 266315
rect 469394 266285 469406 266315
rect 469406 266285 469412 266315
rect 469436 266285 469458 266315
rect 469458 266285 469470 266315
rect 469470 266285 469492 266315
rect 469516 266285 469522 266315
rect 469522 266285 469534 266315
rect 469534 266285 469572 266315
rect 469036 266273 469092 266285
rect 469116 266273 469172 266285
rect 469196 266273 469252 266285
rect 469276 266273 469332 266285
rect 469356 266273 469412 266285
rect 469436 266273 469492 266285
rect 469516 266273 469572 266285
rect 469036 266259 469074 266273
rect 469074 266259 469086 266273
rect 469086 266259 469092 266273
rect 469116 266259 469138 266273
rect 469138 266259 469150 266273
rect 469150 266259 469172 266273
rect 469196 266259 469202 266273
rect 469202 266259 469214 266273
rect 469214 266259 469252 266273
rect 469276 266259 469278 266273
rect 469278 266259 469330 266273
rect 469330 266259 469332 266273
rect 469356 266259 469394 266273
rect 469394 266259 469406 266273
rect 469406 266259 469412 266273
rect 469436 266259 469458 266273
rect 469458 266259 469470 266273
rect 469470 266259 469492 266273
rect 469516 266259 469522 266273
rect 469522 266259 469534 266273
rect 469534 266259 469572 266273
rect 469036 266221 469074 266235
rect 469074 266221 469086 266235
rect 469086 266221 469092 266235
rect 469116 266221 469138 266235
rect 469138 266221 469150 266235
rect 469150 266221 469172 266235
rect 469196 266221 469202 266235
rect 469202 266221 469214 266235
rect 469214 266221 469252 266235
rect 469276 266221 469278 266235
rect 469278 266221 469330 266235
rect 469330 266221 469332 266235
rect 469356 266221 469394 266235
rect 469394 266221 469406 266235
rect 469406 266221 469412 266235
rect 469436 266221 469458 266235
rect 469458 266221 469470 266235
rect 469470 266221 469492 266235
rect 469516 266221 469522 266235
rect 469522 266221 469534 266235
rect 469534 266221 469572 266235
rect 469036 266209 469092 266221
rect 469116 266209 469172 266221
rect 469196 266209 469252 266221
rect 469276 266209 469332 266221
rect 469356 266209 469412 266221
rect 469436 266209 469492 266221
rect 469516 266209 469572 266221
rect 469036 266179 469074 266209
rect 469074 266179 469086 266209
rect 469086 266179 469092 266209
rect 469116 266179 469138 266209
rect 469138 266179 469150 266209
rect 469150 266179 469172 266209
rect 469196 266179 469202 266209
rect 469202 266179 469214 266209
rect 469214 266179 469252 266209
rect 469276 266179 469278 266209
rect 469278 266179 469330 266209
rect 469330 266179 469332 266209
rect 469356 266179 469394 266209
rect 469394 266179 469406 266209
rect 469406 266179 469412 266209
rect 469436 266179 469458 266209
rect 469458 266179 469470 266209
rect 469470 266179 469492 266209
rect 469516 266179 469522 266209
rect 469522 266179 469534 266209
rect 469534 266179 469572 266209
rect 469036 266145 469092 266155
rect 469116 266145 469172 266155
rect 469196 266145 469252 266155
rect 469276 266145 469332 266155
rect 469356 266145 469412 266155
rect 469436 266145 469492 266155
rect 469516 266145 469572 266155
rect 469036 266099 469074 266145
rect 469074 266099 469086 266145
rect 469086 266099 469092 266145
rect 469116 266099 469138 266145
rect 469138 266099 469150 266145
rect 469150 266099 469172 266145
rect 469196 266099 469202 266145
rect 469202 266099 469214 266145
rect 469214 266099 469252 266145
rect 469276 266099 469278 266145
rect 469278 266099 469330 266145
rect 469330 266099 469332 266145
rect 469356 266099 469394 266145
rect 469394 266099 469406 266145
rect 469406 266099 469412 266145
rect 469436 266099 469458 266145
rect 469458 266099 469470 266145
rect 469470 266099 469492 266145
rect 469516 266099 469522 266145
rect 469522 266099 469534 266145
rect 469534 266099 469572 266145
rect 470276 265262 470314 265308
rect 470314 265262 470326 265308
rect 470326 265262 470332 265308
rect 470356 265262 470378 265308
rect 470378 265262 470390 265308
rect 470390 265262 470412 265308
rect 470436 265262 470442 265308
rect 470442 265262 470454 265308
rect 470454 265262 470492 265308
rect 470516 265262 470518 265308
rect 470518 265262 470570 265308
rect 470570 265262 470572 265308
rect 470596 265262 470634 265308
rect 470634 265262 470646 265308
rect 470646 265262 470652 265308
rect 470676 265262 470698 265308
rect 470698 265262 470710 265308
rect 470710 265262 470732 265308
rect 470756 265262 470762 265308
rect 470762 265262 470774 265308
rect 470774 265262 470812 265308
rect 470276 265252 470332 265262
rect 470356 265252 470412 265262
rect 470436 265252 470492 265262
rect 470516 265252 470572 265262
rect 470596 265252 470652 265262
rect 470676 265252 470732 265262
rect 470756 265252 470812 265262
rect 470276 265198 470314 265228
rect 470314 265198 470326 265228
rect 470326 265198 470332 265228
rect 470356 265198 470378 265228
rect 470378 265198 470390 265228
rect 470390 265198 470412 265228
rect 470436 265198 470442 265228
rect 470442 265198 470454 265228
rect 470454 265198 470492 265228
rect 470516 265198 470518 265228
rect 470518 265198 470570 265228
rect 470570 265198 470572 265228
rect 470596 265198 470634 265228
rect 470634 265198 470646 265228
rect 470646 265198 470652 265228
rect 470676 265198 470698 265228
rect 470698 265198 470710 265228
rect 470710 265198 470732 265228
rect 470756 265198 470762 265228
rect 470762 265198 470774 265228
rect 470774 265198 470812 265228
rect 470276 265186 470332 265198
rect 470356 265186 470412 265198
rect 470436 265186 470492 265198
rect 470516 265186 470572 265198
rect 470596 265186 470652 265198
rect 470676 265186 470732 265198
rect 470756 265186 470812 265198
rect 470276 265172 470314 265186
rect 470314 265172 470326 265186
rect 470326 265172 470332 265186
rect 470356 265172 470378 265186
rect 470378 265172 470390 265186
rect 470390 265172 470412 265186
rect 470436 265172 470442 265186
rect 470442 265172 470454 265186
rect 470454 265172 470492 265186
rect 470516 265172 470518 265186
rect 470518 265172 470570 265186
rect 470570 265172 470572 265186
rect 470596 265172 470634 265186
rect 470634 265172 470646 265186
rect 470646 265172 470652 265186
rect 470676 265172 470698 265186
rect 470698 265172 470710 265186
rect 470710 265172 470732 265186
rect 470756 265172 470762 265186
rect 470762 265172 470774 265186
rect 470774 265172 470812 265186
rect 470276 265134 470314 265148
rect 470314 265134 470326 265148
rect 470326 265134 470332 265148
rect 470356 265134 470378 265148
rect 470378 265134 470390 265148
rect 470390 265134 470412 265148
rect 470436 265134 470442 265148
rect 470442 265134 470454 265148
rect 470454 265134 470492 265148
rect 470516 265134 470518 265148
rect 470518 265134 470570 265148
rect 470570 265134 470572 265148
rect 470596 265134 470634 265148
rect 470634 265134 470646 265148
rect 470646 265134 470652 265148
rect 470676 265134 470698 265148
rect 470698 265134 470710 265148
rect 470710 265134 470732 265148
rect 470756 265134 470762 265148
rect 470762 265134 470774 265148
rect 470774 265134 470812 265148
rect 470276 265122 470332 265134
rect 470356 265122 470412 265134
rect 470436 265122 470492 265134
rect 470516 265122 470572 265134
rect 470596 265122 470652 265134
rect 470676 265122 470732 265134
rect 470756 265122 470812 265134
rect 470276 265092 470314 265122
rect 470314 265092 470326 265122
rect 470326 265092 470332 265122
rect 470356 265092 470378 265122
rect 470378 265092 470390 265122
rect 470390 265092 470412 265122
rect 470436 265092 470442 265122
rect 470442 265092 470454 265122
rect 470454 265092 470492 265122
rect 470516 265092 470518 265122
rect 470518 265092 470570 265122
rect 470570 265092 470572 265122
rect 470596 265092 470634 265122
rect 470634 265092 470646 265122
rect 470646 265092 470652 265122
rect 470676 265092 470698 265122
rect 470698 265092 470710 265122
rect 470710 265092 470732 265122
rect 470756 265092 470762 265122
rect 470762 265092 470774 265122
rect 470774 265092 470812 265122
rect 470276 265058 470332 265068
rect 470356 265058 470412 265068
rect 470436 265058 470492 265068
rect 470516 265058 470572 265068
rect 470596 265058 470652 265068
rect 470676 265058 470732 265068
rect 470756 265058 470812 265068
rect 470276 265012 470314 265058
rect 470314 265012 470326 265058
rect 470326 265012 470332 265058
rect 470356 265012 470378 265058
rect 470378 265012 470390 265058
rect 470390 265012 470412 265058
rect 470436 265012 470442 265058
rect 470442 265012 470454 265058
rect 470454 265012 470492 265058
rect 470516 265012 470518 265058
rect 470518 265012 470570 265058
rect 470570 265012 470572 265058
rect 470596 265012 470634 265058
rect 470634 265012 470646 265058
rect 470646 265012 470652 265058
rect 470676 265012 470698 265058
rect 470698 265012 470710 265058
rect 470710 265012 470732 265058
rect 470756 265012 470762 265058
rect 470762 265012 470774 265058
rect 470774 265012 470812 265058
rect 479062 265920 479118 265976
rect 476486 264968 476542 265024
rect 479522 264968 479578 265024
rect 482834 264968 482890 265024
rect 488722 265512 488778 265568
rect 485686 264968 485742 265024
rect 535458 444760 535514 444816
rect 535458 443400 535514 443456
rect 535458 442040 535514 442096
rect 535458 440680 535514 440736
rect 535458 439320 535514 439376
rect 535458 437960 535514 438016
rect 535458 436600 535514 436656
rect 535458 435240 535514 435296
rect 535458 433880 535514 433936
rect 535458 432520 535514 432576
rect 536746 424360 536802 424416
rect 535458 409264 535514 409320
rect 535458 406544 535514 406600
rect 535458 404504 535514 404560
rect 535458 403144 535514 403200
rect 536378 401648 536434 401704
rect 536286 400288 536342 400344
rect 535458 399064 535514 399120
rect 536102 397432 536158 397488
rect 535458 396344 535514 396400
rect 535458 372816 535514 372872
rect 535458 371456 535514 371512
rect 535458 368736 535514 368792
rect 535458 367376 535514 367432
rect 535458 366016 535514 366072
rect 535458 361936 535514 361992
rect 535918 360576 535974 360632
rect 535458 336776 535514 336832
rect 535458 331336 535514 331392
rect 535458 329976 535514 330032
rect 535458 325896 535514 325952
rect 535458 300772 535460 300792
rect 535460 300772 535512 300792
rect 535512 300772 535514 300792
rect 535458 300736 535514 300772
rect 535458 299412 535460 299432
rect 535460 299412 535512 299432
rect 535512 299412 535514 299432
rect 535458 299376 535514 299412
rect 535458 298052 535460 298072
rect 535460 298052 535512 298072
rect 535512 298052 535514 298072
rect 535458 298016 535514 298052
rect 535458 296656 535514 296712
rect 535550 295296 535606 295352
rect 535458 293936 535514 293992
rect 535550 292576 535606 292632
rect 535458 291216 535514 291272
rect 535458 289876 535514 289912
rect 535458 289856 535460 289876
rect 535460 289856 535512 289876
rect 535512 289856 535514 289876
rect 535458 288496 535514 288552
rect 536010 328616 536066 328672
rect 536194 388320 536250 388376
rect 536194 359216 536250 359272
rect 541714 445032 541770 445088
rect 544198 445032 544254 445088
rect 541714 409264 541770 409320
rect 544290 409264 544346 409320
rect 536746 395936 536802 395992
rect 547326 404912 547382 404968
rect 544474 373360 544530 373416
rect 536562 364656 536618 364712
rect 536470 363296 536526 363352
rect 536378 324536 536434 324592
rect 541714 373088 541770 373144
rect 536746 352416 536802 352472
rect 536654 327256 536710 327312
rect 541714 339496 541770 339552
rect 544198 339496 544254 339552
rect 536746 323176 536802 323232
rect 536746 316376 536802 316432
rect 544198 303728 544254 303784
rect 541714 303592 541770 303648
rect 547326 303592 547382 303648
rect 536746 287136 536802 287192
rect 547326 300056 547382 300112
rect 580170 300056 580226 300112
rect 580170 298696 580226 298752
rect 538678 245520 538734 245576
rect 580170 205672 580226 205728
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect 470266 451483 470822 451484
rect 470266 451419 470272 451483
rect 470336 451419 470352 451483
rect 470416 451419 470432 451483
rect 470496 451419 470512 451483
rect 470576 451419 470592 451483
rect 470656 451419 470672 451483
rect 470736 451419 470752 451483
rect 470816 451419 470822 451483
rect 470266 451403 470822 451419
rect 470266 451339 470272 451403
rect 470336 451339 470352 451403
rect 470416 451339 470432 451403
rect 470496 451339 470512 451403
rect 470576 451339 470592 451403
rect 470656 451339 470672 451403
rect 470736 451339 470752 451403
rect 470816 451339 470822 451403
rect 470266 451323 470822 451339
rect 470266 451259 470272 451323
rect 470336 451259 470352 451323
rect 470416 451259 470432 451323
rect 470496 451259 470512 451323
rect 470576 451259 470592 451323
rect 470656 451259 470672 451323
rect 470736 451259 470752 451323
rect 470816 451259 470822 451323
rect 470266 451243 470822 451259
rect 470266 451179 470272 451243
rect 470336 451179 470352 451243
rect 470416 451179 470432 451243
rect 470496 451179 470512 451243
rect 470576 451179 470592 451243
rect 470656 451179 470672 451243
rect 470736 451179 470752 451243
rect 470816 451179 470822 451243
rect 470266 451178 470822 451179
rect 469026 450397 469582 450398
rect 469026 450333 469032 450397
rect 469096 450333 469112 450397
rect 469176 450333 469192 450397
rect 469256 450333 469272 450397
rect 469336 450333 469352 450397
rect 469416 450333 469432 450397
rect 469496 450333 469512 450397
rect 469576 450333 469582 450397
rect 469026 450317 469582 450333
rect 469026 450253 469032 450317
rect 469096 450253 469112 450317
rect 469176 450253 469192 450317
rect 469256 450253 469272 450317
rect 469336 450253 469352 450317
rect 469416 450253 469432 450317
rect 469496 450253 469512 450317
rect 469576 450253 469582 450317
rect 469026 450237 469582 450253
rect 469026 450173 469032 450237
rect 469096 450173 469112 450237
rect 469176 450173 469192 450237
rect 469256 450173 469272 450237
rect 469336 450173 469352 450237
rect 469416 450173 469432 450237
rect 469496 450173 469512 450237
rect 469576 450173 469582 450237
rect 477838 450258 477904 450261
rect 481155 450260 481221 450261
rect 478454 450258 478460 450260
rect 477838 450256 478460 450258
rect 477838 450200 477843 450256
rect 477899 450200 478460 450256
rect 477838 450198 478460 450200
rect 477838 450195 477904 450198
rect 478454 450196 478460 450198
rect 478524 450196 478530 450260
rect 481155 450256 481220 450260
rect 481155 450200 481160 450256
rect 481216 450200 481220 450256
rect 481155 450196 481220 450200
rect 481284 450258 481290 450260
rect 481284 450198 481312 450258
rect 481284 450196 481290 450198
rect 484158 450196 484164 450260
rect 484228 450258 484234 450260
rect 484472 450258 484538 450261
rect 484228 450256 484538 450258
rect 484228 450200 484477 450256
rect 484533 450200 484538 450256
rect 484228 450198 484538 450200
rect 484228 450196 484234 450198
rect 481155 450195 481221 450196
rect 484472 450195 484538 450198
rect 487788 450260 487854 450261
rect 487788 450256 487844 450260
rect 487908 450258 487914 450260
rect 487788 450200 487793 450256
rect 487788 450196 487844 450200
rect 487908 450198 487945 450258
rect 487908 450196 487914 450198
rect 487788 450195 487854 450196
rect 469026 450157 469582 450173
rect 469026 450093 469032 450157
rect 469096 450093 469112 450157
rect 469176 450093 469192 450157
rect 469256 450093 469272 450157
rect 469336 450093 469352 450157
rect 469416 450093 469432 450157
rect 469496 450093 469512 450157
rect 469576 450093 469582 450157
rect 469026 450092 469582 450093
rect -960 449428 480 449668
rect 473670 449652 473676 449716
rect 473740 449714 473746 449716
rect 474089 449714 474155 449717
rect 473740 449712 474155 449714
rect 473740 449656 474094 449712
rect 474150 449656 474155 449712
rect 473740 449654 474155 449656
rect 473740 449652 473746 449654
rect 474089 449651 474155 449654
rect 470266 449312 470822 449313
rect 470266 449248 470272 449312
rect 470336 449248 470352 449312
rect 470416 449248 470432 449312
rect 470496 449248 470512 449312
rect 470576 449248 470592 449312
rect 470656 449248 470672 449312
rect 470736 449248 470752 449312
rect 470816 449248 470822 449312
rect 470266 449232 470822 449248
rect 470266 449168 470272 449232
rect 470336 449168 470352 449232
rect 470416 449168 470432 449232
rect 470496 449168 470512 449232
rect 470576 449168 470592 449232
rect 470656 449168 470672 449232
rect 470736 449168 470752 449232
rect 470816 449168 470822 449232
rect 470266 449152 470822 449168
rect 470266 449088 470272 449152
rect 470336 449088 470352 449152
rect 470416 449088 470432 449152
rect 470496 449088 470512 449152
rect 470576 449088 470592 449152
rect 470656 449088 470672 449152
rect 470736 449088 470752 449152
rect 470816 449088 470822 449152
rect 470266 449072 470822 449088
rect 470266 449008 470272 449072
rect 470336 449008 470352 449072
rect 470416 449008 470432 449072
rect 470496 449008 470512 449072
rect 470576 449008 470592 449072
rect 470656 449008 470672 449072
rect 470736 449008 470752 449072
rect 470816 449008 470822 449072
rect 470266 449007 470822 449008
rect 541566 445028 541572 445092
rect 541636 445090 541642 445092
rect 541709 445090 541775 445093
rect 541636 445088 541775 445090
rect 541636 445032 541714 445088
rect 541770 445032 541775 445088
rect 541636 445030 541775 445032
rect 541636 445028 541642 445030
rect 541709 445027 541775 445030
rect 544193 445090 544259 445093
rect 544326 445090 544332 445092
rect 544193 445088 544332 445090
rect 544193 445032 544198 445088
rect 544254 445032 544332 445088
rect 544193 445030 544332 445032
rect 544193 445027 544259 445030
rect 544326 445028 544332 445030
rect 544396 445028 544402 445092
rect 535453 444818 535519 444821
rect 535453 444816 538108 444818
rect 535453 444760 535458 444816
rect 535514 444760 538108 444816
rect 535453 444758 538108 444760
rect 535453 444755 535519 444758
rect 583520 444668 584960 444908
rect 535453 443458 535519 443461
rect 535453 443456 538108 443458
rect 535453 443400 535458 443456
rect 535514 443400 538108 443456
rect 535453 443398 538108 443400
rect 535453 443395 535519 443398
rect 535453 442098 535519 442101
rect 535453 442096 538108 442098
rect 535453 442040 535458 442096
rect 535514 442040 538108 442096
rect 535453 442038 538108 442040
rect 535453 442035 535519 442038
rect 535453 440738 535519 440741
rect 535453 440736 538108 440738
rect 535453 440680 535458 440736
rect 535514 440680 538108 440736
rect 535453 440678 538108 440680
rect 535453 440675 535519 440678
rect 535453 439378 535519 439381
rect 535453 439376 538108 439378
rect 535453 439320 535458 439376
rect 535514 439320 538108 439376
rect 535453 439318 538108 439320
rect 535453 439315 535519 439318
rect 535453 438018 535519 438021
rect 535453 438016 538108 438018
rect 535453 437960 535458 438016
rect 535514 437960 538108 438016
rect 535453 437958 538108 437960
rect 535453 437955 535519 437958
rect -960 436508 480 436748
rect 535453 436658 535519 436661
rect 535453 436656 538108 436658
rect 535453 436600 535458 436656
rect 535514 436600 538108 436656
rect 535453 436598 538108 436600
rect 535453 436595 535519 436598
rect 535453 435298 535519 435301
rect 535453 435296 538108 435298
rect 535453 435240 535458 435296
rect 535514 435240 538108 435296
rect 535453 435238 538108 435240
rect 535453 435235 535519 435238
rect 549294 434754 549300 434756
rect 547860 434694 549300 434754
rect 549294 434692 549300 434694
rect 549364 434692 549370 434756
rect 535453 433938 535519 433941
rect 535453 433936 538108 433938
rect 535453 433880 535458 433936
rect 535514 433880 538108 433936
rect 535453 433878 538108 433880
rect 535453 433875 535519 433878
rect 470266 433084 470822 433085
rect 470266 433020 470272 433084
rect 470336 433020 470352 433084
rect 470416 433020 470432 433084
rect 470496 433020 470512 433084
rect 470576 433020 470592 433084
rect 470656 433020 470672 433084
rect 470736 433020 470752 433084
rect 470816 433020 470822 433084
rect 470266 433004 470822 433020
rect 470266 432940 470272 433004
rect 470336 432940 470352 433004
rect 470416 432940 470432 433004
rect 470496 432940 470512 433004
rect 470576 432940 470592 433004
rect 470656 432940 470672 433004
rect 470736 432940 470752 433004
rect 470816 432940 470822 433004
rect 470266 432924 470822 432940
rect 470266 432860 470272 432924
rect 470336 432860 470352 432924
rect 470416 432860 470432 432924
rect 470496 432860 470512 432924
rect 470576 432860 470592 432924
rect 470656 432860 470672 432924
rect 470736 432860 470752 432924
rect 470816 432860 470822 432924
rect 470266 432844 470822 432860
rect 470266 432780 470272 432844
rect 470336 432780 470352 432844
rect 470416 432780 470432 432844
rect 470496 432780 470512 432844
rect 470576 432780 470592 432844
rect 470656 432780 470672 432844
rect 470736 432780 470752 432844
rect 470816 432780 470822 432844
rect 470266 432779 470822 432780
rect 535453 432578 535519 432581
rect 535453 432576 538108 432578
rect 535453 432520 535458 432576
rect 535514 432520 538108 432576
rect 535453 432518 538108 432520
rect 535453 432515 535519 432518
rect 483565 432308 483631 432309
rect 483565 432306 483612 432308
rect 483520 432304 483612 432306
rect 483520 432248 483570 432304
rect 483520 432246 483612 432248
rect 483565 432244 483612 432246
rect 483676 432244 483682 432308
rect 483565 432243 483631 432244
rect 481265 432172 481331 432173
rect 481214 432108 481220 432172
rect 481284 432170 481331 432172
rect 481284 432168 481376 432170
rect 481326 432112 481376 432168
rect 481284 432110 481376 432112
rect 481284 432108 481331 432110
rect 481265 432107 481331 432108
rect 469026 431997 469582 431998
rect 469026 431933 469032 431997
rect 469096 431933 469112 431997
rect 469176 431933 469192 431997
rect 469256 431933 469272 431997
rect 469336 431933 469352 431997
rect 469416 431933 469432 431997
rect 469496 431933 469512 431997
rect 469576 431933 469582 431997
rect 469026 431917 469582 431933
rect 469026 431853 469032 431917
rect 469096 431853 469112 431917
rect 469176 431853 469192 431917
rect 469256 431853 469272 431917
rect 469336 431853 469352 431917
rect 469416 431853 469432 431917
rect 469496 431853 469512 431917
rect 469576 431853 469582 431917
rect 469026 431837 469582 431853
rect 469026 431773 469032 431837
rect 469096 431773 469112 431837
rect 469176 431773 469192 431837
rect 469256 431773 469272 431837
rect 469336 431773 469352 431837
rect 469416 431773 469432 431837
rect 469496 431773 469512 431837
rect 469576 431773 469582 431837
rect 473670 431836 473676 431900
rect 473740 431898 473746 431900
rect 474273 431898 474339 431901
rect 473740 431896 474339 431898
rect 473740 431840 474278 431896
rect 474334 431840 474339 431896
rect 473740 431838 474339 431840
rect 473740 431836 473746 431838
rect 474273 431835 474339 431838
rect 487654 431836 487660 431900
rect 487724 431898 487730 431900
rect 488073 431898 488139 431901
rect 487724 431896 488139 431898
rect 487724 431840 488078 431896
rect 488134 431840 488139 431896
rect 487724 431838 488139 431840
rect 487724 431836 487730 431838
rect 488073 431835 488139 431838
rect 469026 431757 469582 431773
rect 469026 431693 469032 431757
rect 469096 431693 469112 431757
rect 469176 431693 469192 431757
rect 469256 431693 469272 431757
rect 469336 431693 469352 431757
rect 469416 431693 469432 431757
rect 469496 431693 469512 431757
rect 469576 431693 469582 431757
rect 469026 431692 469582 431693
rect 478097 431626 478163 431629
rect 478454 431626 478460 431628
rect 478097 431624 478460 431626
rect 478097 431568 478102 431624
rect 478158 431568 478460 431624
rect 478097 431566 478460 431568
rect 478097 431563 478163 431566
rect 478454 431564 478460 431566
rect 478524 431564 478530 431628
rect 583520 431476 584960 431716
rect 470266 430912 470822 430913
rect 470266 430848 470272 430912
rect 470336 430848 470352 430912
rect 470416 430848 470432 430912
rect 470496 430848 470512 430912
rect 470576 430848 470592 430912
rect 470656 430848 470672 430912
rect 470736 430848 470752 430912
rect 470816 430848 470822 430912
rect 470266 430832 470822 430848
rect 470266 430768 470272 430832
rect 470336 430768 470352 430832
rect 470416 430768 470432 430832
rect 470496 430768 470512 430832
rect 470576 430768 470592 430832
rect 470656 430768 470672 430832
rect 470736 430768 470752 430832
rect 470816 430768 470822 430832
rect 470266 430752 470822 430768
rect 470266 430688 470272 430752
rect 470336 430688 470352 430752
rect 470416 430688 470432 430752
rect 470496 430688 470512 430752
rect 470576 430688 470592 430752
rect 470656 430688 470672 430752
rect 470736 430688 470752 430752
rect 470816 430688 470822 430752
rect 470266 430672 470822 430688
rect 470266 430608 470272 430672
rect 470336 430608 470352 430672
rect 470416 430608 470432 430672
rect 470496 430608 470512 430672
rect 470576 430608 470592 430672
rect 470656 430608 470672 430672
rect 470736 430608 470752 430672
rect 470816 430608 470822 430672
rect 470266 430607 470822 430608
rect 478965 427954 479031 427957
rect 480110 427954 480116 427956
rect 478965 427952 480116 427954
rect 478965 427896 478970 427952
rect 479026 427896 480116 427952
rect 478965 427894 480116 427896
rect 478965 427891 479031 427894
rect 480110 427892 480116 427894
rect 480180 427892 480186 427956
rect 485773 427954 485839 427957
rect 486550 427954 486556 427956
rect 485773 427952 486556 427954
rect 485773 427896 485778 427952
rect 485834 427896 486556 427952
rect 485773 427894 486556 427896
rect 485773 427891 485839 427894
rect 486550 427892 486556 427894
rect 486620 427892 486626 427956
rect 536741 424418 536807 424421
rect 538078 424418 538138 431188
rect 536741 424416 538138 424418
rect 536741 424360 536746 424416
rect 536802 424388 538138 424416
rect 536802 424360 538108 424388
rect 536741 424358 538108 424360
rect 536741 424355 536807 424358
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 470266 412084 470822 412085
rect 470266 412020 470272 412084
rect 470336 412020 470352 412084
rect 470416 412020 470432 412084
rect 470496 412020 470512 412084
rect 470576 412020 470592 412084
rect 470656 412020 470672 412084
rect 470736 412020 470752 412084
rect 470816 412020 470822 412084
rect 470266 412004 470822 412020
rect 470266 411940 470272 412004
rect 470336 411940 470352 412004
rect 470416 411940 470432 412004
rect 470496 411940 470512 412004
rect 470576 411940 470592 412004
rect 470656 411940 470672 412004
rect 470736 411940 470752 412004
rect 470816 411940 470822 412004
rect 470266 411924 470822 411940
rect 470266 411860 470272 411924
rect 470336 411860 470352 411924
rect 470416 411860 470432 411924
rect 470496 411860 470512 411924
rect 470576 411860 470592 411924
rect 470656 411860 470672 411924
rect 470736 411860 470752 411924
rect 470816 411860 470822 411924
rect 470266 411844 470822 411860
rect 470266 411780 470272 411844
rect 470336 411780 470352 411844
rect 470416 411780 470432 411844
rect 470496 411780 470512 411844
rect 470576 411780 470592 411844
rect 470656 411780 470672 411844
rect 470736 411780 470752 411844
rect 470816 411780 470822 411844
rect 470266 411779 470822 411780
rect 469026 410998 469582 410999
rect 469026 410934 469032 410998
rect 469096 410934 469112 410998
rect 469176 410934 469192 410998
rect 469256 410934 469272 410998
rect 469336 410934 469352 410998
rect 469416 410934 469432 410998
rect 469496 410934 469512 410998
rect 469576 410934 469582 410998
rect 473721 410956 473787 410957
rect 469026 410918 469582 410934
rect 469026 410854 469032 410918
rect 469096 410854 469112 410918
rect 469176 410854 469192 410918
rect 469256 410854 469272 410918
rect 469336 410854 469352 410918
rect 469416 410854 469432 410918
rect 469496 410854 469512 410918
rect 469576 410854 469582 410918
rect 473670 410892 473676 410956
rect 473740 410954 473787 410956
rect 473740 410952 473832 410954
rect 473782 410896 473832 410952
rect 473740 410894 473832 410896
rect 473740 410892 473787 410894
rect 473721 410891 473787 410892
rect 469026 410838 469582 410854
rect 469026 410774 469032 410838
rect 469096 410774 469112 410838
rect 469176 410774 469192 410838
rect 469256 410774 469272 410838
rect 469336 410774 469352 410838
rect 469416 410774 469432 410838
rect 469496 410774 469512 410838
rect 469576 410774 469582 410838
rect 469026 410758 469582 410774
rect 469026 410694 469032 410758
rect 469096 410694 469112 410758
rect 469176 410694 469192 410758
rect 469256 410694 469272 410758
rect 469336 410694 469352 410758
rect 469416 410694 469432 410758
rect 469496 410694 469512 410758
rect 469576 410694 469582 410758
rect 469026 410693 469582 410694
rect -960 410396 480 410636
rect 484117 410412 484183 410413
rect 484117 410410 484164 410412
rect 484072 410408 484164 410410
rect 484072 410352 484122 410408
rect 484072 410350 484164 410352
rect 484117 410348 484164 410350
rect 484228 410348 484234 410412
rect 484117 410347 484183 410348
rect 478413 410140 478479 410141
rect 481357 410140 481423 410141
rect 487797 410140 487863 410141
rect 478413 410138 478460 410140
rect 478368 410136 478460 410138
rect 478368 410080 478418 410136
rect 478368 410078 478460 410080
rect 478413 410076 478460 410078
rect 478524 410076 478530 410140
rect 481357 410138 481404 410140
rect 481312 410136 481404 410138
rect 481312 410080 481362 410136
rect 481312 410078 481404 410080
rect 481357 410076 481404 410078
rect 481468 410076 481474 410140
rect 487797 410138 487844 410140
rect 487756 410136 487844 410138
rect 487908 410138 487914 410140
rect 488390 410138 488396 410140
rect 487756 410080 487802 410136
rect 487756 410078 487844 410080
rect 487797 410076 487844 410078
rect 487908 410078 488396 410138
rect 487908 410076 487914 410078
rect 488390 410076 488396 410078
rect 488460 410076 488466 410140
rect 478413 410075 478479 410076
rect 481357 410075 481423 410076
rect 487797 410075 487863 410076
rect 470266 409912 470822 409913
rect 470266 409848 470272 409912
rect 470336 409848 470352 409912
rect 470416 409848 470432 409912
rect 470496 409848 470512 409912
rect 470576 409848 470592 409912
rect 470656 409848 470672 409912
rect 470736 409848 470752 409912
rect 470816 409848 470822 409912
rect 470266 409832 470822 409848
rect 470266 409768 470272 409832
rect 470336 409768 470352 409832
rect 470416 409768 470432 409832
rect 470496 409768 470512 409832
rect 470576 409768 470592 409832
rect 470656 409768 470672 409832
rect 470736 409768 470752 409832
rect 470816 409768 470822 409832
rect 470266 409752 470822 409768
rect 470266 409688 470272 409752
rect 470336 409688 470352 409752
rect 470416 409688 470432 409752
rect 470496 409688 470512 409752
rect 470576 409688 470592 409752
rect 470656 409688 470672 409752
rect 470736 409688 470752 409752
rect 470816 409688 470822 409752
rect 470266 409672 470822 409688
rect 470266 409608 470272 409672
rect 470336 409608 470352 409672
rect 470416 409608 470432 409672
rect 470496 409608 470512 409672
rect 470576 409608 470592 409672
rect 470656 409608 470672 409672
rect 470736 409608 470752 409672
rect 470816 409608 470822 409672
rect 470266 409607 470822 409608
rect 535453 409322 535519 409325
rect 535453 409320 538138 409322
rect 535453 409264 535458 409320
rect 535514 409264 538138 409320
rect 535453 409262 538138 409264
rect 535453 409259 535519 409262
rect 538078 408816 538138 409262
rect 541566 409260 541572 409324
rect 541636 409322 541642 409324
rect 541709 409322 541775 409325
rect 544285 409324 544351 409325
rect 544285 409322 544332 409324
rect 541636 409320 541775 409322
rect 541636 409264 541714 409320
rect 541770 409264 541775 409320
rect 541636 409262 541775 409264
rect 544240 409320 544332 409322
rect 544240 409264 544290 409320
rect 544240 409262 544332 409264
rect 541636 409260 541642 409262
rect 541709 409259 541775 409262
rect 544285 409260 544332 409262
rect 544396 409260 544402 409324
rect 544285 409259 544351 409260
rect 480110 407492 480116 407556
rect 480180 407554 480186 407556
rect 480180 407494 538138 407554
rect 480180 407492 480186 407494
rect 538078 407456 538138 407494
rect 481817 407146 481883 407149
rect 482870 407146 482876 407148
rect 481817 407144 482876 407146
rect 481817 407088 481822 407144
rect 481878 407088 482876 407144
rect 481817 407086 482876 407088
rect 481817 407083 481883 407086
rect 482870 407084 482876 407086
rect 482940 407084 482946 407148
rect 485129 407146 485195 407149
rect 485630 407146 485636 407148
rect 485129 407144 485636 407146
rect 485129 407088 485134 407144
rect 485190 407088 485636 407144
rect 485129 407086 485636 407088
rect 485129 407083 485195 407086
rect 485630 407084 485636 407086
rect 485700 407084 485706 407148
rect 535453 406602 535519 406605
rect 535453 406600 538138 406602
rect 535453 406544 535458 406600
rect 535514 406544 538138 406600
rect 535453 406542 538138 406544
rect 535453 406539 535519 406542
rect 538078 406096 538138 406542
rect 547321 404970 547387 404973
rect 583520 404970 584960 405060
rect 547321 404968 584960 404970
rect 547321 404912 547326 404968
rect 547382 404912 584960 404968
rect 547321 404910 584960 404912
rect 547321 404907 547387 404910
rect 583520 404820 584960 404910
rect 535453 404562 535519 404565
rect 538078 404562 538138 404736
rect 535453 404560 538138 404562
rect 535453 404504 535458 404560
rect 535514 404504 538138 404560
rect 535453 404502 538138 404504
rect 535453 404499 535519 404502
rect 535453 403202 535519 403205
rect 538078 403202 538138 403376
rect 535453 403200 538138 403202
rect 535453 403144 535458 403200
rect 535514 403144 538138 403200
rect 535453 403142 538138 403144
rect 535453 403139 535519 403142
rect 536373 401706 536439 401709
rect 538078 401706 538138 402016
rect 536373 401704 538138 401706
rect 536373 401648 536378 401704
rect 536434 401648 538138 401704
rect 536373 401646 538138 401648
rect 536373 401643 536439 401646
rect 536281 400346 536347 400349
rect 538078 400346 538138 400656
rect 536281 400344 538138 400346
rect 536281 400288 536286 400344
rect 536342 400288 538138 400344
rect 536281 400286 538138 400288
rect 536281 400283 536347 400286
rect 535453 399122 535519 399125
rect 538078 399122 538138 399296
rect 535453 399120 538138 399122
rect 535453 399064 535458 399120
rect 535514 399064 538138 399120
rect 535453 399062 538138 399064
rect 535453 399059 535519 399062
rect 547830 398306 547890 398752
rect 549294 398306 549300 398308
rect 547830 398246 549300 398306
rect 549294 398244 549300 398246
rect 549364 398244 549370 398308
rect -960 397340 480 397580
rect 536097 397490 536163 397493
rect 538078 397490 538138 397936
rect 536097 397488 538138 397490
rect 536097 397432 536102 397488
rect 536158 397432 538138 397488
rect 536097 397430 538138 397432
rect 536097 397427 536163 397430
rect 535453 396402 535519 396405
rect 538078 396402 538138 396576
rect 535453 396400 538138 396402
rect 535453 396344 535458 396400
rect 535514 396344 538138 396400
rect 535453 396342 538138 396344
rect 535453 396339 535519 396342
rect 536741 395994 536807 395997
rect 536741 395992 538138 395994
rect 536741 395936 536746 395992
rect 536802 395936 538138 395992
rect 536741 395934 538138 395936
rect 536741 395931 536807 395934
rect 473670 391988 473676 392052
rect 473740 392050 473746 392052
rect 474958 392050 474964 392052
rect 473740 391990 474964 392050
rect 473740 391988 473746 391990
rect 474958 391988 474964 391990
rect 475028 391988 475034 392052
rect 470266 391085 470822 391086
rect 470266 391021 470272 391085
rect 470336 391021 470352 391085
rect 470416 391021 470432 391085
rect 470496 391021 470512 391085
rect 470576 391021 470592 391085
rect 470656 391021 470672 391085
rect 470736 391021 470752 391085
rect 470816 391021 470822 391085
rect 470266 391005 470822 391021
rect 470266 390941 470272 391005
rect 470336 390941 470352 391005
rect 470416 390941 470432 391005
rect 470496 390941 470512 391005
rect 470576 390941 470592 391005
rect 470656 390941 470672 391005
rect 470736 390941 470752 391005
rect 470816 390941 470822 391005
rect 470266 390925 470822 390941
rect 470266 390861 470272 390925
rect 470336 390861 470352 390925
rect 470416 390861 470432 390925
rect 470496 390861 470512 390925
rect 470576 390861 470592 390925
rect 470656 390861 470672 390925
rect 470736 390861 470752 390925
rect 470816 390861 470822 390925
rect 470266 390845 470822 390861
rect 470266 390781 470272 390845
rect 470336 390781 470352 390845
rect 470416 390781 470432 390845
rect 470496 390781 470512 390845
rect 470576 390781 470592 390845
rect 470656 390781 470672 390845
rect 470736 390781 470752 390845
rect 470816 390781 470822 390845
rect 470266 390780 470822 390781
rect 484900 390297 484964 390303
rect 484900 390227 484964 390233
rect 488390 390084 488396 390148
rect 488460 390146 488466 390148
rect 488533 390146 488599 390149
rect 488460 390144 488599 390146
rect 488460 390088 488538 390144
rect 488594 390088 488599 390144
rect 488460 390086 488599 390088
rect 488460 390084 488466 390086
rect 488533 390083 488599 390086
rect 469026 390002 469582 390003
rect 469026 389938 469032 390002
rect 469096 389938 469112 390002
rect 469176 389938 469192 390002
rect 469256 389938 469272 390002
rect 469336 389938 469352 390002
rect 469416 389938 469432 390002
rect 469496 389938 469512 390002
rect 469576 389938 469582 390002
rect 469026 389922 469582 389938
rect 469026 389858 469032 389922
rect 469096 389858 469112 389922
rect 469176 389858 469192 389922
rect 469256 389858 469272 389922
rect 469336 389858 469352 389922
rect 469416 389858 469432 389922
rect 469496 389858 469512 389922
rect 469576 389858 469582 389922
rect 469026 389842 469582 389858
rect 469026 389778 469032 389842
rect 469096 389778 469112 389842
rect 469176 389778 469192 389842
rect 469256 389778 469272 389842
rect 469336 389778 469352 389842
rect 469416 389778 469432 389842
rect 469496 389778 469512 389842
rect 469576 389778 469582 389842
rect 469026 389762 469582 389778
rect 469026 389698 469032 389762
rect 469096 389698 469112 389762
rect 469176 389698 469192 389762
rect 469256 389698 469272 389762
rect 469336 389698 469352 389762
rect 469416 389698 469432 389762
rect 469496 389698 469512 389762
rect 469576 389698 469582 389762
rect 469026 389697 469582 389698
rect 481766 389404 481772 389468
rect 481836 389466 481842 389468
rect 482093 389466 482159 389469
rect 481836 389464 482159 389466
rect 481836 389408 482098 389464
rect 482154 389408 482159 389464
rect 481836 389406 482159 389408
rect 481836 389404 481842 389406
rect 482093 389403 482159 389406
rect 474917 389332 474983 389333
rect 478629 389332 478695 389333
rect 474917 389330 474964 389332
rect 474872 389328 474964 389330
rect 474872 389272 474922 389328
rect 474872 389270 474964 389272
rect 474917 389268 474964 389270
rect 475028 389268 475034 389332
rect 478629 389330 478644 389332
rect 478552 389328 478644 389330
rect 478552 389272 478634 389328
rect 478552 389270 478644 389272
rect 478629 389268 478644 389270
rect 478708 389268 478714 389332
rect 474917 389267 474983 389268
rect 478629 389267 478695 389268
rect 470266 388912 470822 388913
rect 470266 388848 470272 388912
rect 470336 388848 470352 388912
rect 470416 388848 470432 388912
rect 470496 388848 470512 388912
rect 470576 388848 470592 388912
rect 470656 388848 470672 388912
rect 470736 388848 470752 388912
rect 470816 388848 470822 388912
rect 470266 388832 470822 388848
rect 470266 388768 470272 388832
rect 470336 388768 470352 388832
rect 470416 388768 470432 388832
rect 470496 388768 470512 388832
rect 470576 388768 470592 388832
rect 470656 388768 470672 388832
rect 470736 388768 470752 388832
rect 470816 388768 470822 388832
rect 470266 388752 470822 388768
rect 470266 388688 470272 388752
rect 470336 388688 470352 388752
rect 470416 388688 470432 388752
rect 470496 388688 470512 388752
rect 470576 388688 470592 388752
rect 470656 388688 470672 388752
rect 470736 388688 470752 388752
rect 470816 388688 470822 388752
rect 470266 388672 470822 388688
rect 470266 388608 470272 388672
rect 470336 388608 470352 388672
rect 470416 388608 470432 388672
rect 470496 388608 470512 388672
rect 470576 388608 470592 388672
rect 470656 388608 470672 388672
rect 470736 388608 470752 388672
rect 470816 388608 470822 388672
rect 470266 388607 470822 388608
rect 536189 388378 536255 388381
rect 538078 388378 538138 395934
rect 583520 391628 584960 391868
rect 536189 388376 538138 388378
rect 536189 388320 536194 388376
rect 536250 388320 538138 388376
rect 536189 388318 538138 388320
rect 536189 388315 536255 388318
rect 486734 386412 486740 386476
rect 486804 386474 486810 386476
rect 486877 386474 486943 386477
rect 486804 386472 486943 386474
rect 486804 386416 486882 386472
rect 486938 386416 486943 386472
rect 486804 386414 486943 386416
rect 486804 386412 486810 386414
rect 486877 386411 486943 386414
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect 544469 373420 544535 373421
rect 544469 373418 544516 373420
rect 544424 373416 544516 373418
rect 544424 373360 544474 373416
rect 544424 373358 544516 373360
rect 544469 373356 544516 373358
rect 544580 373356 544586 373420
rect 544469 373355 544535 373356
rect 541566 373084 541572 373148
rect 541636 373146 541642 373148
rect 541709 373146 541775 373149
rect 541636 373144 541775 373146
rect 541636 373088 541714 373144
rect 541770 373088 541775 373144
rect 541636 373086 541775 373088
rect 541636 373084 541642 373086
rect 541709 373083 541775 373086
rect 535453 372874 535519 372877
rect 535453 372872 538108 372874
rect 535453 372816 535458 372872
rect 535514 372816 538108 372872
rect 535453 372814 538108 372816
rect 535453 372811 535519 372814
rect 535453 371514 535519 371517
rect 535453 371512 538108 371514
rect -960 371228 480 371468
rect 535453 371456 535458 371512
rect 535514 371456 538108 371512
rect 535453 371454 538108 371456
rect 535453 371451 535519 371454
rect 482870 370092 482876 370156
rect 482940 370154 482946 370156
rect 482940 370094 538108 370154
rect 482940 370092 482946 370094
rect 535453 368794 535519 368797
rect 535453 368792 538108 368794
rect 535453 368736 535458 368792
rect 535514 368736 538108 368792
rect 535453 368734 538108 368736
rect 535453 368731 535519 368734
rect 535453 367434 535519 367437
rect 535453 367432 538108 367434
rect 535453 367376 535458 367432
rect 535514 367376 538108 367432
rect 535453 367374 538108 367376
rect 535453 367371 535519 367374
rect 535453 366074 535519 366077
rect 535453 366072 538108 366074
rect 535453 366016 535458 366072
rect 535514 366016 538108 366072
rect 535453 366014 538108 366016
rect 535453 366011 535519 366014
rect 583520 364972 584960 365212
rect 536557 364714 536623 364717
rect 536557 364712 538108 364714
rect 536557 364656 536562 364712
rect 536618 364656 538108 364712
rect 536557 364654 538108 364656
rect 536557 364651 536623 364654
rect 536465 363354 536531 363357
rect 536465 363352 538108 363354
rect 536465 363296 536470 363352
rect 536526 363296 538108 363352
rect 536465 363294 538108 363296
rect 536465 363291 536531 363294
rect 549294 362810 549300 362812
rect 547860 362750 549300 362810
rect 549294 362748 549300 362750
rect 549364 362748 549370 362812
rect 535453 361994 535519 361997
rect 535453 361992 538108 361994
rect 535453 361936 535458 361992
rect 535514 361936 538108 361992
rect 535453 361934 538108 361936
rect 535453 361931 535519 361934
rect 535913 360634 535979 360637
rect 535913 360632 538108 360634
rect 535913 360576 535918 360632
rect 535974 360576 538108 360632
rect 535913 360574 538108 360576
rect 535913 360571 535979 360574
rect 536189 359274 536255 359277
rect 536189 359272 538108 359274
rect 536189 359216 536194 359272
rect 536250 359244 538108 359272
rect 536250 359216 538138 359244
rect 536189 359214 538138 359216
rect 536189 359211 536255 359214
rect -960 358308 480 358548
rect 470266 358485 470822 358486
rect 470266 358421 470272 358485
rect 470336 358421 470352 358485
rect 470416 358421 470432 358485
rect 470496 358421 470512 358485
rect 470576 358421 470592 358485
rect 470656 358421 470672 358485
rect 470736 358421 470752 358485
rect 470816 358421 470822 358485
rect 470266 358405 470822 358421
rect 470266 358341 470272 358405
rect 470336 358341 470352 358405
rect 470416 358341 470432 358405
rect 470496 358341 470512 358405
rect 470576 358341 470592 358405
rect 470656 358341 470672 358405
rect 470736 358341 470752 358405
rect 470816 358341 470822 358405
rect 470266 358325 470822 358341
rect 470266 358261 470272 358325
rect 470336 358261 470352 358325
rect 470416 358261 470432 358325
rect 470496 358261 470512 358325
rect 470576 358261 470592 358325
rect 470656 358261 470672 358325
rect 470736 358261 470752 358325
rect 470816 358261 470822 358325
rect 470266 358245 470822 358261
rect 470266 358181 470272 358245
rect 470336 358181 470352 358245
rect 470416 358181 470432 358245
rect 470496 358181 470512 358245
rect 470576 358181 470592 358245
rect 470656 358181 470672 358245
rect 470736 358181 470752 358245
rect 470816 358181 470822 358245
rect 470266 358180 470822 358181
rect 478638 357988 478644 358052
rect 478708 358050 478714 358052
rect 478873 358050 478939 358053
rect 481817 358052 481883 358053
rect 484945 358052 485011 358053
rect 478708 358048 478939 358050
rect 478708 357992 478878 358048
rect 478934 357992 478939 358048
rect 478708 357990 478939 357992
rect 478708 357988 478714 357990
rect 478873 357987 478939 357990
rect 481766 357988 481772 358052
rect 481836 358050 481883 358052
rect 481836 358048 481928 358050
rect 481878 357992 481928 358048
rect 481836 357990 481928 357992
rect 481836 357988 481883 357990
rect 484894 357988 484900 358052
rect 484964 358050 485011 358052
rect 488349 358052 488415 358053
rect 488349 358050 488396 358052
rect 484964 358048 485056 358050
rect 485006 357992 485056 358048
rect 484964 357990 485056 357992
rect 488304 358048 488396 358050
rect 488304 357992 488354 358048
rect 488304 357990 488396 357992
rect 484964 357988 485011 357990
rect 481817 357987 481883 357988
rect 484945 357987 485011 357988
rect 488349 357988 488396 357990
rect 488460 357988 488466 358052
rect 488349 357987 488415 357988
rect 475009 357508 475075 357509
rect 474958 357444 474964 357508
rect 475028 357506 475075 357508
rect 475028 357504 475120 357506
rect 475070 357448 475120 357504
rect 475028 357446 475120 357448
rect 475028 357444 475075 357446
rect 475009 357443 475075 357444
rect 469026 357399 469582 357400
rect 469026 357335 469032 357399
rect 469096 357335 469112 357399
rect 469176 357335 469192 357399
rect 469256 357335 469272 357399
rect 469336 357335 469352 357399
rect 469416 357335 469432 357399
rect 469496 357335 469512 357399
rect 469576 357335 469582 357399
rect 469026 357319 469582 357335
rect 469026 357255 469032 357319
rect 469096 357255 469112 357319
rect 469176 357255 469192 357319
rect 469256 357255 469272 357319
rect 469336 357255 469352 357319
rect 469416 357255 469432 357319
rect 469496 357255 469512 357319
rect 469576 357255 469582 357319
rect 469026 357239 469582 357255
rect 469026 357175 469032 357239
rect 469096 357175 469112 357239
rect 469176 357175 469192 357239
rect 469256 357175 469272 357239
rect 469336 357175 469352 357239
rect 469416 357175 469432 357239
rect 469496 357175 469512 357239
rect 469576 357175 469582 357239
rect 469026 357159 469582 357175
rect 469026 357095 469032 357159
rect 469096 357095 469112 357159
rect 469176 357095 469192 357159
rect 469256 357095 469272 357159
rect 469336 357095 469352 357159
rect 469416 357095 469432 357159
rect 469496 357095 469512 357159
rect 469576 357095 469582 357159
rect 469026 357094 469582 357095
rect 470266 356312 470822 356313
rect 470266 356248 470272 356312
rect 470336 356248 470352 356312
rect 470416 356248 470432 356312
rect 470496 356248 470512 356312
rect 470576 356248 470592 356312
rect 470656 356248 470672 356312
rect 470736 356248 470752 356312
rect 470816 356248 470822 356312
rect 470266 356232 470822 356248
rect 470266 356168 470272 356232
rect 470336 356168 470352 356232
rect 470416 356168 470432 356232
rect 470496 356168 470512 356232
rect 470576 356168 470592 356232
rect 470656 356168 470672 356232
rect 470736 356168 470752 356232
rect 470816 356168 470822 356232
rect 470266 356152 470822 356168
rect 470266 356088 470272 356152
rect 470336 356088 470352 356152
rect 470416 356088 470432 356152
rect 470496 356088 470512 356152
rect 470576 356088 470592 356152
rect 470656 356088 470672 356152
rect 470736 356088 470752 356152
rect 470816 356088 470822 356152
rect 470266 356072 470822 356088
rect 470266 356008 470272 356072
rect 470336 356008 470352 356072
rect 470416 356008 470432 356072
rect 470496 356008 470512 356072
rect 470576 356008 470592 356072
rect 470656 356008 470672 356072
rect 470736 356008 470752 356072
rect 470816 356008 470822 356072
rect 470266 356007 470822 356008
rect 536741 352474 536807 352477
rect 538078 352474 538138 359214
rect 536741 352472 538138 352474
rect 536741 352416 536746 352472
rect 536802 352444 538138 352472
rect 536802 352416 538108 352444
rect 536741 352414 538108 352416
rect 536741 352411 536807 352414
rect 544326 351868 544332 351932
rect 544396 351930 544402 351932
rect 583520 351930 584960 352020
rect 544396 351870 584960 351930
rect 544396 351868 544402 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 473670 343708 473676 343772
rect 473740 343770 473746 343772
rect 474958 343770 474964 343772
rect 473740 343710 474964 343770
rect 473740 343708 473746 343710
rect 474958 343708 474964 343710
rect 475028 343708 475034 343772
rect 470266 342484 470822 342485
rect 470266 342420 470272 342484
rect 470336 342420 470352 342484
rect 470416 342420 470432 342484
rect 470496 342420 470512 342484
rect 470576 342420 470592 342484
rect 470656 342420 470672 342484
rect 470736 342420 470752 342484
rect 470816 342420 470822 342484
rect 470266 342404 470822 342420
rect 470266 342340 470272 342404
rect 470336 342340 470352 342404
rect 470416 342340 470432 342404
rect 470496 342340 470512 342404
rect 470576 342340 470592 342404
rect 470656 342340 470672 342404
rect 470736 342340 470752 342404
rect 470816 342340 470822 342404
rect 470266 342324 470822 342340
rect 470266 342260 470272 342324
rect 470336 342260 470352 342324
rect 470416 342260 470432 342324
rect 470496 342260 470512 342324
rect 470576 342260 470592 342324
rect 470656 342260 470672 342324
rect 470736 342260 470752 342324
rect 470816 342260 470822 342324
rect 470266 342244 470822 342260
rect 470266 342180 470272 342244
rect 470336 342180 470352 342244
rect 470416 342180 470432 342244
rect 470496 342180 470512 342244
rect 470576 342180 470592 342244
rect 470656 342180 470672 342244
rect 470736 342180 470752 342244
rect 470816 342180 470822 342244
rect 470266 342179 470822 342180
rect 469026 341397 469582 341398
rect 469026 341333 469032 341397
rect 469096 341333 469112 341397
rect 469176 341333 469192 341397
rect 469256 341333 469272 341397
rect 469336 341333 469352 341397
rect 469416 341333 469432 341397
rect 469496 341333 469512 341397
rect 469576 341333 469582 341397
rect 469026 341317 469582 341333
rect 469026 341253 469032 341317
rect 469096 341253 469112 341317
rect 469176 341253 469192 341317
rect 469256 341253 469272 341317
rect 469336 341253 469352 341317
rect 469416 341253 469432 341317
rect 469496 341253 469512 341317
rect 469576 341253 469582 341317
rect 469026 341237 469582 341253
rect 469026 341173 469032 341237
rect 469096 341173 469112 341237
rect 469176 341173 469192 341237
rect 469256 341173 469272 341237
rect 469336 341173 469352 341237
rect 469416 341173 469432 341237
rect 469496 341173 469512 341237
rect 469576 341173 469582 341237
rect 469026 341157 469582 341173
rect 469026 341093 469032 341157
rect 469096 341093 469112 341157
rect 469176 341093 469192 341157
rect 469256 341093 469272 341157
rect 469336 341093 469352 341157
rect 469416 341093 469432 341157
rect 469496 341093 469512 341157
rect 469576 341093 469582 341157
rect 469026 341092 469582 341093
rect 477910 341050 477976 341053
rect 478454 341050 478460 341052
rect 477910 341048 478460 341050
rect 477910 340992 477915 341048
rect 477971 340992 478460 341048
rect 477910 340990 478460 340992
rect 477910 340987 477976 340990
rect 478454 340988 478460 340990
rect 478524 340988 478530 341052
rect 481227 341050 481293 341053
rect 481398 341050 481404 341052
rect 481227 341048 481404 341050
rect 481227 340992 481232 341048
rect 481288 340992 481404 341048
rect 481227 340990 481404 340992
rect 481227 340987 481293 340990
rect 481398 340988 481404 340990
rect 481468 340988 481474 341052
rect 484158 340988 484164 341052
rect 484228 341050 484234 341052
rect 484393 341050 484459 341053
rect 484228 341048 484459 341050
rect 484228 340992 484398 341048
rect 484454 340992 484459 341048
rect 484228 340990 484459 340992
rect 484228 340988 484234 340990
rect 484393 340987 484459 340990
rect 487889 341050 487955 341053
rect 488022 341050 488028 341052
rect 487889 341048 488028 341050
rect 487889 340992 487894 341048
rect 487950 340992 488028 341048
rect 487889 340990 488028 340992
rect 487889 340987 487955 340990
rect 488022 340988 488028 340990
rect 488092 340988 488098 341052
rect 473670 340444 473676 340508
rect 473740 340506 473746 340508
rect 474549 340506 474615 340509
rect 473740 340504 474615 340506
rect 473740 340448 474554 340504
rect 474610 340448 474615 340504
rect 473740 340446 474615 340448
rect 473740 340444 473746 340446
rect 474549 340443 474615 340446
rect 470266 340312 470822 340313
rect 470266 340248 470272 340312
rect 470336 340248 470352 340312
rect 470416 340248 470432 340312
rect 470496 340248 470512 340312
rect 470576 340248 470592 340312
rect 470656 340248 470672 340312
rect 470736 340248 470752 340312
rect 470816 340248 470822 340312
rect 470266 340232 470822 340248
rect 470266 340168 470272 340232
rect 470336 340168 470352 340232
rect 470416 340168 470432 340232
rect 470496 340168 470512 340232
rect 470576 340168 470592 340232
rect 470656 340168 470672 340232
rect 470736 340168 470752 340232
rect 470816 340168 470822 340232
rect 470266 340152 470822 340168
rect 470266 340088 470272 340152
rect 470336 340088 470352 340152
rect 470416 340088 470432 340152
rect 470496 340088 470512 340152
rect 470576 340088 470592 340152
rect 470656 340088 470672 340152
rect 470736 340088 470752 340152
rect 470816 340088 470822 340152
rect 470266 340072 470822 340088
rect 470266 340008 470272 340072
rect 470336 340008 470352 340072
rect 470416 340008 470432 340072
rect 470496 340008 470512 340072
rect 470576 340008 470592 340072
rect 470656 340008 470672 340072
rect 470736 340008 470752 340072
rect 470816 340008 470822 340072
rect 470266 340007 470822 340008
rect 541566 339492 541572 339556
rect 541636 339554 541642 339556
rect 541709 339554 541775 339557
rect 541636 339552 541775 339554
rect 541636 339496 541714 339552
rect 541770 339496 541775 339552
rect 541636 339494 541775 339496
rect 541636 339492 541642 339494
rect 541709 339491 541775 339494
rect 544193 339554 544259 339557
rect 544326 339554 544332 339556
rect 544193 339552 544332 339554
rect 544193 339496 544198 339552
rect 544254 339496 544332 339552
rect 544193 339494 544332 339496
rect 544193 339491 544259 339494
rect 544326 339492 544332 339494
rect 544396 339492 544402 339556
rect 583520 338452 584960 338692
rect 535453 336834 535519 336837
rect 535453 336832 538108 336834
rect 535453 336776 535458 336832
rect 535514 336776 538108 336832
rect 535453 336774 538108 336776
rect 535453 336771 535519 336774
rect 486550 335412 486556 335476
rect 486620 335474 486626 335476
rect 486620 335414 538108 335474
rect 486620 335412 486626 335414
rect 485630 334052 485636 334116
rect 485700 334114 485706 334116
rect 485700 334054 538108 334114
rect 485700 334052 485706 334054
rect 486734 332692 486740 332756
rect 486804 332754 486810 332756
rect 486804 332694 538108 332754
rect 486804 332692 486810 332694
rect -960 332196 480 332436
rect 535453 331394 535519 331397
rect 535453 331392 538108 331394
rect 535453 331336 535458 331392
rect 535514 331336 538108 331392
rect 535453 331334 538108 331336
rect 535453 331331 535519 331334
rect 535453 330034 535519 330037
rect 535453 330032 538108 330034
rect 535453 329976 535458 330032
rect 535514 329976 538108 330032
rect 535453 329974 538108 329976
rect 535453 329971 535519 329974
rect 536005 328674 536071 328677
rect 536005 328672 538108 328674
rect 536005 328616 536010 328672
rect 536066 328616 538108 328672
rect 536005 328614 538108 328616
rect 536005 328611 536071 328614
rect 536649 327314 536715 327317
rect 536649 327312 538108 327314
rect 536649 327256 536654 327312
rect 536710 327256 538108 327312
rect 536649 327254 538108 327256
rect 536649 327251 536715 327254
rect 549294 326770 549300 326772
rect 547860 326710 549300 326770
rect 549294 326708 549300 326710
rect 549364 326708 549370 326772
rect 535453 325954 535519 325957
rect 535453 325952 538108 325954
rect 535453 325896 535458 325952
rect 535514 325896 538108 325952
rect 535453 325894 538108 325896
rect 535453 325891 535519 325894
rect 583520 325124 584960 325364
rect 536373 324594 536439 324597
rect 536373 324592 538108 324594
rect 536373 324536 536378 324592
rect 536434 324536 538108 324592
rect 536373 324534 538108 324536
rect 536373 324531 536439 324534
rect 536741 323234 536807 323237
rect 536741 323232 538108 323234
rect 536741 323176 536746 323232
rect 536802 323204 538108 323232
rect 536802 323176 538138 323204
rect 536741 323174 538138 323176
rect 536741 323171 536807 323174
rect 470266 322484 470822 322485
rect 470266 322420 470272 322484
rect 470336 322420 470352 322484
rect 470416 322420 470432 322484
rect 470496 322420 470512 322484
rect 470576 322420 470592 322484
rect 470656 322420 470672 322484
rect 470736 322420 470752 322484
rect 470816 322420 470822 322484
rect 470266 322404 470822 322420
rect 470266 322340 470272 322404
rect 470336 322340 470352 322404
rect 470416 322340 470432 322404
rect 470496 322340 470512 322404
rect 470576 322340 470592 322404
rect 470656 322340 470672 322404
rect 470736 322340 470752 322404
rect 470816 322340 470822 322404
rect 470266 322324 470822 322340
rect 470266 322260 470272 322324
rect 470336 322260 470352 322324
rect 470416 322260 470432 322324
rect 470496 322260 470512 322324
rect 470576 322260 470592 322324
rect 470656 322260 470672 322324
rect 470736 322260 470752 322324
rect 470816 322260 470822 322324
rect 470266 322244 470822 322260
rect 470266 322180 470272 322244
rect 470336 322180 470352 322244
rect 470416 322180 470432 322244
rect 470496 322180 470512 322244
rect 470576 322180 470592 322244
rect 470656 322180 470672 322244
rect 470736 322180 470752 322244
rect 470816 322180 470822 322244
rect 470266 322179 470822 322180
rect 469026 321397 469582 321398
rect 469026 321333 469032 321397
rect 469096 321333 469112 321397
rect 469176 321333 469192 321397
rect 469256 321333 469272 321397
rect 469336 321333 469352 321397
rect 469416 321333 469432 321397
rect 469496 321333 469512 321397
rect 469576 321333 469582 321397
rect 469026 321317 469582 321333
rect 469026 321253 469032 321317
rect 469096 321253 469112 321317
rect 469176 321253 469192 321317
rect 469256 321253 469272 321317
rect 469336 321253 469352 321317
rect 469416 321253 469432 321317
rect 469496 321253 469512 321317
rect 469576 321253 469582 321317
rect 473670 321268 473676 321332
rect 473740 321330 473746 321332
rect 474273 321330 474339 321333
rect 473740 321328 474339 321330
rect 473740 321272 474278 321328
rect 474334 321272 474339 321328
rect 473740 321270 474339 321272
rect 473740 321268 473746 321270
rect 474273 321267 474339 321270
rect 484158 321268 484164 321332
rect 484228 321330 484234 321332
rect 484577 321330 484643 321333
rect 484228 321328 484643 321330
rect 484228 321272 484582 321328
rect 484638 321272 484643 321328
rect 484228 321270 484643 321272
rect 484228 321268 484234 321270
rect 484577 321267 484643 321270
rect 469026 321237 469582 321253
rect 469026 321173 469032 321237
rect 469096 321173 469112 321237
rect 469176 321173 469192 321237
rect 469256 321173 469272 321237
rect 469336 321173 469352 321237
rect 469416 321173 469432 321237
rect 469496 321173 469512 321237
rect 469576 321173 469582 321237
rect 469026 321157 469582 321173
rect 469026 321093 469032 321157
rect 469096 321093 469112 321157
rect 469176 321093 469192 321157
rect 469256 321093 469272 321157
rect 469336 321093 469352 321157
rect 469416 321093 469432 321157
rect 469496 321093 469512 321157
rect 469576 321093 469582 321157
rect 469026 321092 469582 321093
rect 488022 320996 488028 321060
rect 488092 321058 488098 321060
rect 488165 321058 488231 321061
rect 488092 321056 488231 321058
rect 488092 321000 488170 321056
rect 488226 321000 488231 321056
rect 488092 320998 488231 321000
rect 488092 320996 488098 320998
rect 488165 320995 488231 320998
rect 478137 320922 478203 320925
rect 481541 320924 481607 320925
rect 478638 320922 478644 320924
rect 478137 320920 478644 320922
rect 478137 320864 478142 320920
rect 478198 320864 478644 320920
rect 478137 320862 478644 320864
rect 478137 320859 478203 320862
rect 478638 320860 478644 320862
rect 478708 320860 478714 320924
rect 481541 320922 481588 320924
rect 481496 320920 481588 320922
rect 481496 320864 481546 320920
rect 481496 320862 481588 320864
rect 481541 320860 481588 320862
rect 481652 320860 481658 320924
rect 481541 320859 481607 320860
rect 470266 320312 470822 320313
rect 470266 320248 470272 320312
rect 470336 320248 470352 320312
rect 470416 320248 470432 320312
rect 470496 320248 470512 320312
rect 470576 320248 470592 320312
rect 470656 320248 470672 320312
rect 470736 320248 470752 320312
rect 470816 320248 470822 320312
rect 470266 320232 470822 320248
rect 470266 320168 470272 320232
rect 470336 320168 470352 320232
rect 470416 320168 470432 320232
rect 470496 320168 470512 320232
rect 470576 320168 470592 320232
rect 470656 320168 470672 320232
rect 470736 320168 470752 320232
rect 470816 320168 470822 320232
rect 470266 320152 470822 320168
rect 470266 320088 470272 320152
rect 470336 320088 470352 320152
rect 470416 320088 470432 320152
rect 470496 320088 470512 320152
rect 470576 320088 470592 320152
rect 470656 320088 470672 320152
rect 470736 320088 470752 320152
rect 470816 320088 470822 320152
rect 470266 320072 470822 320088
rect 470266 320008 470272 320072
rect 470336 320008 470352 320072
rect 470416 320008 470432 320072
rect 470496 320008 470512 320072
rect 470576 320008 470592 320072
rect 470656 320008 470672 320072
rect 470736 320008 470752 320072
rect 470816 320008 470822 320072
rect 470266 320007 470822 320008
rect -960 319140 480 319380
rect 536741 316434 536807 316437
rect 538078 316434 538138 323174
rect 536741 316432 538138 316434
rect 536741 316376 536746 316432
rect 536802 316404 538138 316432
rect 536802 316376 538108 316404
rect 536741 316374 538108 316376
rect 536741 316371 536807 316374
rect 583520 311932 584960 312172
rect 470266 307084 470822 307085
rect 470266 307020 470272 307084
rect 470336 307020 470352 307084
rect 470416 307020 470432 307084
rect 470496 307020 470512 307084
rect 470576 307020 470592 307084
rect 470656 307020 470672 307084
rect 470736 307020 470752 307084
rect 470816 307020 470822 307084
rect 470266 307004 470822 307020
rect 470266 306940 470272 307004
rect 470336 306940 470352 307004
rect 470416 306940 470432 307004
rect 470496 306940 470512 307004
rect 470576 306940 470592 307004
rect 470656 306940 470672 307004
rect 470736 306940 470752 307004
rect 470816 306940 470822 307004
rect 470266 306924 470822 306940
rect 470266 306860 470272 306924
rect 470336 306860 470352 306924
rect 470416 306860 470432 306924
rect 470496 306860 470512 306924
rect 470576 306860 470592 306924
rect 470656 306860 470672 306924
rect 470736 306860 470752 306924
rect 470816 306860 470822 306924
rect 470266 306844 470822 306860
rect 470266 306780 470272 306844
rect 470336 306780 470352 306844
rect 470416 306780 470432 306844
rect 470496 306780 470512 306844
rect 470576 306780 470592 306844
rect 470656 306780 470672 306844
rect 470736 306780 470752 306844
rect 470816 306780 470822 306844
rect 470266 306779 470822 306780
rect -960 306084 480 306324
rect 487654 306308 487660 306372
rect 487724 306308 487730 306372
rect 487529 306234 487595 306237
rect 487662 306234 487722 306308
rect 487529 306232 487722 306234
rect 487529 306176 487534 306232
rect 487590 306176 487722 306232
rect 487529 306174 487722 306176
rect 487529 306171 487595 306174
rect 480999 306098 481065 306101
rect 481582 306098 481588 306100
rect 480999 306096 481588 306098
rect 480999 306040 481004 306096
rect 481060 306040 481588 306096
rect 480999 306038 481588 306040
rect 480999 306035 481065 306038
rect 481582 306036 481588 306038
rect 481652 306036 481658 306100
rect 469026 305999 469582 306000
rect 469026 305935 469032 305999
rect 469096 305935 469112 305999
rect 469176 305935 469192 305999
rect 469256 305935 469272 305999
rect 469336 305935 469352 305999
rect 469416 305935 469432 305999
rect 469496 305935 469512 305999
rect 469576 305935 469582 305999
rect 473721 305964 473787 305965
rect 469026 305919 469582 305935
rect 469026 305855 469032 305919
rect 469096 305855 469112 305919
rect 469176 305855 469192 305919
rect 469256 305855 469272 305919
rect 469336 305855 469352 305919
rect 469416 305855 469432 305919
rect 469496 305855 469512 305919
rect 469576 305855 469582 305919
rect 473670 305900 473676 305964
rect 473740 305962 473787 305964
rect 473740 305960 473832 305962
rect 473782 305904 473832 305960
rect 473740 305902 473832 305904
rect 473740 305900 473787 305902
rect 473721 305899 473787 305900
rect 469026 305839 469582 305855
rect 469026 305775 469032 305839
rect 469096 305775 469112 305839
rect 469176 305775 469192 305839
rect 469256 305775 469272 305839
rect 469336 305775 469352 305839
rect 469416 305775 469432 305839
rect 469496 305775 469512 305839
rect 469576 305775 469582 305839
rect 469026 305759 469582 305775
rect 469026 305695 469032 305759
rect 469096 305695 469112 305759
rect 469176 305695 469192 305759
rect 469256 305695 469272 305759
rect 469336 305695 469352 305759
rect 469416 305695 469432 305759
rect 469496 305695 469512 305759
rect 469576 305695 469582 305759
rect 469026 305694 469582 305695
rect 477734 305690 477800 305693
rect 478822 305690 478828 305692
rect 477734 305688 478828 305690
rect 477734 305632 477739 305688
rect 477795 305632 478828 305688
rect 477734 305630 478828 305632
rect 477734 305627 477800 305630
rect 478822 305628 478828 305630
rect 478892 305628 478898 305692
rect 484117 305556 484183 305557
rect 484117 305554 484164 305556
rect 484072 305552 484164 305554
rect 484072 305496 484122 305552
rect 484072 305494 484164 305496
rect 484117 305492 484164 305494
rect 484228 305492 484234 305556
rect 484117 305491 484183 305492
rect 470266 304912 470822 304913
rect 470266 304848 470272 304912
rect 470336 304848 470352 304912
rect 470416 304848 470432 304912
rect 470496 304848 470512 304912
rect 470576 304848 470592 304912
rect 470656 304848 470672 304912
rect 470736 304848 470752 304912
rect 470816 304848 470822 304912
rect 470266 304832 470822 304848
rect 470266 304768 470272 304832
rect 470336 304768 470352 304832
rect 470416 304768 470432 304832
rect 470496 304768 470512 304832
rect 470576 304768 470592 304832
rect 470656 304768 470672 304832
rect 470736 304768 470752 304832
rect 470816 304768 470822 304832
rect 470266 304752 470822 304768
rect 470266 304688 470272 304752
rect 470336 304688 470352 304752
rect 470416 304688 470432 304752
rect 470496 304688 470512 304752
rect 470576 304688 470592 304752
rect 470656 304688 470672 304752
rect 470736 304688 470752 304752
rect 470816 304688 470822 304752
rect 470266 304672 470822 304688
rect 470266 304608 470272 304672
rect 470336 304608 470352 304672
rect 470416 304608 470432 304672
rect 470496 304608 470512 304672
rect 470576 304608 470592 304672
rect 470656 304608 470672 304672
rect 470736 304608 470752 304672
rect 470816 304608 470822 304672
rect 470266 304607 470822 304608
rect 544193 303786 544259 303789
rect 544326 303786 544332 303788
rect 544193 303784 544332 303786
rect 544193 303728 544198 303784
rect 544254 303728 544332 303784
rect 544193 303726 544332 303728
rect 544193 303723 544259 303726
rect 544326 303724 544332 303726
rect 544396 303724 544402 303788
rect 541566 303588 541572 303652
rect 541636 303650 541642 303652
rect 541709 303650 541775 303653
rect 547321 303650 547387 303653
rect 541636 303648 547387 303650
rect 541636 303592 541714 303648
rect 541770 303592 547326 303648
rect 547382 303592 547387 303648
rect 541636 303590 547387 303592
rect 541636 303588 541642 303590
rect 541709 303587 541775 303590
rect 547321 303587 547387 303590
rect 535453 300794 535519 300797
rect 535453 300792 538108 300794
rect 535453 300736 535458 300792
rect 535514 300736 538108 300792
rect 535453 300734 538108 300736
rect 535453 300731 535519 300734
rect 547321 300114 547387 300117
rect 580165 300114 580231 300117
rect 547321 300112 580231 300114
rect 547321 300056 547326 300112
rect 547382 300056 580170 300112
rect 580226 300056 580231 300112
rect 547321 300054 580231 300056
rect 547321 300051 547387 300054
rect 580165 300051 580231 300054
rect 535453 299434 535519 299437
rect 535453 299432 538108 299434
rect 535453 299376 535458 299432
rect 535514 299376 538108 299432
rect 535453 299374 538108 299376
rect 535453 299371 535519 299374
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 535453 298074 535519 298077
rect 535453 298072 538108 298074
rect 535453 298016 535458 298072
rect 535514 298016 538108 298072
rect 535453 298014 538108 298016
rect 535453 298011 535519 298014
rect 535453 296714 535519 296717
rect 535453 296712 538108 296714
rect 535453 296656 535458 296712
rect 535514 296656 538108 296712
rect 535453 296654 538108 296656
rect 535453 296651 535519 296654
rect 535545 295354 535611 295357
rect 535545 295352 538108 295354
rect 535545 295296 535550 295352
rect 535606 295296 538108 295352
rect 535545 295294 538108 295296
rect 535545 295291 535611 295294
rect 535453 293994 535519 293997
rect 535453 293992 538108 293994
rect 535453 293936 535458 293992
rect 535514 293936 538108 293992
rect 535453 293934 538108 293936
rect 535453 293931 535519 293934
rect -960 293028 480 293268
rect 535545 292634 535611 292637
rect 535545 292632 538108 292634
rect 535545 292576 535550 292632
rect 535606 292576 538108 292632
rect 535545 292574 538108 292576
rect 535545 292571 535611 292574
rect 535453 291274 535519 291277
rect 535453 291272 538108 291274
rect 535453 291216 535458 291272
rect 535514 291216 538108 291272
rect 535453 291214 538108 291216
rect 535453 291211 535519 291214
rect 549294 290730 549300 290732
rect 547860 290670 549300 290730
rect 549294 290668 549300 290670
rect 549364 290668 549370 290732
rect 535453 289914 535519 289917
rect 535453 289912 538108 289914
rect 535453 289856 535458 289912
rect 535514 289856 538108 289912
rect 535453 289854 538108 289856
rect 535453 289851 535519 289854
rect 473670 289716 473676 289780
rect 473740 289778 473746 289780
rect 476062 289778 476068 289780
rect 473740 289718 476068 289778
rect 473740 289716 473746 289718
rect 476062 289716 476068 289718
rect 476132 289716 476138 289780
rect 484158 289716 484164 289780
rect 484228 289778 484234 289780
rect 485814 289778 485820 289780
rect 484228 289718 485820 289778
rect 484228 289716 484234 289718
rect 485814 289716 485820 289718
rect 485884 289716 485890 289780
rect 535453 288554 535519 288557
rect 535453 288552 538108 288554
rect 535453 288496 535458 288552
rect 535514 288496 538108 288552
rect 535453 288494 538108 288496
rect 535453 288491 535519 288494
rect 470266 287485 470822 287486
rect 470266 287421 470272 287485
rect 470336 287421 470352 287485
rect 470416 287421 470432 287485
rect 470496 287421 470512 287485
rect 470576 287421 470592 287485
rect 470656 287421 470672 287485
rect 470736 287421 470752 287485
rect 470816 287421 470822 287485
rect 470266 287405 470822 287421
rect 470266 287341 470272 287405
rect 470336 287341 470352 287405
rect 470416 287341 470432 287405
rect 470496 287341 470512 287405
rect 470576 287341 470592 287405
rect 470656 287341 470672 287405
rect 470736 287341 470752 287405
rect 470816 287341 470822 287405
rect 470266 287325 470822 287341
rect 470266 287261 470272 287325
rect 470336 287261 470352 287325
rect 470416 287261 470432 287325
rect 470496 287261 470512 287325
rect 470576 287261 470592 287325
rect 470656 287261 470672 287325
rect 470736 287261 470752 287325
rect 470816 287261 470822 287325
rect 470266 287245 470822 287261
rect 470266 287181 470272 287245
rect 470336 287181 470352 287245
rect 470416 287181 470432 287245
rect 470496 287181 470512 287245
rect 470576 287181 470592 287245
rect 470656 287181 470672 287245
rect 470736 287181 470752 287245
rect 470816 287181 470822 287245
rect 470266 287180 470822 287181
rect 536741 287194 536807 287197
rect 536741 287192 538108 287194
rect 536741 287136 536746 287192
rect 536802 287164 538108 287192
rect 536802 287136 538138 287164
rect 536741 287134 538138 287136
rect 536741 287131 536807 287134
rect 478628 286922 478694 286925
rect 478822 286922 478828 286924
rect 478628 286920 478828 286922
rect 478628 286864 478633 286920
rect 478689 286864 478828 286920
rect 478628 286862 478828 286864
rect 478628 286859 478694 286862
rect 478822 286860 478828 286862
rect 478892 286860 478898 286924
rect 488574 286724 488580 286788
rect 488644 286724 488650 286788
rect 488582 286653 488642 286724
rect 474916 286650 474982 286653
rect 476062 286650 476068 286652
rect 474916 286648 476068 286650
rect 474916 286592 474921 286648
rect 474977 286592 476068 286648
rect 474916 286590 476068 286592
rect 474916 286587 474982 286590
rect 476062 286588 476068 286590
rect 476132 286588 476138 286652
rect 488582 286648 488691 286653
rect 488582 286592 488630 286648
rect 488686 286592 488691 286648
rect 488582 286590 488691 286592
rect 488625 286587 488691 286590
rect 469026 286400 469582 286401
rect 469026 286336 469032 286400
rect 469096 286336 469112 286400
rect 469176 286336 469192 286400
rect 469256 286336 469272 286400
rect 469336 286336 469352 286400
rect 469416 286336 469432 286400
rect 469496 286336 469512 286400
rect 469576 286336 469582 286400
rect 469026 286320 469582 286336
rect 469026 286256 469032 286320
rect 469096 286256 469112 286320
rect 469176 286256 469192 286320
rect 469256 286256 469272 286320
rect 469336 286256 469352 286320
rect 469416 286256 469432 286320
rect 469496 286256 469512 286320
rect 469576 286256 469582 286320
rect 469026 286240 469582 286256
rect 469026 286176 469032 286240
rect 469096 286176 469112 286240
rect 469176 286176 469192 286240
rect 469256 286176 469272 286240
rect 469336 286176 469352 286240
rect 469416 286176 469432 286240
rect 469496 286176 469512 286240
rect 469576 286176 469582 286240
rect 469026 286160 469582 286176
rect 469026 286096 469032 286160
rect 469096 286096 469112 286160
rect 469176 286096 469192 286160
rect 469256 286096 469272 286160
rect 469336 286096 469352 286160
rect 469416 286096 469432 286160
rect 469496 286096 469512 286160
rect 469576 286096 469582 286160
rect 469026 286095 469582 286096
rect 482340 285836 482406 285837
rect 485865 285836 485931 285837
rect 482318 285834 482324 285836
rect 482213 285774 482324 285834
rect 482388 285834 482406 285836
rect 482870 285834 482876 285836
rect 482388 285832 482876 285834
rect 482401 285776 482876 285832
rect 482318 285772 482324 285774
rect 482388 285774 482876 285776
rect 482388 285772 482406 285774
rect 482870 285772 482876 285774
rect 482940 285772 482946 285836
rect 485814 285772 485820 285836
rect 485884 285834 485931 285836
rect 485884 285832 485976 285834
rect 485926 285776 485976 285832
rect 485884 285774 485976 285776
rect 485884 285772 485931 285774
rect 482340 285771 482406 285772
rect 485865 285771 485931 285772
rect 470266 285312 470822 285313
rect 470266 285248 470272 285312
rect 470336 285248 470352 285312
rect 470416 285248 470432 285312
rect 470496 285248 470512 285312
rect 470576 285248 470592 285312
rect 470656 285248 470672 285312
rect 470736 285248 470752 285312
rect 470816 285248 470822 285312
rect 470266 285232 470822 285248
rect 470266 285168 470272 285232
rect 470336 285168 470352 285232
rect 470416 285168 470432 285232
rect 470496 285168 470512 285232
rect 470576 285168 470592 285232
rect 470656 285168 470672 285232
rect 470736 285168 470752 285232
rect 470816 285168 470822 285232
rect 470266 285152 470822 285168
rect 470266 285088 470272 285152
rect 470336 285088 470352 285152
rect 470416 285088 470432 285152
rect 470496 285088 470512 285152
rect 470576 285088 470592 285152
rect 470656 285088 470672 285152
rect 470736 285088 470752 285152
rect 470816 285088 470822 285152
rect 470266 285072 470822 285088
rect 470266 285008 470272 285072
rect 470336 285008 470352 285072
rect 470416 285008 470432 285072
rect 470496 285008 470512 285072
rect 470576 285008 470592 285072
rect 470656 285008 470672 285072
rect 470736 285008 470752 285072
rect 470816 285008 470822 285072
rect 470266 285007 470822 285008
rect 538078 280364 538138 287134
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect 470266 267485 470822 267486
rect 470266 267421 470272 267485
rect 470336 267421 470352 267485
rect 470416 267421 470432 267485
rect 470496 267421 470512 267485
rect 470576 267421 470592 267485
rect 470656 267421 470672 267485
rect 470736 267421 470752 267485
rect 470816 267421 470822 267485
rect 470266 267405 470822 267421
rect 470266 267341 470272 267405
rect 470336 267341 470352 267405
rect 470416 267341 470432 267405
rect 470496 267341 470512 267405
rect 470576 267341 470592 267405
rect 470656 267341 470672 267405
rect 470736 267341 470752 267405
rect 470816 267341 470822 267405
rect 470266 267325 470822 267341
rect -960 267052 480 267292
rect 470266 267261 470272 267325
rect 470336 267261 470352 267325
rect 470416 267261 470432 267325
rect 470496 267261 470512 267325
rect 470576 267261 470592 267325
rect 470656 267261 470672 267325
rect 470736 267261 470752 267325
rect 470816 267261 470822 267325
rect 470266 267245 470822 267261
rect 470266 267181 470272 267245
rect 470336 267181 470352 267245
rect 470416 267181 470432 267245
rect 470496 267181 470512 267245
rect 470576 267181 470592 267245
rect 470656 267181 470672 267245
rect 470736 267181 470752 267245
rect 470816 267181 470822 267245
rect 470266 267180 470822 267181
rect 469026 266399 469582 266400
rect 469026 266335 469032 266399
rect 469096 266335 469112 266399
rect 469176 266335 469192 266399
rect 469256 266335 469272 266399
rect 469336 266335 469352 266399
rect 469416 266335 469432 266399
rect 469496 266335 469512 266399
rect 469576 266335 469582 266399
rect 469026 266319 469582 266335
rect 469026 266255 469032 266319
rect 469096 266255 469112 266319
rect 469176 266255 469192 266319
rect 469256 266255 469272 266319
rect 469336 266255 469352 266319
rect 469416 266255 469432 266319
rect 469496 266255 469512 266319
rect 469576 266255 469582 266319
rect 469026 266239 469582 266255
rect 469026 266175 469032 266239
rect 469096 266175 469112 266239
rect 469176 266175 469192 266239
rect 469256 266175 469272 266239
rect 469336 266175 469352 266239
rect 469416 266175 469432 266239
rect 469496 266175 469512 266239
rect 469576 266175 469582 266239
rect 469026 266159 469582 266175
rect 469026 266095 469032 266159
rect 469096 266095 469112 266159
rect 469176 266095 469192 266159
rect 469256 266095 469272 266159
rect 469336 266095 469352 266159
rect 469416 266095 469432 266159
rect 469496 266095 469512 266159
rect 469576 266095 469582 266159
rect 469026 266094 469582 266095
rect 479057 265980 479123 265981
rect 479006 265978 479012 265980
rect 478966 265918 479012 265978
rect 479076 265976 479123 265980
rect 479118 265920 479123 265976
rect 479006 265916 479012 265918
rect 479076 265916 479123 265920
rect 479057 265915 479123 265916
rect 488717 265570 488783 265573
rect 489126 265570 489132 265572
rect 488717 265568 489132 265570
rect 488717 265512 488722 265568
rect 488778 265512 489132 265568
rect 488717 265510 489132 265512
rect 488717 265507 488783 265510
rect 489126 265508 489132 265510
rect 489196 265508 489202 265572
rect 470266 265312 470822 265313
rect 470266 265248 470272 265312
rect 470336 265248 470352 265312
rect 470416 265248 470432 265312
rect 470496 265248 470512 265312
rect 470576 265248 470592 265312
rect 470656 265248 470672 265312
rect 470736 265248 470752 265312
rect 470816 265248 470822 265312
rect 470266 265232 470822 265248
rect 470266 265168 470272 265232
rect 470336 265168 470352 265232
rect 470416 265168 470432 265232
rect 470496 265168 470512 265232
rect 470576 265168 470592 265232
rect 470656 265168 470672 265232
rect 470736 265168 470752 265232
rect 470816 265168 470822 265232
rect 470266 265152 470822 265168
rect 470266 265088 470272 265152
rect 470336 265088 470352 265152
rect 470416 265088 470432 265152
rect 470496 265088 470512 265152
rect 470576 265088 470592 265152
rect 470656 265088 470672 265152
rect 470736 265088 470752 265152
rect 470816 265088 470822 265152
rect 470266 265072 470822 265088
rect 470266 265008 470272 265072
rect 470336 265008 470352 265072
rect 470416 265008 470432 265072
rect 470496 265008 470512 265072
rect 470576 265008 470592 265072
rect 470656 265008 470672 265072
rect 470736 265008 470752 265072
rect 470816 265008 470822 265072
rect 476481 265028 476547 265029
rect 476430 265026 476436 265028
rect 470266 265007 470822 265008
rect 476354 264966 476436 265026
rect 476500 265026 476547 265028
rect 477350 265026 477356 265028
rect 476500 265024 477356 265026
rect 476542 264968 477356 265024
rect 476430 264964 476436 264966
rect 476500 264966 477356 264968
rect 476500 264964 476547 264966
rect 477350 264964 477356 264966
rect 477420 264964 477426 265028
rect 479517 265026 479583 265029
rect 482829 265028 482895 265029
rect 480110 265026 480116 265028
rect 479517 265024 480116 265026
rect 479517 264968 479522 265024
rect 479578 264968 480116 265024
rect 479517 264966 480116 264968
rect 476481 264963 476547 264964
rect 479517 264963 479583 264966
rect 480110 264964 480116 264966
rect 480180 264964 480186 265028
rect 482829 265026 482876 265028
rect 482784 265024 482876 265026
rect 482784 264968 482834 265024
rect 482784 264966 482876 264968
rect 482829 264964 482876 264966
rect 482940 264964 482946 265028
rect 485681 265026 485747 265029
rect 485814 265026 485820 265028
rect 485681 265024 485820 265026
rect 485681 264968 485686 265024
rect 485742 264968 485820 265024
rect 485681 264966 485820 264968
rect 482829 264963 482895 264964
rect 485681 264963 485747 264966
rect 485814 264964 485820 264966
rect 485884 265026 485890 265028
rect 486366 265026 486372 265028
rect 485884 264966 486372 265026
rect 485884 264964 485890 264966
rect 486366 264964 486372 264966
rect 486436 264964 486442 265028
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 538673 245578 538739 245581
rect 583520 245578 584960 245668
rect 538673 245576 584960 245578
rect 538673 245520 538678 245576
rect 538734 245520 584960 245576
rect 538673 245518 584960 245520
rect 538673 245515 538739 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 489126 165820 489132 165884
rect 489196 165882 489202 165884
rect 583520 165882 584960 165972
rect 489196 165822 584960 165882
rect 489196 165820 489202 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 486366 125972 486372 126036
rect 486436 126034 486442 126036
rect 583520 126034 584960 126124
rect 486436 125974 584960 126034
rect 486436 125972 486442 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 482870 86124 482876 86188
rect 482940 86186 482946 86188
rect 583520 86186 584960 86276
rect 482940 86126 584960 86186
rect 482940 86124 482946 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 480110 46276 480116 46340
rect 480180 46338 480186 46340
rect 583520 46338 584960 46428
rect 480180 46278 584960 46338
rect 480180 46276 480186 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 549294 19756 549300 19820
rect 549364 19818 549370 19820
rect 583520 19818 584960 19908
rect 549364 19758 584960 19818
rect 549364 19756 549370 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 477350 6564 477356 6628
rect 477420 6626 477426 6628
rect 583520 6626 584960 6716
rect 477420 6566 584960 6626
rect 477420 6564 477426 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 470272 451479 470336 451483
rect 470272 451423 470276 451479
rect 470276 451423 470332 451479
rect 470332 451423 470336 451479
rect 470272 451419 470336 451423
rect 470352 451479 470416 451483
rect 470352 451423 470356 451479
rect 470356 451423 470412 451479
rect 470412 451423 470416 451479
rect 470352 451419 470416 451423
rect 470432 451479 470496 451483
rect 470432 451423 470436 451479
rect 470436 451423 470492 451479
rect 470492 451423 470496 451479
rect 470432 451419 470496 451423
rect 470512 451479 470576 451483
rect 470512 451423 470516 451479
rect 470516 451423 470572 451479
rect 470572 451423 470576 451479
rect 470512 451419 470576 451423
rect 470592 451479 470656 451483
rect 470592 451423 470596 451479
rect 470596 451423 470652 451479
rect 470652 451423 470656 451479
rect 470592 451419 470656 451423
rect 470672 451479 470736 451483
rect 470672 451423 470676 451479
rect 470676 451423 470732 451479
rect 470732 451423 470736 451479
rect 470672 451419 470736 451423
rect 470752 451479 470816 451483
rect 470752 451423 470756 451479
rect 470756 451423 470812 451479
rect 470812 451423 470816 451479
rect 470752 451419 470816 451423
rect 470272 451399 470336 451403
rect 470272 451343 470276 451399
rect 470276 451343 470332 451399
rect 470332 451343 470336 451399
rect 470272 451339 470336 451343
rect 470352 451399 470416 451403
rect 470352 451343 470356 451399
rect 470356 451343 470412 451399
rect 470412 451343 470416 451399
rect 470352 451339 470416 451343
rect 470432 451399 470496 451403
rect 470432 451343 470436 451399
rect 470436 451343 470492 451399
rect 470492 451343 470496 451399
rect 470432 451339 470496 451343
rect 470512 451399 470576 451403
rect 470512 451343 470516 451399
rect 470516 451343 470572 451399
rect 470572 451343 470576 451399
rect 470512 451339 470576 451343
rect 470592 451399 470656 451403
rect 470592 451343 470596 451399
rect 470596 451343 470652 451399
rect 470652 451343 470656 451399
rect 470592 451339 470656 451343
rect 470672 451399 470736 451403
rect 470672 451343 470676 451399
rect 470676 451343 470732 451399
rect 470732 451343 470736 451399
rect 470672 451339 470736 451343
rect 470752 451399 470816 451403
rect 470752 451343 470756 451399
rect 470756 451343 470812 451399
rect 470812 451343 470816 451399
rect 470752 451339 470816 451343
rect 470272 451319 470336 451323
rect 470272 451263 470276 451319
rect 470276 451263 470332 451319
rect 470332 451263 470336 451319
rect 470272 451259 470336 451263
rect 470352 451319 470416 451323
rect 470352 451263 470356 451319
rect 470356 451263 470412 451319
rect 470412 451263 470416 451319
rect 470352 451259 470416 451263
rect 470432 451319 470496 451323
rect 470432 451263 470436 451319
rect 470436 451263 470492 451319
rect 470492 451263 470496 451319
rect 470432 451259 470496 451263
rect 470512 451319 470576 451323
rect 470512 451263 470516 451319
rect 470516 451263 470572 451319
rect 470572 451263 470576 451319
rect 470512 451259 470576 451263
rect 470592 451319 470656 451323
rect 470592 451263 470596 451319
rect 470596 451263 470652 451319
rect 470652 451263 470656 451319
rect 470592 451259 470656 451263
rect 470672 451319 470736 451323
rect 470672 451263 470676 451319
rect 470676 451263 470732 451319
rect 470732 451263 470736 451319
rect 470672 451259 470736 451263
rect 470752 451319 470816 451323
rect 470752 451263 470756 451319
rect 470756 451263 470812 451319
rect 470812 451263 470816 451319
rect 470752 451259 470816 451263
rect 470272 451239 470336 451243
rect 470272 451183 470276 451239
rect 470276 451183 470332 451239
rect 470332 451183 470336 451239
rect 470272 451179 470336 451183
rect 470352 451239 470416 451243
rect 470352 451183 470356 451239
rect 470356 451183 470412 451239
rect 470412 451183 470416 451239
rect 470352 451179 470416 451183
rect 470432 451239 470496 451243
rect 470432 451183 470436 451239
rect 470436 451183 470492 451239
rect 470492 451183 470496 451239
rect 470432 451179 470496 451183
rect 470512 451239 470576 451243
rect 470512 451183 470516 451239
rect 470516 451183 470572 451239
rect 470572 451183 470576 451239
rect 470512 451179 470576 451183
rect 470592 451239 470656 451243
rect 470592 451183 470596 451239
rect 470596 451183 470652 451239
rect 470652 451183 470656 451239
rect 470592 451179 470656 451183
rect 470672 451239 470736 451243
rect 470672 451183 470676 451239
rect 470676 451183 470732 451239
rect 470732 451183 470736 451239
rect 470672 451179 470736 451183
rect 470752 451239 470816 451243
rect 470752 451183 470756 451239
rect 470756 451183 470812 451239
rect 470812 451183 470816 451239
rect 470752 451179 470816 451183
rect 469032 450393 469096 450397
rect 469032 450337 469036 450393
rect 469036 450337 469092 450393
rect 469092 450337 469096 450393
rect 469032 450333 469096 450337
rect 469112 450393 469176 450397
rect 469112 450337 469116 450393
rect 469116 450337 469172 450393
rect 469172 450337 469176 450393
rect 469112 450333 469176 450337
rect 469192 450393 469256 450397
rect 469192 450337 469196 450393
rect 469196 450337 469252 450393
rect 469252 450337 469256 450393
rect 469192 450333 469256 450337
rect 469272 450393 469336 450397
rect 469272 450337 469276 450393
rect 469276 450337 469332 450393
rect 469332 450337 469336 450393
rect 469272 450333 469336 450337
rect 469352 450393 469416 450397
rect 469352 450337 469356 450393
rect 469356 450337 469412 450393
rect 469412 450337 469416 450393
rect 469352 450333 469416 450337
rect 469432 450393 469496 450397
rect 469432 450337 469436 450393
rect 469436 450337 469492 450393
rect 469492 450337 469496 450393
rect 469432 450333 469496 450337
rect 469512 450393 469576 450397
rect 469512 450337 469516 450393
rect 469516 450337 469572 450393
rect 469572 450337 469576 450393
rect 469512 450333 469576 450337
rect 469032 450313 469096 450317
rect 469032 450257 469036 450313
rect 469036 450257 469092 450313
rect 469092 450257 469096 450313
rect 469032 450253 469096 450257
rect 469112 450313 469176 450317
rect 469112 450257 469116 450313
rect 469116 450257 469172 450313
rect 469172 450257 469176 450313
rect 469112 450253 469176 450257
rect 469192 450313 469256 450317
rect 469192 450257 469196 450313
rect 469196 450257 469252 450313
rect 469252 450257 469256 450313
rect 469192 450253 469256 450257
rect 469272 450313 469336 450317
rect 469272 450257 469276 450313
rect 469276 450257 469332 450313
rect 469332 450257 469336 450313
rect 469272 450253 469336 450257
rect 469352 450313 469416 450317
rect 469352 450257 469356 450313
rect 469356 450257 469412 450313
rect 469412 450257 469416 450313
rect 469352 450253 469416 450257
rect 469432 450313 469496 450317
rect 469432 450257 469436 450313
rect 469436 450257 469492 450313
rect 469492 450257 469496 450313
rect 469432 450253 469496 450257
rect 469512 450313 469576 450317
rect 469512 450257 469516 450313
rect 469516 450257 469572 450313
rect 469572 450257 469576 450313
rect 469512 450253 469576 450257
rect 469032 450233 469096 450237
rect 469032 450177 469036 450233
rect 469036 450177 469092 450233
rect 469092 450177 469096 450233
rect 469032 450173 469096 450177
rect 469112 450233 469176 450237
rect 469112 450177 469116 450233
rect 469116 450177 469172 450233
rect 469172 450177 469176 450233
rect 469112 450173 469176 450177
rect 469192 450233 469256 450237
rect 469192 450177 469196 450233
rect 469196 450177 469252 450233
rect 469252 450177 469256 450233
rect 469192 450173 469256 450177
rect 469272 450233 469336 450237
rect 469272 450177 469276 450233
rect 469276 450177 469332 450233
rect 469332 450177 469336 450233
rect 469272 450173 469336 450177
rect 469352 450233 469416 450237
rect 469352 450177 469356 450233
rect 469356 450177 469412 450233
rect 469412 450177 469416 450233
rect 469352 450173 469416 450177
rect 469432 450233 469496 450237
rect 469432 450177 469436 450233
rect 469436 450177 469492 450233
rect 469492 450177 469496 450233
rect 469432 450173 469496 450177
rect 469512 450233 469576 450237
rect 469512 450177 469516 450233
rect 469516 450177 469572 450233
rect 469572 450177 469576 450233
rect 469512 450173 469576 450177
rect 478460 450196 478524 450260
rect 481220 450196 481284 450260
rect 484164 450196 484228 450260
rect 487844 450256 487908 450260
rect 487844 450200 487849 450256
rect 487849 450200 487908 450256
rect 487844 450196 487908 450200
rect 469032 450153 469096 450157
rect 469032 450097 469036 450153
rect 469036 450097 469092 450153
rect 469092 450097 469096 450153
rect 469032 450093 469096 450097
rect 469112 450153 469176 450157
rect 469112 450097 469116 450153
rect 469116 450097 469172 450153
rect 469172 450097 469176 450153
rect 469112 450093 469176 450097
rect 469192 450153 469256 450157
rect 469192 450097 469196 450153
rect 469196 450097 469252 450153
rect 469252 450097 469256 450153
rect 469192 450093 469256 450097
rect 469272 450153 469336 450157
rect 469272 450097 469276 450153
rect 469276 450097 469332 450153
rect 469332 450097 469336 450153
rect 469272 450093 469336 450097
rect 469352 450153 469416 450157
rect 469352 450097 469356 450153
rect 469356 450097 469412 450153
rect 469412 450097 469416 450153
rect 469352 450093 469416 450097
rect 469432 450153 469496 450157
rect 469432 450097 469436 450153
rect 469436 450097 469492 450153
rect 469492 450097 469496 450153
rect 469432 450093 469496 450097
rect 469512 450153 469576 450157
rect 469512 450097 469516 450153
rect 469516 450097 469572 450153
rect 469572 450097 469576 450153
rect 469512 450093 469576 450097
rect 473676 449652 473740 449716
rect 470272 449308 470336 449312
rect 470272 449252 470276 449308
rect 470276 449252 470332 449308
rect 470332 449252 470336 449308
rect 470272 449248 470336 449252
rect 470352 449308 470416 449312
rect 470352 449252 470356 449308
rect 470356 449252 470412 449308
rect 470412 449252 470416 449308
rect 470352 449248 470416 449252
rect 470432 449308 470496 449312
rect 470432 449252 470436 449308
rect 470436 449252 470492 449308
rect 470492 449252 470496 449308
rect 470432 449248 470496 449252
rect 470512 449308 470576 449312
rect 470512 449252 470516 449308
rect 470516 449252 470572 449308
rect 470572 449252 470576 449308
rect 470512 449248 470576 449252
rect 470592 449308 470656 449312
rect 470592 449252 470596 449308
rect 470596 449252 470652 449308
rect 470652 449252 470656 449308
rect 470592 449248 470656 449252
rect 470672 449308 470736 449312
rect 470672 449252 470676 449308
rect 470676 449252 470732 449308
rect 470732 449252 470736 449308
rect 470672 449248 470736 449252
rect 470752 449308 470816 449312
rect 470752 449252 470756 449308
rect 470756 449252 470812 449308
rect 470812 449252 470816 449308
rect 470752 449248 470816 449252
rect 470272 449228 470336 449232
rect 470272 449172 470276 449228
rect 470276 449172 470332 449228
rect 470332 449172 470336 449228
rect 470272 449168 470336 449172
rect 470352 449228 470416 449232
rect 470352 449172 470356 449228
rect 470356 449172 470412 449228
rect 470412 449172 470416 449228
rect 470352 449168 470416 449172
rect 470432 449228 470496 449232
rect 470432 449172 470436 449228
rect 470436 449172 470492 449228
rect 470492 449172 470496 449228
rect 470432 449168 470496 449172
rect 470512 449228 470576 449232
rect 470512 449172 470516 449228
rect 470516 449172 470572 449228
rect 470572 449172 470576 449228
rect 470512 449168 470576 449172
rect 470592 449228 470656 449232
rect 470592 449172 470596 449228
rect 470596 449172 470652 449228
rect 470652 449172 470656 449228
rect 470592 449168 470656 449172
rect 470672 449228 470736 449232
rect 470672 449172 470676 449228
rect 470676 449172 470732 449228
rect 470732 449172 470736 449228
rect 470672 449168 470736 449172
rect 470752 449228 470816 449232
rect 470752 449172 470756 449228
rect 470756 449172 470812 449228
rect 470812 449172 470816 449228
rect 470752 449168 470816 449172
rect 470272 449148 470336 449152
rect 470272 449092 470276 449148
rect 470276 449092 470332 449148
rect 470332 449092 470336 449148
rect 470272 449088 470336 449092
rect 470352 449148 470416 449152
rect 470352 449092 470356 449148
rect 470356 449092 470412 449148
rect 470412 449092 470416 449148
rect 470352 449088 470416 449092
rect 470432 449148 470496 449152
rect 470432 449092 470436 449148
rect 470436 449092 470492 449148
rect 470492 449092 470496 449148
rect 470432 449088 470496 449092
rect 470512 449148 470576 449152
rect 470512 449092 470516 449148
rect 470516 449092 470572 449148
rect 470572 449092 470576 449148
rect 470512 449088 470576 449092
rect 470592 449148 470656 449152
rect 470592 449092 470596 449148
rect 470596 449092 470652 449148
rect 470652 449092 470656 449148
rect 470592 449088 470656 449092
rect 470672 449148 470736 449152
rect 470672 449092 470676 449148
rect 470676 449092 470732 449148
rect 470732 449092 470736 449148
rect 470672 449088 470736 449092
rect 470752 449148 470816 449152
rect 470752 449092 470756 449148
rect 470756 449092 470812 449148
rect 470812 449092 470816 449148
rect 470752 449088 470816 449092
rect 470272 449068 470336 449072
rect 470272 449012 470276 449068
rect 470276 449012 470332 449068
rect 470332 449012 470336 449068
rect 470272 449008 470336 449012
rect 470352 449068 470416 449072
rect 470352 449012 470356 449068
rect 470356 449012 470412 449068
rect 470412 449012 470416 449068
rect 470352 449008 470416 449012
rect 470432 449068 470496 449072
rect 470432 449012 470436 449068
rect 470436 449012 470492 449068
rect 470492 449012 470496 449068
rect 470432 449008 470496 449012
rect 470512 449068 470576 449072
rect 470512 449012 470516 449068
rect 470516 449012 470572 449068
rect 470572 449012 470576 449068
rect 470512 449008 470576 449012
rect 470592 449068 470656 449072
rect 470592 449012 470596 449068
rect 470596 449012 470652 449068
rect 470652 449012 470656 449068
rect 470592 449008 470656 449012
rect 470672 449068 470736 449072
rect 470672 449012 470676 449068
rect 470676 449012 470732 449068
rect 470732 449012 470736 449068
rect 470672 449008 470736 449012
rect 470752 449068 470816 449072
rect 470752 449012 470756 449068
rect 470756 449012 470812 449068
rect 470812 449012 470816 449068
rect 470752 449008 470816 449012
rect 541572 445028 541636 445092
rect 544332 445028 544396 445092
rect 549300 434692 549364 434756
rect 470272 433080 470336 433084
rect 470272 433024 470276 433080
rect 470276 433024 470332 433080
rect 470332 433024 470336 433080
rect 470272 433020 470336 433024
rect 470352 433080 470416 433084
rect 470352 433024 470356 433080
rect 470356 433024 470412 433080
rect 470412 433024 470416 433080
rect 470352 433020 470416 433024
rect 470432 433080 470496 433084
rect 470432 433024 470436 433080
rect 470436 433024 470492 433080
rect 470492 433024 470496 433080
rect 470432 433020 470496 433024
rect 470512 433080 470576 433084
rect 470512 433024 470516 433080
rect 470516 433024 470572 433080
rect 470572 433024 470576 433080
rect 470512 433020 470576 433024
rect 470592 433080 470656 433084
rect 470592 433024 470596 433080
rect 470596 433024 470652 433080
rect 470652 433024 470656 433080
rect 470592 433020 470656 433024
rect 470672 433080 470736 433084
rect 470672 433024 470676 433080
rect 470676 433024 470732 433080
rect 470732 433024 470736 433080
rect 470672 433020 470736 433024
rect 470752 433080 470816 433084
rect 470752 433024 470756 433080
rect 470756 433024 470812 433080
rect 470812 433024 470816 433080
rect 470752 433020 470816 433024
rect 470272 433000 470336 433004
rect 470272 432944 470276 433000
rect 470276 432944 470332 433000
rect 470332 432944 470336 433000
rect 470272 432940 470336 432944
rect 470352 433000 470416 433004
rect 470352 432944 470356 433000
rect 470356 432944 470412 433000
rect 470412 432944 470416 433000
rect 470352 432940 470416 432944
rect 470432 433000 470496 433004
rect 470432 432944 470436 433000
rect 470436 432944 470492 433000
rect 470492 432944 470496 433000
rect 470432 432940 470496 432944
rect 470512 433000 470576 433004
rect 470512 432944 470516 433000
rect 470516 432944 470572 433000
rect 470572 432944 470576 433000
rect 470512 432940 470576 432944
rect 470592 433000 470656 433004
rect 470592 432944 470596 433000
rect 470596 432944 470652 433000
rect 470652 432944 470656 433000
rect 470592 432940 470656 432944
rect 470672 433000 470736 433004
rect 470672 432944 470676 433000
rect 470676 432944 470732 433000
rect 470732 432944 470736 433000
rect 470672 432940 470736 432944
rect 470752 433000 470816 433004
rect 470752 432944 470756 433000
rect 470756 432944 470812 433000
rect 470812 432944 470816 433000
rect 470752 432940 470816 432944
rect 470272 432920 470336 432924
rect 470272 432864 470276 432920
rect 470276 432864 470332 432920
rect 470332 432864 470336 432920
rect 470272 432860 470336 432864
rect 470352 432920 470416 432924
rect 470352 432864 470356 432920
rect 470356 432864 470412 432920
rect 470412 432864 470416 432920
rect 470352 432860 470416 432864
rect 470432 432920 470496 432924
rect 470432 432864 470436 432920
rect 470436 432864 470492 432920
rect 470492 432864 470496 432920
rect 470432 432860 470496 432864
rect 470512 432920 470576 432924
rect 470512 432864 470516 432920
rect 470516 432864 470572 432920
rect 470572 432864 470576 432920
rect 470512 432860 470576 432864
rect 470592 432920 470656 432924
rect 470592 432864 470596 432920
rect 470596 432864 470652 432920
rect 470652 432864 470656 432920
rect 470592 432860 470656 432864
rect 470672 432920 470736 432924
rect 470672 432864 470676 432920
rect 470676 432864 470732 432920
rect 470732 432864 470736 432920
rect 470672 432860 470736 432864
rect 470752 432920 470816 432924
rect 470752 432864 470756 432920
rect 470756 432864 470812 432920
rect 470812 432864 470816 432920
rect 470752 432860 470816 432864
rect 470272 432840 470336 432844
rect 470272 432784 470276 432840
rect 470276 432784 470332 432840
rect 470332 432784 470336 432840
rect 470272 432780 470336 432784
rect 470352 432840 470416 432844
rect 470352 432784 470356 432840
rect 470356 432784 470412 432840
rect 470412 432784 470416 432840
rect 470352 432780 470416 432784
rect 470432 432840 470496 432844
rect 470432 432784 470436 432840
rect 470436 432784 470492 432840
rect 470492 432784 470496 432840
rect 470432 432780 470496 432784
rect 470512 432840 470576 432844
rect 470512 432784 470516 432840
rect 470516 432784 470572 432840
rect 470572 432784 470576 432840
rect 470512 432780 470576 432784
rect 470592 432840 470656 432844
rect 470592 432784 470596 432840
rect 470596 432784 470652 432840
rect 470652 432784 470656 432840
rect 470592 432780 470656 432784
rect 470672 432840 470736 432844
rect 470672 432784 470676 432840
rect 470676 432784 470732 432840
rect 470732 432784 470736 432840
rect 470672 432780 470736 432784
rect 470752 432840 470816 432844
rect 470752 432784 470756 432840
rect 470756 432784 470812 432840
rect 470812 432784 470816 432840
rect 470752 432780 470816 432784
rect 483612 432304 483676 432308
rect 483612 432248 483626 432304
rect 483626 432248 483676 432304
rect 483612 432244 483676 432248
rect 481220 432168 481284 432172
rect 481220 432112 481270 432168
rect 481270 432112 481284 432168
rect 481220 432108 481284 432112
rect 469032 431993 469096 431997
rect 469032 431937 469036 431993
rect 469036 431937 469092 431993
rect 469092 431937 469096 431993
rect 469032 431933 469096 431937
rect 469112 431993 469176 431997
rect 469112 431937 469116 431993
rect 469116 431937 469172 431993
rect 469172 431937 469176 431993
rect 469112 431933 469176 431937
rect 469192 431993 469256 431997
rect 469192 431937 469196 431993
rect 469196 431937 469252 431993
rect 469252 431937 469256 431993
rect 469192 431933 469256 431937
rect 469272 431993 469336 431997
rect 469272 431937 469276 431993
rect 469276 431937 469332 431993
rect 469332 431937 469336 431993
rect 469272 431933 469336 431937
rect 469352 431993 469416 431997
rect 469352 431937 469356 431993
rect 469356 431937 469412 431993
rect 469412 431937 469416 431993
rect 469352 431933 469416 431937
rect 469432 431993 469496 431997
rect 469432 431937 469436 431993
rect 469436 431937 469492 431993
rect 469492 431937 469496 431993
rect 469432 431933 469496 431937
rect 469512 431993 469576 431997
rect 469512 431937 469516 431993
rect 469516 431937 469572 431993
rect 469572 431937 469576 431993
rect 469512 431933 469576 431937
rect 469032 431913 469096 431917
rect 469032 431857 469036 431913
rect 469036 431857 469092 431913
rect 469092 431857 469096 431913
rect 469032 431853 469096 431857
rect 469112 431913 469176 431917
rect 469112 431857 469116 431913
rect 469116 431857 469172 431913
rect 469172 431857 469176 431913
rect 469112 431853 469176 431857
rect 469192 431913 469256 431917
rect 469192 431857 469196 431913
rect 469196 431857 469252 431913
rect 469252 431857 469256 431913
rect 469192 431853 469256 431857
rect 469272 431913 469336 431917
rect 469272 431857 469276 431913
rect 469276 431857 469332 431913
rect 469332 431857 469336 431913
rect 469272 431853 469336 431857
rect 469352 431913 469416 431917
rect 469352 431857 469356 431913
rect 469356 431857 469412 431913
rect 469412 431857 469416 431913
rect 469352 431853 469416 431857
rect 469432 431913 469496 431917
rect 469432 431857 469436 431913
rect 469436 431857 469492 431913
rect 469492 431857 469496 431913
rect 469432 431853 469496 431857
rect 469512 431913 469576 431917
rect 469512 431857 469516 431913
rect 469516 431857 469572 431913
rect 469572 431857 469576 431913
rect 469512 431853 469576 431857
rect 469032 431833 469096 431837
rect 469032 431777 469036 431833
rect 469036 431777 469092 431833
rect 469092 431777 469096 431833
rect 469032 431773 469096 431777
rect 469112 431833 469176 431837
rect 469112 431777 469116 431833
rect 469116 431777 469172 431833
rect 469172 431777 469176 431833
rect 469112 431773 469176 431777
rect 469192 431833 469256 431837
rect 469192 431777 469196 431833
rect 469196 431777 469252 431833
rect 469252 431777 469256 431833
rect 469192 431773 469256 431777
rect 469272 431833 469336 431837
rect 469272 431777 469276 431833
rect 469276 431777 469332 431833
rect 469332 431777 469336 431833
rect 469272 431773 469336 431777
rect 469352 431833 469416 431837
rect 469352 431777 469356 431833
rect 469356 431777 469412 431833
rect 469412 431777 469416 431833
rect 469352 431773 469416 431777
rect 469432 431833 469496 431837
rect 469432 431777 469436 431833
rect 469436 431777 469492 431833
rect 469492 431777 469496 431833
rect 469432 431773 469496 431777
rect 469512 431833 469576 431837
rect 469512 431777 469516 431833
rect 469516 431777 469572 431833
rect 469572 431777 469576 431833
rect 469512 431773 469576 431777
rect 473676 431836 473740 431900
rect 487660 431836 487724 431900
rect 469032 431753 469096 431757
rect 469032 431697 469036 431753
rect 469036 431697 469092 431753
rect 469092 431697 469096 431753
rect 469032 431693 469096 431697
rect 469112 431753 469176 431757
rect 469112 431697 469116 431753
rect 469116 431697 469172 431753
rect 469172 431697 469176 431753
rect 469112 431693 469176 431697
rect 469192 431753 469256 431757
rect 469192 431697 469196 431753
rect 469196 431697 469252 431753
rect 469252 431697 469256 431753
rect 469192 431693 469256 431697
rect 469272 431753 469336 431757
rect 469272 431697 469276 431753
rect 469276 431697 469332 431753
rect 469332 431697 469336 431753
rect 469272 431693 469336 431697
rect 469352 431753 469416 431757
rect 469352 431697 469356 431753
rect 469356 431697 469412 431753
rect 469412 431697 469416 431753
rect 469352 431693 469416 431697
rect 469432 431753 469496 431757
rect 469432 431697 469436 431753
rect 469436 431697 469492 431753
rect 469492 431697 469496 431753
rect 469432 431693 469496 431697
rect 469512 431753 469576 431757
rect 469512 431697 469516 431753
rect 469516 431697 469572 431753
rect 469572 431697 469576 431753
rect 469512 431693 469576 431697
rect 478460 431564 478524 431628
rect 470272 430908 470336 430912
rect 470272 430852 470276 430908
rect 470276 430852 470332 430908
rect 470332 430852 470336 430908
rect 470272 430848 470336 430852
rect 470352 430908 470416 430912
rect 470352 430852 470356 430908
rect 470356 430852 470412 430908
rect 470412 430852 470416 430908
rect 470352 430848 470416 430852
rect 470432 430908 470496 430912
rect 470432 430852 470436 430908
rect 470436 430852 470492 430908
rect 470492 430852 470496 430908
rect 470432 430848 470496 430852
rect 470512 430908 470576 430912
rect 470512 430852 470516 430908
rect 470516 430852 470572 430908
rect 470572 430852 470576 430908
rect 470512 430848 470576 430852
rect 470592 430908 470656 430912
rect 470592 430852 470596 430908
rect 470596 430852 470652 430908
rect 470652 430852 470656 430908
rect 470592 430848 470656 430852
rect 470672 430908 470736 430912
rect 470672 430852 470676 430908
rect 470676 430852 470732 430908
rect 470732 430852 470736 430908
rect 470672 430848 470736 430852
rect 470752 430908 470816 430912
rect 470752 430852 470756 430908
rect 470756 430852 470812 430908
rect 470812 430852 470816 430908
rect 470752 430848 470816 430852
rect 470272 430828 470336 430832
rect 470272 430772 470276 430828
rect 470276 430772 470332 430828
rect 470332 430772 470336 430828
rect 470272 430768 470336 430772
rect 470352 430828 470416 430832
rect 470352 430772 470356 430828
rect 470356 430772 470412 430828
rect 470412 430772 470416 430828
rect 470352 430768 470416 430772
rect 470432 430828 470496 430832
rect 470432 430772 470436 430828
rect 470436 430772 470492 430828
rect 470492 430772 470496 430828
rect 470432 430768 470496 430772
rect 470512 430828 470576 430832
rect 470512 430772 470516 430828
rect 470516 430772 470572 430828
rect 470572 430772 470576 430828
rect 470512 430768 470576 430772
rect 470592 430828 470656 430832
rect 470592 430772 470596 430828
rect 470596 430772 470652 430828
rect 470652 430772 470656 430828
rect 470592 430768 470656 430772
rect 470672 430828 470736 430832
rect 470672 430772 470676 430828
rect 470676 430772 470732 430828
rect 470732 430772 470736 430828
rect 470672 430768 470736 430772
rect 470752 430828 470816 430832
rect 470752 430772 470756 430828
rect 470756 430772 470812 430828
rect 470812 430772 470816 430828
rect 470752 430768 470816 430772
rect 470272 430748 470336 430752
rect 470272 430692 470276 430748
rect 470276 430692 470332 430748
rect 470332 430692 470336 430748
rect 470272 430688 470336 430692
rect 470352 430748 470416 430752
rect 470352 430692 470356 430748
rect 470356 430692 470412 430748
rect 470412 430692 470416 430748
rect 470352 430688 470416 430692
rect 470432 430748 470496 430752
rect 470432 430692 470436 430748
rect 470436 430692 470492 430748
rect 470492 430692 470496 430748
rect 470432 430688 470496 430692
rect 470512 430748 470576 430752
rect 470512 430692 470516 430748
rect 470516 430692 470572 430748
rect 470572 430692 470576 430748
rect 470512 430688 470576 430692
rect 470592 430748 470656 430752
rect 470592 430692 470596 430748
rect 470596 430692 470652 430748
rect 470652 430692 470656 430748
rect 470592 430688 470656 430692
rect 470672 430748 470736 430752
rect 470672 430692 470676 430748
rect 470676 430692 470732 430748
rect 470732 430692 470736 430748
rect 470672 430688 470736 430692
rect 470752 430748 470816 430752
rect 470752 430692 470756 430748
rect 470756 430692 470812 430748
rect 470812 430692 470816 430748
rect 470752 430688 470816 430692
rect 470272 430668 470336 430672
rect 470272 430612 470276 430668
rect 470276 430612 470332 430668
rect 470332 430612 470336 430668
rect 470272 430608 470336 430612
rect 470352 430668 470416 430672
rect 470352 430612 470356 430668
rect 470356 430612 470412 430668
rect 470412 430612 470416 430668
rect 470352 430608 470416 430612
rect 470432 430668 470496 430672
rect 470432 430612 470436 430668
rect 470436 430612 470492 430668
rect 470492 430612 470496 430668
rect 470432 430608 470496 430612
rect 470512 430668 470576 430672
rect 470512 430612 470516 430668
rect 470516 430612 470572 430668
rect 470572 430612 470576 430668
rect 470512 430608 470576 430612
rect 470592 430668 470656 430672
rect 470592 430612 470596 430668
rect 470596 430612 470652 430668
rect 470652 430612 470656 430668
rect 470592 430608 470656 430612
rect 470672 430668 470736 430672
rect 470672 430612 470676 430668
rect 470676 430612 470732 430668
rect 470732 430612 470736 430668
rect 470672 430608 470736 430612
rect 470752 430668 470816 430672
rect 470752 430612 470756 430668
rect 470756 430612 470812 430668
rect 470812 430612 470816 430668
rect 470752 430608 470816 430612
rect 480116 427892 480180 427956
rect 486556 427892 486620 427956
rect 470272 412080 470336 412084
rect 470272 412024 470276 412080
rect 470276 412024 470332 412080
rect 470332 412024 470336 412080
rect 470272 412020 470336 412024
rect 470352 412080 470416 412084
rect 470352 412024 470356 412080
rect 470356 412024 470412 412080
rect 470412 412024 470416 412080
rect 470352 412020 470416 412024
rect 470432 412080 470496 412084
rect 470432 412024 470436 412080
rect 470436 412024 470492 412080
rect 470492 412024 470496 412080
rect 470432 412020 470496 412024
rect 470512 412080 470576 412084
rect 470512 412024 470516 412080
rect 470516 412024 470572 412080
rect 470572 412024 470576 412080
rect 470512 412020 470576 412024
rect 470592 412080 470656 412084
rect 470592 412024 470596 412080
rect 470596 412024 470652 412080
rect 470652 412024 470656 412080
rect 470592 412020 470656 412024
rect 470672 412080 470736 412084
rect 470672 412024 470676 412080
rect 470676 412024 470732 412080
rect 470732 412024 470736 412080
rect 470672 412020 470736 412024
rect 470752 412080 470816 412084
rect 470752 412024 470756 412080
rect 470756 412024 470812 412080
rect 470812 412024 470816 412080
rect 470752 412020 470816 412024
rect 470272 412000 470336 412004
rect 470272 411944 470276 412000
rect 470276 411944 470332 412000
rect 470332 411944 470336 412000
rect 470272 411940 470336 411944
rect 470352 412000 470416 412004
rect 470352 411944 470356 412000
rect 470356 411944 470412 412000
rect 470412 411944 470416 412000
rect 470352 411940 470416 411944
rect 470432 412000 470496 412004
rect 470432 411944 470436 412000
rect 470436 411944 470492 412000
rect 470492 411944 470496 412000
rect 470432 411940 470496 411944
rect 470512 412000 470576 412004
rect 470512 411944 470516 412000
rect 470516 411944 470572 412000
rect 470572 411944 470576 412000
rect 470512 411940 470576 411944
rect 470592 412000 470656 412004
rect 470592 411944 470596 412000
rect 470596 411944 470652 412000
rect 470652 411944 470656 412000
rect 470592 411940 470656 411944
rect 470672 412000 470736 412004
rect 470672 411944 470676 412000
rect 470676 411944 470732 412000
rect 470732 411944 470736 412000
rect 470672 411940 470736 411944
rect 470752 412000 470816 412004
rect 470752 411944 470756 412000
rect 470756 411944 470812 412000
rect 470812 411944 470816 412000
rect 470752 411940 470816 411944
rect 470272 411920 470336 411924
rect 470272 411864 470276 411920
rect 470276 411864 470332 411920
rect 470332 411864 470336 411920
rect 470272 411860 470336 411864
rect 470352 411920 470416 411924
rect 470352 411864 470356 411920
rect 470356 411864 470412 411920
rect 470412 411864 470416 411920
rect 470352 411860 470416 411864
rect 470432 411920 470496 411924
rect 470432 411864 470436 411920
rect 470436 411864 470492 411920
rect 470492 411864 470496 411920
rect 470432 411860 470496 411864
rect 470512 411920 470576 411924
rect 470512 411864 470516 411920
rect 470516 411864 470572 411920
rect 470572 411864 470576 411920
rect 470512 411860 470576 411864
rect 470592 411920 470656 411924
rect 470592 411864 470596 411920
rect 470596 411864 470652 411920
rect 470652 411864 470656 411920
rect 470592 411860 470656 411864
rect 470672 411920 470736 411924
rect 470672 411864 470676 411920
rect 470676 411864 470732 411920
rect 470732 411864 470736 411920
rect 470672 411860 470736 411864
rect 470752 411920 470816 411924
rect 470752 411864 470756 411920
rect 470756 411864 470812 411920
rect 470812 411864 470816 411920
rect 470752 411860 470816 411864
rect 470272 411840 470336 411844
rect 470272 411784 470276 411840
rect 470276 411784 470332 411840
rect 470332 411784 470336 411840
rect 470272 411780 470336 411784
rect 470352 411840 470416 411844
rect 470352 411784 470356 411840
rect 470356 411784 470412 411840
rect 470412 411784 470416 411840
rect 470352 411780 470416 411784
rect 470432 411840 470496 411844
rect 470432 411784 470436 411840
rect 470436 411784 470492 411840
rect 470492 411784 470496 411840
rect 470432 411780 470496 411784
rect 470512 411840 470576 411844
rect 470512 411784 470516 411840
rect 470516 411784 470572 411840
rect 470572 411784 470576 411840
rect 470512 411780 470576 411784
rect 470592 411840 470656 411844
rect 470592 411784 470596 411840
rect 470596 411784 470652 411840
rect 470652 411784 470656 411840
rect 470592 411780 470656 411784
rect 470672 411840 470736 411844
rect 470672 411784 470676 411840
rect 470676 411784 470732 411840
rect 470732 411784 470736 411840
rect 470672 411780 470736 411784
rect 470752 411840 470816 411844
rect 470752 411784 470756 411840
rect 470756 411784 470812 411840
rect 470812 411784 470816 411840
rect 470752 411780 470816 411784
rect 469032 410994 469096 410998
rect 469032 410938 469036 410994
rect 469036 410938 469092 410994
rect 469092 410938 469096 410994
rect 469032 410934 469096 410938
rect 469112 410994 469176 410998
rect 469112 410938 469116 410994
rect 469116 410938 469172 410994
rect 469172 410938 469176 410994
rect 469112 410934 469176 410938
rect 469192 410994 469256 410998
rect 469192 410938 469196 410994
rect 469196 410938 469252 410994
rect 469252 410938 469256 410994
rect 469192 410934 469256 410938
rect 469272 410994 469336 410998
rect 469272 410938 469276 410994
rect 469276 410938 469332 410994
rect 469332 410938 469336 410994
rect 469272 410934 469336 410938
rect 469352 410994 469416 410998
rect 469352 410938 469356 410994
rect 469356 410938 469412 410994
rect 469412 410938 469416 410994
rect 469352 410934 469416 410938
rect 469432 410994 469496 410998
rect 469432 410938 469436 410994
rect 469436 410938 469492 410994
rect 469492 410938 469496 410994
rect 469432 410934 469496 410938
rect 469512 410994 469576 410998
rect 469512 410938 469516 410994
rect 469516 410938 469572 410994
rect 469572 410938 469576 410994
rect 469512 410934 469576 410938
rect 469032 410914 469096 410918
rect 469032 410858 469036 410914
rect 469036 410858 469092 410914
rect 469092 410858 469096 410914
rect 469032 410854 469096 410858
rect 469112 410914 469176 410918
rect 469112 410858 469116 410914
rect 469116 410858 469172 410914
rect 469172 410858 469176 410914
rect 469112 410854 469176 410858
rect 469192 410914 469256 410918
rect 469192 410858 469196 410914
rect 469196 410858 469252 410914
rect 469252 410858 469256 410914
rect 469192 410854 469256 410858
rect 469272 410914 469336 410918
rect 469272 410858 469276 410914
rect 469276 410858 469332 410914
rect 469332 410858 469336 410914
rect 469272 410854 469336 410858
rect 469352 410914 469416 410918
rect 469352 410858 469356 410914
rect 469356 410858 469412 410914
rect 469412 410858 469416 410914
rect 469352 410854 469416 410858
rect 469432 410914 469496 410918
rect 469432 410858 469436 410914
rect 469436 410858 469492 410914
rect 469492 410858 469496 410914
rect 469432 410854 469496 410858
rect 469512 410914 469576 410918
rect 469512 410858 469516 410914
rect 469516 410858 469572 410914
rect 469572 410858 469576 410914
rect 469512 410854 469576 410858
rect 473676 410952 473740 410956
rect 473676 410896 473726 410952
rect 473726 410896 473740 410952
rect 473676 410892 473740 410896
rect 469032 410834 469096 410838
rect 469032 410778 469036 410834
rect 469036 410778 469092 410834
rect 469092 410778 469096 410834
rect 469032 410774 469096 410778
rect 469112 410834 469176 410838
rect 469112 410778 469116 410834
rect 469116 410778 469172 410834
rect 469172 410778 469176 410834
rect 469112 410774 469176 410778
rect 469192 410834 469256 410838
rect 469192 410778 469196 410834
rect 469196 410778 469252 410834
rect 469252 410778 469256 410834
rect 469192 410774 469256 410778
rect 469272 410834 469336 410838
rect 469272 410778 469276 410834
rect 469276 410778 469332 410834
rect 469332 410778 469336 410834
rect 469272 410774 469336 410778
rect 469352 410834 469416 410838
rect 469352 410778 469356 410834
rect 469356 410778 469412 410834
rect 469412 410778 469416 410834
rect 469352 410774 469416 410778
rect 469432 410834 469496 410838
rect 469432 410778 469436 410834
rect 469436 410778 469492 410834
rect 469492 410778 469496 410834
rect 469432 410774 469496 410778
rect 469512 410834 469576 410838
rect 469512 410778 469516 410834
rect 469516 410778 469572 410834
rect 469572 410778 469576 410834
rect 469512 410774 469576 410778
rect 469032 410754 469096 410758
rect 469032 410698 469036 410754
rect 469036 410698 469092 410754
rect 469092 410698 469096 410754
rect 469032 410694 469096 410698
rect 469112 410754 469176 410758
rect 469112 410698 469116 410754
rect 469116 410698 469172 410754
rect 469172 410698 469176 410754
rect 469112 410694 469176 410698
rect 469192 410754 469256 410758
rect 469192 410698 469196 410754
rect 469196 410698 469252 410754
rect 469252 410698 469256 410754
rect 469192 410694 469256 410698
rect 469272 410754 469336 410758
rect 469272 410698 469276 410754
rect 469276 410698 469332 410754
rect 469332 410698 469336 410754
rect 469272 410694 469336 410698
rect 469352 410754 469416 410758
rect 469352 410698 469356 410754
rect 469356 410698 469412 410754
rect 469412 410698 469416 410754
rect 469352 410694 469416 410698
rect 469432 410754 469496 410758
rect 469432 410698 469436 410754
rect 469436 410698 469492 410754
rect 469492 410698 469496 410754
rect 469432 410694 469496 410698
rect 469512 410754 469576 410758
rect 469512 410698 469516 410754
rect 469516 410698 469572 410754
rect 469572 410698 469576 410754
rect 469512 410694 469576 410698
rect 484164 410408 484228 410412
rect 484164 410352 484178 410408
rect 484178 410352 484228 410408
rect 484164 410348 484228 410352
rect 478460 410136 478524 410140
rect 478460 410080 478474 410136
rect 478474 410080 478524 410136
rect 478460 410076 478524 410080
rect 481404 410136 481468 410140
rect 481404 410080 481418 410136
rect 481418 410080 481468 410136
rect 481404 410076 481468 410080
rect 487844 410136 487908 410140
rect 487844 410080 487858 410136
rect 487858 410080 487908 410136
rect 487844 410076 487908 410080
rect 488396 410076 488460 410140
rect 470272 409908 470336 409912
rect 470272 409852 470276 409908
rect 470276 409852 470332 409908
rect 470332 409852 470336 409908
rect 470272 409848 470336 409852
rect 470352 409908 470416 409912
rect 470352 409852 470356 409908
rect 470356 409852 470412 409908
rect 470412 409852 470416 409908
rect 470352 409848 470416 409852
rect 470432 409908 470496 409912
rect 470432 409852 470436 409908
rect 470436 409852 470492 409908
rect 470492 409852 470496 409908
rect 470432 409848 470496 409852
rect 470512 409908 470576 409912
rect 470512 409852 470516 409908
rect 470516 409852 470572 409908
rect 470572 409852 470576 409908
rect 470512 409848 470576 409852
rect 470592 409908 470656 409912
rect 470592 409852 470596 409908
rect 470596 409852 470652 409908
rect 470652 409852 470656 409908
rect 470592 409848 470656 409852
rect 470672 409908 470736 409912
rect 470672 409852 470676 409908
rect 470676 409852 470732 409908
rect 470732 409852 470736 409908
rect 470672 409848 470736 409852
rect 470752 409908 470816 409912
rect 470752 409852 470756 409908
rect 470756 409852 470812 409908
rect 470812 409852 470816 409908
rect 470752 409848 470816 409852
rect 470272 409828 470336 409832
rect 470272 409772 470276 409828
rect 470276 409772 470332 409828
rect 470332 409772 470336 409828
rect 470272 409768 470336 409772
rect 470352 409828 470416 409832
rect 470352 409772 470356 409828
rect 470356 409772 470412 409828
rect 470412 409772 470416 409828
rect 470352 409768 470416 409772
rect 470432 409828 470496 409832
rect 470432 409772 470436 409828
rect 470436 409772 470492 409828
rect 470492 409772 470496 409828
rect 470432 409768 470496 409772
rect 470512 409828 470576 409832
rect 470512 409772 470516 409828
rect 470516 409772 470572 409828
rect 470572 409772 470576 409828
rect 470512 409768 470576 409772
rect 470592 409828 470656 409832
rect 470592 409772 470596 409828
rect 470596 409772 470652 409828
rect 470652 409772 470656 409828
rect 470592 409768 470656 409772
rect 470672 409828 470736 409832
rect 470672 409772 470676 409828
rect 470676 409772 470732 409828
rect 470732 409772 470736 409828
rect 470672 409768 470736 409772
rect 470752 409828 470816 409832
rect 470752 409772 470756 409828
rect 470756 409772 470812 409828
rect 470812 409772 470816 409828
rect 470752 409768 470816 409772
rect 470272 409748 470336 409752
rect 470272 409692 470276 409748
rect 470276 409692 470332 409748
rect 470332 409692 470336 409748
rect 470272 409688 470336 409692
rect 470352 409748 470416 409752
rect 470352 409692 470356 409748
rect 470356 409692 470412 409748
rect 470412 409692 470416 409748
rect 470352 409688 470416 409692
rect 470432 409748 470496 409752
rect 470432 409692 470436 409748
rect 470436 409692 470492 409748
rect 470492 409692 470496 409748
rect 470432 409688 470496 409692
rect 470512 409748 470576 409752
rect 470512 409692 470516 409748
rect 470516 409692 470572 409748
rect 470572 409692 470576 409748
rect 470512 409688 470576 409692
rect 470592 409748 470656 409752
rect 470592 409692 470596 409748
rect 470596 409692 470652 409748
rect 470652 409692 470656 409748
rect 470592 409688 470656 409692
rect 470672 409748 470736 409752
rect 470672 409692 470676 409748
rect 470676 409692 470732 409748
rect 470732 409692 470736 409748
rect 470672 409688 470736 409692
rect 470752 409748 470816 409752
rect 470752 409692 470756 409748
rect 470756 409692 470812 409748
rect 470812 409692 470816 409748
rect 470752 409688 470816 409692
rect 470272 409668 470336 409672
rect 470272 409612 470276 409668
rect 470276 409612 470332 409668
rect 470332 409612 470336 409668
rect 470272 409608 470336 409612
rect 470352 409668 470416 409672
rect 470352 409612 470356 409668
rect 470356 409612 470412 409668
rect 470412 409612 470416 409668
rect 470352 409608 470416 409612
rect 470432 409668 470496 409672
rect 470432 409612 470436 409668
rect 470436 409612 470492 409668
rect 470492 409612 470496 409668
rect 470432 409608 470496 409612
rect 470512 409668 470576 409672
rect 470512 409612 470516 409668
rect 470516 409612 470572 409668
rect 470572 409612 470576 409668
rect 470512 409608 470576 409612
rect 470592 409668 470656 409672
rect 470592 409612 470596 409668
rect 470596 409612 470652 409668
rect 470652 409612 470656 409668
rect 470592 409608 470656 409612
rect 470672 409668 470736 409672
rect 470672 409612 470676 409668
rect 470676 409612 470732 409668
rect 470732 409612 470736 409668
rect 470672 409608 470736 409612
rect 470752 409668 470816 409672
rect 470752 409612 470756 409668
rect 470756 409612 470812 409668
rect 470812 409612 470816 409668
rect 470752 409608 470816 409612
rect 541572 409260 541636 409324
rect 544332 409320 544396 409324
rect 544332 409264 544346 409320
rect 544346 409264 544396 409320
rect 544332 409260 544396 409264
rect 480116 407492 480180 407556
rect 482876 407084 482940 407148
rect 485636 407084 485700 407148
rect 549300 398244 549364 398308
rect 473676 391988 473740 392052
rect 474964 391988 475028 392052
rect 470272 391081 470336 391085
rect 470272 391025 470276 391081
rect 470276 391025 470332 391081
rect 470332 391025 470336 391081
rect 470272 391021 470336 391025
rect 470352 391081 470416 391085
rect 470352 391025 470356 391081
rect 470356 391025 470412 391081
rect 470412 391025 470416 391081
rect 470352 391021 470416 391025
rect 470432 391081 470496 391085
rect 470432 391025 470436 391081
rect 470436 391025 470492 391081
rect 470492 391025 470496 391081
rect 470432 391021 470496 391025
rect 470512 391081 470576 391085
rect 470512 391025 470516 391081
rect 470516 391025 470572 391081
rect 470572 391025 470576 391081
rect 470512 391021 470576 391025
rect 470592 391081 470656 391085
rect 470592 391025 470596 391081
rect 470596 391025 470652 391081
rect 470652 391025 470656 391081
rect 470592 391021 470656 391025
rect 470672 391081 470736 391085
rect 470672 391025 470676 391081
rect 470676 391025 470732 391081
rect 470732 391025 470736 391081
rect 470672 391021 470736 391025
rect 470752 391081 470816 391085
rect 470752 391025 470756 391081
rect 470756 391025 470812 391081
rect 470812 391025 470816 391081
rect 470752 391021 470816 391025
rect 470272 391001 470336 391005
rect 470272 390945 470276 391001
rect 470276 390945 470332 391001
rect 470332 390945 470336 391001
rect 470272 390941 470336 390945
rect 470352 391001 470416 391005
rect 470352 390945 470356 391001
rect 470356 390945 470412 391001
rect 470412 390945 470416 391001
rect 470352 390941 470416 390945
rect 470432 391001 470496 391005
rect 470432 390945 470436 391001
rect 470436 390945 470492 391001
rect 470492 390945 470496 391001
rect 470432 390941 470496 390945
rect 470512 391001 470576 391005
rect 470512 390945 470516 391001
rect 470516 390945 470572 391001
rect 470572 390945 470576 391001
rect 470512 390941 470576 390945
rect 470592 391001 470656 391005
rect 470592 390945 470596 391001
rect 470596 390945 470652 391001
rect 470652 390945 470656 391001
rect 470592 390941 470656 390945
rect 470672 391001 470736 391005
rect 470672 390945 470676 391001
rect 470676 390945 470732 391001
rect 470732 390945 470736 391001
rect 470672 390941 470736 390945
rect 470752 391001 470816 391005
rect 470752 390945 470756 391001
rect 470756 390945 470812 391001
rect 470812 390945 470816 391001
rect 470752 390941 470816 390945
rect 470272 390921 470336 390925
rect 470272 390865 470276 390921
rect 470276 390865 470332 390921
rect 470332 390865 470336 390921
rect 470272 390861 470336 390865
rect 470352 390921 470416 390925
rect 470352 390865 470356 390921
rect 470356 390865 470412 390921
rect 470412 390865 470416 390921
rect 470352 390861 470416 390865
rect 470432 390921 470496 390925
rect 470432 390865 470436 390921
rect 470436 390865 470492 390921
rect 470492 390865 470496 390921
rect 470432 390861 470496 390865
rect 470512 390921 470576 390925
rect 470512 390865 470516 390921
rect 470516 390865 470572 390921
rect 470572 390865 470576 390921
rect 470512 390861 470576 390865
rect 470592 390921 470656 390925
rect 470592 390865 470596 390921
rect 470596 390865 470652 390921
rect 470652 390865 470656 390921
rect 470592 390861 470656 390865
rect 470672 390921 470736 390925
rect 470672 390865 470676 390921
rect 470676 390865 470732 390921
rect 470732 390865 470736 390921
rect 470672 390861 470736 390865
rect 470752 390921 470816 390925
rect 470752 390865 470756 390921
rect 470756 390865 470812 390921
rect 470812 390865 470816 390921
rect 470752 390861 470816 390865
rect 470272 390841 470336 390845
rect 470272 390785 470276 390841
rect 470276 390785 470332 390841
rect 470332 390785 470336 390841
rect 470272 390781 470336 390785
rect 470352 390841 470416 390845
rect 470352 390785 470356 390841
rect 470356 390785 470412 390841
rect 470412 390785 470416 390841
rect 470352 390781 470416 390785
rect 470432 390841 470496 390845
rect 470432 390785 470436 390841
rect 470436 390785 470492 390841
rect 470492 390785 470496 390841
rect 470432 390781 470496 390785
rect 470512 390841 470576 390845
rect 470512 390785 470516 390841
rect 470516 390785 470572 390841
rect 470572 390785 470576 390841
rect 470512 390781 470576 390785
rect 470592 390841 470656 390845
rect 470592 390785 470596 390841
rect 470596 390785 470652 390841
rect 470652 390785 470656 390841
rect 470592 390781 470656 390785
rect 470672 390841 470736 390845
rect 470672 390785 470676 390841
rect 470676 390785 470732 390841
rect 470732 390785 470736 390841
rect 470672 390781 470736 390785
rect 470752 390841 470816 390845
rect 470752 390785 470756 390841
rect 470756 390785 470812 390841
rect 470812 390785 470816 390841
rect 470752 390781 470816 390785
rect 484900 390233 484964 390297
rect 488396 390084 488460 390148
rect 469032 389998 469096 390002
rect 469032 389942 469036 389998
rect 469036 389942 469092 389998
rect 469092 389942 469096 389998
rect 469032 389938 469096 389942
rect 469112 389998 469176 390002
rect 469112 389942 469116 389998
rect 469116 389942 469172 389998
rect 469172 389942 469176 389998
rect 469112 389938 469176 389942
rect 469192 389998 469256 390002
rect 469192 389942 469196 389998
rect 469196 389942 469252 389998
rect 469252 389942 469256 389998
rect 469192 389938 469256 389942
rect 469272 389998 469336 390002
rect 469272 389942 469276 389998
rect 469276 389942 469332 389998
rect 469332 389942 469336 389998
rect 469272 389938 469336 389942
rect 469352 389998 469416 390002
rect 469352 389942 469356 389998
rect 469356 389942 469412 389998
rect 469412 389942 469416 389998
rect 469352 389938 469416 389942
rect 469432 389998 469496 390002
rect 469432 389942 469436 389998
rect 469436 389942 469492 389998
rect 469492 389942 469496 389998
rect 469432 389938 469496 389942
rect 469512 389998 469576 390002
rect 469512 389942 469516 389998
rect 469516 389942 469572 389998
rect 469572 389942 469576 389998
rect 469512 389938 469576 389942
rect 469032 389918 469096 389922
rect 469032 389862 469036 389918
rect 469036 389862 469092 389918
rect 469092 389862 469096 389918
rect 469032 389858 469096 389862
rect 469112 389918 469176 389922
rect 469112 389862 469116 389918
rect 469116 389862 469172 389918
rect 469172 389862 469176 389918
rect 469112 389858 469176 389862
rect 469192 389918 469256 389922
rect 469192 389862 469196 389918
rect 469196 389862 469252 389918
rect 469252 389862 469256 389918
rect 469192 389858 469256 389862
rect 469272 389918 469336 389922
rect 469272 389862 469276 389918
rect 469276 389862 469332 389918
rect 469332 389862 469336 389918
rect 469272 389858 469336 389862
rect 469352 389918 469416 389922
rect 469352 389862 469356 389918
rect 469356 389862 469412 389918
rect 469412 389862 469416 389918
rect 469352 389858 469416 389862
rect 469432 389918 469496 389922
rect 469432 389862 469436 389918
rect 469436 389862 469492 389918
rect 469492 389862 469496 389918
rect 469432 389858 469496 389862
rect 469512 389918 469576 389922
rect 469512 389862 469516 389918
rect 469516 389862 469572 389918
rect 469572 389862 469576 389918
rect 469512 389858 469576 389862
rect 469032 389838 469096 389842
rect 469032 389782 469036 389838
rect 469036 389782 469092 389838
rect 469092 389782 469096 389838
rect 469032 389778 469096 389782
rect 469112 389838 469176 389842
rect 469112 389782 469116 389838
rect 469116 389782 469172 389838
rect 469172 389782 469176 389838
rect 469112 389778 469176 389782
rect 469192 389838 469256 389842
rect 469192 389782 469196 389838
rect 469196 389782 469252 389838
rect 469252 389782 469256 389838
rect 469192 389778 469256 389782
rect 469272 389838 469336 389842
rect 469272 389782 469276 389838
rect 469276 389782 469332 389838
rect 469332 389782 469336 389838
rect 469272 389778 469336 389782
rect 469352 389838 469416 389842
rect 469352 389782 469356 389838
rect 469356 389782 469412 389838
rect 469412 389782 469416 389838
rect 469352 389778 469416 389782
rect 469432 389838 469496 389842
rect 469432 389782 469436 389838
rect 469436 389782 469492 389838
rect 469492 389782 469496 389838
rect 469432 389778 469496 389782
rect 469512 389838 469576 389842
rect 469512 389782 469516 389838
rect 469516 389782 469572 389838
rect 469572 389782 469576 389838
rect 469512 389778 469576 389782
rect 469032 389758 469096 389762
rect 469032 389702 469036 389758
rect 469036 389702 469092 389758
rect 469092 389702 469096 389758
rect 469032 389698 469096 389702
rect 469112 389758 469176 389762
rect 469112 389702 469116 389758
rect 469116 389702 469172 389758
rect 469172 389702 469176 389758
rect 469112 389698 469176 389702
rect 469192 389758 469256 389762
rect 469192 389702 469196 389758
rect 469196 389702 469252 389758
rect 469252 389702 469256 389758
rect 469192 389698 469256 389702
rect 469272 389758 469336 389762
rect 469272 389702 469276 389758
rect 469276 389702 469332 389758
rect 469332 389702 469336 389758
rect 469272 389698 469336 389702
rect 469352 389758 469416 389762
rect 469352 389702 469356 389758
rect 469356 389702 469412 389758
rect 469412 389702 469416 389758
rect 469352 389698 469416 389702
rect 469432 389758 469496 389762
rect 469432 389702 469436 389758
rect 469436 389702 469492 389758
rect 469492 389702 469496 389758
rect 469432 389698 469496 389702
rect 469512 389758 469576 389762
rect 469512 389702 469516 389758
rect 469516 389702 469572 389758
rect 469572 389702 469576 389758
rect 469512 389698 469576 389702
rect 481772 389404 481836 389468
rect 474964 389328 475028 389332
rect 474964 389272 474978 389328
rect 474978 389272 475028 389328
rect 474964 389268 475028 389272
rect 478644 389328 478708 389332
rect 478644 389272 478690 389328
rect 478690 389272 478708 389328
rect 478644 389268 478708 389272
rect 470272 388908 470336 388912
rect 470272 388852 470276 388908
rect 470276 388852 470332 388908
rect 470332 388852 470336 388908
rect 470272 388848 470336 388852
rect 470352 388908 470416 388912
rect 470352 388852 470356 388908
rect 470356 388852 470412 388908
rect 470412 388852 470416 388908
rect 470352 388848 470416 388852
rect 470432 388908 470496 388912
rect 470432 388852 470436 388908
rect 470436 388852 470492 388908
rect 470492 388852 470496 388908
rect 470432 388848 470496 388852
rect 470512 388908 470576 388912
rect 470512 388852 470516 388908
rect 470516 388852 470572 388908
rect 470572 388852 470576 388908
rect 470512 388848 470576 388852
rect 470592 388908 470656 388912
rect 470592 388852 470596 388908
rect 470596 388852 470652 388908
rect 470652 388852 470656 388908
rect 470592 388848 470656 388852
rect 470672 388908 470736 388912
rect 470672 388852 470676 388908
rect 470676 388852 470732 388908
rect 470732 388852 470736 388908
rect 470672 388848 470736 388852
rect 470752 388908 470816 388912
rect 470752 388852 470756 388908
rect 470756 388852 470812 388908
rect 470812 388852 470816 388908
rect 470752 388848 470816 388852
rect 470272 388828 470336 388832
rect 470272 388772 470276 388828
rect 470276 388772 470332 388828
rect 470332 388772 470336 388828
rect 470272 388768 470336 388772
rect 470352 388828 470416 388832
rect 470352 388772 470356 388828
rect 470356 388772 470412 388828
rect 470412 388772 470416 388828
rect 470352 388768 470416 388772
rect 470432 388828 470496 388832
rect 470432 388772 470436 388828
rect 470436 388772 470492 388828
rect 470492 388772 470496 388828
rect 470432 388768 470496 388772
rect 470512 388828 470576 388832
rect 470512 388772 470516 388828
rect 470516 388772 470572 388828
rect 470572 388772 470576 388828
rect 470512 388768 470576 388772
rect 470592 388828 470656 388832
rect 470592 388772 470596 388828
rect 470596 388772 470652 388828
rect 470652 388772 470656 388828
rect 470592 388768 470656 388772
rect 470672 388828 470736 388832
rect 470672 388772 470676 388828
rect 470676 388772 470732 388828
rect 470732 388772 470736 388828
rect 470672 388768 470736 388772
rect 470752 388828 470816 388832
rect 470752 388772 470756 388828
rect 470756 388772 470812 388828
rect 470812 388772 470816 388828
rect 470752 388768 470816 388772
rect 470272 388748 470336 388752
rect 470272 388692 470276 388748
rect 470276 388692 470332 388748
rect 470332 388692 470336 388748
rect 470272 388688 470336 388692
rect 470352 388748 470416 388752
rect 470352 388692 470356 388748
rect 470356 388692 470412 388748
rect 470412 388692 470416 388748
rect 470352 388688 470416 388692
rect 470432 388748 470496 388752
rect 470432 388692 470436 388748
rect 470436 388692 470492 388748
rect 470492 388692 470496 388748
rect 470432 388688 470496 388692
rect 470512 388748 470576 388752
rect 470512 388692 470516 388748
rect 470516 388692 470572 388748
rect 470572 388692 470576 388748
rect 470512 388688 470576 388692
rect 470592 388748 470656 388752
rect 470592 388692 470596 388748
rect 470596 388692 470652 388748
rect 470652 388692 470656 388748
rect 470592 388688 470656 388692
rect 470672 388748 470736 388752
rect 470672 388692 470676 388748
rect 470676 388692 470732 388748
rect 470732 388692 470736 388748
rect 470672 388688 470736 388692
rect 470752 388748 470816 388752
rect 470752 388692 470756 388748
rect 470756 388692 470812 388748
rect 470812 388692 470816 388748
rect 470752 388688 470816 388692
rect 470272 388668 470336 388672
rect 470272 388612 470276 388668
rect 470276 388612 470332 388668
rect 470332 388612 470336 388668
rect 470272 388608 470336 388612
rect 470352 388668 470416 388672
rect 470352 388612 470356 388668
rect 470356 388612 470412 388668
rect 470412 388612 470416 388668
rect 470352 388608 470416 388612
rect 470432 388668 470496 388672
rect 470432 388612 470436 388668
rect 470436 388612 470492 388668
rect 470492 388612 470496 388668
rect 470432 388608 470496 388612
rect 470512 388668 470576 388672
rect 470512 388612 470516 388668
rect 470516 388612 470572 388668
rect 470572 388612 470576 388668
rect 470512 388608 470576 388612
rect 470592 388668 470656 388672
rect 470592 388612 470596 388668
rect 470596 388612 470652 388668
rect 470652 388612 470656 388668
rect 470592 388608 470656 388612
rect 470672 388668 470736 388672
rect 470672 388612 470676 388668
rect 470676 388612 470732 388668
rect 470732 388612 470736 388668
rect 470672 388608 470736 388612
rect 470752 388668 470816 388672
rect 470752 388612 470756 388668
rect 470756 388612 470812 388668
rect 470812 388612 470816 388668
rect 470752 388608 470816 388612
rect 486740 386412 486804 386476
rect 544516 373416 544580 373420
rect 544516 373360 544530 373416
rect 544530 373360 544580 373416
rect 544516 373356 544580 373360
rect 541572 373084 541636 373148
rect 482876 370092 482940 370156
rect 549300 362748 549364 362812
rect 470272 358481 470336 358485
rect 470272 358425 470276 358481
rect 470276 358425 470332 358481
rect 470332 358425 470336 358481
rect 470272 358421 470336 358425
rect 470352 358481 470416 358485
rect 470352 358425 470356 358481
rect 470356 358425 470412 358481
rect 470412 358425 470416 358481
rect 470352 358421 470416 358425
rect 470432 358481 470496 358485
rect 470432 358425 470436 358481
rect 470436 358425 470492 358481
rect 470492 358425 470496 358481
rect 470432 358421 470496 358425
rect 470512 358481 470576 358485
rect 470512 358425 470516 358481
rect 470516 358425 470572 358481
rect 470572 358425 470576 358481
rect 470512 358421 470576 358425
rect 470592 358481 470656 358485
rect 470592 358425 470596 358481
rect 470596 358425 470652 358481
rect 470652 358425 470656 358481
rect 470592 358421 470656 358425
rect 470672 358481 470736 358485
rect 470672 358425 470676 358481
rect 470676 358425 470732 358481
rect 470732 358425 470736 358481
rect 470672 358421 470736 358425
rect 470752 358481 470816 358485
rect 470752 358425 470756 358481
rect 470756 358425 470812 358481
rect 470812 358425 470816 358481
rect 470752 358421 470816 358425
rect 470272 358401 470336 358405
rect 470272 358345 470276 358401
rect 470276 358345 470332 358401
rect 470332 358345 470336 358401
rect 470272 358341 470336 358345
rect 470352 358401 470416 358405
rect 470352 358345 470356 358401
rect 470356 358345 470412 358401
rect 470412 358345 470416 358401
rect 470352 358341 470416 358345
rect 470432 358401 470496 358405
rect 470432 358345 470436 358401
rect 470436 358345 470492 358401
rect 470492 358345 470496 358401
rect 470432 358341 470496 358345
rect 470512 358401 470576 358405
rect 470512 358345 470516 358401
rect 470516 358345 470572 358401
rect 470572 358345 470576 358401
rect 470512 358341 470576 358345
rect 470592 358401 470656 358405
rect 470592 358345 470596 358401
rect 470596 358345 470652 358401
rect 470652 358345 470656 358401
rect 470592 358341 470656 358345
rect 470672 358401 470736 358405
rect 470672 358345 470676 358401
rect 470676 358345 470732 358401
rect 470732 358345 470736 358401
rect 470672 358341 470736 358345
rect 470752 358401 470816 358405
rect 470752 358345 470756 358401
rect 470756 358345 470812 358401
rect 470812 358345 470816 358401
rect 470752 358341 470816 358345
rect 470272 358321 470336 358325
rect 470272 358265 470276 358321
rect 470276 358265 470332 358321
rect 470332 358265 470336 358321
rect 470272 358261 470336 358265
rect 470352 358321 470416 358325
rect 470352 358265 470356 358321
rect 470356 358265 470412 358321
rect 470412 358265 470416 358321
rect 470352 358261 470416 358265
rect 470432 358321 470496 358325
rect 470432 358265 470436 358321
rect 470436 358265 470492 358321
rect 470492 358265 470496 358321
rect 470432 358261 470496 358265
rect 470512 358321 470576 358325
rect 470512 358265 470516 358321
rect 470516 358265 470572 358321
rect 470572 358265 470576 358321
rect 470512 358261 470576 358265
rect 470592 358321 470656 358325
rect 470592 358265 470596 358321
rect 470596 358265 470652 358321
rect 470652 358265 470656 358321
rect 470592 358261 470656 358265
rect 470672 358321 470736 358325
rect 470672 358265 470676 358321
rect 470676 358265 470732 358321
rect 470732 358265 470736 358321
rect 470672 358261 470736 358265
rect 470752 358321 470816 358325
rect 470752 358265 470756 358321
rect 470756 358265 470812 358321
rect 470812 358265 470816 358321
rect 470752 358261 470816 358265
rect 470272 358241 470336 358245
rect 470272 358185 470276 358241
rect 470276 358185 470332 358241
rect 470332 358185 470336 358241
rect 470272 358181 470336 358185
rect 470352 358241 470416 358245
rect 470352 358185 470356 358241
rect 470356 358185 470412 358241
rect 470412 358185 470416 358241
rect 470352 358181 470416 358185
rect 470432 358241 470496 358245
rect 470432 358185 470436 358241
rect 470436 358185 470492 358241
rect 470492 358185 470496 358241
rect 470432 358181 470496 358185
rect 470512 358241 470576 358245
rect 470512 358185 470516 358241
rect 470516 358185 470572 358241
rect 470572 358185 470576 358241
rect 470512 358181 470576 358185
rect 470592 358241 470656 358245
rect 470592 358185 470596 358241
rect 470596 358185 470652 358241
rect 470652 358185 470656 358241
rect 470592 358181 470656 358185
rect 470672 358241 470736 358245
rect 470672 358185 470676 358241
rect 470676 358185 470732 358241
rect 470732 358185 470736 358241
rect 470672 358181 470736 358185
rect 470752 358241 470816 358245
rect 470752 358185 470756 358241
rect 470756 358185 470812 358241
rect 470812 358185 470816 358241
rect 470752 358181 470816 358185
rect 478644 357988 478708 358052
rect 481772 358048 481836 358052
rect 481772 357992 481822 358048
rect 481822 357992 481836 358048
rect 481772 357988 481836 357992
rect 484900 358048 484964 358052
rect 484900 357992 484950 358048
rect 484950 357992 484964 358048
rect 484900 357988 484964 357992
rect 488396 358048 488460 358052
rect 488396 357992 488410 358048
rect 488410 357992 488460 358048
rect 488396 357988 488460 357992
rect 474964 357504 475028 357508
rect 474964 357448 475014 357504
rect 475014 357448 475028 357504
rect 474964 357444 475028 357448
rect 469032 357395 469096 357399
rect 469032 357339 469036 357395
rect 469036 357339 469092 357395
rect 469092 357339 469096 357395
rect 469032 357335 469096 357339
rect 469112 357395 469176 357399
rect 469112 357339 469116 357395
rect 469116 357339 469172 357395
rect 469172 357339 469176 357395
rect 469112 357335 469176 357339
rect 469192 357395 469256 357399
rect 469192 357339 469196 357395
rect 469196 357339 469252 357395
rect 469252 357339 469256 357395
rect 469192 357335 469256 357339
rect 469272 357395 469336 357399
rect 469272 357339 469276 357395
rect 469276 357339 469332 357395
rect 469332 357339 469336 357395
rect 469272 357335 469336 357339
rect 469352 357395 469416 357399
rect 469352 357339 469356 357395
rect 469356 357339 469412 357395
rect 469412 357339 469416 357395
rect 469352 357335 469416 357339
rect 469432 357395 469496 357399
rect 469432 357339 469436 357395
rect 469436 357339 469492 357395
rect 469492 357339 469496 357395
rect 469432 357335 469496 357339
rect 469512 357395 469576 357399
rect 469512 357339 469516 357395
rect 469516 357339 469572 357395
rect 469572 357339 469576 357395
rect 469512 357335 469576 357339
rect 469032 357315 469096 357319
rect 469032 357259 469036 357315
rect 469036 357259 469092 357315
rect 469092 357259 469096 357315
rect 469032 357255 469096 357259
rect 469112 357315 469176 357319
rect 469112 357259 469116 357315
rect 469116 357259 469172 357315
rect 469172 357259 469176 357315
rect 469112 357255 469176 357259
rect 469192 357315 469256 357319
rect 469192 357259 469196 357315
rect 469196 357259 469252 357315
rect 469252 357259 469256 357315
rect 469192 357255 469256 357259
rect 469272 357315 469336 357319
rect 469272 357259 469276 357315
rect 469276 357259 469332 357315
rect 469332 357259 469336 357315
rect 469272 357255 469336 357259
rect 469352 357315 469416 357319
rect 469352 357259 469356 357315
rect 469356 357259 469412 357315
rect 469412 357259 469416 357315
rect 469352 357255 469416 357259
rect 469432 357315 469496 357319
rect 469432 357259 469436 357315
rect 469436 357259 469492 357315
rect 469492 357259 469496 357315
rect 469432 357255 469496 357259
rect 469512 357315 469576 357319
rect 469512 357259 469516 357315
rect 469516 357259 469572 357315
rect 469572 357259 469576 357315
rect 469512 357255 469576 357259
rect 469032 357235 469096 357239
rect 469032 357179 469036 357235
rect 469036 357179 469092 357235
rect 469092 357179 469096 357235
rect 469032 357175 469096 357179
rect 469112 357235 469176 357239
rect 469112 357179 469116 357235
rect 469116 357179 469172 357235
rect 469172 357179 469176 357235
rect 469112 357175 469176 357179
rect 469192 357235 469256 357239
rect 469192 357179 469196 357235
rect 469196 357179 469252 357235
rect 469252 357179 469256 357235
rect 469192 357175 469256 357179
rect 469272 357235 469336 357239
rect 469272 357179 469276 357235
rect 469276 357179 469332 357235
rect 469332 357179 469336 357235
rect 469272 357175 469336 357179
rect 469352 357235 469416 357239
rect 469352 357179 469356 357235
rect 469356 357179 469412 357235
rect 469412 357179 469416 357235
rect 469352 357175 469416 357179
rect 469432 357235 469496 357239
rect 469432 357179 469436 357235
rect 469436 357179 469492 357235
rect 469492 357179 469496 357235
rect 469432 357175 469496 357179
rect 469512 357235 469576 357239
rect 469512 357179 469516 357235
rect 469516 357179 469572 357235
rect 469572 357179 469576 357235
rect 469512 357175 469576 357179
rect 469032 357155 469096 357159
rect 469032 357099 469036 357155
rect 469036 357099 469092 357155
rect 469092 357099 469096 357155
rect 469032 357095 469096 357099
rect 469112 357155 469176 357159
rect 469112 357099 469116 357155
rect 469116 357099 469172 357155
rect 469172 357099 469176 357155
rect 469112 357095 469176 357099
rect 469192 357155 469256 357159
rect 469192 357099 469196 357155
rect 469196 357099 469252 357155
rect 469252 357099 469256 357155
rect 469192 357095 469256 357099
rect 469272 357155 469336 357159
rect 469272 357099 469276 357155
rect 469276 357099 469332 357155
rect 469332 357099 469336 357155
rect 469272 357095 469336 357099
rect 469352 357155 469416 357159
rect 469352 357099 469356 357155
rect 469356 357099 469412 357155
rect 469412 357099 469416 357155
rect 469352 357095 469416 357099
rect 469432 357155 469496 357159
rect 469432 357099 469436 357155
rect 469436 357099 469492 357155
rect 469492 357099 469496 357155
rect 469432 357095 469496 357099
rect 469512 357155 469576 357159
rect 469512 357099 469516 357155
rect 469516 357099 469572 357155
rect 469572 357099 469576 357155
rect 469512 357095 469576 357099
rect 470272 356308 470336 356312
rect 470272 356252 470276 356308
rect 470276 356252 470332 356308
rect 470332 356252 470336 356308
rect 470272 356248 470336 356252
rect 470352 356308 470416 356312
rect 470352 356252 470356 356308
rect 470356 356252 470412 356308
rect 470412 356252 470416 356308
rect 470352 356248 470416 356252
rect 470432 356308 470496 356312
rect 470432 356252 470436 356308
rect 470436 356252 470492 356308
rect 470492 356252 470496 356308
rect 470432 356248 470496 356252
rect 470512 356308 470576 356312
rect 470512 356252 470516 356308
rect 470516 356252 470572 356308
rect 470572 356252 470576 356308
rect 470512 356248 470576 356252
rect 470592 356308 470656 356312
rect 470592 356252 470596 356308
rect 470596 356252 470652 356308
rect 470652 356252 470656 356308
rect 470592 356248 470656 356252
rect 470672 356308 470736 356312
rect 470672 356252 470676 356308
rect 470676 356252 470732 356308
rect 470732 356252 470736 356308
rect 470672 356248 470736 356252
rect 470752 356308 470816 356312
rect 470752 356252 470756 356308
rect 470756 356252 470812 356308
rect 470812 356252 470816 356308
rect 470752 356248 470816 356252
rect 470272 356228 470336 356232
rect 470272 356172 470276 356228
rect 470276 356172 470332 356228
rect 470332 356172 470336 356228
rect 470272 356168 470336 356172
rect 470352 356228 470416 356232
rect 470352 356172 470356 356228
rect 470356 356172 470412 356228
rect 470412 356172 470416 356228
rect 470352 356168 470416 356172
rect 470432 356228 470496 356232
rect 470432 356172 470436 356228
rect 470436 356172 470492 356228
rect 470492 356172 470496 356228
rect 470432 356168 470496 356172
rect 470512 356228 470576 356232
rect 470512 356172 470516 356228
rect 470516 356172 470572 356228
rect 470572 356172 470576 356228
rect 470512 356168 470576 356172
rect 470592 356228 470656 356232
rect 470592 356172 470596 356228
rect 470596 356172 470652 356228
rect 470652 356172 470656 356228
rect 470592 356168 470656 356172
rect 470672 356228 470736 356232
rect 470672 356172 470676 356228
rect 470676 356172 470732 356228
rect 470732 356172 470736 356228
rect 470672 356168 470736 356172
rect 470752 356228 470816 356232
rect 470752 356172 470756 356228
rect 470756 356172 470812 356228
rect 470812 356172 470816 356228
rect 470752 356168 470816 356172
rect 470272 356148 470336 356152
rect 470272 356092 470276 356148
rect 470276 356092 470332 356148
rect 470332 356092 470336 356148
rect 470272 356088 470336 356092
rect 470352 356148 470416 356152
rect 470352 356092 470356 356148
rect 470356 356092 470412 356148
rect 470412 356092 470416 356148
rect 470352 356088 470416 356092
rect 470432 356148 470496 356152
rect 470432 356092 470436 356148
rect 470436 356092 470492 356148
rect 470492 356092 470496 356148
rect 470432 356088 470496 356092
rect 470512 356148 470576 356152
rect 470512 356092 470516 356148
rect 470516 356092 470572 356148
rect 470572 356092 470576 356148
rect 470512 356088 470576 356092
rect 470592 356148 470656 356152
rect 470592 356092 470596 356148
rect 470596 356092 470652 356148
rect 470652 356092 470656 356148
rect 470592 356088 470656 356092
rect 470672 356148 470736 356152
rect 470672 356092 470676 356148
rect 470676 356092 470732 356148
rect 470732 356092 470736 356148
rect 470672 356088 470736 356092
rect 470752 356148 470816 356152
rect 470752 356092 470756 356148
rect 470756 356092 470812 356148
rect 470812 356092 470816 356148
rect 470752 356088 470816 356092
rect 470272 356068 470336 356072
rect 470272 356012 470276 356068
rect 470276 356012 470332 356068
rect 470332 356012 470336 356068
rect 470272 356008 470336 356012
rect 470352 356068 470416 356072
rect 470352 356012 470356 356068
rect 470356 356012 470412 356068
rect 470412 356012 470416 356068
rect 470352 356008 470416 356012
rect 470432 356068 470496 356072
rect 470432 356012 470436 356068
rect 470436 356012 470492 356068
rect 470492 356012 470496 356068
rect 470432 356008 470496 356012
rect 470512 356068 470576 356072
rect 470512 356012 470516 356068
rect 470516 356012 470572 356068
rect 470572 356012 470576 356068
rect 470512 356008 470576 356012
rect 470592 356068 470656 356072
rect 470592 356012 470596 356068
rect 470596 356012 470652 356068
rect 470652 356012 470656 356068
rect 470592 356008 470656 356012
rect 470672 356068 470736 356072
rect 470672 356012 470676 356068
rect 470676 356012 470732 356068
rect 470732 356012 470736 356068
rect 470672 356008 470736 356012
rect 470752 356068 470816 356072
rect 470752 356012 470756 356068
rect 470756 356012 470812 356068
rect 470812 356012 470816 356068
rect 470752 356008 470816 356012
rect 544332 351868 544396 351932
rect 473676 343708 473740 343772
rect 474964 343708 475028 343772
rect 470272 342480 470336 342484
rect 470272 342424 470276 342480
rect 470276 342424 470332 342480
rect 470332 342424 470336 342480
rect 470272 342420 470336 342424
rect 470352 342480 470416 342484
rect 470352 342424 470356 342480
rect 470356 342424 470412 342480
rect 470412 342424 470416 342480
rect 470352 342420 470416 342424
rect 470432 342480 470496 342484
rect 470432 342424 470436 342480
rect 470436 342424 470492 342480
rect 470492 342424 470496 342480
rect 470432 342420 470496 342424
rect 470512 342480 470576 342484
rect 470512 342424 470516 342480
rect 470516 342424 470572 342480
rect 470572 342424 470576 342480
rect 470512 342420 470576 342424
rect 470592 342480 470656 342484
rect 470592 342424 470596 342480
rect 470596 342424 470652 342480
rect 470652 342424 470656 342480
rect 470592 342420 470656 342424
rect 470672 342480 470736 342484
rect 470672 342424 470676 342480
rect 470676 342424 470732 342480
rect 470732 342424 470736 342480
rect 470672 342420 470736 342424
rect 470752 342480 470816 342484
rect 470752 342424 470756 342480
rect 470756 342424 470812 342480
rect 470812 342424 470816 342480
rect 470752 342420 470816 342424
rect 470272 342400 470336 342404
rect 470272 342344 470276 342400
rect 470276 342344 470332 342400
rect 470332 342344 470336 342400
rect 470272 342340 470336 342344
rect 470352 342400 470416 342404
rect 470352 342344 470356 342400
rect 470356 342344 470412 342400
rect 470412 342344 470416 342400
rect 470352 342340 470416 342344
rect 470432 342400 470496 342404
rect 470432 342344 470436 342400
rect 470436 342344 470492 342400
rect 470492 342344 470496 342400
rect 470432 342340 470496 342344
rect 470512 342400 470576 342404
rect 470512 342344 470516 342400
rect 470516 342344 470572 342400
rect 470572 342344 470576 342400
rect 470512 342340 470576 342344
rect 470592 342400 470656 342404
rect 470592 342344 470596 342400
rect 470596 342344 470652 342400
rect 470652 342344 470656 342400
rect 470592 342340 470656 342344
rect 470672 342400 470736 342404
rect 470672 342344 470676 342400
rect 470676 342344 470732 342400
rect 470732 342344 470736 342400
rect 470672 342340 470736 342344
rect 470752 342400 470816 342404
rect 470752 342344 470756 342400
rect 470756 342344 470812 342400
rect 470812 342344 470816 342400
rect 470752 342340 470816 342344
rect 470272 342320 470336 342324
rect 470272 342264 470276 342320
rect 470276 342264 470332 342320
rect 470332 342264 470336 342320
rect 470272 342260 470336 342264
rect 470352 342320 470416 342324
rect 470352 342264 470356 342320
rect 470356 342264 470412 342320
rect 470412 342264 470416 342320
rect 470352 342260 470416 342264
rect 470432 342320 470496 342324
rect 470432 342264 470436 342320
rect 470436 342264 470492 342320
rect 470492 342264 470496 342320
rect 470432 342260 470496 342264
rect 470512 342320 470576 342324
rect 470512 342264 470516 342320
rect 470516 342264 470572 342320
rect 470572 342264 470576 342320
rect 470512 342260 470576 342264
rect 470592 342320 470656 342324
rect 470592 342264 470596 342320
rect 470596 342264 470652 342320
rect 470652 342264 470656 342320
rect 470592 342260 470656 342264
rect 470672 342320 470736 342324
rect 470672 342264 470676 342320
rect 470676 342264 470732 342320
rect 470732 342264 470736 342320
rect 470672 342260 470736 342264
rect 470752 342320 470816 342324
rect 470752 342264 470756 342320
rect 470756 342264 470812 342320
rect 470812 342264 470816 342320
rect 470752 342260 470816 342264
rect 470272 342240 470336 342244
rect 470272 342184 470276 342240
rect 470276 342184 470332 342240
rect 470332 342184 470336 342240
rect 470272 342180 470336 342184
rect 470352 342240 470416 342244
rect 470352 342184 470356 342240
rect 470356 342184 470412 342240
rect 470412 342184 470416 342240
rect 470352 342180 470416 342184
rect 470432 342240 470496 342244
rect 470432 342184 470436 342240
rect 470436 342184 470492 342240
rect 470492 342184 470496 342240
rect 470432 342180 470496 342184
rect 470512 342240 470576 342244
rect 470512 342184 470516 342240
rect 470516 342184 470572 342240
rect 470572 342184 470576 342240
rect 470512 342180 470576 342184
rect 470592 342240 470656 342244
rect 470592 342184 470596 342240
rect 470596 342184 470652 342240
rect 470652 342184 470656 342240
rect 470592 342180 470656 342184
rect 470672 342240 470736 342244
rect 470672 342184 470676 342240
rect 470676 342184 470732 342240
rect 470732 342184 470736 342240
rect 470672 342180 470736 342184
rect 470752 342240 470816 342244
rect 470752 342184 470756 342240
rect 470756 342184 470812 342240
rect 470812 342184 470816 342240
rect 470752 342180 470816 342184
rect 469032 341393 469096 341397
rect 469032 341337 469036 341393
rect 469036 341337 469092 341393
rect 469092 341337 469096 341393
rect 469032 341333 469096 341337
rect 469112 341393 469176 341397
rect 469112 341337 469116 341393
rect 469116 341337 469172 341393
rect 469172 341337 469176 341393
rect 469112 341333 469176 341337
rect 469192 341393 469256 341397
rect 469192 341337 469196 341393
rect 469196 341337 469252 341393
rect 469252 341337 469256 341393
rect 469192 341333 469256 341337
rect 469272 341393 469336 341397
rect 469272 341337 469276 341393
rect 469276 341337 469332 341393
rect 469332 341337 469336 341393
rect 469272 341333 469336 341337
rect 469352 341393 469416 341397
rect 469352 341337 469356 341393
rect 469356 341337 469412 341393
rect 469412 341337 469416 341393
rect 469352 341333 469416 341337
rect 469432 341393 469496 341397
rect 469432 341337 469436 341393
rect 469436 341337 469492 341393
rect 469492 341337 469496 341393
rect 469432 341333 469496 341337
rect 469512 341393 469576 341397
rect 469512 341337 469516 341393
rect 469516 341337 469572 341393
rect 469572 341337 469576 341393
rect 469512 341333 469576 341337
rect 469032 341313 469096 341317
rect 469032 341257 469036 341313
rect 469036 341257 469092 341313
rect 469092 341257 469096 341313
rect 469032 341253 469096 341257
rect 469112 341313 469176 341317
rect 469112 341257 469116 341313
rect 469116 341257 469172 341313
rect 469172 341257 469176 341313
rect 469112 341253 469176 341257
rect 469192 341313 469256 341317
rect 469192 341257 469196 341313
rect 469196 341257 469252 341313
rect 469252 341257 469256 341313
rect 469192 341253 469256 341257
rect 469272 341313 469336 341317
rect 469272 341257 469276 341313
rect 469276 341257 469332 341313
rect 469332 341257 469336 341313
rect 469272 341253 469336 341257
rect 469352 341313 469416 341317
rect 469352 341257 469356 341313
rect 469356 341257 469412 341313
rect 469412 341257 469416 341313
rect 469352 341253 469416 341257
rect 469432 341313 469496 341317
rect 469432 341257 469436 341313
rect 469436 341257 469492 341313
rect 469492 341257 469496 341313
rect 469432 341253 469496 341257
rect 469512 341313 469576 341317
rect 469512 341257 469516 341313
rect 469516 341257 469572 341313
rect 469572 341257 469576 341313
rect 469512 341253 469576 341257
rect 469032 341233 469096 341237
rect 469032 341177 469036 341233
rect 469036 341177 469092 341233
rect 469092 341177 469096 341233
rect 469032 341173 469096 341177
rect 469112 341233 469176 341237
rect 469112 341177 469116 341233
rect 469116 341177 469172 341233
rect 469172 341177 469176 341233
rect 469112 341173 469176 341177
rect 469192 341233 469256 341237
rect 469192 341177 469196 341233
rect 469196 341177 469252 341233
rect 469252 341177 469256 341233
rect 469192 341173 469256 341177
rect 469272 341233 469336 341237
rect 469272 341177 469276 341233
rect 469276 341177 469332 341233
rect 469332 341177 469336 341233
rect 469272 341173 469336 341177
rect 469352 341233 469416 341237
rect 469352 341177 469356 341233
rect 469356 341177 469412 341233
rect 469412 341177 469416 341233
rect 469352 341173 469416 341177
rect 469432 341233 469496 341237
rect 469432 341177 469436 341233
rect 469436 341177 469492 341233
rect 469492 341177 469496 341233
rect 469432 341173 469496 341177
rect 469512 341233 469576 341237
rect 469512 341177 469516 341233
rect 469516 341177 469572 341233
rect 469572 341177 469576 341233
rect 469512 341173 469576 341177
rect 469032 341153 469096 341157
rect 469032 341097 469036 341153
rect 469036 341097 469092 341153
rect 469092 341097 469096 341153
rect 469032 341093 469096 341097
rect 469112 341153 469176 341157
rect 469112 341097 469116 341153
rect 469116 341097 469172 341153
rect 469172 341097 469176 341153
rect 469112 341093 469176 341097
rect 469192 341153 469256 341157
rect 469192 341097 469196 341153
rect 469196 341097 469252 341153
rect 469252 341097 469256 341153
rect 469192 341093 469256 341097
rect 469272 341153 469336 341157
rect 469272 341097 469276 341153
rect 469276 341097 469332 341153
rect 469332 341097 469336 341153
rect 469272 341093 469336 341097
rect 469352 341153 469416 341157
rect 469352 341097 469356 341153
rect 469356 341097 469412 341153
rect 469412 341097 469416 341153
rect 469352 341093 469416 341097
rect 469432 341153 469496 341157
rect 469432 341097 469436 341153
rect 469436 341097 469492 341153
rect 469492 341097 469496 341153
rect 469432 341093 469496 341097
rect 469512 341153 469576 341157
rect 469512 341097 469516 341153
rect 469516 341097 469572 341153
rect 469572 341097 469576 341153
rect 469512 341093 469576 341097
rect 478460 340988 478524 341052
rect 481404 340988 481468 341052
rect 484164 340988 484228 341052
rect 488028 340988 488092 341052
rect 473676 340444 473740 340508
rect 470272 340308 470336 340312
rect 470272 340252 470276 340308
rect 470276 340252 470332 340308
rect 470332 340252 470336 340308
rect 470272 340248 470336 340252
rect 470352 340308 470416 340312
rect 470352 340252 470356 340308
rect 470356 340252 470412 340308
rect 470412 340252 470416 340308
rect 470352 340248 470416 340252
rect 470432 340308 470496 340312
rect 470432 340252 470436 340308
rect 470436 340252 470492 340308
rect 470492 340252 470496 340308
rect 470432 340248 470496 340252
rect 470512 340308 470576 340312
rect 470512 340252 470516 340308
rect 470516 340252 470572 340308
rect 470572 340252 470576 340308
rect 470512 340248 470576 340252
rect 470592 340308 470656 340312
rect 470592 340252 470596 340308
rect 470596 340252 470652 340308
rect 470652 340252 470656 340308
rect 470592 340248 470656 340252
rect 470672 340308 470736 340312
rect 470672 340252 470676 340308
rect 470676 340252 470732 340308
rect 470732 340252 470736 340308
rect 470672 340248 470736 340252
rect 470752 340308 470816 340312
rect 470752 340252 470756 340308
rect 470756 340252 470812 340308
rect 470812 340252 470816 340308
rect 470752 340248 470816 340252
rect 470272 340228 470336 340232
rect 470272 340172 470276 340228
rect 470276 340172 470332 340228
rect 470332 340172 470336 340228
rect 470272 340168 470336 340172
rect 470352 340228 470416 340232
rect 470352 340172 470356 340228
rect 470356 340172 470412 340228
rect 470412 340172 470416 340228
rect 470352 340168 470416 340172
rect 470432 340228 470496 340232
rect 470432 340172 470436 340228
rect 470436 340172 470492 340228
rect 470492 340172 470496 340228
rect 470432 340168 470496 340172
rect 470512 340228 470576 340232
rect 470512 340172 470516 340228
rect 470516 340172 470572 340228
rect 470572 340172 470576 340228
rect 470512 340168 470576 340172
rect 470592 340228 470656 340232
rect 470592 340172 470596 340228
rect 470596 340172 470652 340228
rect 470652 340172 470656 340228
rect 470592 340168 470656 340172
rect 470672 340228 470736 340232
rect 470672 340172 470676 340228
rect 470676 340172 470732 340228
rect 470732 340172 470736 340228
rect 470672 340168 470736 340172
rect 470752 340228 470816 340232
rect 470752 340172 470756 340228
rect 470756 340172 470812 340228
rect 470812 340172 470816 340228
rect 470752 340168 470816 340172
rect 470272 340148 470336 340152
rect 470272 340092 470276 340148
rect 470276 340092 470332 340148
rect 470332 340092 470336 340148
rect 470272 340088 470336 340092
rect 470352 340148 470416 340152
rect 470352 340092 470356 340148
rect 470356 340092 470412 340148
rect 470412 340092 470416 340148
rect 470352 340088 470416 340092
rect 470432 340148 470496 340152
rect 470432 340092 470436 340148
rect 470436 340092 470492 340148
rect 470492 340092 470496 340148
rect 470432 340088 470496 340092
rect 470512 340148 470576 340152
rect 470512 340092 470516 340148
rect 470516 340092 470572 340148
rect 470572 340092 470576 340148
rect 470512 340088 470576 340092
rect 470592 340148 470656 340152
rect 470592 340092 470596 340148
rect 470596 340092 470652 340148
rect 470652 340092 470656 340148
rect 470592 340088 470656 340092
rect 470672 340148 470736 340152
rect 470672 340092 470676 340148
rect 470676 340092 470732 340148
rect 470732 340092 470736 340148
rect 470672 340088 470736 340092
rect 470752 340148 470816 340152
rect 470752 340092 470756 340148
rect 470756 340092 470812 340148
rect 470812 340092 470816 340148
rect 470752 340088 470816 340092
rect 470272 340068 470336 340072
rect 470272 340012 470276 340068
rect 470276 340012 470332 340068
rect 470332 340012 470336 340068
rect 470272 340008 470336 340012
rect 470352 340068 470416 340072
rect 470352 340012 470356 340068
rect 470356 340012 470412 340068
rect 470412 340012 470416 340068
rect 470352 340008 470416 340012
rect 470432 340068 470496 340072
rect 470432 340012 470436 340068
rect 470436 340012 470492 340068
rect 470492 340012 470496 340068
rect 470432 340008 470496 340012
rect 470512 340068 470576 340072
rect 470512 340012 470516 340068
rect 470516 340012 470572 340068
rect 470572 340012 470576 340068
rect 470512 340008 470576 340012
rect 470592 340068 470656 340072
rect 470592 340012 470596 340068
rect 470596 340012 470652 340068
rect 470652 340012 470656 340068
rect 470592 340008 470656 340012
rect 470672 340068 470736 340072
rect 470672 340012 470676 340068
rect 470676 340012 470732 340068
rect 470732 340012 470736 340068
rect 470672 340008 470736 340012
rect 470752 340068 470816 340072
rect 470752 340012 470756 340068
rect 470756 340012 470812 340068
rect 470812 340012 470816 340068
rect 470752 340008 470816 340012
rect 541572 339492 541636 339556
rect 544332 339492 544396 339556
rect 486556 335412 486620 335476
rect 485636 334052 485700 334116
rect 486740 332692 486804 332756
rect 549300 326708 549364 326772
rect 470272 322480 470336 322484
rect 470272 322424 470276 322480
rect 470276 322424 470332 322480
rect 470332 322424 470336 322480
rect 470272 322420 470336 322424
rect 470352 322480 470416 322484
rect 470352 322424 470356 322480
rect 470356 322424 470412 322480
rect 470412 322424 470416 322480
rect 470352 322420 470416 322424
rect 470432 322480 470496 322484
rect 470432 322424 470436 322480
rect 470436 322424 470492 322480
rect 470492 322424 470496 322480
rect 470432 322420 470496 322424
rect 470512 322480 470576 322484
rect 470512 322424 470516 322480
rect 470516 322424 470572 322480
rect 470572 322424 470576 322480
rect 470512 322420 470576 322424
rect 470592 322480 470656 322484
rect 470592 322424 470596 322480
rect 470596 322424 470652 322480
rect 470652 322424 470656 322480
rect 470592 322420 470656 322424
rect 470672 322480 470736 322484
rect 470672 322424 470676 322480
rect 470676 322424 470732 322480
rect 470732 322424 470736 322480
rect 470672 322420 470736 322424
rect 470752 322480 470816 322484
rect 470752 322424 470756 322480
rect 470756 322424 470812 322480
rect 470812 322424 470816 322480
rect 470752 322420 470816 322424
rect 470272 322400 470336 322404
rect 470272 322344 470276 322400
rect 470276 322344 470332 322400
rect 470332 322344 470336 322400
rect 470272 322340 470336 322344
rect 470352 322400 470416 322404
rect 470352 322344 470356 322400
rect 470356 322344 470412 322400
rect 470412 322344 470416 322400
rect 470352 322340 470416 322344
rect 470432 322400 470496 322404
rect 470432 322344 470436 322400
rect 470436 322344 470492 322400
rect 470492 322344 470496 322400
rect 470432 322340 470496 322344
rect 470512 322400 470576 322404
rect 470512 322344 470516 322400
rect 470516 322344 470572 322400
rect 470572 322344 470576 322400
rect 470512 322340 470576 322344
rect 470592 322400 470656 322404
rect 470592 322344 470596 322400
rect 470596 322344 470652 322400
rect 470652 322344 470656 322400
rect 470592 322340 470656 322344
rect 470672 322400 470736 322404
rect 470672 322344 470676 322400
rect 470676 322344 470732 322400
rect 470732 322344 470736 322400
rect 470672 322340 470736 322344
rect 470752 322400 470816 322404
rect 470752 322344 470756 322400
rect 470756 322344 470812 322400
rect 470812 322344 470816 322400
rect 470752 322340 470816 322344
rect 470272 322320 470336 322324
rect 470272 322264 470276 322320
rect 470276 322264 470332 322320
rect 470332 322264 470336 322320
rect 470272 322260 470336 322264
rect 470352 322320 470416 322324
rect 470352 322264 470356 322320
rect 470356 322264 470412 322320
rect 470412 322264 470416 322320
rect 470352 322260 470416 322264
rect 470432 322320 470496 322324
rect 470432 322264 470436 322320
rect 470436 322264 470492 322320
rect 470492 322264 470496 322320
rect 470432 322260 470496 322264
rect 470512 322320 470576 322324
rect 470512 322264 470516 322320
rect 470516 322264 470572 322320
rect 470572 322264 470576 322320
rect 470512 322260 470576 322264
rect 470592 322320 470656 322324
rect 470592 322264 470596 322320
rect 470596 322264 470652 322320
rect 470652 322264 470656 322320
rect 470592 322260 470656 322264
rect 470672 322320 470736 322324
rect 470672 322264 470676 322320
rect 470676 322264 470732 322320
rect 470732 322264 470736 322320
rect 470672 322260 470736 322264
rect 470752 322320 470816 322324
rect 470752 322264 470756 322320
rect 470756 322264 470812 322320
rect 470812 322264 470816 322320
rect 470752 322260 470816 322264
rect 470272 322240 470336 322244
rect 470272 322184 470276 322240
rect 470276 322184 470332 322240
rect 470332 322184 470336 322240
rect 470272 322180 470336 322184
rect 470352 322240 470416 322244
rect 470352 322184 470356 322240
rect 470356 322184 470412 322240
rect 470412 322184 470416 322240
rect 470352 322180 470416 322184
rect 470432 322240 470496 322244
rect 470432 322184 470436 322240
rect 470436 322184 470492 322240
rect 470492 322184 470496 322240
rect 470432 322180 470496 322184
rect 470512 322240 470576 322244
rect 470512 322184 470516 322240
rect 470516 322184 470572 322240
rect 470572 322184 470576 322240
rect 470512 322180 470576 322184
rect 470592 322240 470656 322244
rect 470592 322184 470596 322240
rect 470596 322184 470652 322240
rect 470652 322184 470656 322240
rect 470592 322180 470656 322184
rect 470672 322240 470736 322244
rect 470672 322184 470676 322240
rect 470676 322184 470732 322240
rect 470732 322184 470736 322240
rect 470672 322180 470736 322184
rect 470752 322240 470816 322244
rect 470752 322184 470756 322240
rect 470756 322184 470812 322240
rect 470812 322184 470816 322240
rect 470752 322180 470816 322184
rect 469032 321393 469096 321397
rect 469032 321337 469036 321393
rect 469036 321337 469092 321393
rect 469092 321337 469096 321393
rect 469032 321333 469096 321337
rect 469112 321393 469176 321397
rect 469112 321337 469116 321393
rect 469116 321337 469172 321393
rect 469172 321337 469176 321393
rect 469112 321333 469176 321337
rect 469192 321393 469256 321397
rect 469192 321337 469196 321393
rect 469196 321337 469252 321393
rect 469252 321337 469256 321393
rect 469192 321333 469256 321337
rect 469272 321393 469336 321397
rect 469272 321337 469276 321393
rect 469276 321337 469332 321393
rect 469332 321337 469336 321393
rect 469272 321333 469336 321337
rect 469352 321393 469416 321397
rect 469352 321337 469356 321393
rect 469356 321337 469412 321393
rect 469412 321337 469416 321393
rect 469352 321333 469416 321337
rect 469432 321393 469496 321397
rect 469432 321337 469436 321393
rect 469436 321337 469492 321393
rect 469492 321337 469496 321393
rect 469432 321333 469496 321337
rect 469512 321393 469576 321397
rect 469512 321337 469516 321393
rect 469516 321337 469572 321393
rect 469572 321337 469576 321393
rect 469512 321333 469576 321337
rect 469032 321313 469096 321317
rect 469032 321257 469036 321313
rect 469036 321257 469092 321313
rect 469092 321257 469096 321313
rect 469032 321253 469096 321257
rect 469112 321313 469176 321317
rect 469112 321257 469116 321313
rect 469116 321257 469172 321313
rect 469172 321257 469176 321313
rect 469112 321253 469176 321257
rect 469192 321313 469256 321317
rect 469192 321257 469196 321313
rect 469196 321257 469252 321313
rect 469252 321257 469256 321313
rect 469192 321253 469256 321257
rect 469272 321313 469336 321317
rect 469272 321257 469276 321313
rect 469276 321257 469332 321313
rect 469332 321257 469336 321313
rect 469272 321253 469336 321257
rect 469352 321313 469416 321317
rect 469352 321257 469356 321313
rect 469356 321257 469412 321313
rect 469412 321257 469416 321313
rect 469352 321253 469416 321257
rect 469432 321313 469496 321317
rect 469432 321257 469436 321313
rect 469436 321257 469492 321313
rect 469492 321257 469496 321313
rect 469432 321253 469496 321257
rect 469512 321313 469576 321317
rect 469512 321257 469516 321313
rect 469516 321257 469572 321313
rect 469572 321257 469576 321313
rect 469512 321253 469576 321257
rect 473676 321268 473740 321332
rect 484164 321268 484228 321332
rect 469032 321233 469096 321237
rect 469032 321177 469036 321233
rect 469036 321177 469092 321233
rect 469092 321177 469096 321233
rect 469032 321173 469096 321177
rect 469112 321233 469176 321237
rect 469112 321177 469116 321233
rect 469116 321177 469172 321233
rect 469172 321177 469176 321233
rect 469112 321173 469176 321177
rect 469192 321233 469256 321237
rect 469192 321177 469196 321233
rect 469196 321177 469252 321233
rect 469252 321177 469256 321233
rect 469192 321173 469256 321177
rect 469272 321233 469336 321237
rect 469272 321177 469276 321233
rect 469276 321177 469332 321233
rect 469332 321177 469336 321233
rect 469272 321173 469336 321177
rect 469352 321233 469416 321237
rect 469352 321177 469356 321233
rect 469356 321177 469412 321233
rect 469412 321177 469416 321233
rect 469352 321173 469416 321177
rect 469432 321233 469496 321237
rect 469432 321177 469436 321233
rect 469436 321177 469492 321233
rect 469492 321177 469496 321233
rect 469432 321173 469496 321177
rect 469512 321233 469576 321237
rect 469512 321177 469516 321233
rect 469516 321177 469572 321233
rect 469572 321177 469576 321233
rect 469512 321173 469576 321177
rect 469032 321153 469096 321157
rect 469032 321097 469036 321153
rect 469036 321097 469092 321153
rect 469092 321097 469096 321153
rect 469032 321093 469096 321097
rect 469112 321153 469176 321157
rect 469112 321097 469116 321153
rect 469116 321097 469172 321153
rect 469172 321097 469176 321153
rect 469112 321093 469176 321097
rect 469192 321153 469256 321157
rect 469192 321097 469196 321153
rect 469196 321097 469252 321153
rect 469252 321097 469256 321153
rect 469192 321093 469256 321097
rect 469272 321153 469336 321157
rect 469272 321097 469276 321153
rect 469276 321097 469332 321153
rect 469332 321097 469336 321153
rect 469272 321093 469336 321097
rect 469352 321153 469416 321157
rect 469352 321097 469356 321153
rect 469356 321097 469412 321153
rect 469412 321097 469416 321153
rect 469352 321093 469416 321097
rect 469432 321153 469496 321157
rect 469432 321097 469436 321153
rect 469436 321097 469492 321153
rect 469492 321097 469496 321153
rect 469432 321093 469496 321097
rect 469512 321153 469576 321157
rect 469512 321097 469516 321153
rect 469516 321097 469572 321153
rect 469572 321097 469576 321153
rect 469512 321093 469576 321097
rect 488028 320996 488092 321060
rect 478644 320860 478708 320924
rect 481588 320920 481652 320924
rect 481588 320864 481602 320920
rect 481602 320864 481652 320920
rect 481588 320860 481652 320864
rect 470272 320308 470336 320312
rect 470272 320252 470276 320308
rect 470276 320252 470332 320308
rect 470332 320252 470336 320308
rect 470272 320248 470336 320252
rect 470352 320308 470416 320312
rect 470352 320252 470356 320308
rect 470356 320252 470412 320308
rect 470412 320252 470416 320308
rect 470352 320248 470416 320252
rect 470432 320308 470496 320312
rect 470432 320252 470436 320308
rect 470436 320252 470492 320308
rect 470492 320252 470496 320308
rect 470432 320248 470496 320252
rect 470512 320308 470576 320312
rect 470512 320252 470516 320308
rect 470516 320252 470572 320308
rect 470572 320252 470576 320308
rect 470512 320248 470576 320252
rect 470592 320308 470656 320312
rect 470592 320252 470596 320308
rect 470596 320252 470652 320308
rect 470652 320252 470656 320308
rect 470592 320248 470656 320252
rect 470672 320308 470736 320312
rect 470672 320252 470676 320308
rect 470676 320252 470732 320308
rect 470732 320252 470736 320308
rect 470672 320248 470736 320252
rect 470752 320308 470816 320312
rect 470752 320252 470756 320308
rect 470756 320252 470812 320308
rect 470812 320252 470816 320308
rect 470752 320248 470816 320252
rect 470272 320228 470336 320232
rect 470272 320172 470276 320228
rect 470276 320172 470332 320228
rect 470332 320172 470336 320228
rect 470272 320168 470336 320172
rect 470352 320228 470416 320232
rect 470352 320172 470356 320228
rect 470356 320172 470412 320228
rect 470412 320172 470416 320228
rect 470352 320168 470416 320172
rect 470432 320228 470496 320232
rect 470432 320172 470436 320228
rect 470436 320172 470492 320228
rect 470492 320172 470496 320228
rect 470432 320168 470496 320172
rect 470512 320228 470576 320232
rect 470512 320172 470516 320228
rect 470516 320172 470572 320228
rect 470572 320172 470576 320228
rect 470512 320168 470576 320172
rect 470592 320228 470656 320232
rect 470592 320172 470596 320228
rect 470596 320172 470652 320228
rect 470652 320172 470656 320228
rect 470592 320168 470656 320172
rect 470672 320228 470736 320232
rect 470672 320172 470676 320228
rect 470676 320172 470732 320228
rect 470732 320172 470736 320228
rect 470672 320168 470736 320172
rect 470752 320228 470816 320232
rect 470752 320172 470756 320228
rect 470756 320172 470812 320228
rect 470812 320172 470816 320228
rect 470752 320168 470816 320172
rect 470272 320148 470336 320152
rect 470272 320092 470276 320148
rect 470276 320092 470332 320148
rect 470332 320092 470336 320148
rect 470272 320088 470336 320092
rect 470352 320148 470416 320152
rect 470352 320092 470356 320148
rect 470356 320092 470412 320148
rect 470412 320092 470416 320148
rect 470352 320088 470416 320092
rect 470432 320148 470496 320152
rect 470432 320092 470436 320148
rect 470436 320092 470492 320148
rect 470492 320092 470496 320148
rect 470432 320088 470496 320092
rect 470512 320148 470576 320152
rect 470512 320092 470516 320148
rect 470516 320092 470572 320148
rect 470572 320092 470576 320148
rect 470512 320088 470576 320092
rect 470592 320148 470656 320152
rect 470592 320092 470596 320148
rect 470596 320092 470652 320148
rect 470652 320092 470656 320148
rect 470592 320088 470656 320092
rect 470672 320148 470736 320152
rect 470672 320092 470676 320148
rect 470676 320092 470732 320148
rect 470732 320092 470736 320148
rect 470672 320088 470736 320092
rect 470752 320148 470816 320152
rect 470752 320092 470756 320148
rect 470756 320092 470812 320148
rect 470812 320092 470816 320148
rect 470752 320088 470816 320092
rect 470272 320068 470336 320072
rect 470272 320012 470276 320068
rect 470276 320012 470332 320068
rect 470332 320012 470336 320068
rect 470272 320008 470336 320012
rect 470352 320068 470416 320072
rect 470352 320012 470356 320068
rect 470356 320012 470412 320068
rect 470412 320012 470416 320068
rect 470352 320008 470416 320012
rect 470432 320068 470496 320072
rect 470432 320012 470436 320068
rect 470436 320012 470492 320068
rect 470492 320012 470496 320068
rect 470432 320008 470496 320012
rect 470512 320068 470576 320072
rect 470512 320012 470516 320068
rect 470516 320012 470572 320068
rect 470572 320012 470576 320068
rect 470512 320008 470576 320012
rect 470592 320068 470656 320072
rect 470592 320012 470596 320068
rect 470596 320012 470652 320068
rect 470652 320012 470656 320068
rect 470592 320008 470656 320012
rect 470672 320068 470736 320072
rect 470672 320012 470676 320068
rect 470676 320012 470732 320068
rect 470732 320012 470736 320068
rect 470672 320008 470736 320012
rect 470752 320068 470816 320072
rect 470752 320012 470756 320068
rect 470756 320012 470812 320068
rect 470812 320012 470816 320068
rect 470752 320008 470816 320012
rect 470272 307080 470336 307084
rect 470272 307024 470276 307080
rect 470276 307024 470332 307080
rect 470332 307024 470336 307080
rect 470272 307020 470336 307024
rect 470352 307080 470416 307084
rect 470352 307024 470356 307080
rect 470356 307024 470412 307080
rect 470412 307024 470416 307080
rect 470352 307020 470416 307024
rect 470432 307080 470496 307084
rect 470432 307024 470436 307080
rect 470436 307024 470492 307080
rect 470492 307024 470496 307080
rect 470432 307020 470496 307024
rect 470512 307080 470576 307084
rect 470512 307024 470516 307080
rect 470516 307024 470572 307080
rect 470572 307024 470576 307080
rect 470512 307020 470576 307024
rect 470592 307080 470656 307084
rect 470592 307024 470596 307080
rect 470596 307024 470652 307080
rect 470652 307024 470656 307080
rect 470592 307020 470656 307024
rect 470672 307080 470736 307084
rect 470672 307024 470676 307080
rect 470676 307024 470732 307080
rect 470732 307024 470736 307080
rect 470672 307020 470736 307024
rect 470752 307080 470816 307084
rect 470752 307024 470756 307080
rect 470756 307024 470812 307080
rect 470812 307024 470816 307080
rect 470752 307020 470816 307024
rect 470272 307000 470336 307004
rect 470272 306944 470276 307000
rect 470276 306944 470332 307000
rect 470332 306944 470336 307000
rect 470272 306940 470336 306944
rect 470352 307000 470416 307004
rect 470352 306944 470356 307000
rect 470356 306944 470412 307000
rect 470412 306944 470416 307000
rect 470352 306940 470416 306944
rect 470432 307000 470496 307004
rect 470432 306944 470436 307000
rect 470436 306944 470492 307000
rect 470492 306944 470496 307000
rect 470432 306940 470496 306944
rect 470512 307000 470576 307004
rect 470512 306944 470516 307000
rect 470516 306944 470572 307000
rect 470572 306944 470576 307000
rect 470512 306940 470576 306944
rect 470592 307000 470656 307004
rect 470592 306944 470596 307000
rect 470596 306944 470652 307000
rect 470652 306944 470656 307000
rect 470592 306940 470656 306944
rect 470672 307000 470736 307004
rect 470672 306944 470676 307000
rect 470676 306944 470732 307000
rect 470732 306944 470736 307000
rect 470672 306940 470736 306944
rect 470752 307000 470816 307004
rect 470752 306944 470756 307000
rect 470756 306944 470812 307000
rect 470812 306944 470816 307000
rect 470752 306940 470816 306944
rect 470272 306920 470336 306924
rect 470272 306864 470276 306920
rect 470276 306864 470332 306920
rect 470332 306864 470336 306920
rect 470272 306860 470336 306864
rect 470352 306920 470416 306924
rect 470352 306864 470356 306920
rect 470356 306864 470412 306920
rect 470412 306864 470416 306920
rect 470352 306860 470416 306864
rect 470432 306920 470496 306924
rect 470432 306864 470436 306920
rect 470436 306864 470492 306920
rect 470492 306864 470496 306920
rect 470432 306860 470496 306864
rect 470512 306920 470576 306924
rect 470512 306864 470516 306920
rect 470516 306864 470572 306920
rect 470572 306864 470576 306920
rect 470512 306860 470576 306864
rect 470592 306920 470656 306924
rect 470592 306864 470596 306920
rect 470596 306864 470652 306920
rect 470652 306864 470656 306920
rect 470592 306860 470656 306864
rect 470672 306920 470736 306924
rect 470672 306864 470676 306920
rect 470676 306864 470732 306920
rect 470732 306864 470736 306920
rect 470672 306860 470736 306864
rect 470752 306920 470816 306924
rect 470752 306864 470756 306920
rect 470756 306864 470812 306920
rect 470812 306864 470816 306920
rect 470752 306860 470816 306864
rect 470272 306840 470336 306844
rect 470272 306784 470276 306840
rect 470276 306784 470332 306840
rect 470332 306784 470336 306840
rect 470272 306780 470336 306784
rect 470352 306840 470416 306844
rect 470352 306784 470356 306840
rect 470356 306784 470412 306840
rect 470412 306784 470416 306840
rect 470352 306780 470416 306784
rect 470432 306840 470496 306844
rect 470432 306784 470436 306840
rect 470436 306784 470492 306840
rect 470492 306784 470496 306840
rect 470432 306780 470496 306784
rect 470512 306840 470576 306844
rect 470512 306784 470516 306840
rect 470516 306784 470572 306840
rect 470572 306784 470576 306840
rect 470512 306780 470576 306784
rect 470592 306840 470656 306844
rect 470592 306784 470596 306840
rect 470596 306784 470652 306840
rect 470652 306784 470656 306840
rect 470592 306780 470656 306784
rect 470672 306840 470736 306844
rect 470672 306784 470676 306840
rect 470676 306784 470732 306840
rect 470732 306784 470736 306840
rect 470672 306780 470736 306784
rect 470752 306840 470816 306844
rect 470752 306784 470756 306840
rect 470756 306784 470812 306840
rect 470812 306784 470816 306840
rect 470752 306780 470816 306784
rect 487660 306308 487724 306372
rect 481588 306036 481652 306100
rect 469032 305995 469096 305999
rect 469032 305939 469036 305995
rect 469036 305939 469092 305995
rect 469092 305939 469096 305995
rect 469032 305935 469096 305939
rect 469112 305995 469176 305999
rect 469112 305939 469116 305995
rect 469116 305939 469172 305995
rect 469172 305939 469176 305995
rect 469112 305935 469176 305939
rect 469192 305995 469256 305999
rect 469192 305939 469196 305995
rect 469196 305939 469252 305995
rect 469252 305939 469256 305995
rect 469192 305935 469256 305939
rect 469272 305995 469336 305999
rect 469272 305939 469276 305995
rect 469276 305939 469332 305995
rect 469332 305939 469336 305995
rect 469272 305935 469336 305939
rect 469352 305995 469416 305999
rect 469352 305939 469356 305995
rect 469356 305939 469412 305995
rect 469412 305939 469416 305995
rect 469352 305935 469416 305939
rect 469432 305995 469496 305999
rect 469432 305939 469436 305995
rect 469436 305939 469492 305995
rect 469492 305939 469496 305995
rect 469432 305935 469496 305939
rect 469512 305995 469576 305999
rect 469512 305939 469516 305995
rect 469516 305939 469572 305995
rect 469572 305939 469576 305995
rect 469512 305935 469576 305939
rect 469032 305915 469096 305919
rect 469032 305859 469036 305915
rect 469036 305859 469092 305915
rect 469092 305859 469096 305915
rect 469032 305855 469096 305859
rect 469112 305915 469176 305919
rect 469112 305859 469116 305915
rect 469116 305859 469172 305915
rect 469172 305859 469176 305915
rect 469112 305855 469176 305859
rect 469192 305915 469256 305919
rect 469192 305859 469196 305915
rect 469196 305859 469252 305915
rect 469252 305859 469256 305915
rect 469192 305855 469256 305859
rect 469272 305915 469336 305919
rect 469272 305859 469276 305915
rect 469276 305859 469332 305915
rect 469332 305859 469336 305915
rect 469272 305855 469336 305859
rect 469352 305915 469416 305919
rect 469352 305859 469356 305915
rect 469356 305859 469412 305915
rect 469412 305859 469416 305915
rect 469352 305855 469416 305859
rect 469432 305915 469496 305919
rect 469432 305859 469436 305915
rect 469436 305859 469492 305915
rect 469492 305859 469496 305915
rect 469432 305855 469496 305859
rect 469512 305915 469576 305919
rect 469512 305859 469516 305915
rect 469516 305859 469572 305915
rect 469572 305859 469576 305915
rect 469512 305855 469576 305859
rect 473676 305960 473740 305964
rect 473676 305904 473726 305960
rect 473726 305904 473740 305960
rect 473676 305900 473740 305904
rect 469032 305835 469096 305839
rect 469032 305779 469036 305835
rect 469036 305779 469092 305835
rect 469092 305779 469096 305835
rect 469032 305775 469096 305779
rect 469112 305835 469176 305839
rect 469112 305779 469116 305835
rect 469116 305779 469172 305835
rect 469172 305779 469176 305835
rect 469112 305775 469176 305779
rect 469192 305835 469256 305839
rect 469192 305779 469196 305835
rect 469196 305779 469252 305835
rect 469252 305779 469256 305835
rect 469192 305775 469256 305779
rect 469272 305835 469336 305839
rect 469272 305779 469276 305835
rect 469276 305779 469332 305835
rect 469332 305779 469336 305835
rect 469272 305775 469336 305779
rect 469352 305835 469416 305839
rect 469352 305779 469356 305835
rect 469356 305779 469412 305835
rect 469412 305779 469416 305835
rect 469352 305775 469416 305779
rect 469432 305835 469496 305839
rect 469432 305779 469436 305835
rect 469436 305779 469492 305835
rect 469492 305779 469496 305835
rect 469432 305775 469496 305779
rect 469512 305835 469576 305839
rect 469512 305779 469516 305835
rect 469516 305779 469572 305835
rect 469572 305779 469576 305835
rect 469512 305775 469576 305779
rect 469032 305755 469096 305759
rect 469032 305699 469036 305755
rect 469036 305699 469092 305755
rect 469092 305699 469096 305755
rect 469032 305695 469096 305699
rect 469112 305755 469176 305759
rect 469112 305699 469116 305755
rect 469116 305699 469172 305755
rect 469172 305699 469176 305755
rect 469112 305695 469176 305699
rect 469192 305755 469256 305759
rect 469192 305699 469196 305755
rect 469196 305699 469252 305755
rect 469252 305699 469256 305755
rect 469192 305695 469256 305699
rect 469272 305755 469336 305759
rect 469272 305699 469276 305755
rect 469276 305699 469332 305755
rect 469332 305699 469336 305755
rect 469272 305695 469336 305699
rect 469352 305755 469416 305759
rect 469352 305699 469356 305755
rect 469356 305699 469412 305755
rect 469412 305699 469416 305755
rect 469352 305695 469416 305699
rect 469432 305755 469496 305759
rect 469432 305699 469436 305755
rect 469436 305699 469492 305755
rect 469492 305699 469496 305755
rect 469432 305695 469496 305699
rect 469512 305755 469576 305759
rect 469512 305699 469516 305755
rect 469516 305699 469572 305755
rect 469572 305699 469576 305755
rect 469512 305695 469576 305699
rect 478828 305628 478892 305692
rect 484164 305552 484228 305556
rect 484164 305496 484178 305552
rect 484178 305496 484228 305552
rect 484164 305492 484228 305496
rect 470272 304908 470336 304912
rect 470272 304852 470276 304908
rect 470276 304852 470332 304908
rect 470332 304852 470336 304908
rect 470272 304848 470336 304852
rect 470352 304908 470416 304912
rect 470352 304852 470356 304908
rect 470356 304852 470412 304908
rect 470412 304852 470416 304908
rect 470352 304848 470416 304852
rect 470432 304908 470496 304912
rect 470432 304852 470436 304908
rect 470436 304852 470492 304908
rect 470492 304852 470496 304908
rect 470432 304848 470496 304852
rect 470512 304908 470576 304912
rect 470512 304852 470516 304908
rect 470516 304852 470572 304908
rect 470572 304852 470576 304908
rect 470512 304848 470576 304852
rect 470592 304908 470656 304912
rect 470592 304852 470596 304908
rect 470596 304852 470652 304908
rect 470652 304852 470656 304908
rect 470592 304848 470656 304852
rect 470672 304908 470736 304912
rect 470672 304852 470676 304908
rect 470676 304852 470732 304908
rect 470732 304852 470736 304908
rect 470672 304848 470736 304852
rect 470752 304908 470816 304912
rect 470752 304852 470756 304908
rect 470756 304852 470812 304908
rect 470812 304852 470816 304908
rect 470752 304848 470816 304852
rect 470272 304828 470336 304832
rect 470272 304772 470276 304828
rect 470276 304772 470332 304828
rect 470332 304772 470336 304828
rect 470272 304768 470336 304772
rect 470352 304828 470416 304832
rect 470352 304772 470356 304828
rect 470356 304772 470412 304828
rect 470412 304772 470416 304828
rect 470352 304768 470416 304772
rect 470432 304828 470496 304832
rect 470432 304772 470436 304828
rect 470436 304772 470492 304828
rect 470492 304772 470496 304828
rect 470432 304768 470496 304772
rect 470512 304828 470576 304832
rect 470512 304772 470516 304828
rect 470516 304772 470572 304828
rect 470572 304772 470576 304828
rect 470512 304768 470576 304772
rect 470592 304828 470656 304832
rect 470592 304772 470596 304828
rect 470596 304772 470652 304828
rect 470652 304772 470656 304828
rect 470592 304768 470656 304772
rect 470672 304828 470736 304832
rect 470672 304772 470676 304828
rect 470676 304772 470732 304828
rect 470732 304772 470736 304828
rect 470672 304768 470736 304772
rect 470752 304828 470816 304832
rect 470752 304772 470756 304828
rect 470756 304772 470812 304828
rect 470812 304772 470816 304828
rect 470752 304768 470816 304772
rect 470272 304748 470336 304752
rect 470272 304692 470276 304748
rect 470276 304692 470332 304748
rect 470332 304692 470336 304748
rect 470272 304688 470336 304692
rect 470352 304748 470416 304752
rect 470352 304692 470356 304748
rect 470356 304692 470412 304748
rect 470412 304692 470416 304748
rect 470352 304688 470416 304692
rect 470432 304748 470496 304752
rect 470432 304692 470436 304748
rect 470436 304692 470492 304748
rect 470492 304692 470496 304748
rect 470432 304688 470496 304692
rect 470512 304748 470576 304752
rect 470512 304692 470516 304748
rect 470516 304692 470572 304748
rect 470572 304692 470576 304748
rect 470512 304688 470576 304692
rect 470592 304748 470656 304752
rect 470592 304692 470596 304748
rect 470596 304692 470652 304748
rect 470652 304692 470656 304748
rect 470592 304688 470656 304692
rect 470672 304748 470736 304752
rect 470672 304692 470676 304748
rect 470676 304692 470732 304748
rect 470732 304692 470736 304748
rect 470672 304688 470736 304692
rect 470752 304748 470816 304752
rect 470752 304692 470756 304748
rect 470756 304692 470812 304748
rect 470812 304692 470816 304748
rect 470752 304688 470816 304692
rect 470272 304668 470336 304672
rect 470272 304612 470276 304668
rect 470276 304612 470332 304668
rect 470332 304612 470336 304668
rect 470272 304608 470336 304612
rect 470352 304668 470416 304672
rect 470352 304612 470356 304668
rect 470356 304612 470412 304668
rect 470412 304612 470416 304668
rect 470352 304608 470416 304612
rect 470432 304668 470496 304672
rect 470432 304612 470436 304668
rect 470436 304612 470492 304668
rect 470492 304612 470496 304668
rect 470432 304608 470496 304612
rect 470512 304668 470576 304672
rect 470512 304612 470516 304668
rect 470516 304612 470572 304668
rect 470572 304612 470576 304668
rect 470512 304608 470576 304612
rect 470592 304668 470656 304672
rect 470592 304612 470596 304668
rect 470596 304612 470652 304668
rect 470652 304612 470656 304668
rect 470592 304608 470656 304612
rect 470672 304668 470736 304672
rect 470672 304612 470676 304668
rect 470676 304612 470732 304668
rect 470732 304612 470736 304668
rect 470672 304608 470736 304612
rect 470752 304668 470816 304672
rect 470752 304612 470756 304668
rect 470756 304612 470812 304668
rect 470812 304612 470816 304668
rect 470752 304608 470816 304612
rect 544332 303724 544396 303788
rect 541572 303588 541636 303652
rect 549300 290668 549364 290732
rect 473676 289716 473740 289780
rect 476068 289716 476132 289780
rect 484164 289716 484228 289780
rect 485820 289716 485884 289780
rect 470272 287481 470336 287485
rect 470272 287425 470276 287481
rect 470276 287425 470332 287481
rect 470332 287425 470336 287481
rect 470272 287421 470336 287425
rect 470352 287481 470416 287485
rect 470352 287425 470356 287481
rect 470356 287425 470412 287481
rect 470412 287425 470416 287481
rect 470352 287421 470416 287425
rect 470432 287481 470496 287485
rect 470432 287425 470436 287481
rect 470436 287425 470492 287481
rect 470492 287425 470496 287481
rect 470432 287421 470496 287425
rect 470512 287481 470576 287485
rect 470512 287425 470516 287481
rect 470516 287425 470572 287481
rect 470572 287425 470576 287481
rect 470512 287421 470576 287425
rect 470592 287481 470656 287485
rect 470592 287425 470596 287481
rect 470596 287425 470652 287481
rect 470652 287425 470656 287481
rect 470592 287421 470656 287425
rect 470672 287481 470736 287485
rect 470672 287425 470676 287481
rect 470676 287425 470732 287481
rect 470732 287425 470736 287481
rect 470672 287421 470736 287425
rect 470752 287481 470816 287485
rect 470752 287425 470756 287481
rect 470756 287425 470812 287481
rect 470812 287425 470816 287481
rect 470752 287421 470816 287425
rect 470272 287401 470336 287405
rect 470272 287345 470276 287401
rect 470276 287345 470332 287401
rect 470332 287345 470336 287401
rect 470272 287341 470336 287345
rect 470352 287401 470416 287405
rect 470352 287345 470356 287401
rect 470356 287345 470412 287401
rect 470412 287345 470416 287401
rect 470352 287341 470416 287345
rect 470432 287401 470496 287405
rect 470432 287345 470436 287401
rect 470436 287345 470492 287401
rect 470492 287345 470496 287401
rect 470432 287341 470496 287345
rect 470512 287401 470576 287405
rect 470512 287345 470516 287401
rect 470516 287345 470572 287401
rect 470572 287345 470576 287401
rect 470512 287341 470576 287345
rect 470592 287401 470656 287405
rect 470592 287345 470596 287401
rect 470596 287345 470652 287401
rect 470652 287345 470656 287401
rect 470592 287341 470656 287345
rect 470672 287401 470736 287405
rect 470672 287345 470676 287401
rect 470676 287345 470732 287401
rect 470732 287345 470736 287401
rect 470672 287341 470736 287345
rect 470752 287401 470816 287405
rect 470752 287345 470756 287401
rect 470756 287345 470812 287401
rect 470812 287345 470816 287401
rect 470752 287341 470816 287345
rect 470272 287321 470336 287325
rect 470272 287265 470276 287321
rect 470276 287265 470332 287321
rect 470332 287265 470336 287321
rect 470272 287261 470336 287265
rect 470352 287321 470416 287325
rect 470352 287265 470356 287321
rect 470356 287265 470412 287321
rect 470412 287265 470416 287321
rect 470352 287261 470416 287265
rect 470432 287321 470496 287325
rect 470432 287265 470436 287321
rect 470436 287265 470492 287321
rect 470492 287265 470496 287321
rect 470432 287261 470496 287265
rect 470512 287321 470576 287325
rect 470512 287265 470516 287321
rect 470516 287265 470572 287321
rect 470572 287265 470576 287321
rect 470512 287261 470576 287265
rect 470592 287321 470656 287325
rect 470592 287265 470596 287321
rect 470596 287265 470652 287321
rect 470652 287265 470656 287321
rect 470592 287261 470656 287265
rect 470672 287321 470736 287325
rect 470672 287265 470676 287321
rect 470676 287265 470732 287321
rect 470732 287265 470736 287321
rect 470672 287261 470736 287265
rect 470752 287321 470816 287325
rect 470752 287265 470756 287321
rect 470756 287265 470812 287321
rect 470812 287265 470816 287321
rect 470752 287261 470816 287265
rect 470272 287241 470336 287245
rect 470272 287185 470276 287241
rect 470276 287185 470332 287241
rect 470332 287185 470336 287241
rect 470272 287181 470336 287185
rect 470352 287241 470416 287245
rect 470352 287185 470356 287241
rect 470356 287185 470412 287241
rect 470412 287185 470416 287241
rect 470352 287181 470416 287185
rect 470432 287241 470496 287245
rect 470432 287185 470436 287241
rect 470436 287185 470492 287241
rect 470492 287185 470496 287241
rect 470432 287181 470496 287185
rect 470512 287241 470576 287245
rect 470512 287185 470516 287241
rect 470516 287185 470572 287241
rect 470572 287185 470576 287241
rect 470512 287181 470576 287185
rect 470592 287241 470656 287245
rect 470592 287185 470596 287241
rect 470596 287185 470652 287241
rect 470652 287185 470656 287241
rect 470592 287181 470656 287185
rect 470672 287241 470736 287245
rect 470672 287185 470676 287241
rect 470676 287185 470732 287241
rect 470732 287185 470736 287241
rect 470672 287181 470736 287185
rect 470752 287241 470816 287245
rect 470752 287185 470756 287241
rect 470756 287185 470812 287241
rect 470812 287185 470816 287241
rect 470752 287181 470816 287185
rect 478828 286860 478892 286924
rect 488580 286724 488644 286788
rect 476068 286588 476132 286652
rect 469032 286396 469096 286400
rect 469032 286340 469036 286396
rect 469036 286340 469092 286396
rect 469092 286340 469096 286396
rect 469032 286336 469096 286340
rect 469112 286396 469176 286400
rect 469112 286340 469116 286396
rect 469116 286340 469172 286396
rect 469172 286340 469176 286396
rect 469112 286336 469176 286340
rect 469192 286396 469256 286400
rect 469192 286340 469196 286396
rect 469196 286340 469252 286396
rect 469252 286340 469256 286396
rect 469192 286336 469256 286340
rect 469272 286396 469336 286400
rect 469272 286340 469276 286396
rect 469276 286340 469332 286396
rect 469332 286340 469336 286396
rect 469272 286336 469336 286340
rect 469352 286396 469416 286400
rect 469352 286340 469356 286396
rect 469356 286340 469412 286396
rect 469412 286340 469416 286396
rect 469352 286336 469416 286340
rect 469432 286396 469496 286400
rect 469432 286340 469436 286396
rect 469436 286340 469492 286396
rect 469492 286340 469496 286396
rect 469432 286336 469496 286340
rect 469512 286396 469576 286400
rect 469512 286340 469516 286396
rect 469516 286340 469572 286396
rect 469572 286340 469576 286396
rect 469512 286336 469576 286340
rect 469032 286316 469096 286320
rect 469032 286260 469036 286316
rect 469036 286260 469092 286316
rect 469092 286260 469096 286316
rect 469032 286256 469096 286260
rect 469112 286316 469176 286320
rect 469112 286260 469116 286316
rect 469116 286260 469172 286316
rect 469172 286260 469176 286316
rect 469112 286256 469176 286260
rect 469192 286316 469256 286320
rect 469192 286260 469196 286316
rect 469196 286260 469252 286316
rect 469252 286260 469256 286316
rect 469192 286256 469256 286260
rect 469272 286316 469336 286320
rect 469272 286260 469276 286316
rect 469276 286260 469332 286316
rect 469332 286260 469336 286316
rect 469272 286256 469336 286260
rect 469352 286316 469416 286320
rect 469352 286260 469356 286316
rect 469356 286260 469412 286316
rect 469412 286260 469416 286316
rect 469352 286256 469416 286260
rect 469432 286316 469496 286320
rect 469432 286260 469436 286316
rect 469436 286260 469492 286316
rect 469492 286260 469496 286316
rect 469432 286256 469496 286260
rect 469512 286316 469576 286320
rect 469512 286260 469516 286316
rect 469516 286260 469572 286316
rect 469572 286260 469576 286316
rect 469512 286256 469576 286260
rect 469032 286236 469096 286240
rect 469032 286180 469036 286236
rect 469036 286180 469092 286236
rect 469092 286180 469096 286236
rect 469032 286176 469096 286180
rect 469112 286236 469176 286240
rect 469112 286180 469116 286236
rect 469116 286180 469172 286236
rect 469172 286180 469176 286236
rect 469112 286176 469176 286180
rect 469192 286236 469256 286240
rect 469192 286180 469196 286236
rect 469196 286180 469252 286236
rect 469252 286180 469256 286236
rect 469192 286176 469256 286180
rect 469272 286236 469336 286240
rect 469272 286180 469276 286236
rect 469276 286180 469332 286236
rect 469332 286180 469336 286236
rect 469272 286176 469336 286180
rect 469352 286236 469416 286240
rect 469352 286180 469356 286236
rect 469356 286180 469412 286236
rect 469412 286180 469416 286236
rect 469352 286176 469416 286180
rect 469432 286236 469496 286240
rect 469432 286180 469436 286236
rect 469436 286180 469492 286236
rect 469492 286180 469496 286236
rect 469432 286176 469496 286180
rect 469512 286236 469576 286240
rect 469512 286180 469516 286236
rect 469516 286180 469572 286236
rect 469572 286180 469576 286236
rect 469512 286176 469576 286180
rect 469032 286156 469096 286160
rect 469032 286100 469036 286156
rect 469036 286100 469092 286156
rect 469092 286100 469096 286156
rect 469032 286096 469096 286100
rect 469112 286156 469176 286160
rect 469112 286100 469116 286156
rect 469116 286100 469172 286156
rect 469172 286100 469176 286156
rect 469112 286096 469176 286100
rect 469192 286156 469256 286160
rect 469192 286100 469196 286156
rect 469196 286100 469252 286156
rect 469252 286100 469256 286156
rect 469192 286096 469256 286100
rect 469272 286156 469336 286160
rect 469272 286100 469276 286156
rect 469276 286100 469332 286156
rect 469332 286100 469336 286156
rect 469272 286096 469336 286100
rect 469352 286156 469416 286160
rect 469352 286100 469356 286156
rect 469356 286100 469412 286156
rect 469412 286100 469416 286156
rect 469352 286096 469416 286100
rect 469432 286156 469496 286160
rect 469432 286100 469436 286156
rect 469436 286100 469492 286156
rect 469492 286100 469496 286156
rect 469432 286096 469496 286100
rect 469512 286156 469576 286160
rect 469512 286100 469516 286156
rect 469516 286100 469572 286156
rect 469572 286100 469576 286156
rect 469512 286096 469576 286100
rect 482324 285832 482388 285836
rect 482324 285776 482345 285832
rect 482345 285776 482388 285832
rect 482324 285772 482388 285776
rect 482876 285772 482940 285836
rect 485820 285832 485884 285836
rect 485820 285776 485870 285832
rect 485870 285776 485884 285832
rect 485820 285772 485884 285776
rect 470272 285308 470336 285312
rect 470272 285252 470276 285308
rect 470276 285252 470332 285308
rect 470332 285252 470336 285308
rect 470272 285248 470336 285252
rect 470352 285308 470416 285312
rect 470352 285252 470356 285308
rect 470356 285252 470412 285308
rect 470412 285252 470416 285308
rect 470352 285248 470416 285252
rect 470432 285308 470496 285312
rect 470432 285252 470436 285308
rect 470436 285252 470492 285308
rect 470492 285252 470496 285308
rect 470432 285248 470496 285252
rect 470512 285308 470576 285312
rect 470512 285252 470516 285308
rect 470516 285252 470572 285308
rect 470572 285252 470576 285308
rect 470512 285248 470576 285252
rect 470592 285308 470656 285312
rect 470592 285252 470596 285308
rect 470596 285252 470652 285308
rect 470652 285252 470656 285308
rect 470592 285248 470656 285252
rect 470672 285308 470736 285312
rect 470672 285252 470676 285308
rect 470676 285252 470732 285308
rect 470732 285252 470736 285308
rect 470672 285248 470736 285252
rect 470752 285308 470816 285312
rect 470752 285252 470756 285308
rect 470756 285252 470812 285308
rect 470812 285252 470816 285308
rect 470752 285248 470816 285252
rect 470272 285228 470336 285232
rect 470272 285172 470276 285228
rect 470276 285172 470332 285228
rect 470332 285172 470336 285228
rect 470272 285168 470336 285172
rect 470352 285228 470416 285232
rect 470352 285172 470356 285228
rect 470356 285172 470412 285228
rect 470412 285172 470416 285228
rect 470352 285168 470416 285172
rect 470432 285228 470496 285232
rect 470432 285172 470436 285228
rect 470436 285172 470492 285228
rect 470492 285172 470496 285228
rect 470432 285168 470496 285172
rect 470512 285228 470576 285232
rect 470512 285172 470516 285228
rect 470516 285172 470572 285228
rect 470572 285172 470576 285228
rect 470512 285168 470576 285172
rect 470592 285228 470656 285232
rect 470592 285172 470596 285228
rect 470596 285172 470652 285228
rect 470652 285172 470656 285228
rect 470592 285168 470656 285172
rect 470672 285228 470736 285232
rect 470672 285172 470676 285228
rect 470676 285172 470732 285228
rect 470732 285172 470736 285228
rect 470672 285168 470736 285172
rect 470752 285228 470816 285232
rect 470752 285172 470756 285228
rect 470756 285172 470812 285228
rect 470812 285172 470816 285228
rect 470752 285168 470816 285172
rect 470272 285148 470336 285152
rect 470272 285092 470276 285148
rect 470276 285092 470332 285148
rect 470332 285092 470336 285148
rect 470272 285088 470336 285092
rect 470352 285148 470416 285152
rect 470352 285092 470356 285148
rect 470356 285092 470412 285148
rect 470412 285092 470416 285148
rect 470352 285088 470416 285092
rect 470432 285148 470496 285152
rect 470432 285092 470436 285148
rect 470436 285092 470492 285148
rect 470492 285092 470496 285148
rect 470432 285088 470496 285092
rect 470512 285148 470576 285152
rect 470512 285092 470516 285148
rect 470516 285092 470572 285148
rect 470572 285092 470576 285148
rect 470512 285088 470576 285092
rect 470592 285148 470656 285152
rect 470592 285092 470596 285148
rect 470596 285092 470652 285148
rect 470652 285092 470656 285148
rect 470592 285088 470656 285092
rect 470672 285148 470736 285152
rect 470672 285092 470676 285148
rect 470676 285092 470732 285148
rect 470732 285092 470736 285148
rect 470672 285088 470736 285092
rect 470752 285148 470816 285152
rect 470752 285092 470756 285148
rect 470756 285092 470812 285148
rect 470812 285092 470816 285148
rect 470752 285088 470816 285092
rect 470272 285068 470336 285072
rect 470272 285012 470276 285068
rect 470276 285012 470332 285068
rect 470332 285012 470336 285068
rect 470272 285008 470336 285012
rect 470352 285068 470416 285072
rect 470352 285012 470356 285068
rect 470356 285012 470412 285068
rect 470412 285012 470416 285068
rect 470352 285008 470416 285012
rect 470432 285068 470496 285072
rect 470432 285012 470436 285068
rect 470436 285012 470492 285068
rect 470492 285012 470496 285068
rect 470432 285008 470496 285012
rect 470512 285068 470576 285072
rect 470512 285012 470516 285068
rect 470516 285012 470572 285068
rect 470572 285012 470576 285068
rect 470512 285008 470576 285012
rect 470592 285068 470656 285072
rect 470592 285012 470596 285068
rect 470596 285012 470652 285068
rect 470652 285012 470656 285068
rect 470592 285008 470656 285012
rect 470672 285068 470736 285072
rect 470672 285012 470676 285068
rect 470676 285012 470732 285068
rect 470732 285012 470736 285068
rect 470672 285008 470736 285012
rect 470752 285068 470816 285072
rect 470752 285012 470756 285068
rect 470756 285012 470812 285068
rect 470812 285012 470816 285068
rect 470752 285008 470816 285012
rect 470272 267481 470336 267485
rect 470272 267425 470276 267481
rect 470276 267425 470332 267481
rect 470332 267425 470336 267481
rect 470272 267421 470336 267425
rect 470352 267481 470416 267485
rect 470352 267425 470356 267481
rect 470356 267425 470412 267481
rect 470412 267425 470416 267481
rect 470352 267421 470416 267425
rect 470432 267481 470496 267485
rect 470432 267425 470436 267481
rect 470436 267425 470492 267481
rect 470492 267425 470496 267481
rect 470432 267421 470496 267425
rect 470512 267481 470576 267485
rect 470512 267425 470516 267481
rect 470516 267425 470572 267481
rect 470572 267425 470576 267481
rect 470512 267421 470576 267425
rect 470592 267481 470656 267485
rect 470592 267425 470596 267481
rect 470596 267425 470652 267481
rect 470652 267425 470656 267481
rect 470592 267421 470656 267425
rect 470672 267481 470736 267485
rect 470672 267425 470676 267481
rect 470676 267425 470732 267481
rect 470732 267425 470736 267481
rect 470672 267421 470736 267425
rect 470752 267481 470816 267485
rect 470752 267425 470756 267481
rect 470756 267425 470812 267481
rect 470812 267425 470816 267481
rect 470752 267421 470816 267425
rect 470272 267401 470336 267405
rect 470272 267345 470276 267401
rect 470276 267345 470332 267401
rect 470332 267345 470336 267401
rect 470272 267341 470336 267345
rect 470352 267401 470416 267405
rect 470352 267345 470356 267401
rect 470356 267345 470412 267401
rect 470412 267345 470416 267401
rect 470352 267341 470416 267345
rect 470432 267401 470496 267405
rect 470432 267345 470436 267401
rect 470436 267345 470492 267401
rect 470492 267345 470496 267401
rect 470432 267341 470496 267345
rect 470512 267401 470576 267405
rect 470512 267345 470516 267401
rect 470516 267345 470572 267401
rect 470572 267345 470576 267401
rect 470512 267341 470576 267345
rect 470592 267401 470656 267405
rect 470592 267345 470596 267401
rect 470596 267345 470652 267401
rect 470652 267345 470656 267401
rect 470592 267341 470656 267345
rect 470672 267401 470736 267405
rect 470672 267345 470676 267401
rect 470676 267345 470732 267401
rect 470732 267345 470736 267401
rect 470672 267341 470736 267345
rect 470752 267401 470816 267405
rect 470752 267345 470756 267401
rect 470756 267345 470812 267401
rect 470812 267345 470816 267401
rect 470752 267341 470816 267345
rect 470272 267321 470336 267325
rect 470272 267265 470276 267321
rect 470276 267265 470332 267321
rect 470332 267265 470336 267321
rect 470272 267261 470336 267265
rect 470352 267321 470416 267325
rect 470352 267265 470356 267321
rect 470356 267265 470412 267321
rect 470412 267265 470416 267321
rect 470352 267261 470416 267265
rect 470432 267321 470496 267325
rect 470432 267265 470436 267321
rect 470436 267265 470492 267321
rect 470492 267265 470496 267321
rect 470432 267261 470496 267265
rect 470512 267321 470576 267325
rect 470512 267265 470516 267321
rect 470516 267265 470572 267321
rect 470572 267265 470576 267321
rect 470512 267261 470576 267265
rect 470592 267321 470656 267325
rect 470592 267265 470596 267321
rect 470596 267265 470652 267321
rect 470652 267265 470656 267321
rect 470592 267261 470656 267265
rect 470672 267321 470736 267325
rect 470672 267265 470676 267321
rect 470676 267265 470732 267321
rect 470732 267265 470736 267321
rect 470672 267261 470736 267265
rect 470752 267321 470816 267325
rect 470752 267265 470756 267321
rect 470756 267265 470812 267321
rect 470812 267265 470816 267321
rect 470752 267261 470816 267265
rect 470272 267241 470336 267245
rect 470272 267185 470276 267241
rect 470276 267185 470332 267241
rect 470332 267185 470336 267241
rect 470272 267181 470336 267185
rect 470352 267241 470416 267245
rect 470352 267185 470356 267241
rect 470356 267185 470412 267241
rect 470412 267185 470416 267241
rect 470352 267181 470416 267185
rect 470432 267241 470496 267245
rect 470432 267185 470436 267241
rect 470436 267185 470492 267241
rect 470492 267185 470496 267241
rect 470432 267181 470496 267185
rect 470512 267241 470576 267245
rect 470512 267185 470516 267241
rect 470516 267185 470572 267241
rect 470572 267185 470576 267241
rect 470512 267181 470576 267185
rect 470592 267241 470656 267245
rect 470592 267185 470596 267241
rect 470596 267185 470652 267241
rect 470652 267185 470656 267241
rect 470592 267181 470656 267185
rect 470672 267241 470736 267245
rect 470672 267185 470676 267241
rect 470676 267185 470732 267241
rect 470732 267185 470736 267241
rect 470672 267181 470736 267185
rect 470752 267241 470816 267245
rect 470752 267185 470756 267241
rect 470756 267185 470812 267241
rect 470812 267185 470816 267241
rect 470752 267181 470816 267185
rect 469032 266395 469096 266399
rect 469032 266339 469036 266395
rect 469036 266339 469092 266395
rect 469092 266339 469096 266395
rect 469032 266335 469096 266339
rect 469112 266395 469176 266399
rect 469112 266339 469116 266395
rect 469116 266339 469172 266395
rect 469172 266339 469176 266395
rect 469112 266335 469176 266339
rect 469192 266395 469256 266399
rect 469192 266339 469196 266395
rect 469196 266339 469252 266395
rect 469252 266339 469256 266395
rect 469192 266335 469256 266339
rect 469272 266395 469336 266399
rect 469272 266339 469276 266395
rect 469276 266339 469332 266395
rect 469332 266339 469336 266395
rect 469272 266335 469336 266339
rect 469352 266395 469416 266399
rect 469352 266339 469356 266395
rect 469356 266339 469412 266395
rect 469412 266339 469416 266395
rect 469352 266335 469416 266339
rect 469432 266395 469496 266399
rect 469432 266339 469436 266395
rect 469436 266339 469492 266395
rect 469492 266339 469496 266395
rect 469432 266335 469496 266339
rect 469512 266395 469576 266399
rect 469512 266339 469516 266395
rect 469516 266339 469572 266395
rect 469572 266339 469576 266395
rect 469512 266335 469576 266339
rect 469032 266315 469096 266319
rect 469032 266259 469036 266315
rect 469036 266259 469092 266315
rect 469092 266259 469096 266315
rect 469032 266255 469096 266259
rect 469112 266315 469176 266319
rect 469112 266259 469116 266315
rect 469116 266259 469172 266315
rect 469172 266259 469176 266315
rect 469112 266255 469176 266259
rect 469192 266315 469256 266319
rect 469192 266259 469196 266315
rect 469196 266259 469252 266315
rect 469252 266259 469256 266315
rect 469192 266255 469256 266259
rect 469272 266315 469336 266319
rect 469272 266259 469276 266315
rect 469276 266259 469332 266315
rect 469332 266259 469336 266315
rect 469272 266255 469336 266259
rect 469352 266315 469416 266319
rect 469352 266259 469356 266315
rect 469356 266259 469412 266315
rect 469412 266259 469416 266315
rect 469352 266255 469416 266259
rect 469432 266315 469496 266319
rect 469432 266259 469436 266315
rect 469436 266259 469492 266315
rect 469492 266259 469496 266315
rect 469432 266255 469496 266259
rect 469512 266315 469576 266319
rect 469512 266259 469516 266315
rect 469516 266259 469572 266315
rect 469572 266259 469576 266315
rect 469512 266255 469576 266259
rect 469032 266235 469096 266239
rect 469032 266179 469036 266235
rect 469036 266179 469092 266235
rect 469092 266179 469096 266235
rect 469032 266175 469096 266179
rect 469112 266235 469176 266239
rect 469112 266179 469116 266235
rect 469116 266179 469172 266235
rect 469172 266179 469176 266235
rect 469112 266175 469176 266179
rect 469192 266235 469256 266239
rect 469192 266179 469196 266235
rect 469196 266179 469252 266235
rect 469252 266179 469256 266235
rect 469192 266175 469256 266179
rect 469272 266235 469336 266239
rect 469272 266179 469276 266235
rect 469276 266179 469332 266235
rect 469332 266179 469336 266235
rect 469272 266175 469336 266179
rect 469352 266235 469416 266239
rect 469352 266179 469356 266235
rect 469356 266179 469412 266235
rect 469412 266179 469416 266235
rect 469352 266175 469416 266179
rect 469432 266235 469496 266239
rect 469432 266179 469436 266235
rect 469436 266179 469492 266235
rect 469492 266179 469496 266235
rect 469432 266175 469496 266179
rect 469512 266235 469576 266239
rect 469512 266179 469516 266235
rect 469516 266179 469572 266235
rect 469572 266179 469576 266235
rect 469512 266175 469576 266179
rect 469032 266155 469096 266159
rect 469032 266099 469036 266155
rect 469036 266099 469092 266155
rect 469092 266099 469096 266155
rect 469032 266095 469096 266099
rect 469112 266155 469176 266159
rect 469112 266099 469116 266155
rect 469116 266099 469172 266155
rect 469172 266099 469176 266155
rect 469112 266095 469176 266099
rect 469192 266155 469256 266159
rect 469192 266099 469196 266155
rect 469196 266099 469252 266155
rect 469252 266099 469256 266155
rect 469192 266095 469256 266099
rect 469272 266155 469336 266159
rect 469272 266099 469276 266155
rect 469276 266099 469332 266155
rect 469332 266099 469336 266155
rect 469272 266095 469336 266099
rect 469352 266155 469416 266159
rect 469352 266099 469356 266155
rect 469356 266099 469412 266155
rect 469412 266099 469416 266155
rect 469352 266095 469416 266099
rect 469432 266155 469496 266159
rect 469432 266099 469436 266155
rect 469436 266099 469492 266155
rect 469492 266099 469496 266155
rect 469432 266095 469496 266099
rect 469512 266155 469576 266159
rect 469512 266099 469516 266155
rect 469516 266099 469572 266155
rect 469572 266099 469576 266155
rect 469512 266095 469576 266099
rect 479012 265976 479076 265980
rect 479012 265920 479062 265976
rect 479062 265920 479076 265976
rect 479012 265916 479076 265920
rect 489132 265508 489196 265572
rect 470272 265308 470336 265312
rect 470272 265252 470276 265308
rect 470276 265252 470332 265308
rect 470332 265252 470336 265308
rect 470272 265248 470336 265252
rect 470352 265308 470416 265312
rect 470352 265252 470356 265308
rect 470356 265252 470412 265308
rect 470412 265252 470416 265308
rect 470352 265248 470416 265252
rect 470432 265308 470496 265312
rect 470432 265252 470436 265308
rect 470436 265252 470492 265308
rect 470492 265252 470496 265308
rect 470432 265248 470496 265252
rect 470512 265308 470576 265312
rect 470512 265252 470516 265308
rect 470516 265252 470572 265308
rect 470572 265252 470576 265308
rect 470512 265248 470576 265252
rect 470592 265308 470656 265312
rect 470592 265252 470596 265308
rect 470596 265252 470652 265308
rect 470652 265252 470656 265308
rect 470592 265248 470656 265252
rect 470672 265308 470736 265312
rect 470672 265252 470676 265308
rect 470676 265252 470732 265308
rect 470732 265252 470736 265308
rect 470672 265248 470736 265252
rect 470752 265308 470816 265312
rect 470752 265252 470756 265308
rect 470756 265252 470812 265308
rect 470812 265252 470816 265308
rect 470752 265248 470816 265252
rect 470272 265228 470336 265232
rect 470272 265172 470276 265228
rect 470276 265172 470332 265228
rect 470332 265172 470336 265228
rect 470272 265168 470336 265172
rect 470352 265228 470416 265232
rect 470352 265172 470356 265228
rect 470356 265172 470412 265228
rect 470412 265172 470416 265228
rect 470352 265168 470416 265172
rect 470432 265228 470496 265232
rect 470432 265172 470436 265228
rect 470436 265172 470492 265228
rect 470492 265172 470496 265228
rect 470432 265168 470496 265172
rect 470512 265228 470576 265232
rect 470512 265172 470516 265228
rect 470516 265172 470572 265228
rect 470572 265172 470576 265228
rect 470512 265168 470576 265172
rect 470592 265228 470656 265232
rect 470592 265172 470596 265228
rect 470596 265172 470652 265228
rect 470652 265172 470656 265228
rect 470592 265168 470656 265172
rect 470672 265228 470736 265232
rect 470672 265172 470676 265228
rect 470676 265172 470732 265228
rect 470732 265172 470736 265228
rect 470672 265168 470736 265172
rect 470752 265228 470816 265232
rect 470752 265172 470756 265228
rect 470756 265172 470812 265228
rect 470812 265172 470816 265228
rect 470752 265168 470816 265172
rect 470272 265148 470336 265152
rect 470272 265092 470276 265148
rect 470276 265092 470332 265148
rect 470332 265092 470336 265148
rect 470272 265088 470336 265092
rect 470352 265148 470416 265152
rect 470352 265092 470356 265148
rect 470356 265092 470412 265148
rect 470412 265092 470416 265148
rect 470352 265088 470416 265092
rect 470432 265148 470496 265152
rect 470432 265092 470436 265148
rect 470436 265092 470492 265148
rect 470492 265092 470496 265148
rect 470432 265088 470496 265092
rect 470512 265148 470576 265152
rect 470512 265092 470516 265148
rect 470516 265092 470572 265148
rect 470572 265092 470576 265148
rect 470512 265088 470576 265092
rect 470592 265148 470656 265152
rect 470592 265092 470596 265148
rect 470596 265092 470652 265148
rect 470652 265092 470656 265148
rect 470592 265088 470656 265092
rect 470672 265148 470736 265152
rect 470672 265092 470676 265148
rect 470676 265092 470732 265148
rect 470732 265092 470736 265148
rect 470672 265088 470736 265092
rect 470752 265148 470816 265152
rect 470752 265092 470756 265148
rect 470756 265092 470812 265148
rect 470812 265092 470816 265148
rect 470752 265088 470816 265092
rect 470272 265068 470336 265072
rect 470272 265012 470276 265068
rect 470276 265012 470332 265068
rect 470332 265012 470336 265068
rect 470272 265008 470336 265012
rect 470352 265068 470416 265072
rect 470352 265012 470356 265068
rect 470356 265012 470412 265068
rect 470412 265012 470416 265068
rect 470352 265008 470416 265012
rect 470432 265068 470496 265072
rect 470432 265012 470436 265068
rect 470436 265012 470492 265068
rect 470492 265012 470496 265068
rect 470432 265008 470496 265012
rect 470512 265068 470576 265072
rect 470512 265012 470516 265068
rect 470516 265012 470572 265068
rect 470572 265012 470576 265068
rect 470512 265008 470576 265012
rect 470592 265068 470656 265072
rect 470592 265012 470596 265068
rect 470596 265012 470652 265068
rect 470652 265012 470656 265068
rect 470592 265008 470656 265012
rect 470672 265068 470736 265072
rect 470672 265012 470676 265068
rect 470676 265012 470732 265068
rect 470732 265012 470736 265068
rect 470672 265008 470736 265012
rect 470752 265068 470816 265072
rect 470752 265012 470756 265068
rect 470756 265012 470812 265068
rect 470812 265012 470816 265068
rect 470752 265008 470816 265012
rect 476436 265024 476500 265028
rect 476436 264968 476486 265024
rect 476486 264968 476500 265024
rect 476436 264964 476500 264968
rect 477356 264964 477420 265028
rect 480116 264964 480180 265028
rect 482876 265024 482940 265028
rect 482876 264968 482890 265024
rect 482890 264968 482940 265024
rect 482876 264964 482940 264968
rect 485820 264964 485884 265028
rect 486372 264964 486436 265028
rect 489132 165820 489196 165884
rect 486372 125972 486436 126036
rect 482876 86124 482940 86188
rect 480116 46276 480180 46340
rect 549300 19756 549364 19820
rect 477356 6564 477420 6628
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 695334 -8106 711002
rect -8726 695098 -8694 695334
rect -8458 695098 -8374 695334
rect -8138 695098 -8106 695334
rect -8726 695014 -8106 695098
rect -8726 694778 -8694 695014
rect -8458 694778 -8374 695014
rect -8138 694778 -8106 695014
rect -8726 659334 -8106 694778
rect -8726 659098 -8694 659334
rect -8458 659098 -8374 659334
rect -8138 659098 -8106 659334
rect -8726 659014 -8106 659098
rect -8726 658778 -8694 659014
rect -8458 658778 -8374 659014
rect -8138 658778 -8106 659014
rect -8726 623334 -8106 658778
rect -8726 623098 -8694 623334
rect -8458 623098 -8374 623334
rect -8138 623098 -8106 623334
rect -8726 623014 -8106 623098
rect -8726 622778 -8694 623014
rect -8458 622778 -8374 623014
rect -8138 622778 -8106 623014
rect -8726 587334 -8106 622778
rect -8726 587098 -8694 587334
rect -8458 587098 -8374 587334
rect -8138 587098 -8106 587334
rect -8726 587014 -8106 587098
rect -8726 586778 -8694 587014
rect -8458 586778 -8374 587014
rect -8138 586778 -8106 587014
rect -8726 551334 -8106 586778
rect -8726 551098 -8694 551334
rect -8458 551098 -8374 551334
rect -8138 551098 -8106 551334
rect -8726 551014 -8106 551098
rect -8726 550778 -8694 551014
rect -8458 550778 -8374 551014
rect -8138 550778 -8106 551014
rect -8726 515334 -8106 550778
rect -8726 515098 -8694 515334
rect -8458 515098 -8374 515334
rect -8138 515098 -8106 515334
rect -8726 515014 -8106 515098
rect -8726 514778 -8694 515014
rect -8458 514778 -8374 515014
rect -8138 514778 -8106 515014
rect -8726 479334 -8106 514778
rect -8726 479098 -8694 479334
rect -8458 479098 -8374 479334
rect -8138 479098 -8106 479334
rect -8726 479014 -8106 479098
rect -8726 478778 -8694 479014
rect -8458 478778 -8374 479014
rect -8138 478778 -8106 479014
rect -8726 443334 -8106 478778
rect -8726 443098 -8694 443334
rect -8458 443098 -8374 443334
rect -8138 443098 -8106 443334
rect -8726 443014 -8106 443098
rect -8726 442778 -8694 443014
rect -8458 442778 -8374 443014
rect -8138 442778 -8106 443014
rect -8726 407334 -8106 442778
rect -8726 407098 -8694 407334
rect -8458 407098 -8374 407334
rect -8138 407098 -8106 407334
rect -8726 407014 -8106 407098
rect -8726 406778 -8694 407014
rect -8458 406778 -8374 407014
rect -8138 406778 -8106 407014
rect -8726 371334 -8106 406778
rect -8726 371098 -8694 371334
rect -8458 371098 -8374 371334
rect -8138 371098 -8106 371334
rect -8726 371014 -8106 371098
rect -8726 370778 -8694 371014
rect -8458 370778 -8374 371014
rect -8138 370778 -8106 371014
rect -8726 335334 -8106 370778
rect -8726 335098 -8694 335334
rect -8458 335098 -8374 335334
rect -8138 335098 -8106 335334
rect -8726 335014 -8106 335098
rect -8726 334778 -8694 335014
rect -8458 334778 -8374 335014
rect -8138 334778 -8106 335014
rect -8726 299334 -8106 334778
rect -8726 299098 -8694 299334
rect -8458 299098 -8374 299334
rect -8138 299098 -8106 299334
rect -8726 299014 -8106 299098
rect -8726 298778 -8694 299014
rect -8458 298778 -8374 299014
rect -8138 298778 -8106 299014
rect -8726 263334 -8106 298778
rect -8726 263098 -8694 263334
rect -8458 263098 -8374 263334
rect -8138 263098 -8106 263334
rect -8726 263014 -8106 263098
rect -8726 262778 -8694 263014
rect -8458 262778 -8374 263014
rect -8138 262778 -8106 263014
rect -8726 227334 -8106 262778
rect -8726 227098 -8694 227334
rect -8458 227098 -8374 227334
rect -8138 227098 -8106 227334
rect -8726 227014 -8106 227098
rect -8726 226778 -8694 227014
rect -8458 226778 -8374 227014
rect -8138 226778 -8106 227014
rect -8726 191334 -8106 226778
rect -8726 191098 -8694 191334
rect -8458 191098 -8374 191334
rect -8138 191098 -8106 191334
rect -8726 191014 -8106 191098
rect -8726 190778 -8694 191014
rect -8458 190778 -8374 191014
rect -8138 190778 -8106 191014
rect -8726 155334 -8106 190778
rect -8726 155098 -8694 155334
rect -8458 155098 -8374 155334
rect -8138 155098 -8106 155334
rect -8726 155014 -8106 155098
rect -8726 154778 -8694 155014
rect -8458 154778 -8374 155014
rect -8138 154778 -8106 155014
rect -8726 119334 -8106 154778
rect -8726 119098 -8694 119334
rect -8458 119098 -8374 119334
rect -8138 119098 -8106 119334
rect -8726 119014 -8106 119098
rect -8726 118778 -8694 119014
rect -8458 118778 -8374 119014
rect -8138 118778 -8106 119014
rect -8726 83334 -8106 118778
rect -8726 83098 -8694 83334
rect -8458 83098 -8374 83334
rect -8138 83098 -8106 83334
rect -8726 83014 -8106 83098
rect -8726 82778 -8694 83014
rect -8458 82778 -8374 83014
rect -8138 82778 -8106 83014
rect -8726 47334 -8106 82778
rect -8726 47098 -8694 47334
rect -8458 47098 -8374 47334
rect -8138 47098 -8106 47334
rect -8726 47014 -8106 47098
rect -8726 46778 -8694 47014
rect -8458 46778 -8374 47014
rect -8138 46778 -8106 47014
rect -8726 11334 -8106 46778
rect -8726 11098 -8694 11334
rect -8458 11098 -8374 11334
rect -8138 11098 -8106 11334
rect -8726 11014 -8106 11098
rect -8726 10778 -8694 11014
rect -8458 10778 -8374 11014
rect -8138 10778 -8106 11014
rect -8726 -7066 -8106 10778
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 694094 -7146 710042
rect -7766 693858 -7734 694094
rect -7498 693858 -7414 694094
rect -7178 693858 -7146 694094
rect -7766 693774 -7146 693858
rect -7766 693538 -7734 693774
rect -7498 693538 -7414 693774
rect -7178 693538 -7146 693774
rect -7766 658094 -7146 693538
rect -7766 657858 -7734 658094
rect -7498 657858 -7414 658094
rect -7178 657858 -7146 658094
rect -7766 657774 -7146 657858
rect -7766 657538 -7734 657774
rect -7498 657538 -7414 657774
rect -7178 657538 -7146 657774
rect -7766 622094 -7146 657538
rect -7766 621858 -7734 622094
rect -7498 621858 -7414 622094
rect -7178 621858 -7146 622094
rect -7766 621774 -7146 621858
rect -7766 621538 -7734 621774
rect -7498 621538 -7414 621774
rect -7178 621538 -7146 621774
rect -7766 586094 -7146 621538
rect -7766 585858 -7734 586094
rect -7498 585858 -7414 586094
rect -7178 585858 -7146 586094
rect -7766 585774 -7146 585858
rect -7766 585538 -7734 585774
rect -7498 585538 -7414 585774
rect -7178 585538 -7146 585774
rect -7766 550094 -7146 585538
rect -7766 549858 -7734 550094
rect -7498 549858 -7414 550094
rect -7178 549858 -7146 550094
rect -7766 549774 -7146 549858
rect -7766 549538 -7734 549774
rect -7498 549538 -7414 549774
rect -7178 549538 -7146 549774
rect -7766 514094 -7146 549538
rect -7766 513858 -7734 514094
rect -7498 513858 -7414 514094
rect -7178 513858 -7146 514094
rect -7766 513774 -7146 513858
rect -7766 513538 -7734 513774
rect -7498 513538 -7414 513774
rect -7178 513538 -7146 513774
rect -7766 478094 -7146 513538
rect -7766 477858 -7734 478094
rect -7498 477858 -7414 478094
rect -7178 477858 -7146 478094
rect -7766 477774 -7146 477858
rect -7766 477538 -7734 477774
rect -7498 477538 -7414 477774
rect -7178 477538 -7146 477774
rect -7766 442094 -7146 477538
rect -7766 441858 -7734 442094
rect -7498 441858 -7414 442094
rect -7178 441858 -7146 442094
rect -7766 441774 -7146 441858
rect -7766 441538 -7734 441774
rect -7498 441538 -7414 441774
rect -7178 441538 -7146 441774
rect -7766 406094 -7146 441538
rect -7766 405858 -7734 406094
rect -7498 405858 -7414 406094
rect -7178 405858 -7146 406094
rect -7766 405774 -7146 405858
rect -7766 405538 -7734 405774
rect -7498 405538 -7414 405774
rect -7178 405538 -7146 405774
rect -7766 370094 -7146 405538
rect -7766 369858 -7734 370094
rect -7498 369858 -7414 370094
rect -7178 369858 -7146 370094
rect -7766 369774 -7146 369858
rect -7766 369538 -7734 369774
rect -7498 369538 -7414 369774
rect -7178 369538 -7146 369774
rect -7766 334094 -7146 369538
rect -7766 333858 -7734 334094
rect -7498 333858 -7414 334094
rect -7178 333858 -7146 334094
rect -7766 333774 -7146 333858
rect -7766 333538 -7734 333774
rect -7498 333538 -7414 333774
rect -7178 333538 -7146 333774
rect -7766 298094 -7146 333538
rect -7766 297858 -7734 298094
rect -7498 297858 -7414 298094
rect -7178 297858 -7146 298094
rect -7766 297774 -7146 297858
rect -7766 297538 -7734 297774
rect -7498 297538 -7414 297774
rect -7178 297538 -7146 297774
rect -7766 262094 -7146 297538
rect -7766 261858 -7734 262094
rect -7498 261858 -7414 262094
rect -7178 261858 -7146 262094
rect -7766 261774 -7146 261858
rect -7766 261538 -7734 261774
rect -7498 261538 -7414 261774
rect -7178 261538 -7146 261774
rect -7766 226094 -7146 261538
rect -7766 225858 -7734 226094
rect -7498 225858 -7414 226094
rect -7178 225858 -7146 226094
rect -7766 225774 -7146 225858
rect -7766 225538 -7734 225774
rect -7498 225538 -7414 225774
rect -7178 225538 -7146 225774
rect -7766 190094 -7146 225538
rect -7766 189858 -7734 190094
rect -7498 189858 -7414 190094
rect -7178 189858 -7146 190094
rect -7766 189774 -7146 189858
rect -7766 189538 -7734 189774
rect -7498 189538 -7414 189774
rect -7178 189538 -7146 189774
rect -7766 154094 -7146 189538
rect -7766 153858 -7734 154094
rect -7498 153858 -7414 154094
rect -7178 153858 -7146 154094
rect -7766 153774 -7146 153858
rect -7766 153538 -7734 153774
rect -7498 153538 -7414 153774
rect -7178 153538 -7146 153774
rect -7766 118094 -7146 153538
rect -7766 117858 -7734 118094
rect -7498 117858 -7414 118094
rect -7178 117858 -7146 118094
rect -7766 117774 -7146 117858
rect -7766 117538 -7734 117774
rect -7498 117538 -7414 117774
rect -7178 117538 -7146 117774
rect -7766 82094 -7146 117538
rect -7766 81858 -7734 82094
rect -7498 81858 -7414 82094
rect -7178 81858 -7146 82094
rect -7766 81774 -7146 81858
rect -7766 81538 -7734 81774
rect -7498 81538 -7414 81774
rect -7178 81538 -7146 81774
rect -7766 46094 -7146 81538
rect -7766 45858 -7734 46094
rect -7498 45858 -7414 46094
rect -7178 45858 -7146 46094
rect -7766 45774 -7146 45858
rect -7766 45538 -7734 45774
rect -7498 45538 -7414 45774
rect -7178 45538 -7146 45774
rect -7766 10094 -7146 45538
rect -7766 9858 -7734 10094
rect -7498 9858 -7414 10094
rect -7178 9858 -7146 10094
rect -7766 9774 -7146 9858
rect -7766 9538 -7734 9774
rect -7498 9538 -7414 9774
rect -7178 9538 -7146 9774
rect -7766 -6106 -7146 9538
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 692854 -6186 709082
rect -6806 692618 -6774 692854
rect -6538 692618 -6454 692854
rect -6218 692618 -6186 692854
rect -6806 692534 -6186 692618
rect -6806 692298 -6774 692534
rect -6538 692298 -6454 692534
rect -6218 692298 -6186 692534
rect -6806 656854 -6186 692298
rect -6806 656618 -6774 656854
rect -6538 656618 -6454 656854
rect -6218 656618 -6186 656854
rect -6806 656534 -6186 656618
rect -6806 656298 -6774 656534
rect -6538 656298 -6454 656534
rect -6218 656298 -6186 656534
rect -6806 620854 -6186 656298
rect -6806 620618 -6774 620854
rect -6538 620618 -6454 620854
rect -6218 620618 -6186 620854
rect -6806 620534 -6186 620618
rect -6806 620298 -6774 620534
rect -6538 620298 -6454 620534
rect -6218 620298 -6186 620534
rect -6806 584854 -6186 620298
rect -6806 584618 -6774 584854
rect -6538 584618 -6454 584854
rect -6218 584618 -6186 584854
rect -6806 584534 -6186 584618
rect -6806 584298 -6774 584534
rect -6538 584298 -6454 584534
rect -6218 584298 -6186 584534
rect -6806 548854 -6186 584298
rect -6806 548618 -6774 548854
rect -6538 548618 -6454 548854
rect -6218 548618 -6186 548854
rect -6806 548534 -6186 548618
rect -6806 548298 -6774 548534
rect -6538 548298 -6454 548534
rect -6218 548298 -6186 548534
rect -6806 512854 -6186 548298
rect -6806 512618 -6774 512854
rect -6538 512618 -6454 512854
rect -6218 512618 -6186 512854
rect -6806 512534 -6186 512618
rect -6806 512298 -6774 512534
rect -6538 512298 -6454 512534
rect -6218 512298 -6186 512534
rect -6806 476854 -6186 512298
rect -6806 476618 -6774 476854
rect -6538 476618 -6454 476854
rect -6218 476618 -6186 476854
rect -6806 476534 -6186 476618
rect -6806 476298 -6774 476534
rect -6538 476298 -6454 476534
rect -6218 476298 -6186 476534
rect -6806 440854 -6186 476298
rect -6806 440618 -6774 440854
rect -6538 440618 -6454 440854
rect -6218 440618 -6186 440854
rect -6806 440534 -6186 440618
rect -6806 440298 -6774 440534
rect -6538 440298 -6454 440534
rect -6218 440298 -6186 440534
rect -6806 404854 -6186 440298
rect -6806 404618 -6774 404854
rect -6538 404618 -6454 404854
rect -6218 404618 -6186 404854
rect -6806 404534 -6186 404618
rect -6806 404298 -6774 404534
rect -6538 404298 -6454 404534
rect -6218 404298 -6186 404534
rect -6806 368854 -6186 404298
rect -6806 368618 -6774 368854
rect -6538 368618 -6454 368854
rect -6218 368618 -6186 368854
rect -6806 368534 -6186 368618
rect -6806 368298 -6774 368534
rect -6538 368298 -6454 368534
rect -6218 368298 -6186 368534
rect -6806 332854 -6186 368298
rect -6806 332618 -6774 332854
rect -6538 332618 -6454 332854
rect -6218 332618 -6186 332854
rect -6806 332534 -6186 332618
rect -6806 332298 -6774 332534
rect -6538 332298 -6454 332534
rect -6218 332298 -6186 332534
rect -6806 296854 -6186 332298
rect -6806 296618 -6774 296854
rect -6538 296618 -6454 296854
rect -6218 296618 -6186 296854
rect -6806 296534 -6186 296618
rect -6806 296298 -6774 296534
rect -6538 296298 -6454 296534
rect -6218 296298 -6186 296534
rect -6806 260854 -6186 296298
rect -6806 260618 -6774 260854
rect -6538 260618 -6454 260854
rect -6218 260618 -6186 260854
rect -6806 260534 -6186 260618
rect -6806 260298 -6774 260534
rect -6538 260298 -6454 260534
rect -6218 260298 -6186 260534
rect -6806 224854 -6186 260298
rect -6806 224618 -6774 224854
rect -6538 224618 -6454 224854
rect -6218 224618 -6186 224854
rect -6806 224534 -6186 224618
rect -6806 224298 -6774 224534
rect -6538 224298 -6454 224534
rect -6218 224298 -6186 224534
rect -6806 188854 -6186 224298
rect -6806 188618 -6774 188854
rect -6538 188618 -6454 188854
rect -6218 188618 -6186 188854
rect -6806 188534 -6186 188618
rect -6806 188298 -6774 188534
rect -6538 188298 -6454 188534
rect -6218 188298 -6186 188534
rect -6806 152854 -6186 188298
rect -6806 152618 -6774 152854
rect -6538 152618 -6454 152854
rect -6218 152618 -6186 152854
rect -6806 152534 -6186 152618
rect -6806 152298 -6774 152534
rect -6538 152298 -6454 152534
rect -6218 152298 -6186 152534
rect -6806 116854 -6186 152298
rect -6806 116618 -6774 116854
rect -6538 116618 -6454 116854
rect -6218 116618 -6186 116854
rect -6806 116534 -6186 116618
rect -6806 116298 -6774 116534
rect -6538 116298 -6454 116534
rect -6218 116298 -6186 116534
rect -6806 80854 -6186 116298
rect -6806 80618 -6774 80854
rect -6538 80618 -6454 80854
rect -6218 80618 -6186 80854
rect -6806 80534 -6186 80618
rect -6806 80298 -6774 80534
rect -6538 80298 -6454 80534
rect -6218 80298 -6186 80534
rect -6806 44854 -6186 80298
rect -6806 44618 -6774 44854
rect -6538 44618 -6454 44854
rect -6218 44618 -6186 44854
rect -6806 44534 -6186 44618
rect -6806 44298 -6774 44534
rect -6538 44298 -6454 44534
rect -6218 44298 -6186 44534
rect -6806 8854 -6186 44298
rect -6806 8618 -6774 8854
rect -6538 8618 -6454 8854
rect -6218 8618 -6186 8854
rect -6806 8534 -6186 8618
rect -6806 8298 -6774 8534
rect -6538 8298 -6454 8534
rect -6218 8298 -6186 8534
rect -6806 -5146 -6186 8298
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 691614 -5226 708122
rect -5846 691378 -5814 691614
rect -5578 691378 -5494 691614
rect -5258 691378 -5226 691614
rect -5846 691294 -5226 691378
rect -5846 691058 -5814 691294
rect -5578 691058 -5494 691294
rect -5258 691058 -5226 691294
rect -5846 655614 -5226 691058
rect -5846 655378 -5814 655614
rect -5578 655378 -5494 655614
rect -5258 655378 -5226 655614
rect -5846 655294 -5226 655378
rect -5846 655058 -5814 655294
rect -5578 655058 -5494 655294
rect -5258 655058 -5226 655294
rect -5846 619614 -5226 655058
rect -5846 619378 -5814 619614
rect -5578 619378 -5494 619614
rect -5258 619378 -5226 619614
rect -5846 619294 -5226 619378
rect -5846 619058 -5814 619294
rect -5578 619058 -5494 619294
rect -5258 619058 -5226 619294
rect -5846 583614 -5226 619058
rect -5846 583378 -5814 583614
rect -5578 583378 -5494 583614
rect -5258 583378 -5226 583614
rect -5846 583294 -5226 583378
rect -5846 583058 -5814 583294
rect -5578 583058 -5494 583294
rect -5258 583058 -5226 583294
rect -5846 547614 -5226 583058
rect -5846 547378 -5814 547614
rect -5578 547378 -5494 547614
rect -5258 547378 -5226 547614
rect -5846 547294 -5226 547378
rect -5846 547058 -5814 547294
rect -5578 547058 -5494 547294
rect -5258 547058 -5226 547294
rect -5846 511614 -5226 547058
rect -5846 511378 -5814 511614
rect -5578 511378 -5494 511614
rect -5258 511378 -5226 511614
rect -5846 511294 -5226 511378
rect -5846 511058 -5814 511294
rect -5578 511058 -5494 511294
rect -5258 511058 -5226 511294
rect -5846 475614 -5226 511058
rect -5846 475378 -5814 475614
rect -5578 475378 -5494 475614
rect -5258 475378 -5226 475614
rect -5846 475294 -5226 475378
rect -5846 475058 -5814 475294
rect -5578 475058 -5494 475294
rect -5258 475058 -5226 475294
rect -5846 439614 -5226 475058
rect -5846 439378 -5814 439614
rect -5578 439378 -5494 439614
rect -5258 439378 -5226 439614
rect -5846 439294 -5226 439378
rect -5846 439058 -5814 439294
rect -5578 439058 -5494 439294
rect -5258 439058 -5226 439294
rect -5846 403614 -5226 439058
rect -5846 403378 -5814 403614
rect -5578 403378 -5494 403614
rect -5258 403378 -5226 403614
rect -5846 403294 -5226 403378
rect -5846 403058 -5814 403294
rect -5578 403058 -5494 403294
rect -5258 403058 -5226 403294
rect -5846 367614 -5226 403058
rect -5846 367378 -5814 367614
rect -5578 367378 -5494 367614
rect -5258 367378 -5226 367614
rect -5846 367294 -5226 367378
rect -5846 367058 -5814 367294
rect -5578 367058 -5494 367294
rect -5258 367058 -5226 367294
rect -5846 331614 -5226 367058
rect -5846 331378 -5814 331614
rect -5578 331378 -5494 331614
rect -5258 331378 -5226 331614
rect -5846 331294 -5226 331378
rect -5846 331058 -5814 331294
rect -5578 331058 -5494 331294
rect -5258 331058 -5226 331294
rect -5846 295614 -5226 331058
rect -5846 295378 -5814 295614
rect -5578 295378 -5494 295614
rect -5258 295378 -5226 295614
rect -5846 295294 -5226 295378
rect -5846 295058 -5814 295294
rect -5578 295058 -5494 295294
rect -5258 295058 -5226 295294
rect -5846 259614 -5226 295058
rect -5846 259378 -5814 259614
rect -5578 259378 -5494 259614
rect -5258 259378 -5226 259614
rect -5846 259294 -5226 259378
rect -5846 259058 -5814 259294
rect -5578 259058 -5494 259294
rect -5258 259058 -5226 259294
rect -5846 223614 -5226 259058
rect -5846 223378 -5814 223614
rect -5578 223378 -5494 223614
rect -5258 223378 -5226 223614
rect -5846 223294 -5226 223378
rect -5846 223058 -5814 223294
rect -5578 223058 -5494 223294
rect -5258 223058 -5226 223294
rect -5846 187614 -5226 223058
rect -5846 187378 -5814 187614
rect -5578 187378 -5494 187614
rect -5258 187378 -5226 187614
rect -5846 187294 -5226 187378
rect -5846 187058 -5814 187294
rect -5578 187058 -5494 187294
rect -5258 187058 -5226 187294
rect -5846 151614 -5226 187058
rect -5846 151378 -5814 151614
rect -5578 151378 -5494 151614
rect -5258 151378 -5226 151614
rect -5846 151294 -5226 151378
rect -5846 151058 -5814 151294
rect -5578 151058 -5494 151294
rect -5258 151058 -5226 151294
rect -5846 115614 -5226 151058
rect -5846 115378 -5814 115614
rect -5578 115378 -5494 115614
rect -5258 115378 -5226 115614
rect -5846 115294 -5226 115378
rect -5846 115058 -5814 115294
rect -5578 115058 -5494 115294
rect -5258 115058 -5226 115294
rect -5846 79614 -5226 115058
rect -5846 79378 -5814 79614
rect -5578 79378 -5494 79614
rect -5258 79378 -5226 79614
rect -5846 79294 -5226 79378
rect -5846 79058 -5814 79294
rect -5578 79058 -5494 79294
rect -5258 79058 -5226 79294
rect -5846 43614 -5226 79058
rect -5846 43378 -5814 43614
rect -5578 43378 -5494 43614
rect -5258 43378 -5226 43614
rect -5846 43294 -5226 43378
rect -5846 43058 -5814 43294
rect -5578 43058 -5494 43294
rect -5258 43058 -5226 43294
rect -5846 7614 -5226 43058
rect -5846 7378 -5814 7614
rect -5578 7378 -5494 7614
rect -5258 7378 -5226 7614
rect -5846 7294 -5226 7378
rect -5846 7058 -5814 7294
rect -5578 7058 -5494 7294
rect -5258 7058 -5226 7294
rect -5846 -4186 -5226 7058
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 690374 -4266 707162
rect -4886 690138 -4854 690374
rect -4618 690138 -4534 690374
rect -4298 690138 -4266 690374
rect -4886 690054 -4266 690138
rect -4886 689818 -4854 690054
rect -4618 689818 -4534 690054
rect -4298 689818 -4266 690054
rect -4886 654374 -4266 689818
rect -4886 654138 -4854 654374
rect -4618 654138 -4534 654374
rect -4298 654138 -4266 654374
rect -4886 654054 -4266 654138
rect -4886 653818 -4854 654054
rect -4618 653818 -4534 654054
rect -4298 653818 -4266 654054
rect -4886 618374 -4266 653818
rect -4886 618138 -4854 618374
rect -4618 618138 -4534 618374
rect -4298 618138 -4266 618374
rect -4886 618054 -4266 618138
rect -4886 617818 -4854 618054
rect -4618 617818 -4534 618054
rect -4298 617818 -4266 618054
rect -4886 582374 -4266 617818
rect -4886 582138 -4854 582374
rect -4618 582138 -4534 582374
rect -4298 582138 -4266 582374
rect -4886 582054 -4266 582138
rect -4886 581818 -4854 582054
rect -4618 581818 -4534 582054
rect -4298 581818 -4266 582054
rect -4886 546374 -4266 581818
rect -4886 546138 -4854 546374
rect -4618 546138 -4534 546374
rect -4298 546138 -4266 546374
rect -4886 546054 -4266 546138
rect -4886 545818 -4854 546054
rect -4618 545818 -4534 546054
rect -4298 545818 -4266 546054
rect -4886 510374 -4266 545818
rect -4886 510138 -4854 510374
rect -4618 510138 -4534 510374
rect -4298 510138 -4266 510374
rect -4886 510054 -4266 510138
rect -4886 509818 -4854 510054
rect -4618 509818 -4534 510054
rect -4298 509818 -4266 510054
rect -4886 474374 -4266 509818
rect -4886 474138 -4854 474374
rect -4618 474138 -4534 474374
rect -4298 474138 -4266 474374
rect -4886 474054 -4266 474138
rect -4886 473818 -4854 474054
rect -4618 473818 -4534 474054
rect -4298 473818 -4266 474054
rect -4886 438374 -4266 473818
rect -4886 438138 -4854 438374
rect -4618 438138 -4534 438374
rect -4298 438138 -4266 438374
rect -4886 438054 -4266 438138
rect -4886 437818 -4854 438054
rect -4618 437818 -4534 438054
rect -4298 437818 -4266 438054
rect -4886 402374 -4266 437818
rect -4886 402138 -4854 402374
rect -4618 402138 -4534 402374
rect -4298 402138 -4266 402374
rect -4886 402054 -4266 402138
rect -4886 401818 -4854 402054
rect -4618 401818 -4534 402054
rect -4298 401818 -4266 402054
rect -4886 366374 -4266 401818
rect -4886 366138 -4854 366374
rect -4618 366138 -4534 366374
rect -4298 366138 -4266 366374
rect -4886 366054 -4266 366138
rect -4886 365818 -4854 366054
rect -4618 365818 -4534 366054
rect -4298 365818 -4266 366054
rect -4886 330374 -4266 365818
rect -4886 330138 -4854 330374
rect -4618 330138 -4534 330374
rect -4298 330138 -4266 330374
rect -4886 330054 -4266 330138
rect -4886 329818 -4854 330054
rect -4618 329818 -4534 330054
rect -4298 329818 -4266 330054
rect -4886 294374 -4266 329818
rect -4886 294138 -4854 294374
rect -4618 294138 -4534 294374
rect -4298 294138 -4266 294374
rect -4886 294054 -4266 294138
rect -4886 293818 -4854 294054
rect -4618 293818 -4534 294054
rect -4298 293818 -4266 294054
rect -4886 258374 -4266 293818
rect -4886 258138 -4854 258374
rect -4618 258138 -4534 258374
rect -4298 258138 -4266 258374
rect -4886 258054 -4266 258138
rect -4886 257818 -4854 258054
rect -4618 257818 -4534 258054
rect -4298 257818 -4266 258054
rect -4886 222374 -4266 257818
rect -4886 222138 -4854 222374
rect -4618 222138 -4534 222374
rect -4298 222138 -4266 222374
rect -4886 222054 -4266 222138
rect -4886 221818 -4854 222054
rect -4618 221818 -4534 222054
rect -4298 221818 -4266 222054
rect -4886 186374 -4266 221818
rect -4886 186138 -4854 186374
rect -4618 186138 -4534 186374
rect -4298 186138 -4266 186374
rect -4886 186054 -4266 186138
rect -4886 185818 -4854 186054
rect -4618 185818 -4534 186054
rect -4298 185818 -4266 186054
rect -4886 150374 -4266 185818
rect -4886 150138 -4854 150374
rect -4618 150138 -4534 150374
rect -4298 150138 -4266 150374
rect -4886 150054 -4266 150138
rect -4886 149818 -4854 150054
rect -4618 149818 -4534 150054
rect -4298 149818 -4266 150054
rect -4886 114374 -4266 149818
rect -4886 114138 -4854 114374
rect -4618 114138 -4534 114374
rect -4298 114138 -4266 114374
rect -4886 114054 -4266 114138
rect -4886 113818 -4854 114054
rect -4618 113818 -4534 114054
rect -4298 113818 -4266 114054
rect -4886 78374 -4266 113818
rect -4886 78138 -4854 78374
rect -4618 78138 -4534 78374
rect -4298 78138 -4266 78374
rect -4886 78054 -4266 78138
rect -4886 77818 -4854 78054
rect -4618 77818 -4534 78054
rect -4298 77818 -4266 78054
rect -4886 42374 -4266 77818
rect -4886 42138 -4854 42374
rect -4618 42138 -4534 42374
rect -4298 42138 -4266 42374
rect -4886 42054 -4266 42138
rect -4886 41818 -4854 42054
rect -4618 41818 -4534 42054
rect -4298 41818 -4266 42054
rect -4886 6374 -4266 41818
rect -4886 6138 -4854 6374
rect -4618 6138 -4534 6374
rect -4298 6138 -4266 6374
rect -4886 6054 -4266 6138
rect -4886 5818 -4854 6054
rect -4618 5818 -4534 6054
rect -4298 5818 -4266 6054
rect -4886 -3226 -4266 5818
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 689134 -3306 706202
rect -3926 688898 -3894 689134
rect -3658 688898 -3574 689134
rect -3338 688898 -3306 689134
rect -3926 688814 -3306 688898
rect -3926 688578 -3894 688814
rect -3658 688578 -3574 688814
rect -3338 688578 -3306 688814
rect -3926 653134 -3306 688578
rect -3926 652898 -3894 653134
rect -3658 652898 -3574 653134
rect -3338 652898 -3306 653134
rect -3926 652814 -3306 652898
rect -3926 652578 -3894 652814
rect -3658 652578 -3574 652814
rect -3338 652578 -3306 652814
rect -3926 617134 -3306 652578
rect -3926 616898 -3894 617134
rect -3658 616898 -3574 617134
rect -3338 616898 -3306 617134
rect -3926 616814 -3306 616898
rect -3926 616578 -3894 616814
rect -3658 616578 -3574 616814
rect -3338 616578 -3306 616814
rect -3926 581134 -3306 616578
rect -3926 580898 -3894 581134
rect -3658 580898 -3574 581134
rect -3338 580898 -3306 581134
rect -3926 580814 -3306 580898
rect -3926 580578 -3894 580814
rect -3658 580578 -3574 580814
rect -3338 580578 -3306 580814
rect -3926 545134 -3306 580578
rect -3926 544898 -3894 545134
rect -3658 544898 -3574 545134
rect -3338 544898 -3306 545134
rect -3926 544814 -3306 544898
rect -3926 544578 -3894 544814
rect -3658 544578 -3574 544814
rect -3338 544578 -3306 544814
rect -3926 509134 -3306 544578
rect -3926 508898 -3894 509134
rect -3658 508898 -3574 509134
rect -3338 508898 -3306 509134
rect -3926 508814 -3306 508898
rect -3926 508578 -3894 508814
rect -3658 508578 -3574 508814
rect -3338 508578 -3306 508814
rect -3926 473134 -3306 508578
rect -3926 472898 -3894 473134
rect -3658 472898 -3574 473134
rect -3338 472898 -3306 473134
rect -3926 472814 -3306 472898
rect -3926 472578 -3894 472814
rect -3658 472578 -3574 472814
rect -3338 472578 -3306 472814
rect -3926 437134 -3306 472578
rect -3926 436898 -3894 437134
rect -3658 436898 -3574 437134
rect -3338 436898 -3306 437134
rect -3926 436814 -3306 436898
rect -3926 436578 -3894 436814
rect -3658 436578 -3574 436814
rect -3338 436578 -3306 436814
rect -3926 401134 -3306 436578
rect -3926 400898 -3894 401134
rect -3658 400898 -3574 401134
rect -3338 400898 -3306 401134
rect -3926 400814 -3306 400898
rect -3926 400578 -3894 400814
rect -3658 400578 -3574 400814
rect -3338 400578 -3306 400814
rect -3926 365134 -3306 400578
rect -3926 364898 -3894 365134
rect -3658 364898 -3574 365134
rect -3338 364898 -3306 365134
rect -3926 364814 -3306 364898
rect -3926 364578 -3894 364814
rect -3658 364578 -3574 364814
rect -3338 364578 -3306 364814
rect -3926 329134 -3306 364578
rect -3926 328898 -3894 329134
rect -3658 328898 -3574 329134
rect -3338 328898 -3306 329134
rect -3926 328814 -3306 328898
rect -3926 328578 -3894 328814
rect -3658 328578 -3574 328814
rect -3338 328578 -3306 328814
rect -3926 293134 -3306 328578
rect -3926 292898 -3894 293134
rect -3658 292898 -3574 293134
rect -3338 292898 -3306 293134
rect -3926 292814 -3306 292898
rect -3926 292578 -3894 292814
rect -3658 292578 -3574 292814
rect -3338 292578 -3306 292814
rect -3926 257134 -3306 292578
rect -3926 256898 -3894 257134
rect -3658 256898 -3574 257134
rect -3338 256898 -3306 257134
rect -3926 256814 -3306 256898
rect -3926 256578 -3894 256814
rect -3658 256578 -3574 256814
rect -3338 256578 -3306 256814
rect -3926 221134 -3306 256578
rect -3926 220898 -3894 221134
rect -3658 220898 -3574 221134
rect -3338 220898 -3306 221134
rect -3926 220814 -3306 220898
rect -3926 220578 -3894 220814
rect -3658 220578 -3574 220814
rect -3338 220578 -3306 220814
rect -3926 185134 -3306 220578
rect -3926 184898 -3894 185134
rect -3658 184898 -3574 185134
rect -3338 184898 -3306 185134
rect -3926 184814 -3306 184898
rect -3926 184578 -3894 184814
rect -3658 184578 -3574 184814
rect -3338 184578 -3306 184814
rect -3926 149134 -3306 184578
rect -3926 148898 -3894 149134
rect -3658 148898 -3574 149134
rect -3338 148898 -3306 149134
rect -3926 148814 -3306 148898
rect -3926 148578 -3894 148814
rect -3658 148578 -3574 148814
rect -3338 148578 -3306 148814
rect -3926 113134 -3306 148578
rect -3926 112898 -3894 113134
rect -3658 112898 -3574 113134
rect -3338 112898 -3306 113134
rect -3926 112814 -3306 112898
rect -3926 112578 -3894 112814
rect -3658 112578 -3574 112814
rect -3338 112578 -3306 112814
rect -3926 77134 -3306 112578
rect -3926 76898 -3894 77134
rect -3658 76898 -3574 77134
rect -3338 76898 -3306 77134
rect -3926 76814 -3306 76898
rect -3926 76578 -3894 76814
rect -3658 76578 -3574 76814
rect -3338 76578 -3306 76814
rect -3926 41134 -3306 76578
rect -3926 40898 -3894 41134
rect -3658 40898 -3574 41134
rect -3338 40898 -3306 41134
rect -3926 40814 -3306 40898
rect -3926 40578 -3894 40814
rect -3658 40578 -3574 40814
rect -3338 40578 -3306 40814
rect -3926 5134 -3306 40578
rect -3926 4898 -3894 5134
rect -3658 4898 -3574 5134
rect -3338 4898 -3306 5134
rect -3926 4814 -3306 4898
rect -3926 4578 -3894 4814
rect -3658 4578 -3574 4814
rect -3338 4578 -3306 4814
rect -3926 -2266 -3306 4578
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 687894 -2346 705242
rect -2966 687658 -2934 687894
rect -2698 687658 -2614 687894
rect -2378 687658 -2346 687894
rect -2966 687574 -2346 687658
rect -2966 687338 -2934 687574
rect -2698 687338 -2614 687574
rect -2378 687338 -2346 687574
rect -2966 651894 -2346 687338
rect -2966 651658 -2934 651894
rect -2698 651658 -2614 651894
rect -2378 651658 -2346 651894
rect -2966 651574 -2346 651658
rect -2966 651338 -2934 651574
rect -2698 651338 -2614 651574
rect -2378 651338 -2346 651574
rect -2966 615894 -2346 651338
rect -2966 615658 -2934 615894
rect -2698 615658 -2614 615894
rect -2378 615658 -2346 615894
rect -2966 615574 -2346 615658
rect -2966 615338 -2934 615574
rect -2698 615338 -2614 615574
rect -2378 615338 -2346 615574
rect -2966 579894 -2346 615338
rect -2966 579658 -2934 579894
rect -2698 579658 -2614 579894
rect -2378 579658 -2346 579894
rect -2966 579574 -2346 579658
rect -2966 579338 -2934 579574
rect -2698 579338 -2614 579574
rect -2378 579338 -2346 579574
rect -2966 543894 -2346 579338
rect -2966 543658 -2934 543894
rect -2698 543658 -2614 543894
rect -2378 543658 -2346 543894
rect -2966 543574 -2346 543658
rect -2966 543338 -2934 543574
rect -2698 543338 -2614 543574
rect -2378 543338 -2346 543574
rect -2966 507894 -2346 543338
rect -2966 507658 -2934 507894
rect -2698 507658 -2614 507894
rect -2378 507658 -2346 507894
rect -2966 507574 -2346 507658
rect -2966 507338 -2934 507574
rect -2698 507338 -2614 507574
rect -2378 507338 -2346 507574
rect -2966 471894 -2346 507338
rect -2966 471658 -2934 471894
rect -2698 471658 -2614 471894
rect -2378 471658 -2346 471894
rect -2966 471574 -2346 471658
rect -2966 471338 -2934 471574
rect -2698 471338 -2614 471574
rect -2378 471338 -2346 471574
rect -2966 435894 -2346 471338
rect -2966 435658 -2934 435894
rect -2698 435658 -2614 435894
rect -2378 435658 -2346 435894
rect -2966 435574 -2346 435658
rect -2966 435338 -2934 435574
rect -2698 435338 -2614 435574
rect -2378 435338 -2346 435574
rect -2966 399894 -2346 435338
rect -2966 399658 -2934 399894
rect -2698 399658 -2614 399894
rect -2378 399658 -2346 399894
rect -2966 399574 -2346 399658
rect -2966 399338 -2934 399574
rect -2698 399338 -2614 399574
rect -2378 399338 -2346 399574
rect -2966 363894 -2346 399338
rect -2966 363658 -2934 363894
rect -2698 363658 -2614 363894
rect -2378 363658 -2346 363894
rect -2966 363574 -2346 363658
rect -2966 363338 -2934 363574
rect -2698 363338 -2614 363574
rect -2378 363338 -2346 363574
rect -2966 327894 -2346 363338
rect -2966 327658 -2934 327894
rect -2698 327658 -2614 327894
rect -2378 327658 -2346 327894
rect -2966 327574 -2346 327658
rect -2966 327338 -2934 327574
rect -2698 327338 -2614 327574
rect -2378 327338 -2346 327574
rect -2966 291894 -2346 327338
rect -2966 291658 -2934 291894
rect -2698 291658 -2614 291894
rect -2378 291658 -2346 291894
rect -2966 291574 -2346 291658
rect -2966 291338 -2934 291574
rect -2698 291338 -2614 291574
rect -2378 291338 -2346 291574
rect -2966 255894 -2346 291338
rect -2966 255658 -2934 255894
rect -2698 255658 -2614 255894
rect -2378 255658 -2346 255894
rect -2966 255574 -2346 255658
rect -2966 255338 -2934 255574
rect -2698 255338 -2614 255574
rect -2378 255338 -2346 255574
rect -2966 219894 -2346 255338
rect -2966 219658 -2934 219894
rect -2698 219658 -2614 219894
rect -2378 219658 -2346 219894
rect -2966 219574 -2346 219658
rect -2966 219338 -2934 219574
rect -2698 219338 -2614 219574
rect -2378 219338 -2346 219574
rect -2966 183894 -2346 219338
rect -2966 183658 -2934 183894
rect -2698 183658 -2614 183894
rect -2378 183658 -2346 183894
rect -2966 183574 -2346 183658
rect -2966 183338 -2934 183574
rect -2698 183338 -2614 183574
rect -2378 183338 -2346 183574
rect -2966 147894 -2346 183338
rect -2966 147658 -2934 147894
rect -2698 147658 -2614 147894
rect -2378 147658 -2346 147894
rect -2966 147574 -2346 147658
rect -2966 147338 -2934 147574
rect -2698 147338 -2614 147574
rect -2378 147338 -2346 147574
rect -2966 111894 -2346 147338
rect -2966 111658 -2934 111894
rect -2698 111658 -2614 111894
rect -2378 111658 -2346 111894
rect -2966 111574 -2346 111658
rect -2966 111338 -2934 111574
rect -2698 111338 -2614 111574
rect -2378 111338 -2346 111574
rect -2966 75894 -2346 111338
rect -2966 75658 -2934 75894
rect -2698 75658 -2614 75894
rect -2378 75658 -2346 75894
rect -2966 75574 -2346 75658
rect -2966 75338 -2934 75574
rect -2698 75338 -2614 75574
rect -2378 75338 -2346 75574
rect -2966 39894 -2346 75338
rect -2966 39658 -2934 39894
rect -2698 39658 -2614 39894
rect -2378 39658 -2346 39894
rect -2966 39574 -2346 39658
rect -2966 39338 -2934 39574
rect -2698 39338 -2614 39574
rect -2378 39338 -2346 39574
rect -2966 3894 -2346 39338
rect -2966 3658 -2934 3894
rect -2698 3658 -2614 3894
rect -2378 3658 -2346 3894
rect -2966 3574 -2346 3658
rect -2966 3338 -2934 3574
rect -2698 3338 -2614 3574
rect -2378 3338 -2346 3574
rect -2966 -1306 -2346 3338
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 686654 -1386 704282
rect -2006 686418 -1974 686654
rect -1738 686418 -1654 686654
rect -1418 686418 -1386 686654
rect -2006 686334 -1386 686418
rect -2006 686098 -1974 686334
rect -1738 686098 -1654 686334
rect -1418 686098 -1386 686334
rect -2006 650654 -1386 686098
rect -2006 650418 -1974 650654
rect -1738 650418 -1654 650654
rect -1418 650418 -1386 650654
rect -2006 650334 -1386 650418
rect -2006 650098 -1974 650334
rect -1738 650098 -1654 650334
rect -1418 650098 -1386 650334
rect -2006 614654 -1386 650098
rect -2006 614418 -1974 614654
rect -1738 614418 -1654 614654
rect -1418 614418 -1386 614654
rect -2006 614334 -1386 614418
rect -2006 614098 -1974 614334
rect -1738 614098 -1654 614334
rect -1418 614098 -1386 614334
rect -2006 578654 -1386 614098
rect -2006 578418 -1974 578654
rect -1738 578418 -1654 578654
rect -1418 578418 -1386 578654
rect -2006 578334 -1386 578418
rect -2006 578098 -1974 578334
rect -1738 578098 -1654 578334
rect -1418 578098 -1386 578334
rect -2006 542654 -1386 578098
rect -2006 542418 -1974 542654
rect -1738 542418 -1654 542654
rect -1418 542418 -1386 542654
rect -2006 542334 -1386 542418
rect -2006 542098 -1974 542334
rect -1738 542098 -1654 542334
rect -1418 542098 -1386 542334
rect -2006 506654 -1386 542098
rect -2006 506418 -1974 506654
rect -1738 506418 -1654 506654
rect -1418 506418 -1386 506654
rect -2006 506334 -1386 506418
rect -2006 506098 -1974 506334
rect -1738 506098 -1654 506334
rect -1418 506098 -1386 506334
rect -2006 470654 -1386 506098
rect -2006 470418 -1974 470654
rect -1738 470418 -1654 470654
rect -1418 470418 -1386 470654
rect -2006 470334 -1386 470418
rect -2006 470098 -1974 470334
rect -1738 470098 -1654 470334
rect -1418 470098 -1386 470334
rect -2006 434654 -1386 470098
rect -2006 434418 -1974 434654
rect -1738 434418 -1654 434654
rect -1418 434418 -1386 434654
rect -2006 434334 -1386 434418
rect -2006 434098 -1974 434334
rect -1738 434098 -1654 434334
rect -1418 434098 -1386 434334
rect -2006 398654 -1386 434098
rect -2006 398418 -1974 398654
rect -1738 398418 -1654 398654
rect -1418 398418 -1386 398654
rect -2006 398334 -1386 398418
rect -2006 398098 -1974 398334
rect -1738 398098 -1654 398334
rect -1418 398098 -1386 398334
rect -2006 362654 -1386 398098
rect -2006 362418 -1974 362654
rect -1738 362418 -1654 362654
rect -1418 362418 -1386 362654
rect -2006 362334 -1386 362418
rect -2006 362098 -1974 362334
rect -1738 362098 -1654 362334
rect -1418 362098 -1386 362334
rect -2006 326654 -1386 362098
rect -2006 326418 -1974 326654
rect -1738 326418 -1654 326654
rect -1418 326418 -1386 326654
rect -2006 326334 -1386 326418
rect -2006 326098 -1974 326334
rect -1738 326098 -1654 326334
rect -1418 326098 -1386 326334
rect -2006 290654 -1386 326098
rect -2006 290418 -1974 290654
rect -1738 290418 -1654 290654
rect -1418 290418 -1386 290654
rect -2006 290334 -1386 290418
rect -2006 290098 -1974 290334
rect -1738 290098 -1654 290334
rect -1418 290098 -1386 290334
rect -2006 254654 -1386 290098
rect -2006 254418 -1974 254654
rect -1738 254418 -1654 254654
rect -1418 254418 -1386 254654
rect -2006 254334 -1386 254418
rect -2006 254098 -1974 254334
rect -1738 254098 -1654 254334
rect -1418 254098 -1386 254334
rect -2006 218654 -1386 254098
rect -2006 218418 -1974 218654
rect -1738 218418 -1654 218654
rect -1418 218418 -1386 218654
rect -2006 218334 -1386 218418
rect -2006 218098 -1974 218334
rect -1738 218098 -1654 218334
rect -1418 218098 -1386 218334
rect -2006 182654 -1386 218098
rect -2006 182418 -1974 182654
rect -1738 182418 -1654 182654
rect -1418 182418 -1386 182654
rect -2006 182334 -1386 182418
rect -2006 182098 -1974 182334
rect -1738 182098 -1654 182334
rect -1418 182098 -1386 182334
rect -2006 146654 -1386 182098
rect -2006 146418 -1974 146654
rect -1738 146418 -1654 146654
rect -1418 146418 -1386 146654
rect -2006 146334 -1386 146418
rect -2006 146098 -1974 146334
rect -1738 146098 -1654 146334
rect -1418 146098 -1386 146334
rect -2006 110654 -1386 146098
rect -2006 110418 -1974 110654
rect -1738 110418 -1654 110654
rect -1418 110418 -1386 110654
rect -2006 110334 -1386 110418
rect -2006 110098 -1974 110334
rect -1738 110098 -1654 110334
rect -1418 110098 -1386 110334
rect -2006 74654 -1386 110098
rect -2006 74418 -1974 74654
rect -1738 74418 -1654 74654
rect -1418 74418 -1386 74654
rect -2006 74334 -1386 74418
rect -2006 74098 -1974 74334
rect -1738 74098 -1654 74334
rect -1418 74098 -1386 74334
rect -2006 38654 -1386 74098
rect -2006 38418 -1974 38654
rect -1738 38418 -1654 38654
rect -1418 38418 -1386 38654
rect -2006 38334 -1386 38418
rect -2006 38098 -1974 38334
rect -1738 38098 -1654 38334
rect -1418 38098 -1386 38334
rect -2006 2654 -1386 38098
rect -2006 2418 -1974 2654
rect -1738 2418 -1654 2654
rect -1418 2418 -1386 2654
rect -2006 2334 -1386 2418
rect -2006 2098 -1974 2334
rect -1738 2098 -1654 2334
rect -1418 2098 -1386 2334
rect -2006 -346 -1386 2098
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 994 704838 1614 711590
rect 994 704602 1026 704838
rect 1262 704602 1346 704838
rect 1582 704602 1614 704838
rect 994 704518 1614 704602
rect 994 704282 1026 704518
rect 1262 704282 1346 704518
rect 1582 704282 1614 704518
rect 994 686654 1614 704282
rect 994 686418 1026 686654
rect 1262 686418 1346 686654
rect 1582 686418 1614 686654
rect 994 686334 1614 686418
rect 994 686098 1026 686334
rect 1262 686098 1346 686334
rect 1582 686098 1614 686334
rect 994 650654 1614 686098
rect 994 650418 1026 650654
rect 1262 650418 1346 650654
rect 1582 650418 1614 650654
rect 994 650334 1614 650418
rect 994 650098 1026 650334
rect 1262 650098 1346 650334
rect 1582 650098 1614 650334
rect 994 614654 1614 650098
rect 994 614418 1026 614654
rect 1262 614418 1346 614654
rect 1582 614418 1614 614654
rect 994 614334 1614 614418
rect 994 614098 1026 614334
rect 1262 614098 1346 614334
rect 1582 614098 1614 614334
rect 994 578654 1614 614098
rect 994 578418 1026 578654
rect 1262 578418 1346 578654
rect 1582 578418 1614 578654
rect 994 578334 1614 578418
rect 994 578098 1026 578334
rect 1262 578098 1346 578334
rect 1582 578098 1614 578334
rect 994 542654 1614 578098
rect 994 542418 1026 542654
rect 1262 542418 1346 542654
rect 1582 542418 1614 542654
rect 994 542334 1614 542418
rect 994 542098 1026 542334
rect 1262 542098 1346 542334
rect 1582 542098 1614 542334
rect 994 506654 1614 542098
rect 994 506418 1026 506654
rect 1262 506418 1346 506654
rect 1582 506418 1614 506654
rect 994 506334 1614 506418
rect 994 506098 1026 506334
rect 1262 506098 1346 506334
rect 1582 506098 1614 506334
rect 994 470654 1614 506098
rect 994 470418 1026 470654
rect 1262 470418 1346 470654
rect 1582 470418 1614 470654
rect 994 470334 1614 470418
rect 994 470098 1026 470334
rect 1262 470098 1346 470334
rect 1582 470098 1614 470334
rect 994 434654 1614 470098
rect 994 434418 1026 434654
rect 1262 434418 1346 434654
rect 1582 434418 1614 434654
rect 994 434334 1614 434418
rect 994 434098 1026 434334
rect 1262 434098 1346 434334
rect 1582 434098 1614 434334
rect 994 398654 1614 434098
rect 994 398418 1026 398654
rect 1262 398418 1346 398654
rect 1582 398418 1614 398654
rect 994 398334 1614 398418
rect 994 398098 1026 398334
rect 1262 398098 1346 398334
rect 1582 398098 1614 398334
rect 994 362654 1614 398098
rect 994 362418 1026 362654
rect 1262 362418 1346 362654
rect 1582 362418 1614 362654
rect 994 362334 1614 362418
rect 994 362098 1026 362334
rect 1262 362098 1346 362334
rect 1582 362098 1614 362334
rect 994 326654 1614 362098
rect 994 326418 1026 326654
rect 1262 326418 1346 326654
rect 1582 326418 1614 326654
rect 994 326334 1614 326418
rect 994 326098 1026 326334
rect 1262 326098 1346 326334
rect 1582 326098 1614 326334
rect 994 290654 1614 326098
rect 994 290418 1026 290654
rect 1262 290418 1346 290654
rect 1582 290418 1614 290654
rect 994 290334 1614 290418
rect 994 290098 1026 290334
rect 1262 290098 1346 290334
rect 1582 290098 1614 290334
rect 994 254654 1614 290098
rect 994 254418 1026 254654
rect 1262 254418 1346 254654
rect 1582 254418 1614 254654
rect 994 254334 1614 254418
rect 994 254098 1026 254334
rect 1262 254098 1346 254334
rect 1582 254098 1614 254334
rect 994 218654 1614 254098
rect 994 218418 1026 218654
rect 1262 218418 1346 218654
rect 1582 218418 1614 218654
rect 994 218334 1614 218418
rect 994 218098 1026 218334
rect 1262 218098 1346 218334
rect 1582 218098 1614 218334
rect 994 182654 1614 218098
rect 994 182418 1026 182654
rect 1262 182418 1346 182654
rect 1582 182418 1614 182654
rect 994 182334 1614 182418
rect 994 182098 1026 182334
rect 1262 182098 1346 182334
rect 1582 182098 1614 182334
rect 994 146654 1614 182098
rect 994 146418 1026 146654
rect 1262 146418 1346 146654
rect 1582 146418 1614 146654
rect 994 146334 1614 146418
rect 994 146098 1026 146334
rect 1262 146098 1346 146334
rect 1582 146098 1614 146334
rect 994 110654 1614 146098
rect 994 110418 1026 110654
rect 1262 110418 1346 110654
rect 1582 110418 1614 110654
rect 994 110334 1614 110418
rect 994 110098 1026 110334
rect 1262 110098 1346 110334
rect 1582 110098 1614 110334
rect 994 74654 1614 110098
rect 994 74418 1026 74654
rect 1262 74418 1346 74654
rect 1582 74418 1614 74654
rect 994 74334 1614 74418
rect 994 74098 1026 74334
rect 1262 74098 1346 74334
rect 1582 74098 1614 74334
rect 994 38654 1614 74098
rect 994 38418 1026 38654
rect 1262 38418 1346 38654
rect 1582 38418 1614 38654
rect 994 38334 1614 38418
rect 994 38098 1026 38334
rect 1262 38098 1346 38334
rect 1582 38098 1614 38334
rect 994 2654 1614 38098
rect 994 2418 1026 2654
rect 1262 2418 1346 2654
rect 1582 2418 1614 2654
rect 994 2334 1614 2418
rect 994 2098 1026 2334
rect 1262 2098 1346 2334
rect 1582 2098 1614 2334
rect 994 -346 1614 2098
rect 994 -582 1026 -346
rect 1262 -582 1346 -346
rect 1582 -582 1614 -346
rect 994 -666 1614 -582
rect 994 -902 1026 -666
rect 1262 -902 1346 -666
rect 1582 -902 1614 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 994 -7654 1614 -902
rect 2234 705798 2854 711590
rect 2234 705562 2266 705798
rect 2502 705562 2586 705798
rect 2822 705562 2854 705798
rect 2234 705478 2854 705562
rect 2234 705242 2266 705478
rect 2502 705242 2586 705478
rect 2822 705242 2854 705478
rect 2234 687894 2854 705242
rect 2234 687658 2266 687894
rect 2502 687658 2586 687894
rect 2822 687658 2854 687894
rect 2234 687574 2854 687658
rect 2234 687338 2266 687574
rect 2502 687338 2586 687574
rect 2822 687338 2854 687574
rect 2234 651894 2854 687338
rect 2234 651658 2266 651894
rect 2502 651658 2586 651894
rect 2822 651658 2854 651894
rect 2234 651574 2854 651658
rect 2234 651338 2266 651574
rect 2502 651338 2586 651574
rect 2822 651338 2854 651574
rect 2234 615894 2854 651338
rect 2234 615658 2266 615894
rect 2502 615658 2586 615894
rect 2822 615658 2854 615894
rect 2234 615574 2854 615658
rect 2234 615338 2266 615574
rect 2502 615338 2586 615574
rect 2822 615338 2854 615574
rect 2234 579894 2854 615338
rect 2234 579658 2266 579894
rect 2502 579658 2586 579894
rect 2822 579658 2854 579894
rect 2234 579574 2854 579658
rect 2234 579338 2266 579574
rect 2502 579338 2586 579574
rect 2822 579338 2854 579574
rect 2234 543894 2854 579338
rect 2234 543658 2266 543894
rect 2502 543658 2586 543894
rect 2822 543658 2854 543894
rect 2234 543574 2854 543658
rect 2234 543338 2266 543574
rect 2502 543338 2586 543574
rect 2822 543338 2854 543574
rect 2234 507894 2854 543338
rect 2234 507658 2266 507894
rect 2502 507658 2586 507894
rect 2822 507658 2854 507894
rect 2234 507574 2854 507658
rect 2234 507338 2266 507574
rect 2502 507338 2586 507574
rect 2822 507338 2854 507574
rect 2234 471894 2854 507338
rect 2234 471658 2266 471894
rect 2502 471658 2586 471894
rect 2822 471658 2854 471894
rect 2234 471574 2854 471658
rect 2234 471338 2266 471574
rect 2502 471338 2586 471574
rect 2822 471338 2854 471574
rect 2234 435894 2854 471338
rect 2234 435658 2266 435894
rect 2502 435658 2586 435894
rect 2822 435658 2854 435894
rect 2234 435574 2854 435658
rect 2234 435338 2266 435574
rect 2502 435338 2586 435574
rect 2822 435338 2854 435574
rect 2234 399894 2854 435338
rect 2234 399658 2266 399894
rect 2502 399658 2586 399894
rect 2822 399658 2854 399894
rect 2234 399574 2854 399658
rect 2234 399338 2266 399574
rect 2502 399338 2586 399574
rect 2822 399338 2854 399574
rect 2234 363894 2854 399338
rect 2234 363658 2266 363894
rect 2502 363658 2586 363894
rect 2822 363658 2854 363894
rect 2234 363574 2854 363658
rect 2234 363338 2266 363574
rect 2502 363338 2586 363574
rect 2822 363338 2854 363574
rect 2234 327894 2854 363338
rect 2234 327658 2266 327894
rect 2502 327658 2586 327894
rect 2822 327658 2854 327894
rect 2234 327574 2854 327658
rect 2234 327338 2266 327574
rect 2502 327338 2586 327574
rect 2822 327338 2854 327574
rect 2234 291894 2854 327338
rect 2234 291658 2266 291894
rect 2502 291658 2586 291894
rect 2822 291658 2854 291894
rect 2234 291574 2854 291658
rect 2234 291338 2266 291574
rect 2502 291338 2586 291574
rect 2822 291338 2854 291574
rect 2234 255894 2854 291338
rect 2234 255658 2266 255894
rect 2502 255658 2586 255894
rect 2822 255658 2854 255894
rect 2234 255574 2854 255658
rect 2234 255338 2266 255574
rect 2502 255338 2586 255574
rect 2822 255338 2854 255574
rect 2234 219894 2854 255338
rect 2234 219658 2266 219894
rect 2502 219658 2586 219894
rect 2822 219658 2854 219894
rect 2234 219574 2854 219658
rect 2234 219338 2266 219574
rect 2502 219338 2586 219574
rect 2822 219338 2854 219574
rect 2234 183894 2854 219338
rect 2234 183658 2266 183894
rect 2502 183658 2586 183894
rect 2822 183658 2854 183894
rect 2234 183574 2854 183658
rect 2234 183338 2266 183574
rect 2502 183338 2586 183574
rect 2822 183338 2854 183574
rect 2234 147894 2854 183338
rect 2234 147658 2266 147894
rect 2502 147658 2586 147894
rect 2822 147658 2854 147894
rect 2234 147574 2854 147658
rect 2234 147338 2266 147574
rect 2502 147338 2586 147574
rect 2822 147338 2854 147574
rect 2234 111894 2854 147338
rect 2234 111658 2266 111894
rect 2502 111658 2586 111894
rect 2822 111658 2854 111894
rect 2234 111574 2854 111658
rect 2234 111338 2266 111574
rect 2502 111338 2586 111574
rect 2822 111338 2854 111574
rect 2234 75894 2854 111338
rect 2234 75658 2266 75894
rect 2502 75658 2586 75894
rect 2822 75658 2854 75894
rect 2234 75574 2854 75658
rect 2234 75338 2266 75574
rect 2502 75338 2586 75574
rect 2822 75338 2854 75574
rect 2234 39894 2854 75338
rect 2234 39658 2266 39894
rect 2502 39658 2586 39894
rect 2822 39658 2854 39894
rect 2234 39574 2854 39658
rect 2234 39338 2266 39574
rect 2502 39338 2586 39574
rect 2822 39338 2854 39574
rect 2234 3894 2854 39338
rect 2234 3658 2266 3894
rect 2502 3658 2586 3894
rect 2822 3658 2854 3894
rect 2234 3574 2854 3658
rect 2234 3338 2266 3574
rect 2502 3338 2586 3574
rect 2822 3338 2854 3574
rect 2234 -1306 2854 3338
rect 2234 -1542 2266 -1306
rect 2502 -1542 2586 -1306
rect 2822 -1542 2854 -1306
rect 2234 -1626 2854 -1542
rect 2234 -1862 2266 -1626
rect 2502 -1862 2586 -1626
rect 2822 -1862 2854 -1626
rect 2234 -7654 2854 -1862
rect 3474 706758 4094 711590
rect 3474 706522 3506 706758
rect 3742 706522 3826 706758
rect 4062 706522 4094 706758
rect 3474 706438 4094 706522
rect 3474 706202 3506 706438
rect 3742 706202 3826 706438
rect 4062 706202 4094 706438
rect 3474 689134 4094 706202
rect 3474 688898 3506 689134
rect 3742 688898 3826 689134
rect 4062 688898 4094 689134
rect 3474 688814 4094 688898
rect 3474 688578 3506 688814
rect 3742 688578 3826 688814
rect 4062 688578 4094 688814
rect 3474 653134 4094 688578
rect 3474 652898 3506 653134
rect 3742 652898 3826 653134
rect 4062 652898 4094 653134
rect 3474 652814 4094 652898
rect 3474 652578 3506 652814
rect 3742 652578 3826 652814
rect 4062 652578 4094 652814
rect 3474 617134 4094 652578
rect 3474 616898 3506 617134
rect 3742 616898 3826 617134
rect 4062 616898 4094 617134
rect 3474 616814 4094 616898
rect 3474 616578 3506 616814
rect 3742 616578 3826 616814
rect 4062 616578 4094 616814
rect 3474 581134 4094 616578
rect 3474 580898 3506 581134
rect 3742 580898 3826 581134
rect 4062 580898 4094 581134
rect 3474 580814 4094 580898
rect 3474 580578 3506 580814
rect 3742 580578 3826 580814
rect 4062 580578 4094 580814
rect 3474 545134 4094 580578
rect 3474 544898 3506 545134
rect 3742 544898 3826 545134
rect 4062 544898 4094 545134
rect 3474 544814 4094 544898
rect 3474 544578 3506 544814
rect 3742 544578 3826 544814
rect 4062 544578 4094 544814
rect 3474 509134 4094 544578
rect 3474 508898 3506 509134
rect 3742 508898 3826 509134
rect 4062 508898 4094 509134
rect 3474 508814 4094 508898
rect 3474 508578 3506 508814
rect 3742 508578 3826 508814
rect 4062 508578 4094 508814
rect 3474 473134 4094 508578
rect 3474 472898 3506 473134
rect 3742 472898 3826 473134
rect 4062 472898 4094 473134
rect 3474 472814 4094 472898
rect 3474 472578 3506 472814
rect 3742 472578 3826 472814
rect 4062 472578 4094 472814
rect 3474 437134 4094 472578
rect 3474 436898 3506 437134
rect 3742 436898 3826 437134
rect 4062 436898 4094 437134
rect 3474 436814 4094 436898
rect 3474 436578 3506 436814
rect 3742 436578 3826 436814
rect 4062 436578 4094 436814
rect 3474 401134 4094 436578
rect 3474 400898 3506 401134
rect 3742 400898 3826 401134
rect 4062 400898 4094 401134
rect 3474 400814 4094 400898
rect 3474 400578 3506 400814
rect 3742 400578 3826 400814
rect 4062 400578 4094 400814
rect 3474 365134 4094 400578
rect 3474 364898 3506 365134
rect 3742 364898 3826 365134
rect 4062 364898 4094 365134
rect 3474 364814 4094 364898
rect 3474 364578 3506 364814
rect 3742 364578 3826 364814
rect 4062 364578 4094 364814
rect 3474 329134 4094 364578
rect 3474 328898 3506 329134
rect 3742 328898 3826 329134
rect 4062 328898 4094 329134
rect 3474 328814 4094 328898
rect 3474 328578 3506 328814
rect 3742 328578 3826 328814
rect 4062 328578 4094 328814
rect 3474 293134 4094 328578
rect 3474 292898 3506 293134
rect 3742 292898 3826 293134
rect 4062 292898 4094 293134
rect 3474 292814 4094 292898
rect 3474 292578 3506 292814
rect 3742 292578 3826 292814
rect 4062 292578 4094 292814
rect 3474 257134 4094 292578
rect 3474 256898 3506 257134
rect 3742 256898 3826 257134
rect 4062 256898 4094 257134
rect 3474 256814 4094 256898
rect 3474 256578 3506 256814
rect 3742 256578 3826 256814
rect 4062 256578 4094 256814
rect 3474 221134 4094 256578
rect 3474 220898 3506 221134
rect 3742 220898 3826 221134
rect 4062 220898 4094 221134
rect 3474 220814 4094 220898
rect 3474 220578 3506 220814
rect 3742 220578 3826 220814
rect 4062 220578 4094 220814
rect 3474 185134 4094 220578
rect 3474 184898 3506 185134
rect 3742 184898 3826 185134
rect 4062 184898 4094 185134
rect 3474 184814 4094 184898
rect 3474 184578 3506 184814
rect 3742 184578 3826 184814
rect 4062 184578 4094 184814
rect 3474 149134 4094 184578
rect 3474 148898 3506 149134
rect 3742 148898 3826 149134
rect 4062 148898 4094 149134
rect 3474 148814 4094 148898
rect 3474 148578 3506 148814
rect 3742 148578 3826 148814
rect 4062 148578 4094 148814
rect 3474 113134 4094 148578
rect 3474 112898 3506 113134
rect 3742 112898 3826 113134
rect 4062 112898 4094 113134
rect 3474 112814 4094 112898
rect 3474 112578 3506 112814
rect 3742 112578 3826 112814
rect 4062 112578 4094 112814
rect 3474 77134 4094 112578
rect 3474 76898 3506 77134
rect 3742 76898 3826 77134
rect 4062 76898 4094 77134
rect 3474 76814 4094 76898
rect 3474 76578 3506 76814
rect 3742 76578 3826 76814
rect 4062 76578 4094 76814
rect 3474 41134 4094 76578
rect 3474 40898 3506 41134
rect 3742 40898 3826 41134
rect 4062 40898 4094 41134
rect 3474 40814 4094 40898
rect 3474 40578 3506 40814
rect 3742 40578 3826 40814
rect 4062 40578 4094 40814
rect 3474 5134 4094 40578
rect 3474 4898 3506 5134
rect 3742 4898 3826 5134
rect 4062 4898 4094 5134
rect 3474 4814 4094 4898
rect 3474 4578 3506 4814
rect 3742 4578 3826 4814
rect 4062 4578 4094 4814
rect 3474 -2266 4094 4578
rect 3474 -2502 3506 -2266
rect 3742 -2502 3826 -2266
rect 4062 -2502 4094 -2266
rect 3474 -2586 4094 -2502
rect 3474 -2822 3506 -2586
rect 3742 -2822 3826 -2586
rect 4062 -2822 4094 -2586
rect 3474 -7654 4094 -2822
rect 4714 707718 5334 711590
rect 4714 707482 4746 707718
rect 4982 707482 5066 707718
rect 5302 707482 5334 707718
rect 4714 707398 5334 707482
rect 4714 707162 4746 707398
rect 4982 707162 5066 707398
rect 5302 707162 5334 707398
rect 4714 690374 5334 707162
rect 4714 690138 4746 690374
rect 4982 690138 5066 690374
rect 5302 690138 5334 690374
rect 4714 690054 5334 690138
rect 4714 689818 4746 690054
rect 4982 689818 5066 690054
rect 5302 689818 5334 690054
rect 4714 654374 5334 689818
rect 4714 654138 4746 654374
rect 4982 654138 5066 654374
rect 5302 654138 5334 654374
rect 4714 654054 5334 654138
rect 4714 653818 4746 654054
rect 4982 653818 5066 654054
rect 5302 653818 5334 654054
rect 4714 618374 5334 653818
rect 4714 618138 4746 618374
rect 4982 618138 5066 618374
rect 5302 618138 5334 618374
rect 4714 618054 5334 618138
rect 4714 617818 4746 618054
rect 4982 617818 5066 618054
rect 5302 617818 5334 618054
rect 4714 582374 5334 617818
rect 4714 582138 4746 582374
rect 4982 582138 5066 582374
rect 5302 582138 5334 582374
rect 4714 582054 5334 582138
rect 4714 581818 4746 582054
rect 4982 581818 5066 582054
rect 5302 581818 5334 582054
rect 4714 546374 5334 581818
rect 4714 546138 4746 546374
rect 4982 546138 5066 546374
rect 5302 546138 5334 546374
rect 4714 546054 5334 546138
rect 4714 545818 4746 546054
rect 4982 545818 5066 546054
rect 5302 545818 5334 546054
rect 4714 510374 5334 545818
rect 4714 510138 4746 510374
rect 4982 510138 5066 510374
rect 5302 510138 5334 510374
rect 4714 510054 5334 510138
rect 4714 509818 4746 510054
rect 4982 509818 5066 510054
rect 5302 509818 5334 510054
rect 4714 474374 5334 509818
rect 4714 474138 4746 474374
rect 4982 474138 5066 474374
rect 5302 474138 5334 474374
rect 4714 474054 5334 474138
rect 4714 473818 4746 474054
rect 4982 473818 5066 474054
rect 5302 473818 5334 474054
rect 4714 438374 5334 473818
rect 4714 438138 4746 438374
rect 4982 438138 5066 438374
rect 5302 438138 5334 438374
rect 4714 438054 5334 438138
rect 4714 437818 4746 438054
rect 4982 437818 5066 438054
rect 5302 437818 5334 438054
rect 4714 402374 5334 437818
rect 4714 402138 4746 402374
rect 4982 402138 5066 402374
rect 5302 402138 5334 402374
rect 4714 402054 5334 402138
rect 4714 401818 4746 402054
rect 4982 401818 5066 402054
rect 5302 401818 5334 402054
rect 4714 366374 5334 401818
rect 4714 366138 4746 366374
rect 4982 366138 5066 366374
rect 5302 366138 5334 366374
rect 4714 366054 5334 366138
rect 4714 365818 4746 366054
rect 4982 365818 5066 366054
rect 5302 365818 5334 366054
rect 4714 330374 5334 365818
rect 4714 330138 4746 330374
rect 4982 330138 5066 330374
rect 5302 330138 5334 330374
rect 4714 330054 5334 330138
rect 4714 329818 4746 330054
rect 4982 329818 5066 330054
rect 5302 329818 5334 330054
rect 4714 294374 5334 329818
rect 4714 294138 4746 294374
rect 4982 294138 5066 294374
rect 5302 294138 5334 294374
rect 4714 294054 5334 294138
rect 4714 293818 4746 294054
rect 4982 293818 5066 294054
rect 5302 293818 5334 294054
rect 4714 258374 5334 293818
rect 4714 258138 4746 258374
rect 4982 258138 5066 258374
rect 5302 258138 5334 258374
rect 4714 258054 5334 258138
rect 4714 257818 4746 258054
rect 4982 257818 5066 258054
rect 5302 257818 5334 258054
rect 4714 222374 5334 257818
rect 4714 222138 4746 222374
rect 4982 222138 5066 222374
rect 5302 222138 5334 222374
rect 4714 222054 5334 222138
rect 4714 221818 4746 222054
rect 4982 221818 5066 222054
rect 5302 221818 5334 222054
rect 4714 186374 5334 221818
rect 4714 186138 4746 186374
rect 4982 186138 5066 186374
rect 5302 186138 5334 186374
rect 4714 186054 5334 186138
rect 4714 185818 4746 186054
rect 4982 185818 5066 186054
rect 5302 185818 5334 186054
rect 4714 150374 5334 185818
rect 4714 150138 4746 150374
rect 4982 150138 5066 150374
rect 5302 150138 5334 150374
rect 4714 150054 5334 150138
rect 4714 149818 4746 150054
rect 4982 149818 5066 150054
rect 5302 149818 5334 150054
rect 4714 114374 5334 149818
rect 4714 114138 4746 114374
rect 4982 114138 5066 114374
rect 5302 114138 5334 114374
rect 4714 114054 5334 114138
rect 4714 113818 4746 114054
rect 4982 113818 5066 114054
rect 5302 113818 5334 114054
rect 4714 78374 5334 113818
rect 4714 78138 4746 78374
rect 4982 78138 5066 78374
rect 5302 78138 5334 78374
rect 4714 78054 5334 78138
rect 4714 77818 4746 78054
rect 4982 77818 5066 78054
rect 5302 77818 5334 78054
rect 4714 42374 5334 77818
rect 4714 42138 4746 42374
rect 4982 42138 5066 42374
rect 5302 42138 5334 42374
rect 4714 42054 5334 42138
rect 4714 41818 4746 42054
rect 4982 41818 5066 42054
rect 5302 41818 5334 42054
rect 4714 6374 5334 41818
rect 4714 6138 4746 6374
rect 4982 6138 5066 6374
rect 5302 6138 5334 6374
rect 4714 6054 5334 6138
rect 4714 5818 4746 6054
rect 4982 5818 5066 6054
rect 5302 5818 5334 6054
rect 4714 -3226 5334 5818
rect 4714 -3462 4746 -3226
rect 4982 -3462 5066 -3226
rect 5302 -3462 5334 -3226
rect 4714 -3546 5334 -3462
rect 4714 -3782 4746 -3546
rect 4982 -3782 5066 -3546
rect 5302 -3782 5334 -3546
rect 4714 -7654 5334 -3782
rect 5954 708678 6574 711590
rect 5954 708442 5986 708678
rect 6222 708442 6306 708678
rect 6542 708442 6574 708678
rect 5954 708358 6574 708442
rect 5954 708122 5986 708358
rect 6222 708122 6306 708358
rect 6542 708122 6574 708358
rect 5954 691614 6574 708122
rect 5954 691378 5986 691614
rect 6222 691378 6306 691614
rect 6542 691378 6574 691614
rect 5954 691294 6574 691378
rect 5954 691058 5986 691294
rect 6222 691058 6306 691294
rect 6542 691058 6574 691294
rect 5954 655614 6574 691058
rect 5954 655378 5986 655614
rect 6222 655378 6306 655614
rect 6542 655378 6574 655614
rect 5954 655294 6574 655378
rect 5954 655058 5986 655294
rect 6222 655058 6306 655294
rect 6542 655058 6574 655294
rect 5954 619614 6574 655058
rect 5954 619378 5986 619614
rect 6222 619378 6306 619614
rect 6542 619378 6574 619614
rect 5954 619294 6574 619378
rect 5954 619058 5986 619294
rect 6222 619058 6306 619294
rect 6542 619058 6574 619294
rect 5954 583614 6574 619058
rect 5954 583378 5986 583614
rect 6222 583378 6306 583614
rect 6542 583378 6574 583614
rect 5954 583294 6574 583378
rect 5954 583058 5986 583294
rect 6222 583058 6306 583294
rect 6542 583058 6574 583294
rect 5954 547614 6574 583058
rect 5954 547378 5986 547614
rect 6222 547378 6306 547614
rect 6542 547378 6574 547614
rect 5954 547294 6574 547378
rect 5954 547058 5986 547294
rect 6222 547058 6306 547294
rect 6542 547058 6574 547294
rect 5954 511614 6574 547058
rect 5954 511378 5986 511614
rect 6222 511378 6306 511614
rect 6542 511378 6574 511614
rect 5954 511294 6574 511378
rect 5954 511058 5986 511294
rect 6222 511058 6306 511294
rect 6542 511058 6574 511294
rect 5954 475614 6574 511058
rect 5954 475378 5986 475614
rect 6222 475378 6306 475614
rect 6542 475378 6574 475614
rect 5954 475294 6574 475378
rect 5954 475058 5986 475294
rect 6222 475058 6306 475294
rect 6542 475058 6574 475294
rect 5954 439614 6574 475058
rect 5954 439378 5986 439614
rect 6222 439378 6306 439614
rect 6542 439378 6574 439614
rect 5954 439294 6574 439378
rect 5954 439058 5986 439294
rect 6222 439058 6306 439294
rect 6542 439058 6574 439294
rect 5954 403614 6574 439058
rect 5954 403378 5986 403614
rect 6222 403378 6306 403614
rect 6542 403378 6574 403614
rect 5954 403294 6574 403378
rect 5954 403058 5986 403294
rect 6222 403058 6306 403294
rect 6542 403058 6574 403294
rect 5954 367614 6574 403058
rect 5954 367378 5986 367614
rect 6222 367378 6306 367614
rect 6542 367378 6574 367614
rect 5954 367294 6574 367378
rect 5954 367058 5986 367294
rect 6222 367058 6306 367294
rect 6542 367058 6574 367294
rect 5954 331614 6574 367058
rect 5954 331378 5986 331614
rect 6222 331378 6306 331614
rect 6542 331378 6574 331614
rect 5954 331294 6574 331378
rect 5954 331058 5986 331294
rect 6222 331058 6306 331294
rect 6542 331058 6574 331294
rect 5954 295614 6574 331058
rect 5954 295378 5986 295614
rect 6222 295378 6306 295614
rect 6542 295378 6574 295614
rect 5954 295294 6574 295378
rect 5954 295058 5986 295294
rect 6222 295058 6306 295294
rect 6542 295058 6574 295294
rect 5954 259614 6574 295058
rect 5954 259378 5986 259614
rect 6222 259378 6306 259614
rect 6542 259378 6574 259614
rect 5954 259294 6574 259378
rect 5954 259058 5986 259294
rect 6222 259058 6306 259294
rect 6542 259058 6574 259294
rect 5954 223614 6574 259058
rect 5954 223378 5986 223614
rect 6222 223378 6306 223614
rect 6542 223378 6574 223614
rect 5954 223294 6574 223378
rect 5954 223058 5986 223294
rect 6222 223058 6306 223294
rect 6542 223058 6574 223294
rect 5954 187614 6574 223058
rect 5954 187378 5986 187614
rect 6222 187378 6306 187614
rect 6542 187378 6574 187614
rect 5954 187294 6574 187378
rect 5954 187058 5986 187294
rect 6222 187058 6306 187294
rect 6542 187058 6574 187294
rect 5954 151614 6574 187058
rect 5954 151378 5986 151614
rect 6222 151378 6306 151614
rect 6542 151378 6574 151614
rect 5954 151294 6574 151378
rect 5954 151058 5986 151294
rect 6222 151058 6306 151294
rect 6542 151058 6574 151294
rect 5954 115614 6574 151058
rect 5954 115378 5986 115614
rect 6222 115378 6306 115614
rect 6542 115378 6574 115614
rect 5954 115294 6574 115378
rect 5954 115058 5986 115294
rect 6222 115058 6306 115294
rect 6542 115058 6574 115294
rect 5954 79614 6574 115058
rect 5954 79378 5986 79614
rect 6222 79378 6306 79614
rect 6542 79378 6574 79614
rect 5954 79294 6574 79378
rect 5954 79058 5986 79294
rect 6222 79058 6306 79294
rect 6542 79058 6574 79294
rect 5954 43614 6574 79058
rect 5954 43378 5986 43614
rect 6222 43378 6306 43614
rect 6542 43378 6574 43614
rect 5954 43294 6574 43378
rect 5954 43058 5986 43294
rect 6222 43058 6306 43294
rect 6542 43058 6574 43294
rect 5954 7614 6574 43058
rect 5954 7378 5986 7614
rect 6222 7378 6306 7614
rect 6542 7378 6574 7614
rect 5954 7294 6574 7378
rect 5954 7058 5986 7294
rect 6222 7058 6306 7294
rect 6542 7058 6574 7294
rect 5954 -4186 6574 7058
rect 5954 -4422 5986 -4186
rect 6222 -4422 6306 -4186
rect 6542 -4422 6574 -4186
rect 5954 -4506 6574 -4422
rect 5954 -4742 5986 -4506
rect 6222 -4742 6306 -4506
rect 6542 -4742 6574 -4506
rect 5954 -7654 6574 -4742
rect 7194 709638 7814 711590
rect 7194 709402 7226 709638
rect 7462 709402 7546 709638
rect 7782 709402 7814 709638
rect 7194 709318 7814 709402
rect 7194 709082 7226 709318
rect 7462 709082 7546 709318
rect 7782 709082 7814 709318
rect 7194 692854 7814 709082
rect 7194 692618 7226 692854
rect 7462 692618 7546 692854
rect 7782 692618 7814 692854
rect 7194 692534 7814 692618
rect 7194 692298 7226 692534
rect 7462 692298 7546 692534
rect 7782 692298 7814 692534
rect 7194 656854 7814 692298
rect 7194 656618 7226 656854
rect 7462 656618 7546 656854
rect 7782 656618 7814 656854
rect 7194 656534 7814 656618
rect 7194 656298 7226 656534
rect 7462 656298 7546 656534
rect 7782 656298 7814 656534
rect 7194 620854 7814 656298
rect 7194 620618 7226 620854
rect 7462 620618 7546 620854
rect 7782 620618 7814 620854
rect 7194 620534 7814 620618
rect 7194 620298 7226 620534
rect 7462 620298 7546 620534
rect 7782 620298 7814 620534
rect 7194 584854 7814 620298
rect 7194 584618 7226 584854
rect 7462 584618 7546 584854
rect 7782 584618 7814 584854
rect 7194 584534 7814 584618
rect 7194 584298 7226 584534
rect 7462 584298 7546 584534
rect 7782 584298 7814 584534
rect 7194 548854 7814 584298
rect 7194 548618 7226 548854
rect 7462 548618 7546 548854
rect 7782 548618 7814 548854
rect 7194 548534 7814 548618
rect 7194 548298 7226 548534
rect 7462 548298 7546 548534
rect 7782 548298 7814 548534
rect 7194 512854 7814 548298
rect 7194 512618 7226 512854
rect 7462 512618 7546 512854
rect 7782 512618 7814 512854
rect 7194 512534 7814 512618
rect 7194 512298 7226 512534
rect 7462 512298 7546 512534
rect 7782 512298 7814 512534
rect 7194 476854 7814 512298
rect 7194 476618 7226 476854
rect 7462 476618 7546 476854
rect 7782 476618 7814 476854
rect 7194 476534 7814 476618
rect 7194 476298 7226 476534
rect 7462 476298 7546 476534
rect 7782 476298 7814 476534
rect 7194 440854 7814 476298
rect 7194 440618 7226 440854
rect 7462 440618 7546 440854
rect 7782 440618 7814 440854
rect 7194 440534 7814 440618
rect 7194 440298 7226 440534
rect 7462 440298 7546 440534
rect 7782 440298 7814 440534
rect 7194 404854 7814 440298
rect 7194 404618 7226 404854
rect 7462 404618 7546 404854
rect 7782 404618 7814 404854
rect 7194 404534 7814 404618
rect 7194 404298 7226 404534
rect 7462 404298 7546 404534
rect 7782 404298 7814 404534
rect 7194 368854 7814 404298
rect 7194 368618 7226 368854
rect 7462 368618 7546 368854
rect 7782 368618 7814 368854
rect 7194 368534 7814 368618
rect 7194 368298 7226 368534
rect 7462 368298 7546 368534
rect 7782 368298 7814 368534
rect 7194 332854 7814 368298
rect 7194 332618 7226 332854
rect 7462 332618 7546 332854
rect 7782 332618 7814 332854
rect 7194 332534 7814 332618
rect 7194 332298 7226 332534
rect 7462 332298 7546 332534
rect 7782 332298 7814 332534
rect 7194 296854 7814 332298
rect 7194 296618 7226 296854
rect 7462 296618 7546 296854
rect 7782 296618 7814 296854
rect 7194 296534 7814 296618
rect 7194 296298 7226 296534
rect 7462 296298 7546 296534
rect 7782 296298 7814 296534
rect 7194 260854 7814 296298
rect 7194 260618 7226 260854
rect 7462 260618 7546 260854
rect 7782 260618 7814 260854
rect 7194 260534 7814 260618
rect 7194 260298 7226 260534
rect 7462 260298 7546 260534
rect 7782 260298 7814 260534
rect 7194 224854 7814 260298
rect 7194 224618 7226 224854
rect 7462 224618 7546 224854
rect 7782 224618 7814 224854
rect 7194 224534 7814 224618
rect 7194 224298 7226 224534
rect 7462 224298 7546 224534
rect 7782 224298 7814 224534
rect 7194 188854 7814 224298
rect 7194 188618 7226 188854
rect 7462 188618 7546 188854
rect 7782 188618 7814 188854
rect 7194 188534 7814 188618
rect 7194 188298 7226 188534
rect 7462 188298 7546 188534
rect 7782 188298 7814 188534
rect 7194 152854 7814 188298
rect 7194 152618 7226 152854
rect 7462 152618 7546 152854
rect 7782 152618 7814 152854
rect 7194 152534 7814 152618
rect 7194 152298 7226 152534
rect 7462 152298 7546 152534
rect 7782 152298 7814 152534
rect 7194 116854 7814 152298
rect 7194 116618 7226 116854
rect 7462 116618 7546 116854
rect 7782 116618 7814 116854
rect 7194 116534 7814 116618
rect 7194 116298 7226 116534
rect 7462 116298 7546 116534
rect 7782 116298 7814 116534
rect 7194 80854 7814 116298
rect 7194 80618 7226 80854
rect 7462 80618 7546 80854
rect 7782 80618 7814 80854
rect 7194 80534 7814 80618
rect 7194 80298 7226 80534
rect 7462 80298 7546 80534
rect 7782 80298 7814 80534
rect 7194 44854 7814 80298
rect 7194 44618 7226 44854
rect 7462 44618 7546 44854
rect 7782 44618 7814 44854
rect 7194 44534 7814 44618
rect 7194 44298 7226 44534
rect 7462 44298 7546 44534
rect 7782 44298 7814 44534
rect 7194 8854 7814 44298
rect 7194 8618 7226 8854
rect 7462 8618 7546 8854
rect 7782 8618 7814 8854
rect 7194 8534 7814 8618
rect 7194 8298 7226 8534
rect 7462 8298 7546 8534
rect 7782 8298 7814 8534
rect 7194 -5146 7814 8298
rect 7194 -5382 7226 -5146
rect 7462 -5382 7546 -5146
rect 7782 -5382 7814 -5146
rect 7194 -5466 7814 -5382
rect 7194 -5702 7226 -5466
rect 7462 -5702 7546 -5466
rect 7782 -5702 7814 -5466
rect 7194 -7654 7814 -5702
rect 8434 710598 9054 711590
rect 8434 710362 8466 710598
rect 8702 710362 8786 710598
rect 9022 710362 9054 710598
rect 8434 710278 9054 710362
rect 8434 710042 8466 710278
rect 8702 710042 8786 710278
rect 9022 710042 9054 710278
rect 8434 694094 9054 710042
rect 8434 693858 8466 694094
rect 8702 693858 8786 694094
rect 9022 693858 9054 694094
rect 8434 693774 9054 693858
rect 8434 693538 8466 693774
rect 8702 693538 8786 693774
rect 9022 693538 9054 693774
rect 8434 658094 9054 693538
rect 8434 657858 8466 658094
rect 8702 657858 8786 658094
rect 9022 657858 9054 658094
rect 8434 657774 9054 657858
rect 8434 657538 8466 657774
rect 8702 657538 8786 657774
rect 9022 657538 9054 657774
rect 8434 622094 9054 657538
rect 8434 621858 8466 622094
rect 8702 621858 8786 622094
rect 9022 621858 9054 622094
rect 8434 621774 9054 621858
rect 8434 621538 8466 621774
rect 8702 621538 8786 621774
rect 9022 621538 9054 621774
rect 8434 586094 9054 621538
rect 8434 585858 8466 586094
rect 8702 585858 8786 586094
rect 9022 585858 9054 586094
rect 8434 585774 9054 585858
rect 8434 585538 8466 585774
rect 8702 585538 8786 585774
rect 9022 585538 9054 585774
rect 8434 550094 9054 585538
rect 8434 549858 8466 550094
rect 8702 549858 8786 550094
rect 9022 549858 9054 550094
rect 8434 549774 9054 549858
rect 8434 549538 8466 549774
rect 8702 549538 8786 549774
rect 9022 549538 9054 549774
rect 8434 514094 9054 549538
rect 8434 513858 8466 514094
rect 8702 513858 8786 514094
rect 9022 513858 9054 514094
rect 8434 513774 9054 513858
rect 8434 513538 8466 513774
rect 8702 513538 8786 513774
rect 9022 513538 9054 513774
rect 8434 478094 9054 513538
rect 8434 477858 8466 478094
rect 8702 477858 8786 478094
rect 9022 477858 9054 478094
rect 8434 477774 9054 477858
rect 8434 477538 8466 477774
rect 8702 477538 8786 477774
rect 9022 477538 9054 477774
rect 8434 442094 9054 477538
rect 8434 441858 8466 442094
rect 8702 441858 8786 442094
rect 9022 441858 9054 442094
rect 8434 441774 9054 441858
rect 8434 441538 8466 441774
rect 8702 441538 8786 441774
rect 9022 441538 9054 441774
rect 8434 406094 9054 441538
rect 8434 405858 8466 406094
rect 8702 405858 8786 406094
rect 9022 405858 9054 406094
rect 8434 405774 9054 405858
rect 8434 405538 8466 405774
rect 8702 405538 8786 405774
rect 9022 405538 9054 405774
rect 8434 370094 9054 405538
rect 8434 369858 8466 370094
rect 8702 369858 8786 370094
rect 9022 369858 9054 370094
rect 8434 369774 9054 369858
rect 8434 369538 8466 369774
rect 8702 369538 8786 369774
rect 9022 369538 9054 369774
rect 8434 334094 9054 369538
rect 8434 333858 8466 334094
rect 8702 333858 8786 334094
rect 9022 333858 9054 334094
rect 8434 333774 9054 333858
rect 8434 333538 8466 333774
rect 8702 333538 8786 333774
rect 9022 333538 9054 333774
rect 8434 298094 9054 333538
rect 8434 297858 8466 298094
rect 8702 297858 8786 298094
rect 9022 297858 9054 298094
rect 8434 297774 9054 297858
rect 8434 297538 8466 297774
rect 8702 297538 8786 297774
rect 9022 297538 9054 297774
rect 8434 262094 9054 297538
rect 8434 261858 8466 262094
rect 8702 261858 8786 262094
rect 9022 261858 9054 262094
rect 8434 261774 9054 261858
rect 8434 261538 8466 261774
rect 8702 261538 8786 261774
rect 9022 261538 9054 261774
rect 8434 226094 9054 261538
rect 8434 225858 8466 226094
rect 8702 225858 8786 226094
rect 9022 225858 9054 226094
rect 8434 225774 9054 225858
rect 8434 225538 8466 225774
rect 8702 225538 8786 225774
rect 9022 225538 9054 225774
rect 8434 190094 9054 225538
rect 8434 189858 8466 190094
rect 8702 189858 8786 190094
rect 9022 189858 9054 190094
rect 8434 189774 9054 189858
rect 8434 189538 8466 189774
rect 8702 189538 8786 189774
rect 9022 189538 9054 189774
rect 8434 154094 9054 189538
rect 8434 153858 8466 154094
rect 8702 153858 8786 154094
rect 9022 153858 9054 154094
rect 8434 153774 9054 153858
rect 8434 153538 8466 153774
rect 8702 153538 8786 153774
rect 9022 153538 9054 153774
rect 8434 118094 9054 153538
rect 8434 117858 8466 118094
rect 8702 117858 8786 118094
rect 9022 117858 9054 118094
rect 8434 117774 9054 117858
rect 8434 117538 8466 117774
rect 8702 117538 8786 117774
rect 9022 117538 9054 117774
rect 8434 82094 9054 117538
rect 8434 81858 8466 82094
rect 8702 81858 8786 82094
rect 9022 81858 9054 82094
rect 8434 81774 9054 81858
rect 8434 81538 8466 81774
rect 8702 81538 8786 81774
rect 9022 81538 9054 81774
rect 8434 46094 9054 81538
rect 8434 45858 8466 46094
rect 8702 45858 8786 46094
rect 9022 45858 9054 46094
rect 8434 45774 9054 45858
rect 8434 45538 8466 45774
rect 8702 45538 8786 45774
rect 9022 45538 9054 45774
rect 8434 10094 9054 45538
rect 8434 9858 8466 10094
rect 8702 9858 8786 10094
rect 9022 9858 9054 10094
rect 8434 9774 9054 9858
rect 8434 9538 8466 9774
rect 8702 9538 8786 9774
rect 9022 9538 9054 9774
rect 8434 -6106 9054 9538
rect 8434 -6342 8466 -6106
rect 8702 -6342 8786 -6106
rect 9022 -6342 9054 -6106
rect 8434 -6426 9054 -6342
rect 8434 -6662 8466 -6426
rect 8702 -6662 8786 -6426
rect 9022 -6662 9054 -6426
rect 8434 -7654 9054 -6662
rect 9674 711558 10294 711590
rect 9674 711322 9706 711558
rect 9942 711322 10026 711558
rect 10262 711322 10294 711558
rect 9674 711238 10294 711322
rect 9674 711002 9706 711238
rect 9942 711002 10026 711238
rect 10262 711002 10294 711238
rect 9674 695334 10294 711002
rect 9674 695098 9706 695334
rect 9942 695098 10026 695334
rect 10262 695098 10294 695334
rect 9674 695014 10294 695098
rect 9674 694778 9706 695014
rect 9942 694778 10026 695014
rect 10262 694778 10294 695014
rect 9674 659334 10294 694778
rect 9674 659098 9706 659334
rect 9942 659098 10026 659334
rect 10262 659098 10294 659334
rect 9674 659014 10294 659098
rect 9674 658778 9706 659014
rect 9942 658778 10026 659014
rect 10262 658778 10294 659014
rect 9674 623334 10294 658778
rect 9674 623098 9706 623334
rect 9942 623098 10026 623334
rect 10262 623098 10294 623334
rect 9674 623014 10294 623098
rect 9674 622778 9706 623014
rect 9942 622778 10026 623014
rect 10262 622778 10294 623014
rect 9674 587334 10294 622778
rect 9674 587098 9706 587334
rect 9942 587098 10026 587334
rect 10262 587098 10294 587334
rect 9674 587014 10294 587098
rect 9674 586778 9706 587014
rect 9942 586778 10026 587014
rect 10262 586778 10294 587014
rect 9674 551334 10294 586778
rect 9674 551098 9706 551334
rect 9942 551098 10026 551334
rect 10262 551098 10294 551334
rect 9674 551014 10294 551098
rect 9674 550778 9706 551014
rect 9942 550778 10026 551014
rect 10262 550778 10294 551014
rect 9674 515334 10294 550778
rect 9674 515098 9706 515334
rect 9942 515098 10026 515334
rect 10262 515098 10294 515334
rect 9674 515014 10294 515098
rect 9674 514778 9706 515014
rect 9942 514778 10026 515014
rect 10262 514778 10294 515014
rect 9674 479334 10294 514778
rect 9674 479098 9706 479334
rect 9942 479098 10026 479334
rect 10262 479098 10294 479334
rect 9674 479014 10294 479098
rect 9674 478778 9706 479014
rect 9942 478778 10026 479014
rect 10262 478778 10294 479014
rect 9674 443334 10294 478778
rect 9674 443098 9706 443334
rect 9942 443098 10026 443334
rect 10262 443098 10294 443334
rect 9674 443014 10294 443098
rect 9674 442778 9706 443014
rect 9942 442778 10026 443014
rect 10262 442778 10294 443014
rect 9674 407334 10294 442778
rect 9674 407098 9706 407334
rect 9942 407098 10026 407334
rect 10262 407098 10294 407334
rect 9674 407014 10294 407098
rect 9674 406778 9706 407014
rect 9942 406778 10026 407014
rect 10262 406778 10294 407014
rect 9674 371334 10294 406778
rect 9674 371098 9706 371334
rect 9942 371098 10026 371334
rect 10262 371098 10294 371334
rect 9674 371014 10294 371098
rect 9674 370778 9706 371014
rect 9942 370778 10026 371014
rect 10262 370778 10294 371014
rect 9674 335334 10294 370778
rect 9674 335098 9706 335334
rect 9942 335098 10026 335334
rect 10262 335098 10294 335334
rect 9674 335014 10294 335098
rect 9674 334778 9706 335014
rect 9942 334778 10026 335014
rect 10262 334778 10294 335014
rect 9674 299334 10294 334778
rect 9674 299098 9706 299334
rect 9942 299098 10026 299334
rect 10262 299098 10294 299334
rect 9674 299014 10294 299098
rect 9674 298778 9706 299014
rect 9942 298778 10026 299014
rect 10262 298778 10294 299014
rect 9674 263334 10294 298778
rect 9674 263098 9706 263334
rect 9942 263098 10026 263334
rect 10262 263098 10294 263334
rect 9674 263014 10294 263098
rect 9674 262778 9706 263014
rect 9942 262778 10026 263014
rect 10262 262778 10294 263014
rect 9674 227334 10294 262778
rect 9674 227098 9706 227334
rect 9942 227098 10026 227334
rect 10262 227098 10294 227334
rect 9674 227014 10294 227098
rect 9674 226778 9706 227014
rect 9942 226778 10026 227014
rect 10262 226778 10294 227014
rect 9674 191334 10294 226778
rect 9674 191098 9706 191334
rect 9942 191098 10026 191334
rect 10262 191098 10294 191334
rect 9674 191014 10294 191098
rect 9674 190778 9706 191014
rect 9942 190778 10026 191014
rect 10262 190778 10294 191014
rect 9674 155334 10294 190778
rect 9674 155098 9706 155334
rect 9942 155098 10026 155334
rect 10262 155098 10294 155334
rect 9674 155014 10294 155098
rect 9674 154778 9706 155014
rect 9942 154778 10026 155014
rect 10262 154778 10294 155014
rect 9674 119334 10294 154778
rect 9674 119098 9706 119334
rect 9942 119098 10026 119334
rect 10262 119098 10294 119334
rect 9674 119014 10294 119098
rect 9674 118778 9706 119014
rect 9942 118778 10026 119014
rect 10262 118778 10294 119014
rect 9674 83334 10294 118778
rect 9674 83098 9706 83334
rect 9942 83098 10026 83334
rect 10262 83098 10294 83334
rect 9674 83014 10294 83098
rect 9674 82778 9706 83014
rect 9942 82778 10026 83014
rect 10262 82778 10294 83014
rect 9674 47334 10294 82778
rect 9674 47098 9706 47334
rect 9942 47098 10026 47334
rect 10262 47098 10294 47334
rect 9674 47014 10294 47098
rect 9674 46778 9706 47014
rect 9942 46778 10026 47014
rect 10262 46778 10294 47014
rect 9674 11334 10294 46778
rect 9674 11098 9706 11334
rect 9942 11098 10026 11334
rect 10262 11098 10294 11334
rect 9674 11014 10294 11098
rect 9674 10778 9706 11014
rect 9942 10778 10026 11014
rect 10262 10778 10294 11014
rect 9674 -7066 10294 10778
rect 9674 -7302 9706 -7066
rect 9942 -7302 10026 -7066
rect 10262 -7302 10294 -7066
rect 9674 -7386 10294 -7302
rect 9674 -7622 9706 -7386
rect 9942 -7622 10026 -7386
rect 10262 -7622 10294 -7386
rect 9674 -7654 10294 -7622
rect 36994 704838 37614 711590
rect 36994 704602 37026 704838
rect 37262 704602 37346 704838
rect 37582 704602 37614 704838
rect 36994 704518 37614 704602
rect 36994 704282 37026 704518
rect 37262 704282 37346 704518
rect 37582 704282 37614 704518
rect 36994 686654 37614 704282
rect 36994 686418 37026 686654
rect 37262 686418 37346 686654
rect 37582 686418 37614 686654
rect 36994 686334 37614 686418
rect 36994 686098 37026 686334
rect 37262 686098 37346 686334
rect 37582 686098 37614 686334
rect 36994 650654 37614 686098
rect 36994 650418 37026 650654
rect 37262 650418 37346 650654
rect 37582 650418 37614 650654
rect 36994 650334 37614 650418
rect 36994 650098 37026 650334
rect 37262 650098 37346 650334
rect 37582 650098 37614 650334
rect 36994 614654 37614 650098
rect 36994 614418 37026 614654
rect 37262 614418 37346 614654
rect 37582 614418 37614 614654
rect 36994 614334 37614 614418
rect 36994 614098 37026 614334
rect 37262 614098 37346 614334
rect 37582 614098 37614 614334
rect 36994 578654 37614 614098
rect 36994 578418 37026 578654
rect 37262 578418 37346 578654
rect 37582 578418 37614 578654
rect 36994 578334 37614 578418
rect 36994 578098 37026 578334
rect 37262 578098 37346 578334
rect 37582 578098 37614 578334
rect 36994 542654 37614 578098
rect 36994 542418 37026 542654
rect 37262 542418 37346 542654
rect 37582 542418 37614 542654
rect 36994 542334 37614 542418
rect 36994 542098 37026 542334
rect 37262 542098 37346 542334
rect 37582 542098 37614 542334
rect 36994 506654 37614 542098
rect 36994 506418 37026 506654
rect 37262 506418 37346 506654
rect 37582 506418 37614 506654
rect 36994 506334 37614 506418
rect 36994 506098 37026 506334
rect 37262 506098 37346 506334
rect 37582 506098 37614 506334
rect 36994 470654 37614 506098
rect 36994 470418 37026 470654
rect 37262 470418 37346 470654
rect 37582 470418 37614 470654
rect 36994 470334 37614 470418
rect 36994 470098 37026 470334
rect 37262 470098 37346 470334
rect 37582 470098 37614 470334
rect 36994 434654 37614 470098
rect 36994 434418 37026 434654
rect 37262 434418 37346 434654
rect 37582 434418 37614 434654
rect 36994 434334 37614 434418
rect 36994 434098 37026 434334
rect 37262 434098 37346 434334
rect 37582 434098 37614 434334
rect 36994 398654 37614 434098
rect 36994 398418 37026 398654
rect 37262 398418 37346 398654
rect 37582 398418 37614 398654
rect 36994 398334 37614 398418
rect 36994 398098 37026 398334
rect 37262 398098 37346 398334
rect 37582 398098 37614 398334
rect 36994 362654 37614 398098
rect 36994 362418 37026 362654
rect 37262 362418 37346 362654
rect 37582 362418 37614 362654
rect 36994 362334 37614 362418
rect 36994 362098 37026 362334
rect 37262 362098 37346 362334
rect 37582 362098 37614 362334
rect 36994 326654 37614 362098
rect 36994 326418 37026 326654
rect 37262 326418 37346 326654
rect 37582 326418 37614 326654
rect 36994 326334 37614 326418
rect 36994 326098 37026 326334
rect 37262 326098 37346 326334
rect 37582 326098 37614 326334
rect 36994 290654 37614 326098
rect 36994 290418 37026 290654
rect 37262 290418 37346 290654
rect 37582 290418 37614 290654
rect 36994 290334 37614 290418
rect 36994 290098 37026 290334
rect 37262 290098 37346 290334
rect 37582 290098 37614 290334
rect 36994 254654 37614 290098
rect 36994 254418 37026 254654
rect 37262 254418 37346 254654
rect 37582 254418 37614 254654
rect 36994 254334 37614 254418
rect 36994 254098 37026 254334
rect 37262 254098 37346 254334
rect 37582 254098 37614 254334
rect 36994 218654 37614 254098
rect 36994 218418 37026 218654
rect 37262 218418 37346 218654
rect 37582 218418 37614 218654
rect 36994 218334 37614 218418
rect 36994 218098 37026 218334
rect 37262 218098 37346 218334
rect 37582 218098 37614 218334
rect 36994 182654 37614 218098
rect 36994 182418 37026 182654
rect 37262 182418 37346 182654
rect 37582 182418 37614 182654
rect 36994 182334 37614 182418
rect 36994 182098 37026 182334
rect 37262 182098 37346 182334
rect 37582 182098 37614 182334
rect 36994 146654 37614 182098
rect 36994 146418 37026 146654
rect 37262 146418 37346 146654
rect 37582 146418 37614 146654
rect 36994 146334 37614 146418
rect 36994 146098 37026 146334
rect 37262 146098 37346 146334
rect 37582 146098 37614 146334
rect 36994 110654 37614 146098
rect 36994 110418 37026 110654
rect 37262 110418 37346 110654
rect 37582 110418 37614 110654
rect 36994 110334 37614 110418
rect 36994 110098 37026 110334
rect 37262 110098 37346 110334
rect 37582 110098 37614 110334
rect 36994 74654 37614 110098
rect 36994 74418 37026 74654
rect 37262 74418 37346 74654
rect 37582 74418 37614 74654
rect 36994 74334 37614 74418
rect 36994 74098 37026 74334
rect 37262 74098 37346 74334
rect 37582 74098 37614 74334
rect 36994 38654 37614 74098
rect 36994 38418 37026 38654
rect 37262 38418 37346 38654
rect 37582 38418 37614 38654
rect 36994 38334 37614 38418
rect 36994 38098 37026 38334
rect 37262 38098 37346 38334
rect 37582 38098 37614 38334
rect 36994 2654 37614 38098
rect 36994 2418 37026 2654
rect 37262 2418 37346 2654
rect 37582 2418 37614 2654
rect 36994 2334 37614 2418
rect 36994 2098 37026 2334
rect 37262 2098 37346 2334
rect 37582 2098 37614 2334
rect 36994 -346 37614 2098
rect 36994 -582 37026 -346
rect 37262 -582 37346 -346
rect 37582 -582 37614 -346
rect 36994 -666 37614 -582
rect 36994 -902 37026 -666
rect 37262 -902 37346 -666
rect 37582 -902 37614 -666
rect 36994 -7654 37614 -902
rect 38234 705798 38854 711590
rect 38234 705562 38266 705798
rect 38502 705562 38586 705798
rect 38822 705562 38854 705798
rect 38234 705478 38854 705562
rect 38234 705242 38266 705478
rect 38502 705242 38586 705478
rect 38822 705242 38854 705478
rect 38234 687894 38854 705242
rect 38234 687658 38266 687894
rect 38502 687658 38586 687894
rect 38822 687658 38854 687894
rect 38234 687574 38854 687658
rect 38234 687338 38266 687574
rect 38502 687338 38586 687574
rect 38822 687338 38854 687574
rect 38234 651894 38854 687338
rect 38234 651658 38266 651894
rect 38502 651658 38586 651894
rect 38822 651658 38854 651894
rect 38234 651574 38854 651658
rect 38234 651338 38266 651574
rect 38502 651338 38586 651574
rect 38822 651338 38854 651574
rect 38234 615894 38854 651338
rect 38234 615658 38266 615894
rect 38502 615658 38586 615894
rect 38822 615658 38854 615894
rect 38234 615574 38854 615658
rect 38234 615338 38266 615574
rect 38502 615338 38586 615574
rect 38822 615338 38854 615574
rect 38234 579894 38854 615338
rect 38234 579658 38266 579894
rect 38502 579658 38586 579894
rect 38822 579658 38854 579894
rect 38234 579574 38854 579658
rect 38234 579338 38266 579574
rect 38502 579338 38586 579574
rect 38822 579338 38854 579574
rect 38234 543894 38854 579338
rect 38234 543658 38266 543894
rect 38502 543658 38586 543894
rect 38822 543658 38854 543894
rect 38234 543574 38854 543658
rect 38234 543338 38266 543574
rect 38502 543338 38586 543574
rect 38822 543338 38854 543574
rect 38234 507894 38854 543338
rect 38234 507658 38266 507894
rect 38502 507658 38586 507894
rect 38822 507658 38854 507894
rect 38234 507574 38854 507658
rect 38234 507338 38266 507574
rect 38502 507338 38586 507574
rect 38822 507338 38854 507574
rect 38234 471894 38854 507338
rect 38234 471658 38266 471894
rect 38502 471658 38586 471894
rect 38822 471658 38854 471894
rect 38234 471574 38854 471658
rect 38234 471338 38266 471574
rect 38502 471338 38586 471574
rect 38822 471338 38854 471574
rect 38234 435894 38854 471338
rect 38234 435658 38266 435894
rect 38502 435658 38586 435894
rect 38822 435658 38854 435894
rect 38234 435574 38854 435658
rect 38234 435338 38266 435574
rect 38502 435338 38586 435574
rect 38822 435338 38854 435574
rect 38234 399894 38854 435338
rect 38234 399658 38266 399894
rect 38502 399658 38586 399894
rect 38822 399658 38854 399894
rect 38234 399574 38854 399658
rect 38234 399338 38266 399574
rect 38502 399338 38586 399574
rect 38822 399338 38854 399574
rect 38234 363894 38854 399338
rect 38234 363658 38266 363894
rect 38502 363658 38586 363894
rect 38822 363658 38854 363894
rect 38234 363574 38854 363658
rect 38234 363338 38266 363574
rect 38502 363338 38586 363574
rect 38822 363338 38854 363574
rect 38234 327894 38854 363338
rect 38234 327658 38266 327894
rect 38502 327658 38586 327894
rect 38822 327658 38854 327894
rect 38234 327574 38854 327658
rect 38234 327338 38266 327574
rect 38502 327338 38586 327574
rect 38822 327338 38854 327574
rect 38234 291894 38854 327338
rect 38234 291658 38266 291894
rect 38502 291658 38586 291894
rect 38822 291658 38854 291894
rect 38234 291574 38854 291658
rect 38234 291338 38266 291574
rect 38502 291338 38586 291574
rect 38822 291338 38854 291574
rect 38234 255894 38854 291338
rect 38234 255658 38266 255894
rect 38502 255658 38586 255894
rect 38822 255658 38854 255894
rect 38234 255574 38854 255658
rect 38234 255338 38266 255574
rect 38502 255338 38586 255574
rect 38822 255338 38854 255574
rect 38234 219894 38854 255338
rect 38234 219658 38266 219894
rect 38502 219658 38586 219894
rect 38822 219658 38854 219894
rect 38234 219574 38854 219658
rect 38234 219338 38266 219574
rect 38502 219338 38586 219574
rect 38822 219338 38854 219574
rect 38234 183894 38854 219338
rect 38234 183658 38266 183894
rect 38502 183658 38586 183894
rect 38822 183658 38854 183894
rect 38234 183574 38854 183658
rect 38234 183338 38266 183574
rect 38502 183338 38586 183574
rect 38822 183338 38854 183574
rect 38234 147894 38854 183338
rect 38234 147658 38266 147894
rect 38502 147658 38586 147894
rect 38822 147658 38854 147894
rect 38234 147574 38854 147658
rect 38234 147338 38266 147574
rect 38502 147338 38586 147574
rect 38822 147338 38854 147574
rect 38234 111894 38854 147338
rect 38234 111658 38266 111894
rect 38502 111658 38586 111894
rect 38822 111658 38854 111894
rect 38234 111574 38854 111658
rect 38234 111338 38266 111574
rect 38502 111338 38586 111574
rect 38822 111338 38854 111574
rect 38234 75894 38854 111338
rect 38234 75658 38266 75894
rect 38502 75658 38586 75894
rect 38822 75658 38854 75894
rect 38234 75574 38854 75658
rect 38234 75338 38266 75574
rect 38502 75338 38586 75574
rect 38822 75338 38854 75574
rect 38234 39894 38854 75338
rect 38234 39658 38266 39894
rect 38502 39658 38586 39894
rect 38822 39658 38854 39894
rect 38234 39574 38854 39658
rect 38234 39338 38266 39574
rect 38502 39338 38586 39574
rect 38822 39338 38854 39574
rect 38234 3894 38854 39338
rect 38234 3658 38266 3894
rect 38502 3658 38586 3894
rect 38822 3658 38854 3894
rect 38234 3574 38854 3658
rect 38234 3338 38266 3574
rect 38502 3338 38586 3574
rect 38822 3338 38854 3574
rect 38234 -1306 38854 3338
rect 38234 -1542 38266 -1306
rect 38502 -1542 38586 -1306
rect 38822 -1542 38854 -1306
rect 38234 -1626 38854 -1542
rect 38234 -1862 38266 -1626
rect 38502 -1862 38586 -1626
rect 38822 -1862 38854 -1626
rect 38234 -7654 38854 -1862
rect 39474 706758 40094 711590
rect 39474 706522 39506 706758
rect 39742 706522 39826 706758
rect 40062 706522 40094 706758
rect 39474 706438 40094 706522
rect 39474 706202 39506 706438
rect 39742 706202 39826 706438
rect 40062 706202 40094 706438
rect 39474 689134 40094 706202
rect 39474 688898 39506 689134
rect 39742 688898 39826 689134
rect 40062 688898 40094 689134
rect 39474 688814 40094 688898
rect 39474 688578 39506 688814
rect 39742 688578 39826 688814
rect 40062 688578 40094 688814
rect 39474 653134 40094 688578
rect 39474 652898 39506 653134
rect 39742 652898 39826 653134
rect 40062 652898 40094 653134
rect 39474 652814 40094 652898
rect 39474 652578 39506 652814
rect 39742 652578 39826 652814
rect 40062 652578 40094 652814
rect 39474 617134 40094 652578
rect 39474 616898 39506 617134
rect 39742 616898 39826 617134
rect 40062 616898 40094 617134
rect 39474 616814 40094 616898
rect 39474 616578 39506 616814
rect 39742 616578 39826 616814
rect 40062 616578 40094 616814
rect 39474 581134 40094 616578
rect 39474 580898 39506 581134
rect 39742 580898 39826 581134
rect 40062 580898 40094 581134
rect 39474 580814 40094 580898
rect 39474 580578 39506 580814
rect 39742 580578 39826 580814
rect 40062 580578 40094 580814
rect 39474 545134 40094 580578
rect 39474 544898 39506 545134
rect 39742 544898 39826 545134
rect 40062 544898 40094 545134
rect 39474 544814 40094 544898
rect 39474 544578 39506 544814
rect 39742 544578 39826 544814
rect 40062 544578 40094 544814
rect 39474 509134 40094 544578
rect 39474 508898 39506 509134
rect 39742 508898 39826 509134
rect 40062 508898 40094 509134
rect 39474 508814 40094 508898
rect 39474 508578 39506 508814
rect 39742 508578 39826 508814
rect 40062 508578 40094 508814
rect 39474 473134 40094 508578
rect 39474 472898 39506 473134
rect 39742 472898 39826 473134
rect 40062 472898 40094 473134
rect 39474 472814 40094 472898
rect 39474 472578 39506 472814
rect 39742 472578 39826 472814
rect 40062 472578 40094 472814
rect 39474 437134 40094 472578
rect 39474 436898 39506 437134
rect 39742 436898 39826 437134
rect 40062 436898 40094 437134
rect 39474 436814 40094 436898
rect 39474 436578 39506 436814
rect 39742 436578 39826 436814
rect 40062 436578 40094 436814
rect 39474 401134 40094 436578
rect 39474 400898 39506 401134
rect 39742 400898 39826 401134
rect 40062 400898 40094 401134
rect 39474 400814 40094 400898
rect 39474 400578 39506 400814
rect 39742 400578 39826 400814
rect 40062 400578 40094 400814
rect 39474 365134 40094 400578
rect 39474 364898 39506 365134
rect 39742 364898 39826 365134
rect 40062 364898 40094 365134
rect 39474 364814 40094 364898
rect 39474 364578 39506 364814
rect 39742 364578 39826 364814
rect 40062 364578 40094 364814
rect 39474 329134 40094 364578
rect 39474 328898 39506 329134
rect 39742 328898 39826 329134
rect 40062 328898 40094 329134
rect 39474 328814 40094 328898
rect 39474 328578 39506 328814
rect 39742 328578 39826 328814
rect 40062 328578 40094 328814
rect 39474 293134 40094 328578
rect 39474 292898 39506 293134
rect 39742 292898 39826 293134
rect 40062 292898 40094 293134
rect 39474 292814 40094 292898
rect 39474 292578 39506 292814
rect 39742 292578 39826 292814
rect 40062 292578 40094 292814
rect 39474 257134 40094 292578
rect 39474 256898 39506 257134
rect 39742 256898 39826 257134
rect 40062 256898 40094 257134
rect 39474 256814 40094 256898
rect 39474 256578 39506 256814
rect 39742 256578 39826 256814
rect 40062 256578 40094 256814
rect 39474 221134 40094 256578
rect 39474 220898 39506 221134
rect 39742 220898 39826 221134
rect 40062 220898 40094 221134
rect 39474 220814 40094 220898
rect 39474 220578 39506 220814
rect 39742 220578 39826 220814
rect 40062 220578 40094 220814
rect 39474 185134 40094 220578
rect 39474 184898 39506 185134
rect 39742 184898 39826 185134
rect 40062 184898 40094 185134
rect 39474 184814 40094 184898
rect 39474 184578 39506 184814
rect 39742 184578 39826 184814
rect 40062 184578 40094 184814
rect 39474 149134 40094 184578
rect 39474 148898 39506 149134
rect 39742 148898 39826 149134
rect 40062 148898 40094 149134
rect 39474 148814 40094 148898
rect 39474 148578 39506 148814
rect 39742 148578 39826 148814
rect 40062 148578 40094 148814
rect 39474 113134 40094 148578
rect 39474 112898 39506 113134
rect 39742 112898 39826 113134
rect 40062 112898 40094 113134
rect 39474 112814 40094 112898
rect 39474 112578 39506 112814
rect 39742 112578 39826 112814
rect 40062 112578 40094 112814
rect 39474 77134 40094 112578
rect 39474 76898 39506 77134
rect 39742 76898 39826 77134
rect 40062 76898 40094 77134
rect 39474 76814 40094 76898
rect 39474 76578 39506 76814
rect 39742 76578 39826 76814
rect 40062 76578 40094 76814
rect 39474 41134 40094 76578
rect 39474 40898 39506 41134
rect 39742 40898 39826 41134
rect 40062 40898 40094 41134
rect 39474 40814 40094 40898
rect 39474 40578 39506 40814
rect 39742 40578 39826 40814
rect 40062 40578 40094 40814
rect 39474 5134 40094 40578
rect 39474 4898 39506 5134
rect 39742 4898 39826 5134
rect 40062 4898 40094 5134
rect 39474 4814 40094 4898
rect 39474 4578 39506 4814
rect 39742 4578 39826 4814
rect 40062 4578 40094 4814
rect 39474 -2266 40094 4578
rect 39474 -2502 39506 -2266
rect 39742 -2502 39826 -2266
rect 40062 -2502 40094 -2266
rect 39474 -2586 40094 -2502
rect 39474 -2822 39506 -2586
rect 39742 -2822 39826 -2586
rect 40062 -2822 40094 -2586
rect 39474 -7654 40094 -2822
rect 40714 707718 41334 711590
rect 40714 707482 40746 707718
rect 40982 707482 41066 707718
rect 41302 707482 41334 707718
rect 40714 707398 41334 707482
rect 40714 707162 40746 707398
rect 40982 707162 41066 707398
rect 41302 707162 41334 707398
rect 40714 690374 41334 707162
rect 40714 690138 40746 690374
rect 40982 690138 41066 690374
rect 41302 690138 41334 690374
rect 40714 690054 41334 690138
rect 40714 689818 40746 690054
rect 40982 689818 41066 690054
rect 41302 689818 41334 690054
rect 40714 654374 41334 689818
rect 40714 654138 40746 654374
rect 40982 654138 41066 654374
rect 41302 654138 41334 654374
rect 40714 654054 41334 654138
rect 40714 653818 40746 654054
rect 40982 653818 41066 654054
rect 41302 653818 41334 654054
rect 40714 618374 41334 653818
rect 40714 618138 40746 618374
rect 40982 618138 41066 618374
rect 41302 618138 41334 618374
rect 40714 618054 41334 618138
rect 40714 617818 40746 618054
rect 40982 617818 41066 618054
rect 41302 617818 41334 618054
rect 40714 582374 41334 617818
rect 40714 582138 40746 582374
rect 40982 582138 41066 582374
rect 41302 582138 41334 582374
rect 40714 582054 41334 582138
rect 40714 581818 40746 582054
rect 40982 581818 41066 582054
rect 41302 581818 41334 582054
rect 40714 546374 41334 581818
rect 40714 546138 40746 546374
rect 40982 546138 41066 546374
rect 41302 546138 41334 546374
rect 40714 546054 41334 546138
rect 40714 545818 40746 546054
rect 40982 545818 41066 546054
rect 41302 545818 41334 546054
rect 40714 510374 41334 545818
rect 40714 510138 40746 510374
rect 40982 510138 41066 510374
rect 41302 510138 41334 510374
rect 40714 510054 41334 510138
rect 40714 509818 40746 510054
rect 40982 509818 41066 510054
rect 41302 509818 41334 510054
rect 40714 474374 41334 509818
rect 40714 474138 40746 474374
rect 40982 474138 41066 474374
rect 41302 474138 41334 474374
rect 40714 474054 41334 474138
rect 40714 473818 40746 474054
rect 40982 473818 41066 474054
rect 41302 473818 41334 474054
rect 40714 438374 41334 473818
rect 40714 438138 40746 438374
rect 40982 438138 41066 438374
rect 41302 438138 41334 438374
rect 40714 438054 41334 438138
rect 40714 437818 40746 438054
rect 40982 437818 41066 438054
rect 41302 437818 41334 438054
rect 40714 402374 41334 437818
rect 40714 402138 40746 402374
rect 40982 402138 41066 402374
rect 41302 402138 41334 402374
rect 40714 402054 41334 402138
rect 40714 401818 40746 402054
rect 40982 401818 41066 402054
rect 41302 401818 41334 402054
rect 40714 366374 41334 401818
rect 40714 366138 40746 366374
rect 40982 366138 41066 366374
rect 41302 366138 41334 366374
rect 40714 366054 41334 366138
rect 40714 365818 40746 366054
rect 40982 365818 41066 366054
rect 41302 365818 41334 366054
rect 40714 330374 41334 365818
rect 40714 330138 40746 330374
rect 40982 330138 41066 330374
rect 41302 330138 41334 330374
rect 40714 330054 41334 330138
rect 40714 329818 40746 330054
rect 40982 329818 41066 330054
rect 41302 329818 41334 330054
rect 40714 294374 41334 329818
rect 40714 294138 40746 294374
rect 40982 294138 41066 294374
rect 41302 294138 41334 294374
rect 40714 294054 41334 294138
rect 40714 293818 40746 294054
rect 40982 293818 41066 294054
rect 41302 293818 41334 294054
rect 40714 258374 41334 293818
rect 40714 258138 40746 258374
rect 40982 258138 41066 258374
rect 41302 258138 41334 258374
rect 40714 258054 41334 258138
rect 40714 257818 40746 258054
rect 40982 257818 41066 258054
rect 41302 257818 41334 258054
rect 40714 222374 41334 257818
rect 40714 222138 40746 222374
rect 40982 222138 41066 222374
rect 41302 222138 41334 222374
rect 40714 222054 41334 222138
rect 40714 221818 40746 222054
rect 40982 221818 41066 222054
rect 41302 221818 41334 222054
rect 40714 186374 41334 221818
rect 40714 186138 40746 186374
rect 40982 186138 41066 186374
rect 41302 186138 41334 186374
rect 40714 186054 41334 186138
rect 40714 185818 40746 186054
rect 40982 185818 41066 186054
rect 41302 185818 41334 186054
rect 40714 150374 41334 185818
rect 40714 150138 40746 150374
rect 40982 150138 41066 150374
rect 41302 150138 41334 150374
rect 40714 150054 41334 150138
rect 40714 149818 40746 150054
rect 40982 149818 41066 150054
rect 41302 149818 41334 150054
rect 40714 114374 41334 149818
rect 40714 114138 40746 114374
rect 40982 114138 41066 114374
rect 41302 114138 41334 114374
rect 40714 114054 41334 114138
rect 40714 113818 40746 114054
rect 40982 113818 41066 114054
rect 41302 113818 41334 114054
rect 40714 78374 41334 113818
rect 40714 78138 40746 78374
rect 40982 78138 41066 78374
rect 41302 78138 41334 78374
rect 40714 78054 41334 78138
rect 40714 77818 40746 78054
rect 40982 77818 41066 78054
rect 41302 77818 41334 78054
rect 40714 42374 41334 77818
rect 40714 42138 40746 42374
rect 40982 42138 41066 42374
rect 41302 42138 41334 42374
rect 40714 42054 41334 42138
rect 40714 41818 40746 42054
rect 40982 41818 41066 42054
rect 41302 41818 41334 42054
rect 40714 6374 41334 41818
rect 40714 6138 40746 6374
rect 40982 6138 41066 6374
rect 41302 6138 41334 6374
rect 40714 6054 41334 6138
rect 40714 5818 40746 6054
rect 40982 5818 41066 6054
rect 41302 5818 41334 6054
rect 40714 -3226 41334 5818
rect 40714 -3462 40746 -3226
rect 40982 -3462 41066 -3226
rect 41302 -3462 41334 -3226
rect 40714 -3546 41334 -3462
rect 40714 -3782 40746 -3546
rect 40982 -3782 41066 -3546
rect 41302 -3782 41334 -3546
rect 40714 -7654 41334 -3782
rect 41954 708678 42574 711590
rect 41954 708442 41986 708678
rect 42222 708442 42306 708678
rect 42542 708442 42574 708678
rect 41954 708358 42574 708442
rect 41954 708122 41986 708358
rect 42222 708122 42306 708358
rect 42542 708122 42574 708358
rect 41954 691614 42574 708122
rect 41954 691378 41986 691614
rect 42222 691378 42306 691614
rect 42542 691378 42574 691614
rect 41954 691294 42574 691378
rect 41954 691058 41986 691294
rect 42222 691058 42306 691294
rect 42542 691058 42574 691294
rect 41954 655614 42574 691058
rect 41954 655378 41986 655614
rect 42222 655378 42306 655614
rect 42542 655378 42574 655614
rect 41954 655294 42574 655378
rect 41954 655058 41986 655294
rect 42222 655058 42306 655294
rect 42542 655058 42574 655294
rect 41954 619614 42574 655058
rect 41954 619378 41986 619614
rect 42222 619378 42306 619614
rect 42542 619378 42574 619614
rect 41954 619294 42574 619378
rect 41954 619058 41986 619294
rect 42222 619058 42306 619294
rect 42542 619058 42574 619294
rect 41954 583614 42574 619058
rect 41954 583378 41986 583614
rect 42222 583378 42306 583614
rect 42542 583378 42574 583614
rect 41954 583294 42574 583378
rect 41954 583058 41986 583294
rect 42222 583058 42306 583294
rect 42542 583058 42574 583294
rect 41954 547614 42574 583058
rect 41954 547378 41986 547614
rect 42222 547378 42306 547614
rect 42542 547378 42574 547614
rect 41954 547294 42574 547378
rect 41954 547058 41986 547294
rect 42222 547058 42306 547294
rect 42542 547058 42574 547294
rect 41954 511614 42574 547058
rect 41954 511378 41986 511614
rect 42222 511378 42306 511614
rect 42542 511378 42574 511614
rect 41954 511294 42574 511378
rect 41954 511058 41986 511294
rect 42222 511058 42306 511294
rect 42542 511058 42574 511294
rect 41954 475614 42574 511058
rect 41954 475378 41986 475614
rect 42222 475378 42306 475614
rect 42542 475378 42574 475614
rect 41954 475294 42574 475378
rect 41954 475058 41986 475294
rect 42222 475058 42306 475294
rect 42542 475058 42574 475294
rect 41954 439614 42574 475058
rect 41954 439378 41986 439614
rect 42222 439378 42306 439614
rect 42542 439378 42574 439614
rect 41954 439294 42574 439378
rect 41954 439058 41986 439294
rect 42222 439058 42306 439294
rect 42542 439058 42574 439294
rect 41954 403614 42574 439058
rect 41954 403378 41986 403614
rect 42222 403378 42306 403614
rect 42542 403378 42574 403614
rect 41954 403294 42574 403378
rect 41954 403058 41986 403294
rect 42222 403058 42306 403294
rect 42542 403058 42574 403294
rect 41954 367614 42574 403058
rect 41954 367378 41986 367614
rect 42222 367378 42306 367614
rect 42542 367378 42574 367614
rect 41954 367294 42574 367378
rect 41954 367058 41986 367294
rect 42222 367058 42306 367294
rect 42542 367058 42574 367294
rect 41954 331614 42574 367058
rect 41954 331378 41986 331614
rect 42222 331378 42306 331614
rect 42542 331378 42574 331614
rect 41954 331294 42574 331378
rect 41954 331058 41986 331294
rect 42222 331058 42306 331294
rect 42542 331058 42574 331294
rect 41954 295614 42574 331058
rect 41954 295378 41986 295614
rect 42222 295378 42306 295614
rect 42542 295378 42574 295614
rect 41954 295294 42574 295378
rect 41954 295058 41986 295294
rect 42222 295058 42306 295294
rect 42542 295058 42574 295294
rect 41954 259614 42574 295058
rect 41954 259378 41986 259614
rect 42222 259378 42306 259614
rect 42542 259378 42574 259614
rect 41954 259294 42574 259378
rect 41954 259058 41986 259294
rect 42222 259058 42306 259294
rect 42542 259058 42574 259294
rect 41954 223614 42574 259058
rect 41954 223378 41986 223614
rect 42222 223378 42306 223614
rect 42542 223378 42574 223614
rect 41954 223294 42574 223378
rect 41954 223058 41986 223294
rect 42222 223058 42306 223294
rect 42542 223058 42574 223294
rect 41954 187614 42574 223058
rect 41954 187378 41986 187614
rect 42222 187378 42306 187614
rect 42542 187378 42574 187614
rect 41954 187294 42574 187378
rect 41954 187058 41986 187294
rect 42222 187058 42306 187294
rect 42542 187058 42574 187294
rect 41954 151614 42574 187058
rect 41954 151378 41986 151614
rect 42222 151378 42306 151614
rect 42542 151378 42574 151614
rect 41954 151294 42574 151378
rect 41954 151058 41986 151294
rect 42222 151058 42306 151294
rect 42542 151058 42574 151294
rect 41954 115614 42574 151058
rect 41954 115378 41986 115614
rect 42222 115378 42306 115614
rect 42542 115378 42574 115614
rect 41954 115294 42574 115378
rect 41954 115058 41986 115294
rect 42222 115058 42306 115294
rect 42542 115058 42574 115294
rect 41954 79614 42574 115058
rect 41954 79378 41986 79614
rect 42222 79378 42306 79614
rect 42542 79378 42574 79614
rect 41954 79294 42574 79378
rect 41954 79058 41986 79294
rect 42222 79058 42306 79294
rect 42542 79058 42574 79294
rect 41954 43614 42574 79058
rect 41954 43378 41986 43614
rect 42222 43378 42306 43614
rect 42542 43378 42574 43614
rect 41954 43294 42574 43378
rect 41954 43058 41986 43294
rect 42222 43058 42306 43294
rect 42542 43058 42574 43294
rect 41954 7614 42574 43058
rect 41954 7378 41986 7614
rect 42222 7378 42306 7614
rect 42542 7378 42574 7614
rect 41954 7294 42574 7378
rect 41954 7058 41986 7294
rect 42222 7058 42306 7294
rect 42542 7058 42574 7294
rect 41954 -4186 42574 7058
rect 41954 -4422 41986 -4186
rect 42222 -4422 42306 -4186
rect 42542 -4422 42574 -4186
rect 41954 -4506 42574 -4422
rect 41954 -4742 41986 -4506
rect 42222 -4742 42306 -4506
rect 42542 -4742 42574 -4506
rect 41954 -7654 42574 -4742
rect 43194 709638 43814 711590
rect 43194 709402 43226 709638
rect 43462 709402 43546 709638
rect 43782 709402 43814 709638
rect 43194 709318 43814 709402
rect 43194 709082 43226 709318
rect 43462 709082 43546 709318
rect 43782 709082 43814 709318
rect 43194 692854 43814 709082
rect 43194 692618 43226 692854
rect 43462 692618 43546 692854
rect 43782 692618 43814 692854
rect 43194 692534 43814 692618
rect 43194 692298 43226 692534
rect 43462 692298 43546 692534
rect 43782 692298 43814 692534
rect 43194 656854 43814 692298
rect 43194 656618 43226 656854
rect 43462 656618 43546 656854
rect 43782 656618 43814 656854
rect 43194 656534 43814 656618
rect 43194 656298 43226 656534
rect 43462 656298 43546 656534
rect 43782 656298 43814 656534
rect 43194 620854 43814 656298
rect 43194 620618 43226 620854
rect 43462 620618 43546 620854
rect 43782 620618 43814 620854
rect 43194 620534 43814 620618
rect 43194 620298 43226 620534
rect 43462 620298 43546 620534
rect 43782 620298 43814 620534
rect 43194 584854 43814 620298
rect 43194 584618 43226 584854
rect 43462 584618 43546 584854
rect 43782 584618 43814 584854
rect 43194 584534 43814 584618
rect 43194 584298 43226 584534
rect 43462 584298 43546 584534
rect 43782 584298 43814 584534
rect 43194 548854 43814 584298
rect 43194 548618 43226 548854
rect 43462 548618 43546 548854
rect 43782 548618 43814 548854
rect 43194 548534 43814 548618
rect 43194 548298 43226 548534
rect 43462 548298 43546 548534
rect 43782 548298 43814 548534
rect 43194 512854 43814 548298
rect 43194 512618 43226 512854
rect 43462 512618 43546 512854
rect 43782 512618 43814 512854
rect 43194 512534 43814 512618
rect 43194 512298 43226 512534
rect 43462 512298 43546 512534
rect 43782 512298 43814 512534
rect 43194 476854 43814 512298
rect 43194 476618 43226 476854
rect 43462 476618 43546 476854
rect 43782 476618 43814 476854
rect 43194 476534 43814 476618
rect 43194 476298 43226 476534
rect 43462 476298 43546 476534
rect 43782 476298 43814 476534
rect 43194 440854 43814 476298
rect 43194 440618 43226 440854
rect 43462 440618 43546 440854
rect 43782 440618 43814 440854
rect 43194 440534 43814 440618
rect 43194 440298 43226 440534
rect 43462 440298 43546 440534
rect 43782 440298 43814 440534
rect 43194 404854 43814 440298
rect 43194 404618 43226 404854
rect 43462 404618 43546 404854
rect 43782 404618 43814 404854
rect 43194 404534 43814 404618
rect 43194 404298 43226 404534
rect 43462 404298 43546 404534
rect 43782 404298 43814 404534
rect 43194 368854 43814 404298
rect 43194 368618 43226 368854
rect 43462 368618 43546 368854
rect 43782 368618 43814 368854
rect 43194 368534 43814 368618
rect 43194 368298 43226 368534
rect 43462 368298 43546 368534
rect 43782 368298 43814 368534
rect 43194 332854 43814 368298
rect 43194 332618 43226 332854
rect 43462 332618 43546 332854
rect 43782 332618 43814 332854
rect 43194 332534 43814 332618
rect 43194 332298 43226 332534
rect 43462 332298 43546 332534
rect 43782 332298 43814 332534
rect 43194 296854 43814 332298
rect 43194 296618 43226 296854
rect 43462 296618 43546 296854
rect 43782 296618 43814 296854
rect 43194 296534 43814 296618
rect 43194 296298 43226 296534
rect 43462 296298 43546 296534
rect 43782 296298 43814 296534
rect 43194 260854 43814 296298
rect 43194 260618 43226 260854
rect 43462 260618 43546 260854
rect 43782 260618 43814 260854
rect 43194 260534 43814 260618
rect 43194 260298 43226 260534
rect 43462 260298 43546 260534
rect 43782 260298 43814 260534
rect 43194 224854 43814 260298
rect 43194 224618 43226 224854
rect 43462 224618 43546 224854
rect 43782 224618 43814 224854
rect 43194 224534 43814 224618
rect 43194 224298 43226 224534
rect 43462 224298 43546 224534
rect 43782 224298 43814 224534
rect 43194 188854 43814 224298
rect 43194 188618 43226 188854
rect 43462 188618 43546 188854
rect 43782 188618 43814 188854
rect 43194 188534 43814 188618
rect 43194 188298 43226 188534
rect 43462 188298 43546 188534
rect 43782 188298 43814 188534
rect 43194 152854 43814 188298
rect 43194 152618 43226 152854
rect 43462 152618 43546 152854
rect 43782 152618 43814 152854
rect 43194 152534 43814 152618
rect 43194 152298 43226 152534
rect 43462 152298 43546 152534
rect 43782 152298 43814 152534
rect 43194 116854 43814 152298
rect 43194 116618 43226 116854
rect 43462 116618 43546 116854
rect 43782 116618 43814 116854
rect 43194 116534 43814 116618
rect 43194 116298 43226 116534
rect 43462 116298 43546 116534
rect 43782 116298 43814 116534
rect 43194 80854 43814 116298
rect 43194 80618 43226 80854
rect 43462 80618 43546 80854
rect 43782 80618 43814 80854
rect 43194 80534 43814 80618
rect 43194 80298 43226 80534
rect 43462 80298 43546 80534
rect 43782 80298 43814 80534
rect 43194 44854 43814 80298
rect 43194 44618 43226 44854
rect 43462 44618 43546 44854
rect 43782 44618 43814 44854
rect 43194 44534 43814 44618
rect 43194 44298 43226 44534
rect 43462 44298 43546 44534
rect 43782 44298 43814 44534
rect 43194 8854 43814 44298
rect 43194 8618 43226 8854
rect 43462 8618 43546 8854
rect 43782 8618 43814 8854
rect 43194 8534 43814 8618
rect 43194 8298 43226 8534
rect 43462 8298 43546 8534
rect 43782 8298 43814 8534
rect 43194 -5146 43814 8298
rect 43194 -5382 43226 -5146
rect 43462 -5382 43546 -5146
rect 43782 -5382 43814 -5146
rect 43194 -5466 43814 -5382
rect 43194 -5702 43226 -5466
rect 43462 -5702 43546 -5466
rect 43782 -5702 43814 -5466
rect 43194 -7654 43814 -5702
rect 44434 710598 45054 711590
rect 44434 710362 44466 710598
rect 44702 710362 44786 710598
rect 45022 710362 45054 710598
rect 44434 710278 45054 710362
rect 44434 710042 44466 710278
rect 44702 710042 44786 710278
rect 45022 710042 45054 710278
rect 44434 694094 45054 710042
rect 44434 693858 44466 694094
rect 44702 693858 44786 694094
rect 45022 693858 45054 694094
rect 44434 693774 45054 693858
rect 44434 693538 44466 693774
rect 44702 693538 44786 693774
rect 45022 693538 45054 693774
rect 44434 658094 45054 693538
rect 44434 657858 44466 658094
rect 44702 657858 44786 658094
rect 45022 657858 45054 658094
rect 44434 657774 45054 657858
rect 44434 657538 44466 657774
rect 44702 657538 44786 657774
rect 45022 657538 45054 657774
rect 44434 622094 45054 657538
rect 44434 621858 44466 622094
rect 44702 621858 44786 622094
rect 45022 621858 45054 622094
rect 44434 621774 45054 621858
rect 44434 621538 44466 621774
rect 44702 621538 44786 621774
rect 45022 621538 45054 621774
rect 44434 586094 45054 621538
rect 44434 585858 44466 586094
rect 44702 585858 44786 586094
rect 45022 585858 45054 586094
rect 44434 585774 45054 585858
rect 44434 585538 44466 585774
rect 44702 585538 44786 585774
rect 45022 585538 45054 585774
rect 44434 550094 45054 585538
rect 44434 549858 44466 550094
rect 44702 549858 44786 550094
rect 45022 549858 45054 550094
rect 44434 549774 45054 549858
rect 44434 549538 44466 549774
rect 44702 549538 44786 549774
rect 45022 549538 45054 549774
rect 44434 514094 45054 549538
rect 44434 513858 44466 514094
rect 44702 513858 44786 514094
rect 45022 513858 45054 514094
rect 44434 513774 45054 513858
rect 44434 513538 44466 513774
rect 44702 513538 44786 513774
rect 45022 513538 45054 513774
rect 44434 478094 45054 513538
rect 44434 477858 44466 478094
rect 44702 477858 44786 478094
rect 45022 477858 45054 478094
rect 44434 477774 45054 477858
rect 44434 477538 44466 477774
rect 44702 477538 44786 477774
rect 45022 477538 45054 477774
rect 44434 442094 45054 477538
rect 44434 441858 44466 442094
rect 44702 441858 44786 442094
rect 45022 441858 45054 442094
rect 44434 441774 45054 441858
rect 44434 441538 44466 441774
rect 44702 441538 44786 441774
rect 45022 441538 45054 441774
rect 44434 406094 45054 441538
rect 44434 405858 44466 406094
rect 44702 405858 44786 406094
rect 45022 405858 45054 406094
rect 44434 405774 45054 405858
rect 44434 405538 44466 405774
rect 44702 405538 44786 405774
rect 45022 405538 45054 405774
rect 44434 370094 45054 405538
rect 44434 369858 44466 370094
rect 44702 369858 44786 370094
rect 45022 369858 45054 370094
rect 44434 369774 45054 369858
rect 44434 369538 44466 369774
rect 44702 369538 44786 369774
rect 45022 369538 45054 369774
rect 44434 334094 45054 369538
rect 44434 333858 44466 334094
rect 44702 333858 44786 334094
rect 45022 333858 45054 334094
rect 44434 333774 45054 333858
rect 44434 333538 44466 333774
rect 44702 333538 44786 333774
rect 45022 333538 45054 333774
rect 44434 298094 45054 333538
rect 44434 297858 44466 298094
rect 44702 297858 44786 298094
rect 45022 297858 45054 298094
rect 44434 297774 45054 297858
rect 44434 297538 44466 297774
rect 44702 297538 44786 297774
rect 45022 297538 45054 297774
rect 44434 262094 45054 297538
rect 44434 261858 44466 262094
rect 44702 261858 44786 262094
rect 45022 261858 45054 262094
rect 44434 261774 45054 261858
rect 44434 261538 44466 261774
rect 44702 261538 44786 261774
rect 45022 261538 45054 261774
rect 44434 226094 45054 261538
rect 44434 225858 44466 226094
rect 44702 225858 44786 226094
rect 45022 225858 45054 226094
rect 44434 225774 45054 225858
rect 44434 225538 44466 225774
rect 44702 225538 44786 225774
rect 45022 225538 45054 225774
rect 44434 190094 45054 225538
rect 44434 189858 44466 190094
rect 44702 189858 44786 190094
rect 45022 189858 45054 190094
rect 44434 189774 45054 189858
rect 44434 189538 44466 189774
rect 44702 189538 44786 189774
rect 45022 189538 45054 189774
rect 44434 154094 45054 189538
rect 44434 153858 44466 154094
rect 44702 153858 44786 154094
rect 45022 153858 45054 154094
rect 44434 153774 45054 153858
rect 44434 153538 44466 153774
rect 44702 153538 44786 153774
rect 45022 153538 45054 153774
rect 44434 118094 45054 153538
rect 44434 117858 44466 118094
rect 44702 117858 44786 118094
rect 45022 117858 45054 118094
rect 44434 117774 45054 117858
rect 44434 117538 44466 117774
rect 44702 117538 44786 117774
rect 45022 117538 45054 117774
rect 44434 82094 45054 117538
rect 44434 81858 44466 82094
rect 44702 81858 44786 82094
rect 45022 81858 45054 82094
rect 44434 81774 45054 81858
rect 44434 81538 44466 81774
rect 44702 81538 44786 81774
rect 45022 81538 45054 81774
rect 44434 46094 45054 81538
rect 44434 45858 44466 46094
rect 44702 45858 44786 46094
rect 45022 45858 45054 46094
rect 44434 45774 45054 45858
rect 44434 45538 44466 45774
rect 44702 45538 44786 45774
rect 45022 45538 45054 45774
rect 44434 10094 45054 45538
rect 44434 9858 44466 10094
rect 44702 9858 44786 10094
rect 45022 9858 45054 10094
rect 44434 9774 45054 9858
rect 44434 9538 44466 9774
rect 44702 9538 44786 9774
rect 45022 9538 45054 9774
rect 44434 -6106 45054 9538
rect 44434 -6342 44466 -6106
rect 44702 -6342 44786 -6106
rect 45022 -6342 45054 -6106
rect 44434 -6426 45054 -6342
rect 44434 -6662 44466 -6426
rect 44702 -6662 44786 -6426
rect 45022 -6662 45054 -6426
rect 44434 -7654 45054 -6662
rect 45674 711558 46294 711590
rect 45674 711322 45706 711558
rect 45942 711322 46026 711558
rect 46262 711322 46294 711558
rect 45674 711238 46294 711322
rect 45674 711002 45706 711238
rect 45942 711002 46026 711238
rect 46262 711002 46294 711238
rect 45674 695334 46294 711002
rect 45674 695098 45706 695334
rect 45942 695098 46026 695334
rect 46262 695098 46294 695334
rect 45674 695014 46294 695098
rect 45674 694778 45706 695014
rect 45942 694778 46026 695014
rect 46262 694778 46294 695014
rect 45674 659334 46294 694778
rect 45674 659098 45706 659334
rect 45942 659098 46026 659334
rect 46262 659098 46294 659334
rect 45674 659014 46294 659098
rect 45674 658778 45706 659014
rect 45942 658778 46026 659014
rect 46262 658778 46294 659014
rect 45674 623334 46294 658778
rect 45674 623098 45706 623334
rect 45942 623098 46026 623334
rect 46262 623098 46294 623334
rect 45674 623014 46294 623098
rect 45674 622778 45706 623014
rect 45942 622778 46026 623014
rect 46262 622778 46294 623014
rect 45674 587334 46294 622778
rect 45674 587098 45706 587334
rect 45942 587098 46026 587334
rect 46262 587098 46294 587334
rect 45674 587014 46294 587098
rect 45674 586778 45706 587014
rect 45942 586778 46026 587014
rect 46262 586778 46294 587014
rect 45674 551334 46294 586778
rect 45674 551098 45706 551334
rect 45942 551098 46026 551334
rect 46262 551098 46294 551334
rect 45674 551014 46294 551098
rect 45674 550778 45706 551014
rect 45942 550778 46026 551014
rect 46262 550778 46294 551014
rect 45674 515334 46294 550778
rect 45674 515098 45706 515334
rect 45942 515098 46026 515334
rect 46262 515098 46294 515334
rect 45674 515014 46294 515098
rect 45674 514778 45706 515014
rect 45942 514778 46026 515014
rect 46262 514778 46294 515014
rect 45674 479334 46294 514778
rect 45674 479098 45706 479334
rect 45942 479098 46026 479334
rect 46262 479098 46294 479334
rect 45674 479014 46294 479098
rect 45674 478778 45706 479014
rect 45942 478778 46026 479014
rect 46262 478778 46294 479014
rect 45674 443334 46294 478778
rect 45674 443098 45706 443334
rect 45942 443098 46026 443334
rect 46262 443098 46294 443334
rect 45674 443014 46294 443098
rect 45674 442778 45706 443014
rect 45942 442778 46026 443014
rect 46262 442778 46294 443014
rect 45674 407334 46294 442778
rect 45674 407098 45706 407334
rect 45942 407098 46026 407334
rect 46262 407098 46294 407334
rect 45674 407014 46294 407098
rect 45674 406778 45706 407014
rect 45942 406778 46026 407014
rect 46262 406778 46294 407014
rect 45674 371334 46294 406778
rect 45674 371098 45706 371334
rect 45942 371098 46026 371334
rect 46262 371098 46294 371334
rect 45674 371014 46294 371098
rect 45674 370778 45706 371014
rect 45942 370778 46026 371014
rect 46262 370778 46294 371014
rect 45674 335334 46294 370778
rect 45674 335098 45706 335334
rect 45942 335098 46026 335334
rect 46262 335098 46294 335334
rect 45674 335014 46294 335098
rect 45674 334778 45706 335014
rect 45942 334778 46026 335014
rect 46262 334778 46294 335014
rect 45674 299334 46294 334778
rect 45674 299098 45706 299334
rect 45942 299098 46026 299334
rect 46262 299098 46294 299334
rect 45674 299014 46294 299098
rect 45674 298778 45706 299014
rect 45942 298778 46026 299014
rect 46262 298778 46294 299014
rect 45674 263334 46294 298778
rect 45674 263098 45706 263334
rect 45942 263098 46026 263334
rect 46262 263098 46294 263334
rect 45674 263014 46294 263098
rect 45674 262778 45706 263014
rect 45942 262778 46026 263014
rect 46262 262778 46294 263014
rect 45674 227334 46294 262778
rect 45674 227098 45706 227334
rect 45942 227098 46026 227334
rect 46262 227098 46294 227334
rect 45674 227014 46294 227098
rect 45674 226778 45706 227014
rect 45942 226778 46026 227014
rect 46262 226778 46294 227014
rect 45674 191334 46294 226778
rect 45674 191098 45706 191334
rect 45942 191098 46026 191334
rect 46262 191098 46294 191334
rect 45674 191014 46294 191098
rect 45674 190778 45706 191014
rect 45942 190778 46026 191014
rect 46262 190778 46294 191014
rect 45674 155334 46294 190778
rect 45674 155098 45706 155334
rect 45942 155098 46026 155334
rect 46262 155098 46294 155334
rect 45674 155014 46294 155098
rect 45674 154778 45706 155014
rect 45942 154778 46026 155014
rect 46262 154778 46294 155014
rect 45674 119334 46294 154778
rect 45674 119098 45706 119334
rect 45942 119098 46026 119334
rect 46262 119098 46294 119334
rect 45674 119014 46294 119098
rect 45674 118778 45706 119014
rect 45942 118778 46026 119014
rect 46262 118778 46294 119014
rect 45674 83334 46294 118778
rect 45674 83098 45706 83334
rect 45942 83098 46026 83334
rect 46262 83098 46294 83334
rect 45674 83014 46294 83098
rect 45674 82778 45706 83014
rect 45942 82778 46026 83014
rect 46262 82778 46294 83014
rect 45674 47334 46294 82778
rect 45674 47098 45706 47334
rect 45942 47098 46026 47334
rect 46262 47098 46294 47334
rect 45674 47014 46294 47098
rect 45674 46778 45706 47014
rect 45942 46778 46026 47014
rect 46262 46778 46294 47014
rect 45674 11334 46294 46778
rect 45674 11098 45706 11334
rect 45942 11098 46026 11334
rect 46262 11098 46294 11334
rect 45674 11014 46294 11098
rect 45674 10778 45706 11014
rect 45942 10778 46026 11014
rect 46262 10778 46294 11014
rect 45674 -7066 46294 10778
rect 45674 -7302 45706 -7066
rect 45942 -7302 46026 -7066
rect 46262 -7302 46294 -7066
rect 45674 -7386 46294 -7302
rect 45674 -7622 45706 -7386
rect 45942 -7622 46026 -7386
rect 46262 -7622 46294 -7386
rect 45674 -7654 46294 -7622
rect 72994 704838 73614 711590
rect 72994 704602 73026 704838
rect 73262 704602 73346 704838
rect 73582 704602 73614 704838
rect 72994 704518 73614 704602
rect 72994 704282 73026 704518
rect 73262 704282 73346 704518
rect 73582 704282 73614 704518
rect 72994 686654 73614 704282
rect 72994 686418 73026 686654
rect 73262 686418 73346 686654
rect 73582 686418 73614 686654
rect 72994 686334 73614 686418
rect 72994 686098 73026 686334
rect 73262 686098 73346 686334
rect 73582 686098 73614 686334
rect 72994 650654 73614 686098
rect 72994 650418 73026 650654
rect 73262 650418 73346 650654
rect 73582 650418 73614 650654
rect 72994 650334 73614 650418
rect 72994 650098 73026 650334
rect 73262 650098 73346 650334
rect 73582 650098 73614 650334
rect 72994 614654 73614 650098
rect 72994 614418 73026 614654
rect 73262 614418 73346 614654
rect 73582 614418 73614 614654
rect 72994 614334 73614 614418
rect 72994 614098 73026 614334
rect 73262 614098 73346 614334
rect 73582 614098 73614 614334
rect 72994 578654 73614 614098
rect 72994 578418 73026 578654
rect 73262 578418 73346 578654
rect 73582 578418 73614 578654
rect 72994 578334 73614 578418
rect 72994 578098 73026 578334
rect 73262 578098 73346 578334
rect 73582 578098 73614 578334
rect 72994 542654 73614 578098
rect 72994 542418 73026 542654
rect 73262 542418 73346 542654
rect 73582 542418 73614 542654
rect 72994 542334 73614 542418
rect 72994 542098 73026 542334
rect 73262 542098 73346 542334
rect 73582 542098 73614 542334
rect 72994 506654 73614 542098
rect 72994 506418 73026 506654
rect 73262 506418 73346 506654
rect 73582 506418 73614 506654
rect 72994 506334 73614 506418
rect 72994 506098 73026 506334
rect 73262 506098 73346 506334
rect 73582 506098 73614 506334
rect 72994 470654 73614 506098
rect 72994 470418 73026 470654
rect 73262 470418 73346 470654
rect 73582 470418 73614 470654
rect 72994 470334 73614 470418
rect 72994 470098 73026 470334
rect 73262 470098 73346 470334
rect 73582 470098 73614 470334
rect 72994 434654 73614 470098
rect 72994 434418 73026 434654
rect 73262 434418 73346 434654
rect 73582 434418 73614 434654
rect 72994 434334 73614 434418
rect 72994 434098 73026 434334
rect 73262 434098 73346 434334
rect 73582 434098 73614 434334
rect 72994 398654 73614 434098
rect 72994 398418 73026 398654
rect 73262 398418 73346 398654
rect 73582 398418 73614 398654
rect 72994 398334 73614 398418
rect 72994 398098 73026 398334
rect 73262 398098 73346 398334
rect 73582 398098 73614 398334
rect 72994 362654 73614 398098
rect 72994 362418 73026 362654
rect 73262 362418 73346 362654
rect 73582 362418 73614 362654
rect 72994 362334 73614 362418
rect 72994 362098 73026 362334
rect 73262 362098 73346 362334
rect 73582 362098 73614 362334
rect 72994 326654 73614 362098
rect 72994 326418 73026 326654
rect 73262 326418 73346 326654
rect 73582 326418 73614 326654
rect 72994 326334 73614 326418
rect 72994 326098 73026 326334
rect 73262 326098 73346 326334
rect 73582 326098 73614 326334
rect 72994 290654 73614 326098
rect 72994 290418 73026 290654
rect 73262 290418 73346 290654
rect 73582 290418 73614 290654
rect 72994 290334 73614 290418
rect 72994 290098 73026 290334
rect 73262 290098 73346 290334
rect 73582 290098 73614 290334
rect 72994 254654 73614 290098
rect 72994 254418 73026 254654
rect 73262 254418 73346 254654
rect 73582 254418 73614 254654
rect 72994 254334 73614 254418
rect 72994 254098 73026 254334
rect 73262 254098 73346 254334
rect 73582 254098 73614 254334
rect 72994 218654 73614 254098
rect 72994 218418 73026 218654
rect 73262 218418 73346 218654
rect 73582 218418 73614 218654
rect 72994 218334 73614 218418
rect 72994 218098 73026 218334
rect 73262 218098 73346 218334
rect 73582 218098 73614 218334
rect 72994 182654 73614 218098
rect 72994 182418 73026 182654
rect 73262 182418 73346 182654
rect 73582 182418 73614 182654
rect 72994 182334 73614 182418
rect 72994 182098 73026 182334
rect 73262 182098 73346 182334
rect 73582 182098 73614 182334
rect 72994 146654 73614 182098
rect 72994 146418 73026 146654
rect 73262 146418 73346 146654
rect 73582 146418 73614 146654
rect 72994 146334 73614 146418
rect 72994 146098 73026 146334
rect 73262 146098 73346 146334
rect 73582 146098 73614 146334
rect 72994 110654 73614 146098
rect 72994 110418 73026 110654
rect 73262 110418 73346 110654
rect 73582 110418 73614 110654
rect 72994 110334 73614 110418
rect 72994 110098 73026 110334
rect 73262 110098 73346 110334
rect 73582 110098 73614 110334
rect 72994 74654 73614 110098
rect 72994 74418 73026 74654
rect 73262 74418 73346 74654
rect 73582 74418 73614 74654
rect 72994 74334 73614 74418
rect 72994 74098 73026 74334
rect 73262 74098 73346 74334
rect 73582 74098 73614 74334
rect 72994 38654 73614 74098
rect 72994 38418 73026 38654
rect 73262 38418 73346 38654
rect 73582 38418 73614 38654
rect 72994 38334 73614 38418
rect 72994 38098 73026 38334
rect 73262 38098 73346 38334
rect 73582 38098 73614 38334
rect 72994 2654 73614 38098
rect 72994 2418 73026 2654
rect 73262 2418 73346 2654
rect 73582 2418 73614 2654
rect 72994 2334 73614 2418
rect 72994 2098 73026 2334
rect 73262 2098 73346 2334
rect 73582 2098 73614 2334
rect 72994 -346 73614 2098
rect 72994 -582 73026 -346
rect 73262 -582 73346 -346
rect 73582 -582 73614 -346
rect 72994 -666 73614 -582
rect 72994 -902 73026 -666
rect 73262 -902 73346 -666
rect 73582 -902 73614 -666
rect 72994 -7654 73614 -902
rect 74234 705798 74854 711590
rect 74234 705562 74266 705798
rect 74502 705562 74586 705798
rect 74822 705562 74854 705798
rect 74234 705478 74854 705562
rect 74234 705242 74266 705478
rect 74502 705242 74586 705478
rect 74822 705242 74854 705478
rect 74234 687894 74854 705242
rect 74234 687658 74266 687894
rect 74502 687658 74586 687894
rect 74822 687658 74854 687894
rect 74234 687574 74854 687658
rect 74234 687338 74266 687574
rect 74502 687338 74586 687574
rect 74822 687338 74854 687574
rect 74234 651894 74854 687338
rect 74234 651658 74266 651894
rect 74502 651658 74586 651894
rect 74822 651658 74854 651894
rect 74234 651574 74854 651658
rect 74234 651338 74266 651574
rect 74502 651338 74586 651574
rect 74822 651338 74854 651574
rect 74234 615894 74854 651338
rect 74234 615658 74266 615894
rect 74502 615658 74586 615894
rect 74822 615658 74854 615894
rect 74234 615574 74854 615658
rect 74234 615338 74266 615574
rect 74502 615338 74586 615574
rect 74822 615338 74854 615574
rect 74234 579894 74854 615338
rect 74234 579658 74266 579894
rect 74502 579658 74586 579894
rect 74822 579658 74854 579894
rect 74234 579574 74854 579658
rect 74234 579338 74266 579574
rect 74502 579338 74586 579574
rect 74822 579338 74854 579574
rect 74234 543894 74854 579338
rect 74234 543658 74266 543894
rect 74502 543658 74586 543894
rect 74822 543658 74854 543894
rect 74234 543574 74854 543658
rect 74234 543338 74266 543574
rect 74502 543338 74586 543574
rect 74822 543338 74854 543574
rect 74234 507894 74854 543338
rect 74234 507658 74266 507894
rect 74502 507658 74586 507894
rect 74822 507658 74854 507894
rect 74234 507574 74854 507658
rect 74234 507338 74266 507574
rect 74502 507338 74586 507574
rect 74822 507338 74854 507574
rect 74234 471894 74854 507338
rect 74234 471658 74266 471894
rect 74502 471658 74586 471894
rect 74822 471658 74854 471894
rect 74234 471574 74854 471658
rect 74234 471338 74266 471574
rect 74502 471338 74586 471574
rect 74822 471338 74854 471574
rect 74234 435894 74854 471338
rect 74234 435658 74266 435894
rect 74502 435658 74586 435894
rect 74822 435658 74854 435894
rect 74234 435574 74854 435658
rect 74234 435338 74266 435574
rect 74502 435338 74586 435574
rect 74822 435338 74854 435574
rect 74234 399894 74854 435338
rect 74234 399658 74266 399894
rect 74502 399658 74586 399894
rect 74822 399658 74854 399894
rect 74234 399574 74854 399658
rect 74234 399338 74266 399574
rect 74502 399338 74586 399574
rect 74822 399338 74854 399574
rect 74234 363894 74854 399338
rect 74234 363658 74266 363894
rect 74502 363658 74586 363894
rect 74822 363658 74854 363894
rect 74234 363574 74854 363658
rect 74234 363338 74266 363574
rect 74502 363338 74586 363574
rect 74822 363338 74854 363574
rect 74234 327894 74854 363338
rect 74234 327658 74266 327894
rect 74502 327658 74586 327894
rect 74822 327658 74854 327894
rect 74234 327574 74854 327658
rect 74234 327338 74266 327574
rect 74502 327338 74586 327574
rect 74822 327338 74854 327574
rect 74234 291894 74854 327338
rect 74234 291658 74266 291894
rect 74502 291658 74586 291894
rect 74822 291658 74854 291894
rect 74234 291574 74854 291658
rect 74234 291338 74266 291574
rect 74502 291338 74586 291574
rect 74822 291338 74854 291574
rect 74234 255894 74854 291338
rect 74234 255658 74266 255894
rect 74502 255658 74586 255894
rect 74822 255658 74854 255894
rect 74234 255574 74854 255658
rect 74234 255338 74266 255574
rect 74502 255338 74586 255574
rect 74822 255338 74854 255574
rect 74234 219894 74854 255338
rect 74234 219658 74266 219894
rect 74502 219658 74586 219894
rect 74822 219658 74854 219894
rect 74234 219574 74854 219658
rect 74234 219338 74266 219574
rect 74502 219338 74586 219574
rect 74822 219338 74854 219574
rect 74234 183894 74854 219338
rect 74234 183658 74266 183894
rect 74502 183658 74586 183894
rect 74822 183658 74854 183894
rect 74234 183574 74854 183658
rect 74234 183338 74266 183574
rect 74502 183338 74586 183574
rect 74822 183338 74854 183574
rect 74234 147894 74854 183338
rect 74234 147658 74266 147894
rect 74502 147658 74586 147894
rect 74822 147658 74854 147894
rect 74234 147574 74854 147658
rect 74234 147338 74266 147574
rect 74502 147338 74586 147574
rect 74822 147338 74854 147574
rect 74234 111894 74854 147338
rect 74234 111658 74266 111894
rect 74502 111658 74586 111894
rect 74822 111658 74854 111894
rect 74234 111574 74854 111658
rect 74234 111338 74266 111574
rect 74502 111338 74586 111574
rect 74822 111338 74854 111574
rect 74234 75894 74854 111338
rect 74234 75658 74266 75894
rect 74502 75658 74586 75894
rect 74822 75658 74854 75894
rect 74234 75574 74854 75658
rect 74234 75338 74266 75574
rect 74502 75338 74586 75574
rect 74822 75338 74854 75574
rect 74234 39894 74854 75338
rect 74234 39658 74266 39894
rect 74502 39658 74586 39894
rect 74822 39658 74854 39894
rect 74234 39574 74854 39658
rect 74234 39338 74266 39574
rect 74502 39338 74586 39574
rect 74822 39338 74854 39574
rect 74234 3894 74854 39338
rect 74234 3658 74266 3894
rect 74502 3658 74586 3894
rect 74822 3658 74854 3894
rect 74234 3574 74854 3658
rect 74234 3338 74266 3574
rect 74502 3338 74586 3574
rect 74822 3338 74854 3574
rect 74234 -1306 74854 3338
rect 74234 -1542 74266 -1306
rect 74502 -1542 74586 -1306
rect 74822 -1542 74854 -1306
rect 74234 -1626 74854 -1542
rect 74234 -1862 74266 -1626
rect 74502 -1862 74586 -1626
rect 74822 -1862 74854 -1626
rect 74234 -7654 74854 -1862
rect 75474 706758 76094 711590
rect 75474 706522 75506 706758
rect 75742 706522 75826 706758
rect 76062 706522 76094 706758
rect 75474 706438 76094 706522
rect 75474 706202 75506 706438
rect 75742 706202 75826 706438
rect 76062 706202 76094 706438
rect 75474 689134 76094 706202
rect 75474 688898 75506 689134
rect 75742 688898 75826 689134
rect 76062 688898 76094 689134
rect 75474 688814 76094 688898
rect 75474 688578 75506 688814
rect 75742 688578 75826 688814
rect 76062 688578 76094 688814
rect 75474 653134 76094 688578
rect 75474 652898 75506 653134
rect 75742 652898 75826 653134
rect 76062 652898 76094 653134
rect 75474 652814 76094 652898
rect 75474 652578 75506 652814
rect 75742 652578 75826 652814
rect 76062 652578 76094 652814
rect 75474 617134 76094 652578
rect 75474 616898 75506 617134
rect 75742 616898 75826 617134
rect 76062 616898 76094 617134
rect 75474 616814 76094 616898
rect 75474 616578 75506 616814
rect 75742 616578 75826 616814
rect 76062 616578 76094 616814
rect 75474 581134 76094 616578
rect 75474 580898 75506 581134
rect 75742 580898 75826 581134
rect 76062 580898 76094 581134
rect 75474 580814 76094 580898
rect 75474 580578 75506 580814
rect 75742 580578 75826 580814
rect 76062 580578 76094 580814
rect 75474 545134 76094 580578
rect 75474 544898 75506 545134
rect 75742 544898 75826 545134
rect 76062 544898 76094 545134
rect 75474 544814 76094 544898
rect 75474 544578 75506 544814
rect 75742 544578 75826 544814
rect 76062 544578 76094 544814
rect 75474 509134 76094 544578
rect 75474 508898 75506 509134
rect 75742 508898 75826 509134
rect 76062 508898 76094 509134
rect 75474 508814 76094 508898
rect 75474 508578 75506 508814
rect 75742 508578 75826 508814
rect 76062 508578 76094 508814
rect 75474 473134 76094 508578
rect 75474 472898 75506 473134
rect 75742 472898 75826 473134
rect 76062 472898 76094 473134
rect 75474 472814 76094 472898
rect 75474 472578 75506 472814
rect 75742 472578 75826 472814
rect 76062 472578 76094 472814
rect 75474 437134 76094 472578
rect 75474 436898 75506 437134
rect 75742 436898 75826 437134
rect 76062 436898 76094 437134
rect 75474 436814 76094 436898
rect 75474 436578 75506 436814
rect 75742 436578 75826 436814
rect 76062 436578 76094 436814
rect 75474 401134 76094 436578
rect 75474 400898 75506 401134
rect 75742 400898 75826 401134
rect 76062 400898 76094 401134
rect 75474 400814 76094 400898
rect 75474 400578 75506 400814
rect 75742 400578 75826 400814
rect 76062 400578 76094 400814
rect 75474 365134 76094 400578
rect 75474 364898 75506 365134
rect 75742 364898 75826 365134
rect 76062 364898 76094 365134
rect 75474 364814 76094 364898
rect 75474 364578 75506 364814
rect 75742 364578 75826 364814
rect 76062 364578 76094 364814
rect 75474 329134 76094 364578
rect 75474 328898 75506 329134
rect 75742 328898 75826 329134
rect 76062 328898 76094 329134
rect 75474 328814 76094 328898
rect 75474 328578 75506 328814
rect 75742 328578 75826 328814
rect 76062 328578 76094 328814
rect 75474 293134 76094 328578
rect 75474 292898 75506 293134
rect 75742 292898 75826 293134
rect 76062 292898 76094 293134
rect 75474 292814 76094 292898
rect 75474 292578 75506 292814
rect 75742 292578 75826 292814
rect 76062 292578 76094 292814
rect 75474 257134 76094 292578
rect 75474 256898 75506 257134
rect 75742 256898 75826 257134
rect 76062 256898 76094 257134
rect 75474 256814 76094 256898
rect 75474 256578 75506 256814
rect 75742 256578 75826 256814
rect 76062 256578 76094 256814
rect 75474 221134 76094 256578
rect 75474 220898 75506 221134
rect 75742 220898 75826 221134
rect 76062 220898 76094 221134
rect 75474 220814 76094 220898
rect 75474 220578 75506 220814
rect 75742 220578 75826 220814
rect 76062 220578 76094 220814
rect 75474 185134 76094 220578
rect 75474 184898 75506 185134
rect 75742 184898 75826 185134
rect 76062 184898 76094 185134
rect 75474 184814 76094 184898
rect 75474 184578 75506 184814
rect 75742 184578 75826 184814
rect 76062 184578 76094 184814
rect 75474 149134 76094 184578
rect 75474 148898 75506 149134
rect 75742 148898 75826 149134
rect 76062 148898 76094 149134
rect 75474 148814 76094 148898
rect 75474 148578 75506 148814
rect 75742 148578 75826 148814
rect 76062 148578 76094 148814
rect 75474 113134 76094 148578
rect 75474 112898 75506 113134
rect 75742 112898 75826 113134
rect 76062 112898 76094 113134
rect 75474 112814 76094 112898
rect 75474 112578 75506 112814
rect 75742 112578 75826 112814
rect 76062 112578 76094 112814
rect 75474 77134 76094 112578
rect 75474 76898 75506 77134
rect 75742 76898 75826 77134
rect 76062 76898 76094 77134
rect 75474 76814 76094 76898
rect 75474 76578 75506 76814
rect 75742 76578 75826 76814
rect 76062 76578 76094 76814
rect 75474 41134 76094 76578
rect 75474 40898 75506 41134
rect 75742 40898 75826 41134
rect 76062 40898 76094 41134
rect 75474 40814 76094 40898
rect 75474 40578 75506 40814
rect 75742 40578 75826 40814
rect 76062 40578 76094 40814
rect 75474 5134 76094 40578
rect 75474 4898 75506 5134
rect 75742 4898 75826 5134
rect 76062 4898 76094 5134
rect 75474 4814 76094 4898
rect 75474 4578 75506 4814
rect 75742 4578 75826 4814
rect 76062 4578 76094 4814
rect 75474 -2266 76094 4578
rect 75474 -2502 75506 -2266
rect 75742 -2502 75826 -2266
rect 76062 -2502 76094 -2266
rect 75474 -2586 76094 -2502
rect 75474 -2822 75506 -2586
rect 75742 -2822 75826 -2586
rect 76062 -2822 76094 -2586
rect 75474 -7654 76094 -2822
rect 76714 707718 77334 711590
rect 76714 707482 76746 707718
rect 76982 707482 77066 707718
rect 77302 707482 77334 707718
rect 76714 707398 77334 707482
rect 76714 707162 76746 707398
rect 76982 707162 77066 707398
rect 77302 707162 77334 707398
rect 76714 690374 77334 707162
rect 76714 690138 76746 690374
rect 76982 690138 77066 690374
rect 77302 690138 77334 690374
rect 76714 690054 77334 690138
rect 76714 689818 76746 690054
rect 76982 689818 77066 690054
rect 77302 689818 77334 690054
rect 76714 654374 77334 689818
rect 76714 654138 76746 654374
rect 76982 654138 77066 654374
rect 77302 654138 77334 654374
rect 76714 654054 77334 654138
rect 76714 653818 76746 654054
rect 76982 653818 77066 654054
rect 77302 653818 77334 654054
rect 76714 618374 77334 653818
rect 76714 618138 76746 618374
rect 76982 618138 77066 618374
rect 77302 618138 77334 618374
rect 76714 618054 77334 618138
rect 76714 617818 76746 618054
rect 76982 617818 77066 618054
rect 77302 617818 77334 618054
rect 76714 582374 77334 617818
rect 76714 582138 76746 582374
rect 76982 582138 77066 582374
rect 77302 582138 77334 582374
rect 76714 582054 77334 582138
rect 76714 581818 76746 582054
rect 76982 581818 77066 582054
rect 77302 581818 77334 582054
rect 76714 546374 77334 581818
rect 76714 546138 76746 546374
rect 76982 546138 77066 546374
rect 77302 546138 77334 546374
rect 76714 546054 77334 546138
rect 76714 545818 76746 546054
rect 76982 545818 77066 546054
rect 77302 545818 77334 546054
rect 76714 510374 77334 545818
rect 76714 510138 76746 510374
rect 76982 510138 77066 510374
rect 77302 510138 77334 510374
rect 76714 510054 77334 510138
rect 76714 509818 76746 510054
rect 76982 509818 77066 510054
rect 77302 509818 77334 510054
rect 76714 474374 77334 509818
rect 76714 474138 76746 474374
rect 76982 474138 77066 474374
rect 77302 474138 77334 474374
rect 76714 474054 77334 474138
rect 76714 473818 76746 474054
rect 76982 473818 77066 474054
rect 77302 473818 77334 474054
rect 76714 438374 77334 473818
rect 76714 438138 76746 438374
rect 76982 438138 77066 438374
rect 77302 438138 77334 438374
rect 76714 438054 77334 438138
rect 76714 437818 76746 438054
rect 76982 437818 77066 438054
rect 77302 437818 77334 438054
rect 76714 402374 77334 437818
rect 76714 402138 76746 402374
rect 76982 402138 77066 402374
rect 77302 402138 77334 402374
rect 76714 402054 77334 402138
rect 76714 401818 76746 402054
rect 76982 401818 77066 402054
rect 77302 401818 77334 402054
rect 76714 366374 77334 401818
rect 76714 366138 76746 366374
rect 76982 366138 77066 366374
rect 77302 366138 77334 366374
rect 76714 366054 77334 366138
rect 76714 365818 76746 366054
rect 76982 365818 77066 366054
rect 77302 365818 77334 366054
rect 76714 330374 77334 365818
rect 76714 330138 76746 330374
rect 76982 330138 77066 330374
rect 77302 330138 77334 330374
rect 76714 330054 77334 330138
rect 76714 329818 76746 330054
rect 76982 329818 77066 330054
rect 77302 329818 77334 330054
rect 76714 294374 77334 329818
rect 76714 294138 76746 294374
rect 76982 294138 77066 294374
rect 77302 294138 77334 294374
rect 76714 294054 77334 294138
rect 76714 293818 76746 294054
rect 76982 293818 77066 294054
rect 77302 293818 77334 294054
rect 76714 258374 77334 293818
rect 76714 258138 76746 258374
rect 76982 258138 77066 258374
rect 77302 258138 77334 258374
rect 76714 258054 77334 258138
rect 76714 257818 76746 258054
rect 76982 257818 77066 258054
rect 77302 257818 77334 258054
rect 76714 222374 77334 257818
rect 76714 222138 76746 222374
rect 76982 222138 77066 222374
rect 77302 222138 77334 222374
rect 76714 222054 77334 222138
rect 76714 221818 76746 222054
rect 76982 221818 77066 222054
rect 77302 221818 77334 222054
rect 76714 186374 77334 221818
rect 76714 186138 76746 186374
rect 76982 186138 77066 186374
rect 77302 186138 77334 186374
rect 76714 186054 77334 186138
rect 76714 185818 76746 186054
rect 76982 185818 77066 186054
rect 77302 185818 77334 186054
rect 76714 150374 77334 185818
rect 76714 150138 76746 150374
rect 76982 150138 77066 150374
rect 77302 150138 77334 150374
rect 76714 150054 77334 150138
rect 76714 149818 76746 150054
rect 76982 149818 77066 150054
rect 77302 149818 77334 150054
rect 76714 114374 77334 149818
rect 76714 114138 76746 114374
rect 76982 114138 77066 114374
rect 77302 114138 77334 114374
rect 76714 114054 77334 114138
rect 76714 113818 76746 114054
rect 76982 113818 77066 114054
rect 77302 113818 77334 114054
rect 76714 78374 77334 113818
rect 76714 78138 76746 78374
rect 76982 78138 77066 78374
rect 77302 78138 77334 78374
rect 76714 78054 77334 78138
rect 76714 77818 76746 78054
rect 76982 77818 77066 78054
rect 77302 77818 77334 78054
rect 76714 42374 77334 77818
rect 76714 42138 76746 42374
rect 76982 42138 77066 42374
rect 77302 42138 77334 42374
rect 76714 42054 77334 42138
rect 76714 41818 76746 42054
rect 76982 41818 77066 42054
rect 77302 41818 77334 42054
rect 76714 6374 77334 41818
rect 76714 6138 76746 6374
rect 76982 6138 77066 6374
rect 77302 6138 77334 6374
rect 76714 6054 77334 6138
rect 76714 5818 76746 6054
rect 76982 5818 77066 6054
rect 77302 5818 77334 6054
rect 76714 -3226 77334 5818
rect 76714 -3462 76746 -3226
rect 76982 -3462 77066 -3226
rect 77302 -3462 77334 -3226
rect 76714 -3546 77334 -3462
rect 76714 -3782 76746 -3546
rect 76982 -3782 77066 -3546
rect 77302 -3782 77334 -3546
rect 76714 -7654 77334 -3782
rect 77954 708678 78574 711590
rect 77954 708442 77986 708678
rect 78222 708442 78306 708678
rect 78542 708442 78574 708678
rect 77954 708358 78574 708442
rect 77954 708122 77986 708358
rect 78222 708122 78306 708358
rect 78542 708122 78574 708358
rect 77954 691614 78574 708122
rect 77954 691378 77986 691614
rect 78222 691378 78306 691614
rect 78542 691378 78574 691614
rect 77954 691294 78574 691378
rect 77954 691058 77986 691294
rect 78222 691058 78306 691294
rect 78542 691058 78574 691294
rect 77954 655614 78574 691058
rect 77954 655378 77986 655614
rect 78222 655378 78306 655614
rect 78542 655378 78574 655614
rect 77954 655294 78574 655378
rect 77954 655058 77986 655294
rect 78222 655058 78306 655294
rect 78542 655058 78574 655294
rect 77954 619614 78574 655058
rect 77954 619378 77986 619614
rect 78222 619378 78306 619614
rect 78542 619378 78574 619614
rect 77954 619294 78574 619378
rect 77954 619058 77986 619294
rect 78222 619058 78306 619294
rect 78542 619058 78574 619294
rect 77954 583614 78574 619058
rect 77954 583378 77986 583614
rect 78222 583378 78306 583614
rect 78542 583378 78574 583614
rect 77954 583294 78574 583378
rect 77954 583058 77986 583294
rect 78222 583058 78306 583294
rect 78542 583058 78574 583294
rect 77954 547614 78574 583058
rect 77954 547378 77986 547614
rect 78222 547378 78306 547614
rect 78542 547378 78574 547614
rect 77954 547294 78574 547378
rect 77954 547058 77986 547294
rect 78222 547058 78306 547294
rect 78542 547058 78574 547294
rect 77954 511614 78574 547058
rect 77954 511378 77986 511614
rect 78222 511378 78306 511614
rect 78542 511378 78574 511614
rect 77954 511294 78574 511378
rect 77954 511058 77986 511294
rect 78222 511058 78306 511294
rect 78542 511058 78574 511294
rect 77954 475614 78574 511058
rect 77954 475378 77986 475614
rect 78222 475378 78306 475614
rect 78542 475378 78574 475614
rect 77954 475294 78574 475378
rect 77954 475058 77986 475294
rect 78222 475058 78306 475294
rect 78542 475058 78574 475294
rect 77954 439614 78574 475058
rect 77954 439378 77986 439614
rect 78222 439378 78306 439614
rect 78542 439378 78574 439614
rect 77954 439294 78574 439378
rect 77954 439058 77986 439294
rect 78222 439058 78306 439294
rect 78542 439058 78574 439294
rect 77954 403614 78574 439058
rect 77954 403378 77986 403614
rect 78222 403378 78306 403614
rect 78542 403378 78574 403614
rect 77954 403294 78574 403378
rect 77954 403058 77986 403294
rect 78222 403058 78306 403294
rect 78542 403058 78574 403294
rect 77954 367614 78574 403058
rect 77954 367378 77986 367614
rect 78222 367378 78306 367614
rect 78542 367378 78574 367614
rect 77954 367294 78574 367378
rect 77954 367058 77986 367294
rect 78222 367058 78306 367294
rect 78542 367058 78574 367294
rect 77954 331614 78574 367058
rect 77954 331378 77986 331614
rect 78222 331378 78306 331614
rect 78542 331378 78574 331614
rect 77954 331294 78574 331378
rect 77954 331058 77986 331294
rect 78222 331058 78306 331294
rect 78542 331058 78574 331294
rect 77954 295614 78574 331058
rect 77954 295378 77986 295614
rect 78222 295378 78306 295614
rect 78542 295378 78574 295614
rect 77954 295294 78574 295378
rect 77954 295058 77986 295294
rect 78222 295058 78306 295294
rect 78542 295058 78574 295294
rect 77954 259614 78574 295058
rect 77954 259378 77986 259614
rect 78222 259378 78306 259614
rect 78542 259378 78574 259614
rect 77954 259294 78574 259378
rect 77954 259058 77986 259294
rect 78222 259058 78306 259294
rect 78542 259058 78574 259294
rect 77954 223614 78574 259058
rect 77954 223378 77986 223614
rect 78222 223378 78306 223614
rect 78542 223378 78574 223614
rect 77954 223294 78574 223378
rect 77954 223058 77986 223294
rect 78222 223058 78306 223294
rect 78542 223058 78574 223294
rect 77954 187614 78574 223058
rect 77954 187378 77986 187614
rect 78222 187378 78306 187614
rect 78542 187378 78574 187614
rect 77954 187294 78574 187378
rect 77954 187058 77986 187294
rect 78222 187058 78306 187294
rect 78542 187058 78574 187294
rect 77954 151614 78574 187058
rect 77954 151378 77986 151614
rect 78222 151378 78306 151614
rect 78542 151378 78574 151614
rect 77954 151294 78574 151378
rect 77954 151058 77986 151294
rect 78222 151058 78306 151294
rect 78542 151058 78574 151294
rect 77954 115614 78574 151058
rect 77954 115378 77986 115614
rect 78222 115378 78306 115614
rect 78542 115378 78574 115614
rect 77954 115294 78574 115378
rect 77954 115058 77986 115294
rect 78222 115058 78306 115294
rect 78542 115058 78574 115294
rect 77954 79614 78574 115058
rect 77954 79378 77986 79614
rect 78222 79378 78306 79614
rect 78542 79378 78574 79614
rect 77954 79294 78574 79378
rect 77954 79058 77986 79294
rect 78222 79058 78306 79294
rect 78542 79058 78574 79294
rect 77954 43614 78574 79058
rect 77954 43378 77986 43614
rect 78222 43378 78306 43614
rect 78542 43378 78574 43614
rect 77954 43294 78574 43378
rect 77954 43058 77986 43294
rect 78222 43058 78306 43294
rect 78542 43058 78574 43294
rect 77954 7614 78574 43058
rect 77954 7378 77986 7614
rect 78222 7378 78306 7614
rect 78542 7378 78574 7614
rect 77954 7294 78574 7378
rect 77954 7058 77986 7294
rect 78222 7058 78306 7294
rect 78542 7058 78574 7294
rect 77954 -4186 78574 7058
rect 77954 -4422 77986 -4186
rect 78222 -4422 78306 -4186
rect 78542 -4422 78574 -4186
rect 77954 -4506 78574 -4422
rect 77954 -4742 77986 -4506
rect 78222 -4742 78306 -4506
rect 78542 -4742 78574 -4506
rect 77954 -7654 78574 -4742
rect 79194 709638 79814 711590
rect 79194 709402 79226 709638
rect 79462 709402 79546 709638
rect 79782 709402 79814 709638
rect 79194 709318 79814 709402
rect 79194 709082 79226 709318
rect 79462 709082 79546 709318
rect 79782 709082 79814 709318
rect 79194 692854 79814 709082
rect 79194 692618 79226 692854
rect 79462 692618 79546 692854
rect 79782 692618 79814 692854
rect 79194 692534 79814 692618
rect 79194 692298 79226 692534
rect 79462 692298 79546 692534
rect 79782 692298 79814 692534
rect 79194 656854 79814 692298
rect 79194 656618 79226 656854
rect 79462 656618 79546 656854
rect 79782 656618 79814 656854
rect 79194 656534 79814 656618
rect 79194 656298 79226 656534
rect 79462 656298 79546 656534
rect 79782 656298 79814 656534
rect 79194 620854 79814 656298
rect 79194 620618 79226 620854
rect 79462 620618 79546 620854
rect 79782 620618 79814 620854
rect 79194 620534 79814 620618
rect 79194 620298 79226 620534
rect 79462 620298 79546 620534
rect 79782 620298 79814 620534
rect 79194 584854 79814 620298
rect 79194 584618 79226 584854
rect 79462 584618 79546 584854
rect 79782 584618 79814 584854
rect 79194 584534 79814 584618
rect 79194 584298 79226 584534
rect 79462 584298 79546 584534
rect 79782 584298 79814 584534
rect 79194 548854 79814 584298
rect 79194 548618 79226 548854
rect 79462 548618 79546 548854
rect 79782 548618 79814 548854
rect 79194 548534 79814 548618
rect 79194 548298 79226 548534
rect 79462 548298 79546 548534
rect 79782 548298 79814 548534
rect 79194 512854 79814 548298
rect 79194 512618 79226 512854
rect 79462 512618 79546 512854
rect 79782 512618 79814 512854
rect 79194 512534 79814 512618
rect 79194 512298 79226 512534
rect 79462 512298 79546 512534
rect 79782 512298 79814 512534
rect 79194 476854 79814 512298
rect 79194 476618 79226 476854
rect 79462 476618 79546 476854
rect 79782 476618 79814 476854
rect 79194 476534 79814 476618
rect 79194 476298 79226 476534
rect 79462 476298 79546 476534
rect 79782 476298 79814 476534
rect 79194 440854 79814 476298
rect 79194 440618 79226 440854
rect 79462 440618 79546 440854
rect 79782 440618 79814 440854
rect 79194 440534 79814 440618
rect 79194 440298 79226 440534
rect 79462 440298 79546 440534
rect 79782 440298 79814 440534
rect 79194 404854 79814 440298
rect 79194 404618 79226 404854
rect 79462 404618 79546 404854
rect 79782 404618 79814 404854
rect 79194 404534 79814 404618
rect 79194 404298 79226 404534
rect 79462 404298 79546 404534
rect 79782 404298 79814 404534
rect 79194 368854 79814 404298
rect 79194 368618 79226 368854
rect 79462 368618 79546 368854
rect 79782 368618 79814 368854
rect 79194 368534 79814 368618
rect 79194 368298 79226 368534
rect 79462 368298 79546 368534
rect 79782 368298 79814 368534
rect 79194 332854 79814 368298
rect 79194 332618 79226 332854
rect 79462 332618 79546 332854
rect 79782 332618 79814 332854
rect 79194 332534 79814 332618
rect 79194 332298 79226 332534
rect 79462 332298 79546 332534
rect 79782 332298 79814 332534
rect 79194 296854 79814 332298
rect 79194 296618 79226 296854
rect 79462 296618 79546 296854
rect 79782 296618 79814 296854
rect 79194 296534 79814 296618
rect 79194 296298 79226 296534
rect 79462 296298 79546 296534
rect 79782 296298 79814 296534
rect 79194 260854 79814 296298
rect 79194 260618 79226 260854
rect 79462 260618 79546 260854
rect 79782 260618 79814 260854
rect 79194 260534 79814 260618
rect 79194 260298 79226 260534
rect 79462 260298 79546 260534
rect 79782 260298 79814 260534
rect 79194 224854 79814 260298
rect 79194 224618 79226 224854
rect 79462 224618 79546 224854
rect 79782 224618 79814 224854
rect 79194 224534 79814 224618
rect 79194 224298 79226 224534
rect 79462 224298 79546 224534
rect 79782 224298 79814 224534
rect 79194 188854 79814 224298
rect 79194 188618 79226 188854
rect 79462 188618 79546 188854
rect 79782 188618 79814 188854
rect 79194 188534 79814 188618
rect 79194 188298 79226 188534
rect 79462 188298 79546 188534
rect 79782 188298 79814 188534
rect 79194 152854 79814 188298
rect 79194 152618 79226 152854
rect 79462 152618 79546 152854
rect 79782 152618 79814 152854
rect 79194 152534 79814 152618
rect 79194 152298 79226 152534
rect 79462 152298 79546 152534
rect 79782 152298 79814 152534
rect 79194 116854 79814 152298
rect 79194 116618 79226 116854
rect 79462 116618 79546 116854
rect 79782 116618 79814 116854
rect 79194 116534 79814 116618
rect 79194 116298 79226 116534
rect 79462 116298 79546 116534
rect 79782 116298 79814 116534
rect 79194 80854 79814 116298
rect 79194 80618 79226 80854
rect 79462 80618 79546 80854
rect 79782 80618 79814 80854
rect 79194 80534 79814 80618
rect 79194 80298 79226 80534
rect 79462 80298 79546 80534
rect 79782 80298 79814 80534
rect 79194 44854 79814 80298
rect 79194 44618 79226 44854
rect 79462 44618 79546 44854
rect 79782 44618 79814 44854
rect 79194 44534 79814 44618
rect 79194 44298 79226 44534
rect 79462 44298 79546 44534
rect 79782 44298 79814 44534
rect 79194 8854 79814 44298
rect 79194 8618 79226 8854
rect 79462 8618 79546 8854
rect 79782 8618 79814 8854
rect 79194 8534 79814 8618
rect 79194 8298 79226 8534
rect 79462 8298 79546 8534
rect 79782 8298 79814 8534
rect 79194 -5146 79814 8298
rect 79194 -5382 79226 -5146
rect 79462 -5382 79546 -5146
rect 79782 -5382 79814 -5146
rect 79194 -5466 79814 -5382
rect 79194 -5702 79226 -5466
rect 79462 -5702 79546 -5466
rect 79782 -5702 79814 -5466
rect 79194 -7654 79814 -5702
rect 80434 710598 81054 711590
rect 80434 710362 80466 710598
rect 80702 710362 80786 710598
rect 81022 710362 81054 710598
rect 80434 710278 81054 710362
rect 80434 710042 80466 710278
rect 80702 710042 80786 710278
rect 81022 710042 81054 710278
rect 80434 694094 81054 710042
rect 80434 693858 80466 694094
rect 80702 693858 80786 694094
rect 81022 693858 81054 694094
rect 80434 693774 81054 693858
rect 80434 693538 80466 693774
rect 80702 693538 80786 693774
rect 81022 693538 81054 693774
rect 80434 658094 81054 693538
rect 80434 657858 80466 658094
rect 80702 657858 80786 658094
rect 81022 657858 81054 658094
rect 80434 657774 81054 657858
rect 80434 657538 80466 657774
rect 80702 657538 80786 657774
rect 81022 657538 81054 657774
rect 80434 622094 81054 657538
rect 80434 621858 80466 622094
rect 80702 621858 80786 622094
rect 81022 621858 81054 622094
rect 80434 621774 81054 621858
rect 80434 621538 80466 621774
rect 80702 621538 80786 621774
rect 81022 621538 81054 621774
rect 80434 586094 81054 621538
rect 80434 585858 80466 586094
rect 80702 585858 80786 586094
rect 81022 585858 81054 586094
rect 80434 585774 81054 585858
rect 80434 585538 80466 585774
rect 80702 585538 80786 585774
rect 81022 585538 81054 585774
rect 80434 550094 81054 585538
rect 80434 549858 80466 550094
rect 80702 549858 80786 550094
rect 81022 549858 81054 550094
rect 80434 549774 81054 549858
rect 80434 549538 80466 549774
rect 80702 549538 80786 549774
rect 81022 549538 81054 549774
rect 80434 514094 81054 549538
rect 80434 513858 80466 514094
rect 80702 513858 80786 514094
rect 81022 513858 81054 514094
rect 80434 513774 81054 513858
rect 80434 513538 80466 513774
rect 80702 513538 80786 513774
rect 81022 513538 81054 513774
rect 80434 478094 81054 513538
rect 80434 477858 80466 478094
rect 80702 477858 80786 478094
rect 81022 477858 81054 478094
rect 80434 477774 81054 477858
rect 80434 477538 80466 477774
rect 80702 477538 80786 477774
rect 81022 477538 81054 477774
rect 80434 442094 81054 477538
rect 80434 441858 80466 442094
rect 80702 441858 80786 442094
rect 81022 441858 81054 442094
rect 80434 441774 81054 441858
rect 80434 441538 80466 441774
rect 80702 441538 80786 441774
rect 81022 441538 81054 441774
rect 80434 406094 81054 441538
rect 80434 405858 80466 406094
rect 80702 405858 80786 406094
rect 81022 405858 81054 406094
rect 80434 405774 81054 405858
rect 80434 405538 80466 405774
rect 80702 405538 80786 405774
rect 81022 405538 81054 405774
rect 80434 370094 81054 405538
rect 80434 369858 80466 370094
rect 80702 369858 80786 370094
rect 81022 369858 81054 370094
rect 80434 369774 81054 369858
rect 80434 369538 80466 369774
rect 80702 369538 80786 369774
rect 81022 369538 81054 369774
rect 80434 334094 81054 369538
rect 80434 333858 80466 334094
rect 80702 333858 80786 334094
rect 81022 333858 81054 334094
rect 80434 333774 81054 333858
rect 80434 333538 80466 333774
rect 80702 333538 80786 333774
rect 81022 333538 81054 333774
rect 80434 298094 81054 333538
rect 80434 297858 80466 298094
rect 80702 297858 80786 298094
rect 81022 297858 81054 298094
rect 80434 297774 81054 297858
rect 80434 297538 80466 297774
rect 80702 297538 80786 297774
rect 81022 297538 81054 297774
rect 80434 262094 81054 297538
rect 80434 261858 80466 262094
rect 80702 261858 80786 262094
rect 81022 261858 81054 262094
rect 80434 261774 81054 261858
rect 80434 261538 80466 261774
rect 80702 261538 80786 261774
rect 81022 261538 81054 261774
rect 80434 226094 81054 261538
rect 80434 225858 80466 226094
rect 80702 225858 80786 226094
rect 81022 225858 81054 226094
rect 80434 225774 81054 225858
rect 80434 225538 80466 225774
rect 80702 225538 80786 225774
rect 81022 225538 81054 225774
rect 80434 190094 81054 225538
rect 80434 189858 80466 190094
rect 80702 189858 80786 190094
rect 81022 189858 81054 190094
rect 80434 189774 81054 189858
rect 80434 189538 80466 189774
rect 80702 189538 80786 189774
rect 81022 189538 81054 189774
rect 80434 154094 81054 189538
rect 80434 153858 80466 154094
rect 80702 153858 80786 154094
rect 81022 153858 81054 154094
rect 80434 153774 81054 153858
rect 80434 153538 80466 153774
rect 80702 153538 80786 153774
rect 81022 153538 81054 153774
rect 80434 118094 81054 153538
rect 80434 117858 80466 118094
rect 80702 117858 80786 118094
rect 81022 117858 81054 118094
rect 80434 117774 81054 117858
rect 80434 117538 80466 117774
rect 80702 117538 80786 117774
rect 81022 117538 81054 117774
rect 80434 82094 81054 117538
rect 80434 81858 80466 82094
rect 80702 81858 80786 82094
rect 81022 81858 81054 82094
rect 80434 81774 81054 81858
rect 80434 81538 80466 81774
rect 80702 81538 80786 81774
rect 81022 81538 81054 81774
rect 80434 46094 81054 81538
rect 80434 45858 80466 46094
rect 80702 45858 80786 46094
rect 81022 45858 81054 46094
rect 80434 45774 81054 45858
rect 80434 45538 80466 45774
rect 80702 45538 80786 45774
rect 81022 45538 81054 45774
rect 80434 10094 81054 45538
rect 80434 9858 80466 10094
rect 80702 9858 80786 10094
rect 81022 9858 81054 10094
rect 80434 9774 81054 9858
rect 80434 9538 80466 9774
rect 80702 9538 80786 9774
rect 81022 9538 81054 9774
rect 80434 -6106 81054 9538
rect 80434 -6342 80466 -6106
rect 80702 -6342 80786 -6106
rect 81022 -6342 81054 -6106
rect 80434 -6426 81054 -6342
rect 80434 -6662 80466 -6426
rect 80702 -6662 80786 -6426
rect 81022 -6662 81054 -6426
rect 80434 -7654 81054 -6662
rect 81674 711558 82294 711590
rect 81674 711322 81706 711558
rect 81942 711322 82026 711558
rect 82262 711322 82294 711558
rect 81674 711238 82294 711322
rect 81674 711002 81706 711238
rect 81942 711002 82026 711238
rect 82262 711002 82294 711238
rect 81674 695334 82294 711002
rect 81674 695098 81706 695334
rect 81942 695098 82026 695334
rect 82262 695098 82294 695334
rect 81674 695014 82294 695098
rect 81674 694778 81706 695014
rect 81942 694778 82026 695014
rect 82262 694778 82294 695014
rect 81674 659334 82294 694778
rect 81674 659098 81706 659334
rect 81942 659098 82026 659334
rect 82262 659098 82294 659334
rect 81674 659014 82294 659098
rect 81674 658778 81706 659014
rect 81942 658778 82026 659014
rect 82262 658778 82294 659014
rect 81674 623334 82294 658778
rect 81674 623098 81706 623334
rect 81942 623098 82026 623334
rect 82262 623098 82294 623334
rect 81674 623014 82294 623098
rect 81674 622778 81706 623014
rect 81942 622778 82026 623014
rect 82262 622778 82294 623014
rect 81674 587334 82294 622778
rect 81674 587098 81706 587334
rect 81942 587098 82026 587334
rect 82262 587098 82294 587334
rect 81674 587014 82294 587098
rect 81674 586778 81706 587014
rect 81942 586778 82026 587014
rect 82262 586778 82294 587014
rect 81674 551334 82294 586778
rect 81674 551098 81706 551334
rect 81942 551098 82026 551334
rect 82262 551098 82294 551334
rect 81674 551014 82294 551098
rect 81674 550778 81706 551014
rect 81942 550778 82026 551014
rect 82262 550778 82294 551014
rect 81674 515334 82294 550778
rect 81674 515098 81706 515334
rect 81942 515098 82026 515334
rect 82262 515098 82294 515334
rect 81674 515014 82294 515098
rect 81674 514778 81706 515014
rect 81942 514778 82026 515014
rect 82262 514778 82294 515014
rect 81674 479334 82294 514778
rect 81674 479098 81706 479334
rect 81942 479098 82026 479334
rect 82262 479098 82294 479334
rect 81674 479014 82294 479098
rect 81674 478778 81706 479014
rect 81942 478778 82026 479014
rect 82262 478778 82294 479014
rect 81674 443334 82294 478778
rect 81674 443098 81706 443334
rect 81942 443098 82026 443334
rect 82262 443098 82294 443334
rect 81674 443014 82294 443098
rect 81674 442778 81706 443014
rect 81942 442778 82026 443014
rect 82262 442778 82294 443014
rect 81674 407334 82294 442778
rect 81674 407098 81706 407334
rect 81942 407098 82026 407334
rect 82262 407098 82294 407334
rect 81674 407014 82294 407098
rect 81674 406778 81706 407014
rect 81942 406778 82026 407014
rect 82262 406778 82294 407014
rect 81674 371334 82294 406778
rect 81674 371098 81706 371334
rect 81942 371098 82026 371334
rect 82262 371098 82294 371334
rect 81674 371014 82294 371098
rect 81674 370778 81706 371014
rect 81942 370778 82026 371014
rect 82262 370778 82294 371014
rect 81674 335334 82294 370778
rect 81674 335098 81706 335334
rect 81942 335098 82026 335334
rect 82262 335098 82294 335334
rect 81674 335014 82294 335098
rect 81674 334778 81706 335014
rect 81942 334778 82026 335014
rect 82262 334778 82294 335014
rect 81674 299334 82294 334778
rect 81674 299098 81706 299334
rect 81942 299098 82026 299334
rect 82262 299098 82294 299334
rect 81674 299014 82294 299098
rect 81674 298778 81706 299014
rect 81942 298778 82026 299014
rect 82262 298778 82294 299014
rect 81674 263334 82294 298778
rect 81674 263098 81706 263334
rect 81942 263098 82026 263334
rect 82262 263098 82294 263334
rect 81674 263014 82294 263098
rect 81674 262778 81706 263014
rect 81942 262778 82026 263014
rect 82262 262778 82294 263014
rect 81674 227334 82294 262778
rect 81674 227098 81706 227334
rect 81942 227098 82026 227334
rect 82262 227098 82294 227334
rect 81674 227014 82294 227098
rect 81674 226778 81706 227014
rect 81942 226778 82026 227014
rect 82262 226778 82294 227014
rect 81674 191334 82294 226778
rect 81674 191098 81706 191334
rect 81942 191098 82026 191334
rect 82262 191098 82294 191334
rect 81674 191014 82294 191098
rect 81674 190778 81706 191014
rect 81942 190778 82026 191014
rect 82262 190778 82294 191014
rect 81674 155334 82294 190778
rect 81674 155098 81706 155334
rect 81942 155098 82026 155334
rect 82262 155098 82294 155334
rect 81674 155014 82294 155098
rect 81674 154778 81706 155014
rect 81942 154778 82026 155014
rect 82262 154778 82294 155014
rect 81674 119334 82294 154778
rect 81674 119098 81706 119334
rect 81942 119098 82026 119334
rect 82262 119098 82294 119334
rect 81674 119014 82294 119098
rect 81674 118778 81706 119014
rect 81942 118778 82026 119014
rect 82262 118778 82294 119014
rect 81674 83334 82294 118778
rect 81674 83098 81706 83334
rect 81942 83098 82026 83334
rect 82262 83098 82294 83334
rect 81674 83014 82294 83098
rect 81674 82778 81706 83014
rect 81942 82778 82026 83014
rect 82262 82778 82294 83014
rect 81674 47334 82294 82778
rect 81674 47098 81706 47334
rect 81942 47098 82026 47334
rect 82262 47098 82294 47334
rect 81674 47014 82294 47098
rect 81674 46778 81706 47014
rect 81942 46778 82026 47014
rect 82262 46778 82294 47014
rect 81674 11334 82294 46778
rect 81674 11098 81706 11334
rect 81942 11098 82026 11334
rect 82262 11098 82294 11334
rect 81674 11014 82294 11098
rect 81674 10778 81706 11014
rect 81942 10778 82026 11014
rect 82262 10778 82294 11014
rect 81674 -7066 82294 10778
rect 81674 -7302 81706 -7066
rect 81942 -7302 82026 -7066
rect 82262 -7302 82294 -7066
rect 81674 -7386 82294 -7302
rect 81674 -7622 81706 -7386
rect 81942 -7622 82026 -7386
rect 82262 -7622 82294 -7386
rect 81674 -7654 82294 -7622
rect 108994 704838 109614 711590
rect 108994 704602 109026 704838
rect 109262 704602 109346 704838
rect 109582 704602 109614 704838
rect 108994 704518 109614 704602
rect 108994 704282 109026 704518
rect 109262 704282 109346 704518
rect 109582 704282 109614 704518
rect 108994 686654 109614 704282
rect 108994 686418 109026 686654
rect 109262 686418 109346 686654
rect 109582 686418 109614 686654
rect 108994 686334 109614 686418
rect 108994 686098 109026 686334
rect 109262 686098 109346 686334
rect 109582 686098 109614 686334
rect 108994 650654 109614 686098
rect 108994 650418 109026 650654
rect 109262 650418 109346 650654
rect 109582 650418 109614 650654
rect 108994 650334 109614 650418
rect 108994 650098 109026 650334
rect 109262 650098 109346 650334
rect 109582 650098 109614 650334
rect 108994 614654 109614 650098
rect 108994 614418 109026 614654
rect 109262 614418 109346 614654
rect 109582 614418 109614 614654
rect 108994 614334 109614 614418
rect 108994 614098 109026 614334
rect 109262 614098 109346 614334
rect 109582 614098 109614 614334
rect 108994 578654 109614 614098
rect 108994 578418 109026 578654
rect 109262 578418 109346 578654
rect 109582 578418 109614 578654
rect 108994 578334 109614 578418
rect 108994 578098 109026 578334
rect 109262 578098 109346 578334
rect 109582 578098 109614 578334
rect 108994 542654 109614 578098
rect 108994 542418 109026 542654
rect 109262 542418 109346 542654
rect 109582 542418 109614 542654
rect 108994 542334 109614 542418
rect 108994 542098 109026 542334
rect 109262 542098 109346 542334
rect 109582 542098 109614 542334
rect 108994 506654 109614 542098
rect 108994 506418 109026 506654
rect 109262 506418 109346 506654
rect 109582 506418 109614 506654
rect 108994 506334 109614 506418
rect 108994 506098 109026 506334
rect 109262 506098 109346 506334
rect 109582 506098 109614 506334
rect 108994 470654 109614 506098
rect 108994 470418 109026 470654
rect 109262 470418 109346 470654
rect 109582 470418 109614 470654
rect 108994 470334 109614 470418
rect 108994 470098 109026 470334
rect 109262 470098 109346 470334
rect 109582 470098 109614 470334
rect 108994 434654 109614 470098
rect 108994 434418 109026 434654
rect 109262 434418 109346 434654
rect 109582 434418 109614 434654
rect 108994 434334 109614 434418
rect 108994 434098 109026 434334
rect 109262 434098 109346 434334
rect 109582 434098 109614 434334
rect 108994 398654 109614 434098
rect 108994 398418 109026 398654
rect 109262 398418 109346 398654
rect 109582 398418 109614 398654
rect 108994 398334 109614 398418
rect 108994 398098 109026 398334
rect 109262 398098 109346 398334
rect 109582 398098 109614 398334
rect 108994 362654 109614 398098
rect 108994 362418 109026 362654
rect 109262 362418 109346 362654
rect 109582 362418 109614 362654
rect 108994 362334 109614 362418
rect 108994 362098 109026 362334
rect 109262 362098 109346 362334
rect 109582 362098 109614 362334
rect 108994 326654 109614 362098
rect 108994 326418 109026 326654
rect 109262 326418 109346 326654
rect 109582 326418 109614 326654
rect 108994 326334 109614 326418
rect 108994 326098 109026 326334
rect 109262 326098 109346 326334
rect 109582 326098 109614 326334
rect 108994 290654 109614 326098
rect 108994 290418 109026 290654
rect 109262 290418 109346 290654
rect 109582 290418 109614 290654
rect 108994 290334 109614 290418
rect 108994 290098 109026 290334
rect 109262 290098 109346 290334
rect 109582 290098 109614 290334
rect 108994 254654 109614 290098
rect 108994 254418 109026 254654
rect 109262 254418 109346 254654
rect 109582 254418 109614 254654
rect 108994 254334 109614 254418
rect 108994 254098 109026 254334
rect 109262 254098 109346 254334
rect 109582 254098 109614 254334
rect 108994 218654 109614 254098
rect 108994 218418 109026 218654
rect 109262 218418 109346 218654
rect 109582 218418 109614 218654
rect 108994 218334 109614 218418
rect 108994 218098 109026 218334
rect 109262 218098 109346 218334
rect 109582 218098 109614 218334
rect 108994 182654 109614 218098
rect 108994 182418 109026 182654
rect 109262 182418 109346 182654
rect 109582 182418 109614 182654
rect 108994 182334 109614 182418
rect 108994 182098 109026 182334
rect 109262 182098 109346 182334
rect 109582 182098 109614 182334
rect 108994 146654 109614 182098
rect 108994 146418 109026 146654
rect 109262 146418 109346 146654
rect 109582 146418 109614 146654
rect 108994 146334 109614 146418
rect 108994 146098 109026 146334
rect 109262 146098 109346 146334
rect 109582 146098 109614 146334
rect 108994 110654 109614 146098
rect 108994 110418 109026 110654
rect 109262 110418 109346 110654
rect 109582 110418 109614 110654
rect 108994 110334 109614 110418
rect 108994 110098 109026 110334
rect 109262 110098 109346 110334
rect 109582 110098 109614 110334
rect 108994 74654 109614 110098
rect 108994 74418 109026 74654
rect 109262 74418 109346 74654
rect 109582 74418 109614 74654
rect 108994 74334 109614 74418
rect 108994 74098 109026 74334
rect 109262 74098 109346 74334
rect 109582 74098 109614 74334
rect 108994 38654 109614 74098
rect 108994 38418 109026 38654
rect 109262 38418 109346 38654
rect 109582 38418 109614 38654
rect 108994 38334 109614 38418
rect 108994 38098 109026 38334
rect 109262 38098 109346 38334
rect 109582 38098 109614 38334
rect 108994 2654 109614 38098
rect 108994 2418 109026 2654
rect 109262 2418 109346 2654
rect 109582 2418 109614 2654
rect 108994 2334 109614 2418
rect 108994 2098 109026 2334
rect 109262 2098 109346 2334
rect 109582 2098 109614 2334
rect 108994 -346 109614 2098
rect 108994 -582 109026 -346
rect 109262 -582 109346 -346
rect 109582 -582 109614 -346
rect 108994 -666 109614 -582
rect 108994 -902 109026 -666
rect 109262 -902 109346 -666
rect 109582 -902 109614 -666
rect 108994 -7654 109614 -902
rect 110234 705798 110854 711590
rect 110234 705562 110266 705798
rect 110502 705562 110586 705798
rect 110822 705562 110854 705798
rect 110234 705478 110854 705562
rect 110234 705242 110266 705478
rect 110502 705242 110586 705478
rect 110822 705242 110854 705478
rect 110234 687894 110854 705242
rect 110234 687658 110266 687894
rect 110502 687658 110586 687894
rect 110822 687658 110854 687894
rect 110234 687574 110854 687658
rect 110234 687338 110266 687574
rect 110502 687338 110586 687574
rect 110822 687338 110854 687574
rect 110234 651894 110854 687338
rect 110234 651658 110266 651894
rect 110502 651658 110586 651894
rect 110822 651658 110854 651894
rect 110234 651574 110854 651658
rect 110234 651338 110266 651574
rect 110502 651338 110586 651574
rect 110822 651338 110854 651574
rect 110234 615894 110854 651338
rect 110234 615658 110266 615894
rect 110502 615658 110586 615894
rect 110822 615658 110854 615894
rect 110234 615574 110854 615658
rect 110234 615338 110266 615574
rect 110502 615338 110586 615574
rect 110822 615338 110854 615574
rect 110234 579894 110854 615338
rect 110234 579658 110266 579894
rect 110502 579658 110586 579894
rect 110822 579658 110854 579894
rect 110234 579574 110854 579658
rect 110234 579338 110266 579574
rect 110502 579338 110586 579574
rect 110822 579338 110854 579574
rect 110234 543894 110854 579338
rect 110234 543658 110266 543894
rect 110502 543658 110586 543894
rect 110822 543658 110854 543894
rect 110234 543574 110854 543658
rect 110234 543338 110266 543574
rect 110502 543338 110586 543574
rect 110822 543338 110854 543574
rect 110234 507894 110854 543338
rect 110234 507658 110266 507894
rect 110502 507658 110586 507894
rect 110822 507658 110854 507894
rect 110234 507574 110854 507658
rect 110234 507338 110266 507574
rect 110502 507338 110586 507574
rect 110822 507338 110854 507574
rect 110234 471894 110854 507338
rect 110234 471658 110266 471894
rect 110502 471658 110586 471894
rect 110822 471658 110854 471894
rect 110234 471574 110854 471658
rect 110234 471338 110266 471574
rect 110502 471338 110586 471574
rect 110822 471338 110854 471574
rect 110234 435894 110854 471338
rect 110234 435658 110266 435894
rect 110502 435658 110586 435894
rect 110822 435658 110854 435894
rect 110234 435574 110854 435658
rect 110234 435338 110266 435574
rect 110502 435338 110586 435574
rect 110822 435338 110854 435574
rect 110234 399894 110854 435338
rect 110234 399658 110266 399894
rect 110502 399658 110586 399894
rect 110822 399658 110854 399894
rect 110234 399574 110854 399658
rect 110234 399338 110266 399574
rect 110502 399338 110586 399574
rect 110822 399338 110854 399574
rect 110234 363894 110854 399338
rect 110234 363658 110266 363894
rect 110502 363658 110586 363894
rect 110822 363658 110854 363894
rect 110234 363574 110854 363658
rect 110234 363338 110266 363574
rect 110502 363338 110586 363574
rect 110822 363338 110854 363574
rect 110234 327894 110854 363338
rect 110234 327658 110266 327894
rect 110502 327658 110586 327894
rect 110822 327658 110854 327894
rect 110234 327574 110854 327658
rect 110234 327338 110266 327574
rect 110502 327338 110586 327574
rect 110822 327338 110854 327574
rect 110234 291894 110854 327338
rect 110234 291658 110266 291894
rect 110502 291658 110586 291894
rect 110822 291658 110854 291894
rect 110234 291574 110854 291658
rect 110234 291338 110266 291574
rect 110502 291338 110586 291574
rect 110822 291338 110854 291574
rect 110234 255894 110854 291338
rect 110234 255658 110266 255894
rect 110502 255658 110586 255894
rect 110822 255658 110854 255894
rect 110234 255574 110854 255658
rect 110234 255338 110266 255574
rect 110502 255338 110586 255574
rect 110822 255338 110854 255574
rect 110234 219894 110854 255338
rect 110234 219658 110266 219894
rect 110502 219658 110586 219894
rect 110822 219658 110854 219894
rect 110234 219574 110854 219658
rect 110234 219338 110266 219574
rect 110502 219338 110586 219574
rect 110822 219338 110854 219574
rect 110234 183894 110854 219338
rect 110234 183658 110266 183894
rect 110502 183658 110586 183894
rect 110822 183658 110854 183894
rect 110234 183574 110854 183658
rect 110234 183338 110266 183574
rect 110502 183338 110586 183574
rect 110822 183338 110854 183574
rect 110234 147894 110854 183338
rect 110234 147658 110266 147894
rect 110502 147658 110586 147894
rect 110822 147658 110854 147894
rect 110234 147574 110854 147658
rect 110234 147338 110266 147574
rect 110502 147338 110586 147574
rect 110822 147338 110854 147574
rect 110234 111894 110854 147338
rect 110234 111658 110266 111894
rect 110502 111658 110586 111894
rect 110822 111658 110854 111894
rect 110234 111574 110854 111658
rect 110234 111338 110266 111574
rect 110502 111338 110586 111574
rect 110822 111338 110854 111574
rect 110234 75894 110854 111338
rect 110234 75658 110266 75894
rect 110502 75658 110586 75894
rect 110822 75658 110854 75894
rect 110234 75574 110854 75658
rect 110234 75338 110266 75574
rect 110502 75338 110586 75574
rect 110822 75338 110854 75574
rect 110234 39894 110854 75338
rect 110234 39658 110266 39894
rect 110502 39658 110586 39894
rect 110822 39658 110854 39894
rect 110234 39574 110854 39658
rect 110234 39338 110266 39574
rect 110502 39338 110586 39574
rect 110822 39338 110854 39574
rect 110234 3894 110854 39338
rect 110234 3658 110266 3894
rect 110502 3658 110586 3894
rect 110822 3658 110854 3894
rect 110234 3574 110854 3658
rect 110234 3338 110266 3574
rect 110502 3338 110586 3574
rect 110822 3338 110854 3574
rect 110234 -1306 110854 3338
rect 110234 -1542 110266 -1306
rect 110502 -1542 110586 -1306
rect 110822 -1542 110854 -1306
rect 110234 -1626 110854 -1542
rect 110234 -1862 110266 -1626
rect 110502 -1862 110586 -1626
rect 110822 -1862 110854 -1626
rect 110234 -7654 110854 -1862
rect 111474 706758 112094 711590
rect 111474 706522 111506 706758
rect 111742 706522 111826 706758
rect 112062 706522 112094 706758
rect 111474 706438 112094 706522
rect 111474 706202 111506 706438
rect 111742 706202 111826 706438
rect 112062 706202 112094 706438
rect 111474 689134 112094 706202
rect 111474 688898 111506 689134
rect 111742 688898 111826 689134
rect 112062 688898 112094 689134
rect 111474 688814 112094 688898
rect 111474 688578 111506 688814
rect 111742 688578 111826 688814
rect 112062 688578 112094 688814
rect 111474 653134 112094 688578
rect 111474 652898 111506 653134
rect 111742 652898 111826 653134
rect 112062 652898 112094 653134
rect 111474 652814 112094 652898
rect 111474 652578 111506 652814
rect 111742 652578 111826 652814
rect 112062 652578 112094 652814
rect 111474 617134 112094 652578
rect 111474 616898 111506 617134
rect 111742 616898 111826 617134
rect 112062 616898 112094 617134
rect 111474 616814 112094 616898
rect 111474 616578 111506 616814
rect 111742 616578 111826 616814
rect 112062 616578 112094 616814
rect 111474 581134 112094 616578
rect 111474 580898 111506 581134
rect 111742 580898 111826 581134
rect 112062 580898 112094 581134
rect 111474 580814 112094 580898
rect 111474 580578 111506 580814
rect 111742 580578 111826 580814
rect 112062 580578 112094 580814
rect 111474 545134 112094 580578
rect 111474 544898 111506 545134
rect 111742 544898 111826 545134
rect 112062 544898 112094 545134
rect 111474 544814 112094 544898
rect 111474 544578 111506 544814
rect 111742 544578 111826 544814
rect 112062 544578 112094 544814
rect 111474 509134 112094 544578
rect 111474 508898 111506 509134
rect 111742 508898 111826 509134
rect 112062 508898 112094 509134
rect 111474 508814 112094 508898
rect 111474 508578 111506 508814
rect 111742 508578 111826 508814
rect 112062 508578 112094 508814
rect 111474 473134 112094 508578
rect 111474 472898 111506 473134
rect 111742 472898 111826 473134
rect 112062 472898 112094 473134
rect 111474 472814 112094 472898
rect 111474 472578 111506 472814
rect 111742 472578 111826 472814
rect 112062 472578 112094 472814
rect 111474 437134 112094 472578
rect 111474 436898 111506 437134
rect 111742 436898 111826 437134
rect 112062 436898 112094 437134
rect 111474 436814 112094 436898
rect 111474 436578 111506 436814
rect 111742 436578 111826 436814
rect 112062 436578 112094 436814
rect 111474 401134 112094 436578
rect 111474 400898 111506 401134
rect 111742 400898 111826 401134
rect 112062 400898 112094 401134
rect 111474 400814 112094 400898
rect 111474 400578 111506 400814
rect 111742 400578 111826 400814
rect 112062 400578 112094 400814
rect 111474 365134 112094 400578
rect 111474 364898 111506 365134
rect 111742 364898 111826 365134
rect 112062 364898 112094 365134
rect 111474 364814 112094 364898
rect 111474 364578 111506 364814
rect 111742 364578 111826 364814
rect 112062 364578 112094 364814
rect 111474 329134 112094 364578
rect 111474 328898 111506 329134
rect 111742 328898 111826 329134
rect 112062 328898 112094 329134
rect 111474 328814 112094 328898
rect 111474 328578 111506 328814
rect 111742 328578 111826 328814
rect 112062 328578 112094 328814
rect 111474 293134 112094 328578
rect 111474 292898 111506 293134
rect 111742 292898 111826 293134
rect 112062 292898 112094 293134
rect 111474 292814 112094 292898
rect 111474 292578 111506 292814
rect 111742 292578 111826 292814
rect 112062 292578 112094 292814
rect 111474 257134 112094 292578
rect 111474 256898 111506 257134
rect 111742 256898 111826 257134
rect 112062 256898 112094 257134
rect 111474 256814 112094 256898
rect 111474 256578 111506 256814
rect 111742 256578 111826 256814
rect 112062 256578 112094 256814
rect 111474 221134 112094 256578
rect 111474 220898 111506 221134
rect 111742 220898 111826 221134
rect 112062 220898 112094 221134
rect 111474 220814 112094 220898
rect 111474 220578 111506 220814
rect 111742 220578 111826 220814
rect 112062 220578 112094 220814
rect 111474 185134 112094 220578
rect 111474 184898 111506 185134
rect 111742 184898 111826 185134
rect 112062 184898 112094 185134
rect 111474 184814 112094 184898
rect 111474 184578 111506 184814
rect 111742 184578 111826 184814
rect 112062 184578 112094 184814
rect 111474 149134 112094 184578
rect 111474 148898 111506 149134
rect 111742 148898 111826 149134
rect 112062 148898 112094 149134
rect 111474 148814 112094 148898
rect 111474 148578 111506 148814
rect 111742 148578 111826 148814
rect 112062 148578 112094 148814
rect 111474 113134 112094 148578
rect 111474 112898 111506 113134
rect 111742 112898 111826 113134
rect 112062 112898 112094 113134
rect 111474 112814 112094 112898
rect 111474 112578 111506 112814
rect 111742 112578 111826 112814
rect 112062 112578 112094 112814
rect 111474 77134 112094 112578
rect 111474 76898 111506 77134
rect 111742 76898 111826 77134
rect 112062 76898 112094 77134
rect 111474 76814 112094 76898
rect 111474 76578 111506 76814
rect 111742 76578 111826 76814
rect 112062 76578 112094 76814
rect 111474 41134 112094 76578
rect 111474 40898 111506 41134
rect 111742 40898 111826 41134
rect 112062 40898 112094 41134
rect 111474 40814 112094 40898
rect 111474 40578 111506 40814
rect 111742 40578 111826 40814
rect 112062 40578 112094 40814
rect 111474 5134 112094 40578
rect 111474 4898 111506 5134
rect 111742 4898 111826 5134
rect 112062 4898 112094 5134
rect 111474 4814 112094 4898
rect 111474 4578 111506 4814
rect 111742 4578 111826 4814
rect 112062 4578 112094 4814
rect 111474 -2266 112094 4578
rect 111474 -2502 111506 -2266
rect 111742 -2502 111826 -2266
rect 112062 -2502 112094 -2266
rect 111474 -2586 112094 -2502
rect 111474 -2822 111506 -2586
rect 111742 -2822 111826 -2586
rect 112062 -2822 112094 -2586
rect 111474 -7654 112094 -2822
rect 112714 707718 113334 711590
rect 112714 707482 112746 707718
rect 112982 707482 113066 707718
rect 113302 707482 113334 707718
rect 112714 707398 113334 707482
rect 112714 707162 112746 707398
rect 112982 707162 113066 707398
rect 113302 707162 113334 707398
rect 112714 690374 113334 707162
rect 112714 690138 112746 690374
rect 112982 690138 113066 690374
rect 113302 690138 113334 690374
rect 112714 690054 113334 690138
rect 112714 689818 112746 690054
rect 112982 689818 113066 690054
rect 113302 689818 113334 690054
rect 112714 654374 113334 689818
rect 112714 654138 112746 654374
rect 112982 654138 113066 654374
rect 113302 654138 113334 654374
rect 112714 654054 113334 654138
rect 112714 653818 112746 654054
rect 112982 653818 113066 654054
rect 113302 653818 113334 654054
rect 112714 618374 113334 653818
rect 112714 618138 112746 618374
rect 112982 618138 113066 618374
rect 113302 618138 113334 618374
rect 112714 618054 113334 618138
rect 112714 617818 112746 618054
rect 112982 617818 113066 618054
rect 113302 617818 113334 618054
rect 112714 582374 113334 617818
rect 112714 582138 112746 582374
rect 112982 582138 113066 582374
rect 113302 582138 113334 582374
rect 112714 582054 113334 582138
rect 112714 581818 112746 582054
rect 112982 581818 113066 582054
rect 113302 581818 113334 582054
rect 112714 546374 113334 581818
rect 112714 546138 112746 546374
rect 112982 546138 113066 546374
rect 113302 546138 113334 546374
rect 112714 546054 113334 546138
rect 112714 545818 112746 546054
rect 112982 545818 113066 546054
rect 113302 545818 113334 546054
rect 112714 510374 113334 545818
rect 112714 510138 112746 510374
rect 112982 510138 113066 510374
rect 113302 510138 113334 510374
rect 112714 510054 113334 510138
rect 112714 509818 112746 510054
rect 112982 509818 113066 510054
rect 113302 509818 113334 510054
rect 112714 474374 113334 509818
rect 112714 474138 112746 474374
rect 112982 474138 113066 474374
rect 113302 474138 113334 474374
rect 112714 474054 113334 474138
rect 112714 473818 112746 474054
rect 112982 473818 113066 474054
rect 113302 473818 113334 474054
rect 112714 438374 113334 473818
rect 112714 438138 112746 438374
rect 112982 438138 113066 438374
rect 113302 438138 113334 438374
rect 112714 438054 113334 438138
rect 112714 437818 112746 438054
rect 112982 437818 113066 438054
rect 113302 437818 113334 438054
rect 112714 402374 113334 437818
rect 112714 402138 112746 402374
rect 112982 402138 113066 402374
rect 113302 402138 113334 402374
rect 112714 402054 113334 402138
rect 112714 401818 112746 402054
rect 112982 401818 113066 402054
rect 113302 401818 113334 402054
rect 112714 366374 113334 401818
rect 112714 366138 112746 366374
rect 112982 366138 113066 366374
rect 113302 366138 113334 366374
rect 112714 366054 113334 366138
rect 112714 365818 112746 366054
rect 112982 365818 113066 366054
rect 113302 365818 113334 366054
rect 112714 330374 113334 365818
rect 112714 330138 112746 330374
rect 112982 330138 113066 330374
rect 113302 330138 113334 330374
rect 112714 330054 113334 330138
rect 112714 329818 112746 330054
rect 112982 329818 113066 330054
rect 113302 329818 113334 330054
rect 112714 294374 113334 329818
rect 112714 294138 112746 294374
rect 112982 294138 113066 294374
rect 113302 294138 113334 294374
rect 112714 294054 113334 294138
rect 112714 293818 112746 294054
rect 112982 293818 113066 294054
rect 113302 293818 113334 294054
rect 112714 258374 113334 293818
rect 112714 258138 112746 258374
rect 112982 258138 113066 258374
rect 113302 258138 113334 258374
rect 112714 258054 113334 258138
rect 112714 257818 112746 258054
rect 112982 257818 113066 258054
rect 113302 257818 113334 258054
rect 112714 222374 113334 257818
rect 112714 222138 112746 222374
rect 112982 222138 113066 222374
rect 113302 222138 113334 222374
rect 112714 222054 113334 222138
rect 112714 221818 112746 222054
rect 112982 221818 113066 222054
rect 113302 221818 113334 222054
rect 112714 186374 113334 221818
rect 112714 186138 112746 186374
rect 112982 186138 113066 186374
rect 113302 186138 113334 186374
rect 112714 186054 113334 186138
rect 112714 185818 112746 186054
rect 112982 185818 113066 186054
rect 113302 185818 113334 186054
rect 112714 150374 113334 185818
rect 112714 150138 112746 150374
rect 112982 150138 113066 150374
rect 113302 150138 113334 150374
rect 112714 150054 113334 150138
rect 112714 149818 112746 150054
rect 112982 149818 113066 150054
rect 113302 149818 113334 150054
rect 112714 114374 113334 149818
rect 112714 114138 112746 114374
rect 112982 114138 113066 114374
rect 113302 114138 113334 114374
rect 112714 114054 113334 114138
rect 112714 113818 112746 114054
rect 112982 113818 113066 114054
rect 113302 113818 113334 114054
rect 112714 78374 113334 113818
rect 112714 78138 112746 78374
rect 112982 78138 113066 78374
rect 113302 78138 113334 78374
rect 112714 78054 113334 78138
rect 112714 77818 112746 78054
rect 112982 77818 113066 78054
rect 113302 77818 113334 78054
rect 112714 42374 113334 77818
rect 112714 42138 112746 42374
rect 112982 42138 113066 42374
rect 113302 42138 113334 42374
rect 112714 42054 113334 42138
rect 112714 41818 112746 42054
rect 112982 41818 113066 42054
rect 113302 41818 113334 42054
rect 112714 6374 113334 41818
rect 112714 6138 112746 6374
rect 112982 6138 113066 6374
rect 113302 6138 113334 6374
rect 112714 6054 113334 6138
rect 112714 5818 112746 6054
rect 112982 5818 113066 6054
rect 113302 5818 113334 6054
rect 112714 -3226 113334 5818
rect 112714 -3462 112746 -3226
rect 112982 -3462 113066 -3226
rect 113302 -3462 113334 -3226
rect 112714 -3546 113334 -3462
rect 112714 -3782 112746 -3546
rect 112982 -3782 113066 -3546
rect 113302 -3782 113334 -3546
rect 112714 -7654 113334 -3782
rect 113954 708678 114574 711590
rect 113954 708442 113986 708678
rect 114222 708442 114306 708678
rect 114542 708442 114574 708678
rect 113954 708358 114574 708442
rect 113954 708122 113986 708358
rect 114222 708122 114306 708358
rect 114542 708122 114574 708358
rect 113954 691614 114574 708122
rect 113954 691378 113986 691614
rect 114222 691378 114306 691614
rect 114542 691378 114574 691614
rect 113954 691294 114574 691378
rect 113954 691058 113986 691294
rect 114222 691058 114306 691294
rect 114542 691058 114574 691294
rect 113954 655614 114574 691058
rect 113954 655378 113986 655614
rect 114222 655378 114306 655614
rect 114542 655378 114574 655614
rect 113954 655294 114574 655378
rect 113954 655058 113986 655294
rect 114222 655058 114306 655294
rect 114542 655058 114574 655294
rect 113954 619614 114574 655058
rect 113954 619378 113986 619614
rect 114222 619378 114306 619614
rect 114542 619378 114574 619614
rect 113954 619294 114574 619378
rect 113954 619058 113986 619294
rect 114222 619058 114306 619294
rect 114542 619058 114574 619294
rect 113954 583614 114574 619058
rect 113954 583378 113986 583614
rect 114222 583378 114306 583614
rect 114542 583378 114574 583614
rect 113954 583294 114574 583378
rect 113954 583058 113986 583294
rect 114222 583058 114306 583294
rect 114542 583058 114574 583294
rect 113954 547614 114574 583058
rect 113954 547378 113986 547614
rect 114222 547378 114306 547614
rect 114542 547378 114574 547614
rect 113954 547294 114574 547378
rect 113954 547058 113986 547294
rect 114222 547058 114306 547294
rect 114542 547058 114574 547294
rect 113954 511614 114574 547058
rect 113954 511378 113986 511614
rect 114222 511378 114306 511614
rect 114542 511378 114574 511614
rect 113954 511294 114574 511378
rect 113954 511058 113986 511294
rect 114222 511058 114306 511294
rect 114542 511058 114574 511294
rect 113954 475614 114574 511058
rect 113954 475378 113986 475614
rect 114222 475378 114306 475614
rect 114542 475378 114574 475614
rect 113954 475294 114574 475378
rect 113954 475058 113986 475294
rect 114222 475058 114306 475294
rect 114542 475058 114574 475294
rect 113954 439614 114574 475058
rect 113954 439378 113986 439614
rect 114222 439378 114306 439614
rect 114542 439378 114574 439614
rect 113954 439294 114574 439378
rect 113954 439058 113986 439294
rect 114222 439058 114306 439294
rect 114542 439058 114574 439294
rect 113954 403614 114574 439058
rect 113954 403378 113986 403614
rect 114222 403378 114306 403614
rect 114542 403378 114574 403614
rect 113954 403294 114574 403378
rect 113954 403058 113986 403294
rect 114222 403058 114306 403294
rect 114542 403058 114574 403294
rect 113954 367614 114574 403058
rect 113954 367378 113986 367614
rect 114222 367378 114306 367614
rect 114542 367378 114574 367614
rect 113954 367294 114574 367378
rect 113954 367058 113986 367294
rect 114222 367058 114306 367294
rect 114542 367058 114574 367294
rect 113954 331614 114574 367058
rect 113954 331378 113986 331614
rect 114222 331378 114306 331614
rect 114542 331378 114574 331614
rect 113954 331294 114574 331378
rect 113954 331058 113986 331294
rect 114222 331058 114306 331294
rect 114542 331058 114574 331294
rect 113954 295614 114574 331058
rect 113954 295378 113986 295614
rect 114222 295378 114306 295614
rect 114542 295378 114574 295614
rect 113954 295294 114574 295378
rect 113954 295058 113986 295294
rect 114222 295058 114306 295294
rect 114542 295058 114574 295294
rect 113954 259614 114574 295058
rect 113954 259378 113986 259614
rect 114222 259378 114306 259614
rect 114542 259378 114574 259614
rect 113954 259294 114574 259378
rect 113954 259058 113986 259294
rect 114222 259058 114306 259294
rect 114542 259058 114574 259294
rect 113954 223614 114574 259058
rect 113954 223378 113986 223614
rect 114222 223378 114306 223614
rect 114542 223378 114574 223614
rect 113954 223294 114574 223378
rect 113954 223058 113986 223294
rect 114222 223058 114306 223294
rect 114542 223058 114574 223294
rect 113954 187614 114574 223058
rect 113954 187378 113986 187614
rect 114222 187378 114306 187614
rect 114542 187378 114574 187614
rect 113954 187294 114574 187378
rect 113954 187058 113986 187294
rect 114222 187058 114306 187294
rect 114542 187058 114574 187294
rect 113954 151614 114574 187058
rect 113954 151378 113986 151614
rect 114222 151378 114306 151614
rect 114542 151378 114574 151614
rect 113954 151294 114574 151378
rect 113954 151058 113986 151294
rect 114222 151058 114306 151294
rect 114542 151058 114574 151294
rect 113954 115614 114574 151058
rect 113954 115378 113986 115614
rect 114222 115378 114306 115614
rect 114542 115378 114574 115614
rect 113954 115294 114574 115378
rect 113954 115058 113986 115294
rect 114222 115058 114306 115294
rect 114542 115058 114574 115294
rect 113954 79614 114574 115058
rect 113954 79378 113986 79614
rect 114222 79378 114306 79614
rect 114542 79378 114574 79614
rect 113954 79294 114574 79378
rect 113954 79058 113986 79294
rect 114222 79058 114306 79294
rect 114542 79058 114574 79294
rect 113954 43614 114574 79058
rect 113954 43378 113986 43614
rect 114222 43378 114306 43614
rect 114542 43378 114574 43614
rect 113954 43294 114574 43378
rect 113954 43058 113986 43294
rect 114222 43058 114306 43294
rect 114542 43058 114574 43294
rect 113954 7614 114574 43058
rect 113954 7378 113986 7614
rect 114222 7378 114306 7614
rect 114542 7378 114574 7614
rect 113954 7294 114574 7378
rect 113954 7058 113986 7294
rect 114222 7058 114306 7294
rect 114542 7058 114574 7294
rect 113954 -4186 114574 7058
rect 113954 -4422 113986 -4186
rect 114222 -4422 114306 -4186
rect 114542 -4422 114574 -4186
rect 113954 -4506 114574 -4422
rect 113954 -4742 113986 -4506
rect 114222 -4742 114306 -4506
rect 114542 -4742 114574 -4506
rect 113954 -7654 114574 -4742
rect 115194 709638 115814 711590
rect 115194 709402 115226 709638
rect 115462 709402 115546 709638
rect 115782 709402 115814 709638
rect 115194 709318 115814 709402
rect 115194 709082 115226 709318
rect 115462 709082 115546 709318
rect 115782 709082 115814 709318
rect 115194 692854 115814 709082
rect 115194 692618 115226 692854
rect 115462 692618 115546 692854
rect 115782 692618 115814 692854
rect 115194 692534 115814 692618
rect 115194 692298 115226 692534
rect 115462 692298 115546 692534
rect 115782 692298 115814 692534
rect 115194 656854 115814 692298
rect 115194 656618 115226 656854
rect 115462 656618 115546 656854
rect 115782 656618 115814 656854
rect 115194 656534 115814 656618
rect 115194 656298 115226 656534
rect 115462 656298 115546 656534
rect 115782 656298 115814 656534
rect 115194 620854 115814 656298
rect 115194 620618 115226 620854
rect 115462 620618 115546 620854
rect 115782 620618 115814 620854
rect 115194 620534 115814 620618
rect 115194 620298 115226 620534
rect 115462 620298 115546 620534
rect 115782 620298 115814 620534
rect 115194 584854 115814 620298
rect 115194 584618 115226 584854
rect 115462 584618 115546 584854
rect 115782 584618 115814 584854
rect 115194 584534 115814 584618
rect 115194 584298 115226 584534
rect 115462 584298 115546 584534
rect 115782 584298 115814 584534
rect 115194 548854 115814 584298
rect 115194 548618 115226 548854
rect 115462 548618 115546 548854
rect 115782 548618 115814 548854
rect 115194 548534 115814 548618
rect 115194 548298 115226 548534
rect 115462 548298 115546 548534
rect 115782 548298 115814 548534
rect 115194 512854 115814 548298
rect 115194 512618 115226 512854
rect 115462 512618 115546 512854
rect 115782 512618 115814 512854
rect 115194 512534 115814 512618
rect 115194 512298 115226 512534
rect 115462 512298 115546 512534
rect 115782 512298 115814 512534
rect 115194 476854 115814 512298
rect 115194 476618 115226 476854
rect 115462 476618 115546 476854
rect 115782 476618 115814 476854
rect 115194 476534 115814 476618
rect 115194 476298 115226 476534
rect 115462 476298 115546 476534
rect 115782 476298 115814 476534
rect 115194 440854 115814 476298
rect 115194 440618 115226 440854
rect 115462 440618 115546 440854
rect 115782 440618 115814 440854
rect 115194 440534 115814 440618
rect 115194 440298 115226 440534
rect 115462 440298 115546 440534
rect 115782 440298 115814 440534
rect 115194 404854 115814 440298
rect 115194 404618 115226 404854
rect 115462 404618 115546 404854
rect 115782 404618 115814 404854
rect 115194 404534 115814 404618
rect 115194 404298 115226 404534
rect 115462 404298 115546 404534
rect 115782 404298 115814 404534
rect 115194 368854 115814 404298
rect 115194 368618 115226 368854
rect 115462 368618 115546 368854
rect 115782 368618 115814 368854
rect 115194 368534 115814 368618
rect 115194 368298 115226 368534
rect 115462 368298 115546 368534
rect 115782 368298 115814 368534
rect 115194 332854 115814 368298
rect 115194 332618 115226 332854
rect 115462 332618 115546 332854
rect 115782 332618 115814 332854
rect 115194 332534 115814 332618
rect 115194 332298 115226 332534
rect 115462 332298 115546 332534
rect 115782 332298 115814 332534
rect 115194 296854 115814 332298
rect 115194 296618 115226 296854
rect 115462 296618 115546 296854
rect 115782 296618 115814 296854
rect 115194 296534 115814 296618
rect 115194 296298 115226 296534
rect 115462 296298 115546 296534
rect 115782 296298 115814 296534
rect 115194 260854 115814 296298
rect 115194 260618 115226 260854
rect 115462 260618 115546 260854
rect 115782 260618 115814 260854
rect 115194 260534 115814 260618
rect 115194 260298 115226 260534
rect 115462 260298 115546 260534
rect 115782 260298 115814 260534
rect 115194 224854 115814 260298
rect 115194 224618 115226 224854
rect 115462 224618 115546 224854
rect 115782 224618 115814 224854
rect 115194 224534 115814 224618
rect 115194 224298 115226 224534
rect 115462 224298 115546 224534
rect 115782 224298 115814 224534
rect 115194 188854 115814 224298
rect 115194 188618 115226 188854
rect 115462 188618 115546 188854
rect 115782 188618 115814 188854
rect 115194 188534 115814 188618
rect 115194 188298 115226 188534
rect 115462 188298 115546 188534
rect 115782 188298 115814 188534
rect 115194 152854 115814 188298
rect 115194 152618 115226 152854
rect 115462 152618 115546 152854
rect 115782 152618 115814 152854
rect 115194 152534 115814 152618
rect 115194 152298 115226 152534
rect 115462 152298 115546 152534
rect 115782 152298 115814 152534
rect 115194 116854 115814 152298
rect 115194 116618 115226 116854
rect 115462 116618 115546 116854
rect 115782 116618 115814 116854
rect 115194 116534 115814 116618
rect 115194 116298 115226 116534
rect 115462 116298 115546 116534
rect 115782 116298 115814 116534
rect 115194 80854 115814 116298
rect 115194 80618 115226 80854
rect 115462 80618 115546 80854
rect 115782 80618 115814 80854
rect 115194 80534 115814 80618
rect 115194 80298 115226 80534
rect 115462 80298 115546 80534
rect 115782 80298 115814 80534
rect 115194 44854 115814 80298
rect 115194 44618 115226 44854
rect 115462 44618 115546 44854
rect 115782 44618 115814 44854
rect 115194 44534 115814 44618
rect 115194 44298 115226 44534
rect 115462 44298 115546 44534
rect 115782 44298 115814 44534
rect 115194 8854 115814 44298
rect 115194 8618 115226 8854
rect 115462 8618 115546 8854
rect 115782 8618 115814 8854
rect 115194 8534 115814 8618
rect 115194 8298 115226 8534
rect 115462 8298 115546 8534
rect 115782 8298 115814 8534
rect 115194 -5146 115814 8298
rect 115194 -5382 115226 -5146
rect 115462 -5382 115546 -5146
rect 115782 -5382 115814 -5146
rect 115194 -5466 115814 -5382
rect 115194 -5702 115226 -5466
rect 115462 -5702 115546 -5466
rect 115782 -5702 115814 -5466
rect 115194 -7654 115814 -5702
rect 116434 710598 117054 711590
rect 116434 710362 116466 710598
rect 116702 710362 116786 710598
rect 117022 710362 117054 710598
rect 116434 710278 117054 710362
rect 116434 710042 116466 710278
rect 116702 710042 116786 710278
rect 117022 710042 117054 710278
rect 116434 694094 117054 710042
rect 116434 693858 116466 694094
rect 116702 693858 116786 694094
rect 117022 693858 117054 694094
rect 116434 693774 117054 693858
rect 116434 693538 116466 693774
rect 116702 693538 116786 693774
rect 117022 693538 117054 693774
rect 116434 658094 117054 693538
rect 116434 657858 116466 658094
rect 116702 657858 116786 658094
rect 117022 657858 117054 658094
rect 116434 657774 117054 657858
rect 116434 657538 116466 657774
rect 116702 657538 116786 657774
rect 117022 657538 117054 657774
rect 116434 622094 117054 657538
rect 116434 621858 116466 622094
rect 116702 621858 116786 622094
rect 117022 621858 117054 622094
rect 116434 621774 117054 621858
rect 116434 621538 116466 621774
rect 116702 621538 116786 621774
rect 117022 621538 117054 621774
rect 116434 586094 117054 621538
rect 116434 585858 116466 586094
rect 116702 585858 116786 586094
rect 117022 585858 117054 586094
rect 116434 585774 117054 585858
rect 116434 585538 116466 585774
rect 116702 585538 116786 585774
rect 117022 585538 117054 585774
rect 116434 550094 117054 585538
rect 116434 549858 116466 550094
rect 116702 549858 116786 550094
rect 117022 549858 117054 550094
rect 116434 549774 117054 549858
rect 116434 549538 116466 549774
rect 116702 549538 116786 549774
rect 117022 549538 117054 549774
rect 116434 514094 117054 549538
rect 116434 513858 116466 514094
rect 116702 513858 116786 514094
rect 117022 513858 117054 514094
rect 116434 513774 117054 513858
rect 116434 513538 116466 513774
rect 116702 513538 116786 513774
rect 117022 513538 117054 513774
rect 116434 478094 117054 513538
rect 116434 477858 116466 478094
rect 116702 477858 116786 478094
rect 117022 477858 117054 478094
rect 116434 477774 117054 477858
rect 116434 477538 116466 477774
rect 116702 477538 116786 477774
rect 117022 477538 117054 477774
rect 116434 442094 117054 477538
rect 116434 441858 116466 442094
rect 116702 441858 116786 442094
rect 117022 441858 117054 442094
rect 116434 441774 117054 441858
rect 116434 441538 116466 441774
rect 116702 441538 116786 441774
rect 117022 441538 117054 441774
rect 116434 406094 117054 441538
rect 116434 405858 116466 406094
rect 116702 405858 116786 406094
rect 117022 405858 117054 406094
rect 116434 405774 117054 405858
rect 116434 405538 116466 405774
rect 116702 405538 116786 405774
rect 117022 405538 117054 405774
rect 116434 370094 117054 405538
rect 116434 369858 116466 370094
rect 116702 369858 116786 370094
rect 117022 369858 117054 370094
rect 116434 369774 117054 369858
rect 116434 369538 116466 369774
rect 116702 369538 116786 369774
rect 117022 369538 117054 369774
rect 116434 334094 117054 369538
rect 116434 333858 116466 334094
rect 116702 333858 116786 334094
rect 117022 333858 117054 334094
rect 116434 333774 117054 333858
rect 116434 333538 116466 333774
rect 116702 333538 116786 333774
rect 117022 333538 117054 333774
rect 116434 298094 117054 333538
rect 116434 297858 116466 298094
rect 116702 297858 116786 298094
rect 117022 297858 117054 298094
rect 116434 297774 117054 297858
rect 116434 297538 116466 297774
rect 116702 297538 116786 297774
rect 117022 297538 117054 297774
rect 116434 262094 117054 297538
rect 116434 261858 116466 262094
rect 116702 261858 116786 262094
rect 117022 261858 117054 262094
rect 116434 261774 117054 261858
rect 116434 261538 116466 261774
rect 116702 261538 116786 261774
rect 117022 261538 117054 261774
rect 116434 226094 117054 261538
rect 116434 225858 116466 226094
rect 116702 225858 116786 226094
rect 117022 225858 117054 226094
rect 116434 225774 117054 225858
rect 116434 225538 116466 225774
rect 116702 225538 116786 225774
rect 117022 225538 117054 225774
rect 116434 190094 117054 225538
rect 116434 189858 116466 190094
rect 116702 189858 116786 190094
rect 117022 189858 117054 190094
rect 116434 189774 117054 189858
rect 116434 189538 116466 189774
rect 116702 189538 116786 189774
rect 117022 189538 117054 189774
rect 116434 154094 117054 189538
rect 116434 153858 116466 154094
rect 116702 153858 116786 154094
rect 117022 153858 117054 154094
rect 116434 153774 117054 153858
rect 116434 153538 116466 153774
rect 116702 153538 116786 153774
rect 117022 153538 117054 153774
rect 116434 118094 117054 153538
rect 116434 117858 116466 118094
rect 116702 117858 116786 118094
rect 117022 117858 117054 118094
rect 116434 117774 117054 117858
rect 116434 117538 116466 117774
rect 116702 117538 116786 117774
rect 117022 117538 117054 117774
rect 116434 82094 117054 117538
rect 116434 81858 116466 82094
rect 116702 81858 116786 82094
rect 117022 81858 117054 82094
rect 116434 81774 117054 81858
rect 116434 81538 116466 81774
rect 116702 81538 116786 81774
rect 117022 81538 117054 81774
rect 116434 46094 117054 81538
rect 116434 45858 116466 46094
rect 116702 45858 116786 46094
rect 117022 45858 117054 46094
rect 116434 45774 117054 45858
rect 116434 45538 116466 45774
rect 116702 45538 116786 45774
rect 117022 45538 117054 45774
rect 116434 10094 117054 45538
rect 116434 9858 116466 10094
rect 116702 9858 116786 10094
rect 117022 9858 117054 10094
rect 116434 9774 117054 9858
rect 116434 9538 116466 9774
rect 116702 9538 116786 9774
rect 117022 9538 117054 9774
rect 116434 -6106 117054 9538
rect 116434 -6342 116466 -6106
rect 116702 -6342 116786 -6106
rect 117022 -6342 117054 -6106
rect 116434 -6426 117054 -6342
rect 116434 -6662 116466 -6426
rect 116702 -6662 116786 -6426
rect 117022 -6662 117054 -6426
rect 116434 -7654 117054 -6662
rect 117674 711558 118294 711590
rect 117674 711322 117706 711558
rect 117942 711322 118026 711558
rect 118262 711322 118294 711558
rect 117674 711238 118294 711322
rect 117674 711002 117706 711238
rect 117942 711002 118026 711238
rect 118262 711002 118294 711238
rect 117674 695334 118294 711002
rect 117674 695098 117706 695334
rect 117942 695098 118026 695334
rect 118262 695098 118294 695334
rect 117674 695014 118294 695098
rect 117674 694778 117706 695014
rect 117942 694778 118026 695014
rect 118262 694778 118294 695014
rect 117674 659334 118294 694778
rect 117674 659098 117706 659334
rect 117942 659098 118026 659334
rect 118262 659098 118294 659334
rect 117674 659014 118294 659098
rect 117674 658778 117706 659014
rect 117942 658778 118026 659014
rect 118262 658778 118294 659014
rect 117674 623334 118294 658778
rect 117674 623098 117706 623334
rect 117942 623098 118026 623334
rect 118262 623098 118294 623334
rect 117674 623014 118294 623098
rect 117674 622778 117706 623014
rect 117942 622778 118026 623014
rect 118262 622778 118294 623014
rect 117674 587334 118294 622778
rect 117674 587098 117706 587334
rect 117942 587098 118026 587334
rect 118262 587098 118294 587334
rect 117674 587014 118294 587098
rect 117674 586778 117706 587014
rect 117942 586778 118026 587014
rect 118262 586778 118294 587014
rect 117674 551334 118294 586778
rect 117674 551098 117706 551334
rect 117942 551098 118026 551334
rect 118262 551098 118294 551334
rect 117674 551014 118294 551098
rect 117674 550778 117706 551014
rect 117942 550778 118026 551014
rect 118262 550778 118294 551014
rect 117674 515334 118294 550778
rect 117674 515098 117706 515334
rect 117942 515098 118026 515334
rect 118262 515098 118294 515334
rect 117674 515014 118294 515098
rect 117674 514778 117706 515014
rect 117942 514778 118026 515014
rect 118262 514778 118294 515014
rect 117674 479334 118294 514778
rect 117674 479098 117706 479334
rect 117942 479098 118026 479334
rect 118262 479098 118294 479334
rect 117674 479014 118294 479098
rect 117674 478778 117706 479014
rect 117942 478778 118026 479014
rect 118262 478778 118294 479014
rect 117674 443334 118294 478778
rect 117674 443098 117706 443334
rect 117942 443098 118026 443334
rect 118262 443098 118294 443334
rect 117674 443014 118294 443098
rect 117674 442778 117706 443014
rect 117942 442778 118026 443014
rect 118262 442778 118294 443014
rect 117674 407334 118294 442778
rect 117674 407098 117706 407334
rect 117942 407098 118026 407334
rect 118262 407098 118294 407334
rect 117674 407014 118294 407098
rect 117674 406778 117706 407014
rect 117942 406778 118026 407014
rect 118262 406778 118294 407014
rect 117674 371334 118294 406778
rect 117674 371098 117706 371334
rect 117942 371098 118026 371334
rect 118262 371098 118294 371334
rect 117674 371014 118294 371098
rect 117674 370778 117706 371014
rect 117942 370778 118026 371014
rect 118262 370778 118294 371014
rect 117674 335334 118294 370778
rect 117674 335098 117706 335334
rect 117942 335098 118026 335334
rect 118262 335098 118294 335334
rect 117674 335014 118294 335098
rect 117674 334778 117706 335014
rect 117942 334778 118026 335014
rect 118262 334778 118294 335014
rect 117674 299334 118294 334778
rect 117674 299098 117706 299334
rect 117942 299098 118026 299334
rect 118262 299098 118294 299334
rect 117674 299014 118294 299098
rect 117674 298778 117706 299014
rect 117942 298778 118026 299014
rect 118262 298778 118294 299014
rect 117674 263334 118294 298778
rect 117674 263098 117706 263334
rect 117942 263098 118026 263334
rect 118262 263098 118294 263334
rect 117674 263014 118294 263098
rect 117674 262778 117706 263014
rect 117942 262778 118026 263014
rect 118262 262778 118294 263014
rect 117674 227334 118294 262778
rect 117674 227098 117706 227334
rect 117942 227098 118026 227334
rect 118262 227098 118294 227334
rect 117674 227014 118294 227098
rect 117674 226778 117706 227014
rect 117942 226778 118026 227014
rect 118262 226778 118294 227014
rect 117674 191334 118294 226778
rect 117674 191098 117706 191334
rect 117942 191098 118026 191334
rect 118262 191098 118294 191334
rect 117674 191014 118294 191098
rect 117674 190778 117706 191014
rect 117942 190778 118026 191014
rect 118262 190778 118294 191014
rect 117674 155334 118294 190778
rect 117674 155098 117706 155334
rect 117942 155098 118026 155334
rect 118262 155098 118294 155334
rect 117674 155014 118294 155098
rect 117674 154778 117706 155014
rect 117942 154778 118026 155014
rect 118262 154778 118294 155014
rect 117674 119334 118294 154778
rect 117674 119098 117706 119334
rect 117942 119098 118026 119334
rect 118262 119098 118294 119334
rect 117674 119014 118294 119098
rect 117674 118778 117706 119014
rect 117942 118778 118026 119014
rect 118262 118778 118294 119014
rect 117674 83334 118294 118778
rect 117674 83098 117706 83334
rect 117942 83098 118026 83334
rect 118262 83098 118294 83334
rect 117674 83014 118294 83098
rect 117674 82778 117706 83014
rect 117942 82778 118026 83014
rect 118262 82778 118294 83014
rect 117674 47334 118294 82778
rect 117674 47098 117706 47334
rect 117942 47098 118026 47334
rect 118262 47098 118294 47334
rect 117674 47014 118294 47098
rect 117674 46778 117706 47014
rect 117942 46778 118026 47014
rect 118262 46778 118294 47014
rect 117674 11334 118294 46778
rect 117674 11098 117706 11334
rect 117942 11098 118026 11334
rect 118262 11098 118294 11334
rect 117674 11014 118294 11098
rect 117674 10778 117706 11014
rect 117942 10778 118026 11014
rect 118262 10778 118294 11014
rect 117674 -7066 118294 10778
rect 117674 -7302 117706 -7066
rect 117942 -7302 118026 -7066
rect 118262 -7302 118294 -7066
rect 117674 -7386 118294 -7302
rect 117674 -7622 117706 -7386
rect 117942 -7622 118026 -7386
rect 118262 -7622 118294 -7386
rect 117674 -7654 118294 -7622
rect 144994 704838 145614 711590
rect 144994 704602 145026 704838
rect 145262 704602 145346 704838
rect 145582 704602 145614 704838
rect 144994 704518 145614 704602
rect 144994 704282 145026 704518
rect 145262 704282 145346 704518
rect 145582 704282 145614 704518
rect 144994 686654 145614 704282
rect 144994 686418 145026 686654
rect 145262 686418 145346 686654
rect 145582 686418 145614 686654
rect 144994 686334 145614 686418
rect 144994 686098 145026 686334
rect 145262 686098 145346 686334
rect 145582 686098 145614 686334
rect 144994 650654 145614 686098
rect 144994 650418 145026 650654
rect 145262 650418 145346 650654
rect 145582 650418 145614 650654
rect 144994 650334 145614 650418
rect 144994 650098 145026 650334
rect 145262 650098 145346 650334
rect 145582 650098 145614 650334
rect 144994 614654 145614 650098
rect 144994 614418 145026 614654
rect 145262 614418 145346 614654
rect 145582 614418 145614 614654
rect 144994 614334 145614 614418
rect 144994 614098 145026 614334
rect 145262 614098 145346 614334
rect 145582 614098 145614 614334
rect 144994 578654 145614 614098
rect 144994 578418 145026 578654
rect 145262 578418 145346 578654
rect 145582 578418 145614 578654
rect 144994 578334 145614 578418
rect 144994 578098 145026 578334
rect 145262 578098 145346 578334
rect 145582 578098 145614 578334
rect 144994 542654 145614 578098
rect 144994 542418 145026 542654
rect 145262 542418 145346 542654
rect 145582 542418 145614 542654
rect 144994 542334 145614 542418
rect 144994 542098 145026 542334
rect 145262 542098 145346 542334
rect 145582 542098 145614 542334
rect 144994 506654 145614 542098
rect 144994 506418 145026 506654
rect 145262 506418 145346 506654
rect 145582 506418 145614 506654
rect 144994 506334 145614 506418
rect 144994 506098 145026 506334
rect 145262 506098 145346 506334
rect 145582 506098 145614 506334
rect 144994 470654 145614 506098
rect 144994 470418 145026 470654
rect 145262 470418 145346 470654
rect 145582 470418 145614 470654
rect 144994 470334 145614 470418
rect 144994 470098 145026 470334
rect 145262 470098 145346 470334
rect 145582 470098 145614 470334
rect 144994 434654 145614 470098
rect 144994 434418 145026 434654
rect 145262 434418 145346 434654
rect 145582 434418 145614 434654
rect 144994 434334 145614 434418
rect 144994 434098 145026 434334
rect 145262 434098 145346 434334
rect 145582 434098 145614 434334
rect 144994 398654 145614 434098
rect 144994 398418 145026 398654
rect 145262 398418 145346 398654
rect 145582 398418 145614 398654
rect 144994 398334 145614 398418
rect 144994 398098 145026 398334
rect 145262 398098 145346 398334
rect 145582 398098 145614 398334
rect 144994 362654 145614 398098
rect 144994 362418 145026 362654
rect 145262 362418 145346 362654
rect 145582 362418 145614 362654
rect 144994 362334 145614 362418
rect 144994 362098 145026 362334
rect 145262 362098 145346 362334
rect 145582 362098 145614 362334
rect 144994 326654 145614 362098
rect 144994 326418 145026 326654
rect 145262 326418 145346 326654
rect 145582 326418 145614 326654
rect 144994 326334 145614 326418
rect 144994 326098 145026 326334
rect 145262 326098 145346 326334
rect 145582 326098 145614 326334
rect 144994 290654 145614 326098
rect 144994 290418 145026 290654
rect 145262 290418 145346 290654
rect 145582 290418 145614 290654
rect 144994 290334 145614 290418
rect 144994 290098 145026 290334
rect 145262 290098 145346 290334
rect 145582 290098 145614 290334
rect 144994 254654 145614 290098
rect 144994 254418 145026 254654
rect 145262 254418 145346 254654
rect 145582 254418 145614 254654
rect 144994 254334 145614 254418
rect 144994 254098 145026 254334
rect 145262 254098 145346 254334
rect 145582 254098 145614 254334
rect 144994 218654 145614 254098
rect 144994 218418 145026 218654
rect 145262 218418 145346 218654
rect 145582 218418 145614 218654
rect 144994 218334 145614 218418
rect 144994 218098 145026 218334
rect 145262 218098 145346 218334
rect 145582 218098 145614 218334
rect 144994 182654 145614 218098
rect 144994 182418 145026 182654
rect 145262 182418 145346 182654
rect 145582 182418 145614 182654
rect 144994 182334 145614 182418
rect 144994 182098 145026 182334
rect 145262 182098 145346 182334
rect 145582 182098 145614 182334
rect 144994 146654 145614 182098
rect 144994 146418 145026 146654
rect 145262 146418 145346 146654
rect 145582 146418 145614 146654
rect 144994 146334 145614 146418
rect 144994 146098 145026 146334
rect 145262 146098 145346 146334
rect 145582 146098 145614 146334
rect 144994 110654 145614 146098
rect 144994 110418 145026 110654
rect 145262 110418 145346 110654
rect 145582 110418 145614 110654
rect 144994 110334 145614 110418
rect 144994 110098 145026 110334
rect 145262 110098 145346 110334
rect 145582 110098 145614 110334
rect 144994 74654 145614 110098
rect 144994 74418 145026 74654
rect 145262 74418 145346 74654
rect 145582 74418 145614 74654
rect 144994 74334 145614 74418
rect 144994 74098 145026 74334
rect 145262 74098 145346 74334
rect 145582 74098 145614 74334
rect 144994 38654 145614 74098
rect 144994 38418 145026 38654
rect 145262 38418 145346 38654
rect 145582 38418 145614 38654
rect 144994 38334 145614 38418
rect 144994 38098 145026 38334
rect 145262 38098 145346 38334
rect 145582 38098 145614 38334
rect 144994 2654 145614 38098
rect 144994 2418 145026 2654
rect 145262 2418 145346 2654
rect 145582 2418 145614 2654
rect 144994 2334 145614 2418
rect 144994 2098 145026 2334
rect 145262 2098 145346 2334
rect 145582 2098 145614 2334
rect 144994 -346 145614 2098
rect 144994 -582 145026 -346
rect 145262 -582 145346 -346
rect 145582 -582 145614 -346
rect 144994 -666 145614 -582
rect 144994 -902 145026 -666
rect 145262 -902 145346 -666
rect 145582 -902 145614 -666
rect 144994 -7654 145614 -902
rect 146234 705798 146854 711590
rect 146234 705562 146266 705798
rect 146502 705562 146586 705798
rect 146822 705562 146854 705798
rect 146234 705478 146854 705562
rect 146234 705242 146266 705478
rect 146502 705242 146586 705478
rect 146822 705242 146854 705478
rect 146234 687894 146854 705242
rect 146234 687658 146266 687894
rect 146502 687658 146586 687894
rect 146822 687658 146854 687894
rect 146234 687574 146854 687658
rect 146234 687338 146266 687574
rect 146502 687338 146586 687574
rect 146822 687338 146854 687574
rect 146234 651894 146854 687338
rect 146234 651658 146266 651894
rect 146502 651658 146586 651894
rect 146822 651658 146854 651894
rect 146234 651574 146854 651658
rect 146234 651338 146266 651574
rect 146502 651338 146586 651574
rect 146822 651338 146854 651574
rect 146234 615894 146854 651338
rect 146234 615658 146266 615894
rect 146502 615658 146586 615894
rect 146822 615658 146854 615894
rect 146234 615574 146854 615658
rect 146234 615338 146266 615574
rect 146502 615338 146586 615574
rect 146822 615338 146854 615574
rect 146234 579894 146854 615338
rect 146234 579658 146266 579894
rect 146502 579658 146586 579894
rect 146822 579658 146854 579894
rect 146234 579574 146854 579658
rect 146234 579338 146266 579574
rect 146502 579338 146586 579574
rect 146822 579338 146854 579574
rect 146234 543894 146854 579338
rect 146234 543658 146266 543894
rect 146502 543658 146586 543894
rect 146822 543658 146854 543894
rect 146234 543574 146854 543658
rect 146234 543338 146266 543574
rect 146502 543338 146586 543574
rect 146822 543338 146854 543574
rect 146234 507894 146854 543338
rect 146234 507658 146266 507894
rect 146502 507658 146586 507894
rect 146822 507658 146854 507894
rect 146234 507574 146854 507658
rect 146234 507338 146266 507574
rect 146502 507338 146586 507574
rect 146822 507338 146854 507574
rect 146234 471894 146854 507338
rect 146234 471658 146266 471894
rect 146502 471658 146586 471894
rect 146822 471658 146854 471894
rect 146234 471574 146854 471658
rect 146234 471338 146266 471574
rect 146502 471338 146586 471574
rect 146822 471338 146854 471574
rect 146234 435894 146854 471338
rect 146234 435658 146266 435894
rect 146502 435658 146586 435894
rect 146822 435658 146854 435894
rect 146234 435574 146854 435658
rect 146234 435338 146266 435574
rect 146502 435338 146586 435574
rect 146822 435338 146854 435574
rect 146234 399894 146854 435338
rect 146234 399658 146266 399894
rect 146502 399658 146586 399894
rect 146822 399658 146854 399894
rect 146234 399574 146854 399658
rect 146234 399338 146266 399574
rect 146502 399338 146586 399574
rect 146822 399338 146854 399574
rect 146234 363894 146854 399338
rect 146234 363658 146266 363894
rect 146502 363658 146586 363894
rect 146822 363658 146854 363894
rect 146234 363574 146854 363658
rect 146234 363338 146266 363574
rect 146502 363338 146586 363574
rect 146822 363338 146854 363574
rect 146234 327894 146854 363338
rect 146234 327658 146266 327894
rect 146502 327658 146586 327894
rect 146822 327658 146854 327894
rect 146234 327574 146854 327658
rect 146234 327338 146266 327574
rect 146502 327338 146586 327574
rect 146822 327338 146854 327574
rect 146234 291894 146854 327338
rect 146234 291658 146266 291894
rect 146502 291658 146586 291894
rect 146822 291658 146854 291894
rect 146234 291574 146854 291658
rect 146234 291338 146266 291574
rect 146502 291338 146586 291574
rect 146822 291338 146854 291574
rect 146234 255894 146854 291338
rect 146234 255658 146266 255894
rect 146502 255658 146586 255894
rect 146822 255658 146854 255894
rect 146234 255574 146854 255658
rect 146234 255338 146266 255574
rect 146502 255338 146586 255574
rect 146822 255338 146854 255574
rect 146234 219894 146854 255338
rect 146234 219658 146266 219894
rect 146502 219658 146586 219894
rect 146822 219658 146854 219894
rect 146234 219574 146854 219658
rect 146234 219338 146266 219574
rect 146502 219338 146586 219574
rect 146822 219338 146854 219574
rect 146234 183894 146854 219338
rect 146234 183658 146266 183894
rect 146502 183658 146586 183894
rect 146822 183658 146854 183894
rect 146234 183574 146854 183658
rect 146234 183338 146266 183574
rect 146502 183338 146586 183574
rect 146822 183338 146854 183574
rect 146234 147894 146854 183338
rect 146234 147658 146266 147894
rect 146502 147658 146586 147894
rect 146822 147658 146854 147894
rect 146234 147574 146854 147658
rect 146234 147338 146266 147574
rect 146502 147338 146586 147574
rect 146822 147338 146854 147574
rect 146234 111894 146854 147338
rect 146234 111658 146266 111894
rect 146502 111658 146586 111894
rect 146822 111658 146854 111894
rect 146234 111574 146854 111658
rect 146234 111338 146266 111574
rect 146502 111338 146586 111574
rect 146822 111338 146854 111574
rect 146234 75894 146854 111338
rect 146234 75658 146266 75894
rect 146502 75658 146586 75894
rect 146822 75658 146854 75894
rect 146234 75574 146854 75658
rect 146234 75338 146266 75574
rect 146502 75338 146586 75574
rect 146822 75338 146854 75574
rect 146234 39894 146854 75338
rect 146234 39658 146266 39894
rect 146502 39658 146586 39894
rect 146822 39658 146854 39894
rect 146234 39574 146854 39658
rect 146234 39338 146266 39574
rect 146502 39338 146586 39574
rect 146822 39338 146854 39574
rect 146234 3894 146854 39338
rect 146234 3658 146266 3894
rect 146502 3658 146586 3894
rect 146822 3658 146854 3894
rect 146234 3574 146854 3658
rect 146234 3338 146266 3574
rect 146502 3338 146586 3574
rect 146822 3338 146854 3574
rect 146234 -1306 146854 3338
rect 146234 -1542 146266 -1306
rect 146502 -1542 146586 -1306
rect 146822 -1542 146854 -1306
rect 146234 -1626 146854 -1542
rect 146234 -1862 146266 -1626
rect 146502 -1862 146586 -1626
rect 146822 -1862 146854 -1626
rect 146234 -7654 146854 -1862
rect 147474 706758 148094 711590
rect 147474 706522 147506 706758
rect 147742 706522 147826 706758
rect 148062 706522 148094 706758
rect 147474 706438 148094 706522
rect 147474 706202 147506 706438
rect 147742 706202 147826 706438
rect 148062 706202 148094 706438
rect 147474 689134 148094 706202
rect 147474 688898 147506 689134
rect 147742 688898 147826 689134
rect 148062 688898 148094 689134
rect 147474 688814 148094 688898
rect 147474 688578 147506 688814
rect 147742 688578 147826 688814
rect 148062 688578 148094 688814
rect 147474 653134 148094 688578
rect 147474 652898 147506 653134
rect 147742 652898 147826 653134
rect 148062 652898 148094 653134
rect 147474 652814 148094 652898
rect 147474 652578 147506 652814
rect 147742 652578 147826 652814
rect 148062 652578 148094 652814
rect 147474 617134 148094 652578
rect 147474 616898 147506 617134
rect 147742 616898 147826 617134
rect 148062 616898 148094 617134
rect 147474 616814 148094 616898
rect 147474 616578 147506 616814
rect 147742 616578 147826 616814
rect 148062 616578 148094 616814
rect 147474 581134 148094 616578
rect 147474 580898 147506 581134
rect 147742 580898 147826 581134
rect 148062 580898 148094 581134
rect 147474 580814 148094 580898
rect 147474 580578 147506 580814
rect 147742 580578 147826 580814
rect 148062 580578 148094 580814
rect 147474 545134 148094 580578
rect 147474 544898 147506 545134
rect 147742 544898 147826 545134
rect 148062 544898 148094 545134
rect 147474 544814 148094 544898
rect 147474 544578 147506 544814
rect 147742 544578 147826 544814
rect 148062 544578 148094 544814
rect 147474 509134 148094 544578
rect 147474 508898 147506 509134
rect 147742 508898 147826 509134
rect 148062 508898 148094 509134
rect 147474 508814 148094 508898
rect 147474 508578 147506 508814
rect 147742 508578 147826 508814
rect 148062 508578 148094 508814
rect 147474 473134 148094 508578
rect 147474 472898 147506 473134
rect 147742 472898 147826 473134
rect 148062 472898 148094 473134
rect 147474 472814 148094 472898
rect 147474 472578 147506 472814
rect 147742 472578 147826 472814
rect 148062 472578 148094 472814
rect 147474 437134 148094 472578
rect 147474 436898 147506 437134
rect 147742 436898 147826 437134
rect 148062 436898 148094 437134
rect 147474 436814 148094 436898
rect 147474 436578 147506 436814
rect 147742 436578 147826 436814
rect 148062 436578 148094 436814
rect 147474 401134 148094 436578
rect 147474 400898 147506 401134
rect 147742 400898 147826 401134
rect 148062 400898 148094 401134
rect 147474 400814 148094 400898
rect 147474 400578 147506 400814
rect 147742 400578 147826 400814
rect 148062 400578 148094 400814
rect 147474 365134 148094 400578
rect 147474 364898 147506 365134
rect 147742 364898 147826 365134
rect 148062 364898 148094 365134
rect 147474 364814 148094 364898
rect 147474 364578 147506 364814
rect 147742 364578 147826 364814
rect 148062 364578 148094 364814
rect 147474 329134 148094 364578
rect 147474 328898 147506 329134
rect 147742 328898 147826 329134
rect 148062 328898 148094 329134
rect 147474 328814 148094 328898
rect 147474 328578 147506 328814
rect 147742 328578 147826 328814
rect 148062 328578 148094 328814
rect 147474 293134 148094 328578
rect 147474 292898 147506 293134
rect 147742 292898 147826 293134
rect 148062 292898 148094 293134
rect 147474 292814 148094 292898
rect 147474 292578 147506 292814
rect 147742 292578 147826 292814
rect 148062 292578 148094 292814
rect 147474 257134 148094 292578
rect 147474 256898 147506 257134
rect 147742 256898 147826 257134
rect 148062 256898 148094 257134
rect 147474 256814 148094 256898
rect 147474 256578 147506 256814
rect 147742 256578 147826 256814
rect 148062 256578 148094 256814
rect 147474 221134 148094 256578
rect 147474 220898 147506 221134
rect 147742 220898 147826 221134
rect 148062 220898 148094 221134
rect 147474 220814 148094 220898
rect 147474 220578 147506 220814
rect 147742 220578 147826 220814
rect 148062 220578 148094 220814
rect 147474 185134 148094 220578
rect 147474 184898 147506 185134
rect 147742 184898 147826 185134
rect 148062 184898 148094 185134
rect 147474 184814 148094 184898
rect 147474 184578 147506 184814
rect 147742 184578 147826 184814
rect 148062 184578 148094 184814
rect 147474 149134 148094 184578
rect 147474 148898 147506 149134
rect 147742 148898 147826 149134
rect 148062 148898 148094 149134
rect 147474 148814 148094 148898
rect 147474 148578 147506 148814
rect 147742 148578 147826 148814
rect 148062 148578 148094 148814
rect 147474 113134 148094 148578
rect 147474 112898 147506 113134
rect 147742 112898 147826 113134
rect 148062 112898 148094 113134
rect 147474 112814 148094 112898
rect 147474 112578 147506 112814
rect 147742 112578 147826 112814
rect 148062 112578 148094 112814
rect 147474 77134 148094 112578
rect 147474 76898 147506 77134
rect 147742 76898 147826 77134
rect 148062 76898 148094 77134
rect 147474 76814 148094 76898
rect 147474 76578 147506 76814
rect 147742 76578 147826 76814
rect 148062 76578 148094 76814
rect 147474 41134 148094 76578
rect 147474 40898 147506 41134
rect 147742 40898 147826 41134
rect 148062 40898 148094 41134
rect 147474 40814 148094 40898
rect 147474 40578 147506 40814
rect 147742 40578 147826 40814
rect 148062 40578 148094 40814
rect 147474 5134 148094 40578
rect 147474 4898 147506 5134
rect 147742 4898 147826 5134
rect 148062 4898 148094 5134
rect 147474 4814 148094 4898
rect 147474 4578 147506 4814
rect 147742 4578 147826 4814
rect 148062 4578 148094 4814
rect 147474 -2266 148094 4578
rect 147474 -2502 147506 -2266
rect 147742 -2502 147826 -2266
rect 148062 -2502 148094 -2266
rect 147474 -2586 148094 -2502
rect 147474 -2822 147506 -2586
rect 147742 -2822 147826 -2586
rect 148062 -2822 148094 -2586
rect 147474 -7654 148094 -2822
rect 148714 707718 149334 711590
rect 148714 707482 148746 707718
rect 148982 707482 149066 707718
rect 149302 707482 149334 707718
rect 148714 707398 149334 707482
rect 148714 707162 148746 707398
rect 148982 707162 149066 707398
rect 149302 707162 149334 707398
rect 148714 690374 149334 707162
rect 148714 690138 148746 690374
rect 148982 690138 149066 690374
rect 149302 690138 149334 690374
rect 148714 690054 149334 690138
rect 148714 689818 148746 690054
rect 148982 689818 149066 690054
rect 149302 689818 149334 690054
rect 148714 654374 149334 689818
rect 148714 654138 148746 654374
rect 148982 654138 149066 654374
rect 149302 654138 149334 654374
rect 148714 654054 149334 654138
rect 148714 653818 148746 654054
rect 148982 653818 149066 654054
rect 149302 653818 149334 654054
rect 148714 618374 149334 653818
rect 148714 618138 148746 618374
rect 148982 618138 149066 618374
rect 149302 618138 149334 618374
rect 148714 618054 149334 618138
rect 148714 617818 148746 618054
rect 148982 617818 149066 618054
rect 149302 617818 149334 618054
rect 148714 582374 149334 617818
rect 148714 582138 148746 582374
rect 148982 582138 149066 582374
rect 149302 582138 149334 582374
rect 148714 582054 149334 582138
rect 148714 581818 148746 582054
rect 148982 581818 149066 582054
rect 149302 581818 149334 582054
rect 148714 546374 149334 581818
rect 148714 546138 148746 546374
rect 148982 546138 149066 546374
rect 149302 546138 149334 546374
rect 148714 546054 149334 546138
rect 148714 545818 148746 546054
rect 148982 545818 149066 546054
rect 149302 545818 149334 546054
rect 148714 510374 149334 545818
rect 148714 510138 148746 510374
rect 148982 510138 149066 510374
rect 149302 510138 149334 510374
rect 148714 510054 149334 510138
rect 148714 509818 148746 510054
rect 148982 509818 149066 510054
rect 149302 509818 149334 510054
rect 148714 474374 149334 509818
rect 148714 474138 148746 474374
rect 148982 474138 149066 474374
rect 149302 474138 149334 474374
rect 148714 474054 149334 474138
rect 148714 473818 148746 474054
rect 148982 473818 149066 474054
rect 149302 473818 149334 474054
rect 148714 438374 149334 473818
rect 148714 438138 148746 438374
rect 148982 438138 149066 438374
rect 149302 438138 149334 438374
rect 148714 438054 149334 438138
rect 148714 437818 148746 438054
rect 148982 437818 149066 438054
rect 149302 437818 149334 438054
rect 148714 402374 149334 437818
rect 148714 402138 148746 402374
rect 148982 402138 149066 402374
rect 149302 402138 149334 402374
rect 148714 402054 149334 402138
rect 148714 401818 148746 402054
rect 148982 401818 149066 402054
rect 149302 401818 149334 402054
rect 148714 366374 149334 401818
rect 148714 366138 148746 366374
rect 148982 366138 149066 366374
rect 149302 366138 149334 366374
rect 148714 366054 149334 366138
rect 148714 365818 148746 366054
rect 148982 365818 149066 366054
rect 149302 365818 149334 366054
rect 148714 330374 149334 365818
rect 148714 330138 148746 330374
rect 148982 330138 149066 330374
rect 149302 330138 149334 330374
rect 148714 330054 149334 330138
rect 148714 329818 148746 330054
rect 148982 329818 149066 330054
rect 149302 329818 149334 330054
rect 148714 294374 149334 329818
rect 148714 294138 148746 294374
rect 148982 294138 149066 294374
rect 149302 294138 149334 294374
rect 148714 294054 149334 294138
rect 148714 293818 148746 294054
rect 148982 293818 149066 294054
rect 149302 293818 149334 294054
rect 148714 258374 149334 293818
rect 148714 258138 148746 258374
rect 148982 258138 149066 258374
rect 149302 258138 149334 258374
rect 148714 258054 149334 258138
rect 148714 257818 148746 258054
rect 148982 257818 149066 258054
rect 149302 257818 149334 258054
rect 148714 222374 149334 257818
rect 148714 222138 148746 222374
rect 148982 222138 149066 222374
rect 149302 222138 149334 222374
rect 148714 222054 149334 222138
rect 148714 221818 148746 222054
rect 148982 221818 149066 222054
rect 149302 221818 149334 222054
rect 148714 186374 149334 221818
rect 148714 186138 148746 186374
rect 148982 186138 149066 186374
rect 149302 186138 149334 186374
rect 148714 186054 149334 186138
rect 148714 185818 148746 186054
rect 148982 185818 149066 186054
rect 149302 185818 149334 186054
rect 148714 150374 149334 185818
rect 148714 150138 148746 150374
rect 148982 150138 149066 150374
rect 149302 150138 149334 150374
rect 148714 150054 149334 150138
rect 148714 149818 148746 150054
rect 148982 149818 149066 150054
rect 149302 149818 149334 150054
rect 148714 114374 149334 149818
rect 148714 114138 148746 114374
rect 148982 114138 149066 114374
rect 149302 114138 149334 114374
rect 148714 114054 149334 114138
rect 148714 113818 148746 114054
rect 148982 113818 149066 114054
rect 149302 113818 149334 114054
rect 148714 78374 149334 113818
rect 148714 78138 148746 78374
rect 148982 78138 149066 78374
rect 149302 78138 149334 78374
rect 148714 78054 149334 78138
rect 148714 77818 148746 78054
rect 148982 77818 149066 78054
rect 149302 77818 149334 78054
rect 148714 42374 149334 77818
rect 148714 42138 148746 42374
rect 148982 42138 149066 42374
rect 149302 42138 149334 42374
rect 148714 42054 149334 42138
rect 148714 41818 148746 42054
rect 148982 41818 149066 42054
rect 149302 41818 149334 42054
rect 148714 6374 149334 41818
rect 148714 6138 148746 6374
rect 148982 6138 149066 6374
rect 149302 6138 149334 6374
rect 148714 6054 149334 6138
rect 148714 5818 148746 6054
rect 148982 5818 149066 6054
rect 149302 5818 149334 6054
rect 148714 -3226 149334 5818
rect 148714 -3462 148746 -3226
rect 148982 -3462 149066 -3226
rect 149302 -3462 149334 -3226
rect 148714 -3546 149334 -3462
rect 148714 -3782 148746 -3546
rect 148982 -3782 149066 -3546
rect 149302 -3782 149334 -3546
rect 148714 -7654 149334 -3782
rect 149954 708678 150574 711590
rect 149954 708442 149986 708678
rect 150222 708442 150306 708678
rect 150542 708442 150574 708678
rect 149954 708358 150574 708442
rect 149954 708122 149986 708358
rect 150222 708122 150306 708358
rect 150542 708122 150574 708358
rect 149954 691614 150574 708122
rect 149954 691378 149986 691614
rect 150222 691378 150306 691614
rect 150542 691378 150574 691614
rect 149954 691294 150574 691378
rect 149954 691058 149986 691294
rect 150222 691058 150306 691294
rect 150542 691058 150574 691294
rect 149954 655614 150574 691058
rect 149954 655378 149986 655614
rect 150222 655378 150306 655614
rect 150542 655378 150574 655614
rect 149954 655294 150574 655378
rect 149954 655058 149986 655294
rect 150222 655058 150306 655294
rect 150542 655058 150574 655294
rect 149954 619614 150574 655058
rect 149954 619378 149986 619614
rect 150222 619378 150306 619614
rect 150542 619378 150574 619614
rect 149954 619294 150574 619378
rect 149954 619058 149986 619294
rect 150222 619058 150306 619294
rect 150542 619058 150574 619294
rect 149954 583614 150574 619058
rect 149954 583378 149986 583614
rect 150222 583378 150306 583614
rect 150542 583378 150574 583614
rect 149954 583294 150574 583378
rect 149954 583058 149986 583294
rect 150222 583058 150306 583294
rect 150542 583058 150574 583294
rect 149954 547614 150574 583058
rect 149954 547378 149986 547614
rect 150222 547378 150306 547614
rect 150542 547378 150574 547614
rect 149954 547294 150574 547378
rect 149954 547058 149986 547294
rect 150222 547058 150306 547294
rect 150542 547058 150574 547294
rect 149954 511614 150574 547058
rect 149954 511378 149986 511614
rect 150222 511378 150306 511614
rect 150542 511378 150574 511614
rect 149954 511294 150574 511378
rect 149954 511058 149986 511294
rect 150222 511058 150306 511294
rect 150542 511058 150574 511294
rect 149954 475614 150574 511058
rect 149954 475378 149986 475614
rect 150222 475378 150306 475614
rect 150542 475378 150574 475614
rect 149954 475294 150574 475378
rect 149954 475058 149986 475294
rect 150222 475058 150306 475294
rect 150542 475058 150574 475294
rect 149954 439614 150574 475058
rect 149954 439378 149986 439614
rect 150222 439378 150306 439614
rect 150542 439378 150574 439614
rect 149954 439294 150574 439378
rect 149954 439058 149986 439294
rect 150222 439058 150306 439294
rect 150542 439058 150574 439294
rect 149954 403614 150574 439058
rect 149954 403378 149986 403614
rect 150222 403378 150306 403614
rect 150542 403378 150574 403614
rect 149954 403294 150574 403378
rect 149954 403058 149986 403294
rect 150222 403058 150306 403294
rect 150542 403058 150574 403294
rect 149954 367614 150574 403058
rect 149954 367378 149986 367614
rect 150222 367378 150306 367614
rect 150542 367378 150574 367614
rect 149954 367294 150574 367378
rect 149954 367058 149986 367294
rect 150222 367058 150306 367294
rect 150542 367058 150574 367294
rect 149954 331614 150574 367058
rect 149954 331378 149986 331614
rect 150222 331378 150306 331614
rect 150542 331378 150574 331614
rect 149954 331294 150574 331378
rect 149954 331058 149986 331294
rect 150222 331058 150306 331294
rect 150542 331058 150574 331294
rect 149954 295614 150574 331058
rect 149954 295378 149986 295614
rect 150222 295378 150306 295614
rect 150542 295378 150574 295614
rect 149954 295294 150574 295378
rect 149954 295058 149986 295294
rect 150222 295058 150306 295294
rect 150542 295058 150574 295294
rect 149954 259614 150574 295058
rect 149954 259378 149986 259614
rect 150222 259378 150306 259614
rect 150542 259378 150574 259614
rect 149954 259294 150574 259378
rect 149954 259058 149986 259294
rect 150222 259058 150306 259294
rect 150542 259058 150574 259294
rect 149954 223614 150574 259058
rect 149954 223378 149986 223614
rect 150222 223378 150306 223614
rect 150542 223378 150574 223614
rect 149954 223294 150574 223378
rect 149954 223058 149986 223294
rect 150222 223058 150306 223294
rect 150542 223058 150574 223294
rect 149954 187614 150574 223058
rect 149954 187378 149986 187614
rect 150222 187378 150306 187614
rect 150542 187378 150574 187614
rect 149954 187294 150574 187378
rect 149954 187058 149986 187294
rect 150222 187058 150306 187294
rect 150542 187058 150574 187294
rect 149954 151614 150574 187058
rect 149954 151378 149986 151614
rect 150222 151378 150306 151614
rect 150542 151378 150574 151614
rect 149954 151294 150574 151378
rect 149954 151058 149986 151294
rect 150222 151058 150306 151294
rect 150542 151058 150574 151294
rect 149954 115614 150574 151058
rect 149954 115378 149986 115614
rect 150222 115378 150306 115614
rect 150542 115378 150574 115614
rect 149954 115294 150574 115378
rect 149954 115058 149986 115294
rect 150222 115058 150306 115294
rect 150542 115058 150574 115294
rect 149954 79614 150574 115058
rect 149954 79378 149986 79614
rect 150222 79378 150306 79614
rect 150542 79378 150574 79614
rect 149954 79294 150574 79378
rect 149954 79058 149986 79294
rect 150222 79058 150306 79294
rect 150542 79058 150574 79294
rect 149954 43614 150574 79058
rect 149954 43378 149986 43614
rect 150222 43378 150306 43614
rect 150542 43378 150574 43614
rect 149954 43294 150574 43378
rect 149954 43058 149986 43294
rect 150222 43058 150306 43294
rect 150542 43058 150574 43294
rect 149954 7614 150574 43058
rect 149954 7378 149986 7614
rect 150222 7378 150306 7614
rect 150542 7378 150574 7614
rect 149954 7294 150574 7378
rect 149954 7058 149986 7294
rect 150222 7058 150306 7294
rect 150542 7058 150574 7294
rect 149954 -4186 150574 7058
rect 149954 -4422 149986 -4186
rect 150222 -4422 150306 -4186
rect 150542 -4422 150574 -4186
rect 149954 -4506 150574 -4422
rect 149954 -4742 149986 -4506
rect 150222 -4742 150306 -4506
rect 150542 -4742 150574 -4506
rect 149954 -7654 150574 -4742
rect 151194 709638 151814 711590
rect 151194 709402 151226 709638
rect 151462 709402 151546 709638
rect 151782 709402 151814 709638
rect 151194 709318 151814 709402
rect 151194 709082 151226 709318
rect 151462 709082 151546 709318
rect 151782 709082 151814 709318
rect 151194 692854 151814 709082
rect 151194 692618 151226 692854
rect 151462 692618 151546 692854
rect 151782 692618 151814 692854
rect 151194 692534 151814 692618
rect 151194 692298 151226 692534
rect 151462 692298 151546 692534
rect 151782 692298 151814 692534
rect 151194 656854 151814 692298
rect 151194 656618 151226 656854
rect 151462 656618 151546 656854
rect 151782 656618 151814 656854
rect 151194 656534 151814 656618
rect 151194 656298 151226 656534
rect 151462 656298 151546 656534
rect 151782 656298 151814 656534
rect 151194 620854 151814 656298
rect 151194 620618 151226 620854
rect 151462 620618 151546 620854
rect 151782 620618 151814 620854
rect 151194 620534 151814 620618
rect 151194 620298 151226 620534
rect 151462 620298 151546 620534
rect 151782 620298 151814 620534
rect 151194 584854 151814 620298
rect 151194 584618 151226 584854
rect 151462 584618 151546 584854
rect 151782 584618 151814 584854
rect 151194 584534 151814 584618
rect 151194 584298 151226 584534
rect 151462 584298 151546 584534
rect 151782 584298 151814 584534
rect 151194 548854 151814 584298
rect 151194 548618 151226 548854
rect 151462 548618 151546 548854
rect 151782 548618 151814 548854
rect 151194 548534 151814 548618
rect 151194 548298 151226 548534
rect 151462 548298 151546 548534
rect 151782 548298 151814 548534
rect 151194 512854 151814 548298
rect 151194 512618 151226 512854
rect 151462 512618 151546 512854
rect 151782 512618 151814 512854
rect 151194 512534 151814 512618
rect 151194 512298 151226 512534
rect 151462 512298 151546 512534
rect 151782 512298 151814 512534
rect 151194 476854 151814 512298
rect 151194 476618 151226 476854
rect 151462 476618 151546 476854
rect 151782 476618 151814 476854
rect 151194 476534 151814 476618
rect 151194 476298 151226 476534
rect 151462 476298 151546 476534
rect 151782 476298 151814 476534
rect 151194 440854 151814 476298
rect 151194 440618 151226 440854
rect 151462 440618 151546 440854
rect 151782 440618 151814 440854
rect 151194 440534 151814 440618
rect 151194 440298 151226 440534
rect 151462 440298 151546 440534
rect 151782 440298 151814 440534
rect 151194 404854 151814 440298
rect 151194 404618 151226 404854
rect 151462 404618 151546 404854
rect 151782 404618 151814 404854
rect 151194 404534 151814 404618
rect 151194 404298 151226 404534
rect 151462 404298 151546 404534
rect 151782 404298 151814 404534
rect 151194 368854 151814 404298
rect 151194 368618 151226 368854
rect 151462 368618 151546 368854
rect 151782 368618 151814 368854
rect 151194 368534 151814 368618
rect 151194 368298 151226 368534
rect 151462 368298 151546 368534
rect 151782 368298 151814 368534
rect 151194 332854 151814 368298
rect 151194 332618 151226 332854
rect 151462 332618 151546 332854
rect 151782 332618 151814 332854
rect 151194 332534 151814 332618
rect 151194 332298 151226 332534
rect 151462 332298 151546 332534
rect 151782 332298 151814 332534
rect 151194 296854 151814 332298
rect 151194 296618 151226 296854
rect 151462 296618 151546 296854
rect 151782 296618 151814 296854
rect 151194 296534 151814 296618
rect 151194 296298 151226 296534
rect 151462 296298 151546 296534
rect 151782 296298 151814 296534
rect 151194 260854 151814 296298
rect 151194 260618 151226 260854
rect 151462 260618 151546 260854
rect 151782 260618 151814 260854
rect 151194 260534 151814 260618
rect 151194 260298 151226 260534
rect 151462 260298 151546 260534
rect 151782 260298 151814 260534
rect 151194 224854 151814 260298
rect 151194 224618 151226 224854
rect 151462 224618 151546 224854
rect 151782 224618 151814 224854
rect 151194 224534 151814 224618
rect 151194 224298 151226 224534
rect 151462 224298 151546 224534
rect 151782 224298 151814 224534
rect 151194 188854 151814 224298
rect 151194 188618 151226 188854
rect 151462 188618 151546 188854
rect 151782 188618 151814 188854
rect 151194 188534 151814 188618
rect 151194 188298 151226 188534
rect 151462 188298 151546 188534
rect 151782 188298 151814 188534
rect 151194 152854 151814 188298
rect 151194 152618 151226 152854
rect 151462 152618 151546 152854
rect 151782 152618 151814 152854
rect 151194 152534 151814 152618
rect 151194 152298 151226 152534
rect 151462 152298 151546 152534
rect 151782 152298 151814 152534
rect 151194 116854 151814 152298
rect 151194 116618 151226 116854
rect 151462 116618 151546 116854
rect 151782 116618 151814 116854
rect 151194 116534 151814 116618
rect 151194 116298 151226 116534
rect 151462 116298 151546 116534
rect 151782 116298 151814 116534
rect 151194 80854 151814 116298
rect 151194 80618 151226 80854
rect 151462 80618 151546 80854
rect 151782 80618 151814 80854
rect 151194 80534 151814 80618
rect 151194 80298 151226 80534
rect 151462 80298 151546 80534
rect 151782 80298 151814 80534
rect 151194 44854 151814 80298
rect 151194 44618 151226 44854
rect 151462 44618 151546 44854
rect 151782 44618 151814 44854
rect 151194 44534 151814 44618
rect 151194 44298 151226 44534
rect 151462 44298 151546 44534
rect 151782 44298 151814 44534
rect 151194 8854 151814 44298
rect 151194 8618 151226 8854
rect 151462 8618 151546 8854
rect 151782 8618 151814 8854
rect 151194 8534 151814 8618
rect 151194 8298 151226 8534
rect 151462 8298 151546 8534
rect 151782 8298 151814 8534
rect 151194 -5146 151814 8298
rect 151194 -5382 151226 -5146
rect 151462 -5382 151546 -5146
rect 151782 -5382 151814 -5146
rect 151194 -5466 151814 -5382
rect 151194 -5702 151226 -5466
rect 151462 -5702 151546 -5466
rect 151782 -5702 151814 -5466
rect 151194 -7654 151814 -5702
rect 152434 710598 153054 711590
rect 152434 710362 152466 710598
rect 152702 710362 152786 710598
rect 153022 710362 153054 710598
rect 152434 710278 153054 710362
rect 152434 710042 152466 710278
rect 152702 710042 152786 710278
rect 153022 710042 153054 710278
rect 152434 694094 153054 710042
rect 152434 693858 152466 694094
rect 152702 693858 152786 694094
rect 153022 693858 153054 694094
rect 152434 693774 153054 693858
rect 152434 693538 152466 693774
rect 152702 693538 152786 693774
rect 153022 693538 153054 693774
rect 152434 658094 153054 693538
rect 152434 657858 152466 658094
rect 152702 657858 152786 658094
rect 153022 657858 153054 658094
rect 152434 657774 153054 657858
rect 152434 657538 152466 657774
rect 152702 657538 152786 657774
rect 153022 657538 153054 657774
rect 152434 622094 153054 657538
rect 152434 621858 152466 622094
rect 152702 621858 152786 622094
rect 153022 621858 153054 622094
rect 152434 621774 153054 621858
rect 152434 621538 152466 621774
rect 152702 621538 152786 621774
rect 153022 621538 153054 621774
rect 152434 586094 153054 621538
rect 152434 585858 152466 586094
rect 152702 585858 152786 586094
rect 153022 585858 153054 586094
rect 152434 585774 153054 585858
rect 152434 585538 152466 585774
rect 152702 585538 152786 585774
rect 153022 585538 153054 585774
rect 152434 550094 153054 585538
rect 152434 549858 152466 550094
rect 152702 549858 152786 550094
rect 153022 549858 153054 550094
rect 152434 549774 153054 549858
rect 152434 549538 152466 549774
rect 152702 549538 152786 549774
rect 153022 549538 153054 549774
rect 152434 514094 153054 549538
rect 152434 513858 152466 514094
rect 152702 513858 152786 514094
rect 153022 513858 153054 514094
rect 152434 513774 153054 513858
rect 152434 513538 152466 513774
rect 152702 513538 152786 513774
rect 153022 513538 153054 513774
rect 152434 478094 153054 513538
rect 152434 477858 152466 478094
rect 152702 477858 152786 478094
rect 153022 477858 153054 478094
rect 152434 477774 153054 477858
rect 152434 477538 152466 477774
rect 152702 477538 152786 477774
rect 153022 477538 153054 477774
rect 152434 442094 153054 477538
rect 152434 441858 152466 442094
rect 152702 441858 152786 442094
rect 153022 441858 153054 442094
rect 152434 441774 153054 441858
rect 152434 441538 152466 441774
rect 152702 441538 152786 441774
rect 153022 441538 153054 441774
rect 152434 406094 153054 441538
rect 152434 405858 152466 406094
rect 152702 405858 152786 406094
rect 153022 405858 153054 406094
rect 152434 405774 153054 405858
rect 152434 405538 152466 405774
rect 152702 405538 152786 405774
rect 153022 405538 153054 405774
rect 152434 370094 153054 405538
rect 152434 369858 152466 370094
rect 152702 369858 152786 370094
rect 153022 369858 153054 370094
rect 152434 369774 153054 369858
rect 152434 369538 152466 369774
rect 152702 369538 152786 369774
rect 153022 369538 153054 369774
rect 152434 334094 153054 369538
rect 152434 333858 152466 334094
rect 152702 333858 152786 334094
rect 153022 333858 153054 334094
rect 152434 333774 153054 333858
rect 152434 333538 152466 333774
rect 152702 333538 152786 333774
rect 153022 333538 153054 333774
rect 152434 298094 153054 333538
rect 152434 297858 152466 298094
rect 152702 297858 152786 298094
rect 153022 297858 153054 298094
rect 152434 297774 153054 297858
rect 152434 297538 152466 297774
rect 152702 297538 152786 297774
rect 153022 297538 153054 297774
rect 152434 262094 153054 297538
rect 152434 261858 152466 262094
rect 152702 261858 152786 262094
rect 153022 261858 153054 262094
rect 152434 261774 153054 261858
rect 152434 261538 152466 261774
rect 152702 261538 152786 261774
rect 153022 261538 153054 261774
rect 152434 226094 153054 261538
rect 152434 225858 152466 226094
rect 152702 225858 152786 226094
rect 153022 225858 153054 226094
rect 152434 225774 153054 225858
rect 152434 225538 152466 225774
rect 152702 225538 152786 225774
rect 153022 225538 153054 225774
rect 152434 190094 153054 225538
rect 152434 189858 152466 190094
rect 152702 189858 152786 190094
rect 153022 189858 153054 190094
rect 152434 189774 153054 189858
rect 152434 189538 152466 189774
rect 152702 189538 152786 189774
rect 153022 189538 153054 189774
rect 152434 154094 153054 189538
rect 152434 153858 152466 154094
rect 152702 153858 152786 154094
rect 153022 153858 153054 154094
rect 152434 153774 153054 153858
rect 152434 153538 152466 153774
rect 152702 153538 152786 153774
rect 153022 153538 153054 153774
rect 152434 118094 153054 153538
rect 152434 117858 152466 118094
rect 152702 117858 152786 118094
rect 153022 117858 153054 118094
rect 152434 117774 153054 117858
rect 152434 117538 152466 117774
rect 152702 117538 152786 117774
rect 153022 117538 153054 117774
rect 152434 82094 153054 117538
rect 152434 81858 152466 82094
rect 152702 81858 152786 82094
rect 153022 81858 153054 82094
rect 152434 81774 153054 81858
rect 152434 81538 152466 81774
rect 152702 81538 152786 81774
rect 153022 81538 153054 81774
rect 152434 46094 153054 81538
rect 152434 45858 152466 46094
rect 152702 45858 152786 46094
rect 153022 45858 153054 46094
rect 152434 45774 153054 45858
rect 152434 45538 152466 45774
rect 152702 45538 152786 45774
rect 153022 45538 153054 45774
rect 152434 10094 153054 45538
rect 152434 9858 152466 10094
rect 152702 9858 152786 10094
rect 153022 9858 153054 10094
rect 152434 9774 153054 9858
rect 152434 9538 152466 9774
rect 152702 9538 152786 9774
rect 153022 9538 153054 9774
rect 152434 -6106 153054 9538
rect 152434 -6342 152466 -6106
rect 152702 -6342 152786 -6106
rect 153022 -6342 153054 -6106
rect 152434 -6426 153054 -6342
rect 152434 -6662 152466 -6426
rect 152702 -6662 152786 -6426
rect 153022 -6662 153054 -6426
rect 152434 -7654 153054 -6662
rect 153674 711558 154294 711590
rect 153674 711322 153706 711558
rect 153942 711322 154026 711558
rect 154262 711322 154294 711558
rect 153674 711238 154294 711322
rect 153674 711002 153706 711238
rect 153942 711002 154026 711238
rect 154262 711002 154294 711238
rect 153674 695334 154294 711002
rect 153674 695098 153706 695334
rect 153942 695098 154026 695334
rect 154262 695098 154294 695334
rect 153674 695014 154294 695098
rect 153674 694778 153706 695014
rect 153942 694778 154026 695014
rect 154262 694778 154294 695014
rect 153674 659334 154294 694778
rect 153674 659098 153706 659334
rect 153942 659098 154026 659334
rect 154262 659098 154294 659334
rect 153674 659014 154294 659098
rect 153674 658778 153706 659014
rect 153942 658778 154026 659014
rect 154262 658778 154294 659014
rect 153674 623334 154294 658778
rect 153674 623098 153706 623334
rect 153942 623098 154026 623334
rect 154262 623098 154294 623334
rect 153674 623014 154294 623098
rect 153674 622778 153706 623014
rect 153942 622778 154026 623014
rect 154262 622778 154294 623014
rect 153674 587334 154294 622778
rect 153674 587098 153706 587334
rect 153942 587098 154026 587334
rect 154262 587098 154294 587334
rect 153674 587014 154294 587098
rect 153674 586778 153706 587014
rect 153942 586778 154026 587014
rect 154262 586778 154294 587014
rect 153674 551334 154294 586778
rect 153674 551098 153706 551334
rect 153942 551098 154026 551334
rect 154262 551098 154294 551334
rect 153674 551014 154294 551098
rect 153674 550778 153706 551014
rect 153942 550778 154026 551014
rect 154262 550778 154294 551014
rect 153674 515334 154294 550778
rect 153674 515098 153706 515334
rect 153942 515098 154026 515334
rect 154262 515098 154294 515334
rect 153674 515014 154294 515098
rect 153674 514778 153706 515014
rect 153942 514778 154026 515014
rect 154262 514778 154294 515014
rect 153674 479334 154294 514778
rect 153674 479098 153706 479334
rect 153942 479098 154026 479334
rect 154262 479098 154294 479334
rect 153674 479014 154294 479098
rect 153674 478778 153706 479014
rect 153942 478778 154026 479014
rect 154262 478778 154294 479014
rect 153674 443334 154294 478778
rect 153674 443098 153706 443334
rect 153942 443098 154026 443334
rect 154262 443098 154294 443334
rect 153674 443014 154294 443098
rect 153674 442778 153706 443014
rect 153942 442778 154026 443014
rect 154262 442778 154294 443014
rect 153674 407334 154294 442778
rect 153674 407098 153706 407334
rect 153942 407098 154026 407334
rect 154262 407098 154294 407334
rect 153674 407014 154294 407098
rect 153674 406778 153706 407014
rect 153942 406778 154026 407014
rect 154262 406778 154294 407014
rect 153674 371334 154294 406778
rect 153674 371098 153706 371334
rect 153942 371098 154026 371334
rect 154262 371098 154294 371334
rect 153674 371014 154294 371098
rect 153674 370778 153706 371014
rect 153942 370778 154026 371014
rect 154262 370778 154294 371014
rect 153674 335334 154294 370778
rect 153674 335098 153706 335334
rect 153942 335098 154026 335334
rect 154262 335098 154294 335334
rect 153674 335014 154294 335098
rect 153674 334778 153706 335014
rect 153942 334778 154026 335014
rect 154262 334778 154294 335014
rect 153674 299334 154294 334778
rect 153674 299098 153706 299334
rect 153942 299098 154026 299334
rect 154262 299098 154294 299334
rect 153674 299014 154294 299098
rect 153674 298778 153706 299014
rect 153942 298778 154026 299014
rect 154262 298778 154294 299014
rect 153674 263334 154294 298778
rect 153674 263098 153706 263334
rect 153942 263098 154026 263334
rect 154262 263098 154294 263334
rect 153674 263014 154294 263098
rect 153674 262778 153706 263014
rect 153942 262778 154026 263014
rect 154262 262778 154294 263014
rect 153674 227334 154294 262778
rect 153674 227098 153706 227334
rect 153942 227098 154026 227334
rect 154262 227098 154294 227334
rect 153674 227014 154294 227098
rect 153674 226778 153706 227014
rect 153942 226778 154026 227014
rect 154262 226778 154294 227014
rect 153674 191334 154294 226778
rect 153674 191098 153706 191334
rect 153942 191098 154026 191334
rect 154262 191098 154294 191334
rect 153674 191014 154294 191098
rect 153674 190778 153706 191014
rect 153942 190778 154026 191014
rect 154262 190778 154294 191014
rect 153674 155334 154294 190778
rect 153674 155098 153706 155334
rect 153942 155098 154026 155334
rect 154262 155098 154294 155334
rect 153674 155014 154294 155098
rect 153674 154778 153706 155014
rect 153942 154778 154026 155014
rect 154262 154778 154294 155014
rect 153674 119334 154294 154778
rect 153674 119098 153706 119334
rect 153942 119098 154026 119334
rect 154262 119098 154294 119334
rect 153674 119014 154294 119098
rect 153674 118778 153706 119014
rect 153942 118778 154026 119014
rect 154262 118778 154294 119014
rect 153674 83334 154294 118778
rect 153674 83098 153706 83334
rect 153942 83098 154026 83334
rect 154262 83098 154294 83334
rect 153674 83014 154294 83098
rect 153674 82778 153706 83014
rect 153942 82778 154026 83014
rect 154262 82778 154294 83014
rect 153674 47334 154294 82778
rect 153674 47098 153706 47334
rect 153942 47098 154026 47334
rect 154262 47098 154294 47334
rect 153674 47014 154294 47098
rect 153674 46778 153706 47014
rect 153942 46778 154026 47014
rect 154262 46778 154294 47014
rect 153674 11334 154294 46778
rect 153674 11098 153706 11334
rect 153942 11098 154026 11334
rect 154262 11098 154294 11334
rect 153674 11014 154294 11098
rect 153674 10778 153706 11014
rect 153942 10778 154026 11014
rect 154262 10778 154294 11014
rect 153674 -7066 154294 10778
rect 153674 -7302 153706 -7066
rect 153942 -7302 154026 -7066
rect 154262 -7302 154294 -7066
rect 153674 -7386 154294 -7302
rect 153674 -7622 153706 -7386
rect 153942 -7622 154026 -7386
rect 154262 -7622 154294 -7386
rect 153674 -7654 154294 -7622
rect 180994 704838 181614 711590
rect 180994 704602 181026 704838
rect 181262 704602 181346 704838
rect 181582 704602 181614 704838
rect 180994 704518 181614 704602
rect 180994 704282 181026 704518
rect 181262 704282 181346 704518
rect 181582 704282 181614 704518
rect 180994 686654 181614 704282
rect 180994 686418 181026 686654
rect 181262 686418 181346 686654
rect 181582 686418 181614 686654
rect 180994 686334 181614 686418
rect 180994 686098 181026 686334
rect 181262 686098 181346 686334
rect 181582 686098 181614 686334
rect 180994 650654 181614 686098
rect 180994 650418 181026 650654
rect 181262 650418 181346 650654
rect 181582 650418 181614 650654
rect 180994 650334 181614 650418
rect 180994 650098 181026 650334
rect 181262 650098 181346 650334
rect 181582 650098 181614 650334
rect 180994 614654 181614 650098
rect 180994 614418 181026 614654
rect 181262 614418 181346 614654
rect 181582 614418 181614 614654
rect 180994 614334 181614 614418
rect 180994 614098 181026 614334
rect 181262 614098 181346 614334
rect 181582 614098 181614 614334
rect 180994 578654 181614 614098
rect 180994 578418 181026 578654
rect 181262 578418 181346 578654
rect 181582 578418 181614 578654
rect 180994 578334 181614 578418
rect 180994 578098 181026 578334
rect 181262 578098 181346 578334
rect 181582 578098 181614 578334
rect 180994 542654 181614 578098
rect 180994 542418 181026 542654
rect 181262 542418 181346 542654
rect 181582 542418 181614 542654
rect 180994 542334 181614 542418
rect 180994 542098 181026 542334
rect 181262 542098 181346 542334
rect 181582 542098 181614 542334
rect 180994 506654 181614 542098
rect 180994 506418 181026 506654
rect 181262 506418 181346 506654
rect 181582 506418 181614 506654
rect 180994 506334 181614 506418
rect 180994 506098 181026 506334
rect 181262 506098 181346 506334
rect 181582 506098 181614 506334
rect 180994 470654 181614 506098
rect 180994 470418 181026 470654
rect 181262 470418 181346 470654
rect 181582 470418 181614 470654
rect 180994 470334 181614 470418
rect 180994 470098 181026 470334
rect 181262 470098 181346 470334
rect 181582 470098 181614 470334
rect 180994 434654 181614 470098
rect 180994 434418 181026 434654
rect 181262 434418 181346 434654
rect 181582 434418 181614 434654
rect 180994 434334 181614 434418
rect 180994 434098 181026 434334
rect 181262 434098 181346 434334
rect 181582 434098 181614 434334
rect 180994 398654 181614 434098
rect 180994 398418 181026 398654
rect 181262 398418 181346 398654
rect 181582 398418 181614 398654
rect 180994 398334 181614 398418
rect 180994 398098 181026 398334
rect 181262 398098 181346 398334
rect 181582 398098 181614 398334
rect 180994 362654 181614 398098
rect 180994 362418 181026 362654
rect 181262 362418 181346 362654
rect 181582 362418 181614 362654
rect 180994 362334 181614 362418
rect 180994 362098 181026 362334
rect 181262 362098 181346 362334
rect 181582 362098 181614 362334
rect 180994 326654 181614 362098
rect 180994 326418 181026 326654
rect 181262 326418 181346 326654
rect 181582 326418 181614 326654
rect 180994 326334 181614 326418
rect 180994 326098 181026 326334
rect 181262 326098 181346 326334
rect 181582 326098 181614 326334
rect 180994 290654 181614 326098
rect 180994 290418 181026 290654
rect 181262 290418 181346 290654
rect 181582 290418 181614 290654
rect 180994 290334 181614 290418
rect 180994 290098 181026 290334
rect 181262 290098 181346 290334
rect 181582 290098 181614 290334
rect 180994 254654 181614 290098
rect 180994 254418 181026 254654
rect 181262 254418 181346 254654
rect 181582 254418 181614 254654
rect 180994 254334 181614 254418
rect 180994 254098 181026 254334
rect 181262 254098 181346 254334
rect 181582 254098 181614 254334
rect 180994 218654 181614 254098
rect 180994 218418 181026 218654
rect 181262 218418 181346 218654
rect 181582 218418 181614 218654
rect 180994 218334 181614 218418
rect 180994 218098 181026 218334
rect 181262 218098 181346 218334
rect 181582 218098 181614 218334
rect 180994 182654 181614 218098
rect 180994 182418 181026 182654
rect 181262 182418 181346 182654
rect 181582 182418 181614 182654
rect 180994 182334 181614 182418
rect 180994 182098 181026 182334
rect 181262 182098 181346 182334
rect 181582 182098 181614 182334
rect 180994 146654 181614 182098
rect 180994 146418 181026 146654
rect 181262 146418 181346 146654
rect 181582 146418 181614 146654
rect 180994 146334 181614 146418
rect 180994 146098 181026 146334
rect 181262 146098 181346 146334
rect 181582 146098 181614 146334
rect 180994 110654 181614 146098
rect 180994 110418 181026 110654
rect 181262 110418 181346 110654
rect 181582 110418 181614 110654
rect 180994 110334 181614 110418
rect 180994 110098 181026 110334
rect 181262 110098 181346 110334
rect 181582 110098 181614 110334
rect 180994 74654 181614 110098
rect 180994 74418 181026 74654
rect 181262 74418 181346 74654
rect 181582 74418 181614 74654
rect 180994 74334 181614 74418
rect 180994 74098 181026 74334
rect 181262 74098 181346 74334
rect 181582 74098 181614 74334
rect 180994 38654 181614 74098
rect 180994 38418 181026 38654
rect 181262 38418 181346 38654
rect 181582 38418 181614 38654
rect 180994 38334 181614 38418
rect 180994 38098 181026 38334
rect 181262 38098 181346 38334
rect 181582 38098 181614 38334
rect 180994 2654 181614 38098
rect 180994 2418 181026 2654
rect 181262 2418 181346 2654
rect 181582 2418 181614 2654
rect 180994 2334 181614 2418
rect 180994 2098 181026 2334
rect 181262 2098 181346 2334
rect 181582 2098 181614 2334
rect 180994 -346 181614 2098
rect 180994 -582 181026 -346
rect 181262 -582 181346 -346
rect 181582 -582 181614 -346
rect 180994 -666 181614 -582
rect 180994 -902 181026 -666
rect 181262 -902 181346 -666
rect 181582 -902 181614 -666
rect 180994 -7654 181614 -902
rect 182234 705798 182854 711590
rect 182234 705562 182266 705798
rect 182502 705562 182586 705798
rect 182822 705562 182854 705798
rect 182234 705478 182854 705562
rect 182234 705242 182266 705478
rect 182502 705242 182586 705478
rect 182822 705242 182854 705478
rect 182234 687894 182854 705242
rect 182234 687658 182266 687894
rect 182502 687658 182586 687894
rect 182822 687658 182854 687894
rect 182234 687574 182854 687658
rect 182234 687338 182266 687574
rect 182502 687338 182586 687574
rect 182822 687338 182854 687574
rect 182234 651894 182854 687338
rect 182234 651658 182266 651894
rect 182502 651658 182586 651894
rect 182822 651658 182854 651894
rect 182234 651574 182854 651658
rect 182234 651338 182266 651574
rect 182502 651338 182586 651574
rect 182822 651338 182854 651574
rect 182234 615894 182854 651338
rect 182234 615658 182266 615894
rect 182502 615658 182586 615894
rect 182822 615658 182854 615894
rect 182234 615574 182854 615658
rect 182234 615338 182266 615574
rect 182502 615338 182586 615574
rect 182822 615338 182854 615574
rect 182234 579894 182854 615338
rect 182234 579658 182266 579894
rect 182502 579658 182586 579894
rect 182822 579658 182854 579894
rect 182234 579574 182854 579658
rect 182234 579338 182266 579574
rect 182502 579338 182586 579574
rect 182822 579338 182854 579574
rect 182234 543894 182854 579338
rect 182234 543658 182266 543894
rect 182502 543658 182586 543894
rect 182822 543658 182854 543894
rect 182234 543574 182854 543658
rect 182234 543338 182266 543574
rect 182502 543338 182586 543574
rect 182822 543338 182854 543574
rect 182234 507894 182854 543338
rect 182234 507658 182266 507894
rect 182502 507658 182586 507894
rect 182822 507658 182854 507894
rect 182234 507574 182854 507658
rect 182234 507338 182266 507574
rect 182502 507338 182586 507574
rect 182822 507338 182854 507574
rect 182234 471894 182854 507338
rect 182234 471658 182266 471894
rect 182502 471658 182586 471894
rect 182822 471658 182854 471894
rect 182234 471574 182854 471658
rect 182234 471338 182266 471574
rect 182502 471338 182586 471574
rect 182822 471338 182854 471574
rect 182234 435894 182854 471338
rect 182234 435658 182266 435894
rect 182502 435658 182586 435894
rect 182822 435658 182854 435894
rect 182234 435574 182854 435658
rect 182234 435338 182266 435574
rect 182502 435338 182586 435574
rect 182822 435338 182854 435574
rect 182234 399894 182854 435338
rect 182234 399658 182266 399894
rect 182502 399658 182586 399894
rect 182822 399658 182854 399894
rect 182234 399574 182854 399658
rect 182234 399338 182266 399574
rect 182502 399338 182586 399574
rect 182822 399338 182854 399574
rect 182234 363894 182854 399338
rect 182234 363658 182266 363894
rect 182502 363658 182586 363894
rect 182822 363658 182854 363894
rect 182234 363574 182854 363658
rect 182234 363338 182266 363574
rect 182502 363338 182586 363574
rect 182822 363338 182854 363574
rect 182234 327894 182854 363338
rect 182234 327658 182266 327894
rect 182502 327658 182586 327894
rect 182822 327658 182854 327894
rect 182234 327574 182854 327658
rect 182234 327338 182266 327574
rect 182502 327338 182586 327574
rect 182822 327338 182854 327574
rect 182234 291894 182854 327338
rect 182234 291658 182266 291894
rect 182502 291658 182586 291894
rect 182822 291658 182854 291894
rect 182234 291574 182854 291658
rect 182234 291338 182266 291574
rect 182502 291338 182586 291574
rect 182822 291338 182854 291574
rect 182234 255894 182854 291338
rect 182234 255658 182266 255894
rect 182502 255658 182586 255894
rect 182822 255658 182854 255894
rect 182234 255574 182854 255658
rect 182234 255338 182266 255574
rect 182502 255338 182586 255574
rect 182822 255338 182854 255574
rect 182234 219894 182854 255338
rect 182234 219658 182266 219894
rect 182502 219658 182586 219894
rect 182822 219658 182854 219894
rect 182234 219574 182854 219658
rect 182234 219338 182266 219574
rect 182502 219338 182586 219574
rect 182822 219338 182854 219574
rect 182234 183894 182854 219338
rect 182234 183658 182266 183894
rect 182502 183658 182586 183894
rect 182822 183658 182854 183894
rect 182234 183574 182854 183658
rect 182234 183338 182266 183574
rect 182502 183338 182586 183574
rect 182822 183338 182854 183574
rect 182234 147894 182854 183338
rect 182234 147658 182266 147894
rect 182502 147658 182586 147894
rect 182822 147658 182854 147894
rect 182234 147574 182854 147658
rect 182234 147338 182266 147574
rect 182502 147338 182586 147574
rect 182822 147338 182854 147574
rect 182234 111894 182854 147338
rect 182234 111658 182266 111894
rect 182502 111658 182586 111894
rect 182822 111658 182854 111894
rect 182234 111574 182854 111658
rect 182234 111338 182266 111574
rect 182502 111338 182586 111574
rect 182822 111338 182854 111574
rect 182234 75894 182854 111338
rect 182234 75658 182266 75894
rect 182502 75658 182586 75894
rect 182822 75658 182854 75894
rect 182234 75574 182854 75658
rect 182234 75338 182266 75574
rect 182502 75338 182586 75574
rect 182822 75338 182854 75574
rect 182234 39894 182854 75338
rect 182234 39658 182266 39894
rect 182502 39658 182586 39894
rect 182822 39658 182854 39894
rect 182234 39574 182854 39658
rect 182234 39338 182266 39574
rect 182502 39338 182586 39574
rect 182822 39338 182854 39574
rect 182234 3894 182854 39338
rect 182234 3658 182266 3894
rect 182502 3658 182586 3894
rect 182822 3658 182854 3894
rect 182234 3574 182854 3658
rect 182234 3338 182266 3574
rect 182502 3338 182586 3574
rect 182822 3338 182854 3574
rect 182234 -1306 182854 3338
rect 182234 -1542 182266 -1306
rect 182502 -1542 182586 -1306
rect 182822 -1542 182854 -1306
rect 182234 -1626 182854 -1542
rect 182234 -1862 182266 -1626
rect 182502 -1862 182586 -1626
rect 182822 -1862 182854 -1626
rect 182234 -7654 182854 -1862
rect 183474 706758 184094 711590
rect 183474 706522 183506 706758
rect 183742 706522 183826 706758
rect 184062 706522 184094 706758
rect 183474 706438 184094 706522
rect 183474 706202 183506 706438
rect 183742 706202 183826 706438
rect 184062 706202 184094 706438
rect 183474 689134 184094 706202
rect 183474 688898 183506 689134
rect 183742 688898 183826 689134
rect 184062 688898 184094 689134
rect 183474 688814 184094 688898
rect 183474 688578 183506 688814
rect 183742 688578 183826 688814
rect 184062 688578 184094 688814
rect 183474 653134 184094 688578
rect 183474 652898 183506 653134
rect 183742 652898 183826 653134
rect 184062 652898 184094 653134
rect 183474 652814 184094 652898
rect 183474 652578 183506 652814
rect 183742 652578 183826 652814
rect 184062 652578 184094 652814
rect 183474 617134 184094 652578
rect 183474 616898 183506 617134
rect 183742 616898 183826 617134
rect 184062 616898 184094 617134
rect 183474 616814 184094 616898
rect 183474 616578 183506 616814
rect 183742 616578 183826 616814
rect 184062 616578 184094 616814
rect 183474 581134 184094 616578
rect 183474 580898 183506 581134
rect 183742 580898 183826 581134
rect 184062 580898 184094 581134
rect 183474 580814 184094 580898
rect 183474 580578 183506 580814
rect 183742 580578 183826 580814
rect 184062 580578 184094 580814
rect 183474 545134 184094 580578
rect 183474 544898 183506 545134
rect 183742 544898 183826 545134
rect 184062 544898 184094 545134
rect 183474 544814 184094 544898
rect 183474 544578 183506 544814
rect 183742 544578 183826 544814
rect 184062 544578 184094 544814
rect 183474 509134 184094 544578
rect 183474 508898 183506 509134
rect 183742 508898 183826 509134
rect 184062 508898 184094 509134
rect 183474 508814 184094 508898
rect 183474 508578 183506 508814
rect 183742 508578 183826 508814
rect 184062 508578 184094 508814
rect 183474 473134 184094 508578
rect 183474 472898 183506 473134
rect 183742 472898 183826 473134
rect 184062 472898 184094 473134
rect 183474 472814 184094 472898
rect 183474 472578 183506 472814
rect 183742 472578 183826 472814
rect 184062 472578 184094 472814
rect 183474 437134 184094 472578
rect 183474 436898 183506 437134
rect 183742 436898 183826 437134
rect 184062 436898 184094 437134
rect 183474 436814 184094 436898
rect 183474 436578 183506 436814
rect 183742 436578 183826 436814
rect 184062 436578 184094 436814
rect 183474 401134 184094 436578
rect 183474 400898 183506 401134
rect 183742 400898 183826 401134
rect 184062 400898 184094 401134
rect 183474 400814 184094 400898
rect 183474 400578 183506 400814
rect 183742 400578 183826 400814
rect 184062 400578 184094 400814
rect 183474 365134 184094 400578
rect 183474 364898 183506 365134
rect 183742 364898 183826 365134
rect 184062 364898 184094 365134
rect 183474 364814 184094 364898
rect 183474 364578 183506 364814
rect 183742 364578 183826 364814
rect 184062 364578 184094 364814
rect 183474 329134 184094 364578
rect 183474 328898 183506 329134
rect 183742 328898 183826 329134
rect 184062 328898 184094 329134
rect 183474 328814 184094 328898
rect 183474 328578 183506 328814
rect 183742 328578 183826 328814
rect 184062 328578 184094 328814
rect 183474 293134 184094 328578
rect 183474 292898 183506 293134
rect 183742 292898 183826 293134
rect 184062 292898 184094 293134
rect 183474 292814 184094 292898
rect 183474 292578 183506 292814
rect 183742 292578 183826 292814
rect 184062 292578 184094 292814
rect 183474 257134 184094 292578
rect 183474 256898 183506 257134
rect 183742 256898 183826 257134
rect 184062 256898 184094 257134
rect 183474 256814 184094 256898
rect 183474 256578 183506 256814
rect 183742 256578 183826 256814
rect 184062 256578 184094 256814
rect 183474 221134 184094 256578
rect 183474 220898 183506 221134
rect 183742 220898 183826 221134
rect 184062 220898 184094 221134
rect 183474 220814 184094 220898
rect 183474 220578 183506 220814
rect 183742 220578 183826 220814
rect 184062 220578 184094 220814
rect 183474 185134 184094 220578
rect 183474 184898 183506 185134
rect 183742 184898 183826 185134
rect 184062 184898 184094 185134
rect 183474 184814 184094 184898
rect 183474 184578 183506 184814
rect 183742 184578 183826 184814
rect 184062 184578 184094 184814
rect 183474 149134 184094 184578
rect 183474 148898 183506 149134
rect 183742 148898 183826 149134
rect 184062 148898 184094 149134
rect 183474 148814 184094 148898
rect 183474 148578 183506 148814
rect 183742 148578 183826 148814
rect 184062 148578 184094 148814
rect 183474 113134 184094 148578
rect 183474 112898 183506 113134
rect 183742 112898 183826 113134
rect 184062 112898 184094 113134
rect 183474 112814 184094 112898
rect 183474 112578 183506 112814
rect 183742 112578 183826 112814
rect 184062 112578 184094 112814
rect 183474 77134 184094 112578
rect 183474 76898 183506 77134
rect 183742 76898 183826 77134
rect 184062 76898 184094 77134
rect 183474 76814 184094 76898
rect 183474 76578 183506 76814
rect 183742 76578 183826 76814
rect 184062 76578 184094 76814
rect 183474 41134 184094 76578
rect 183474 40898 183506 41134
rect 183742 40898 183826 41134
rect 184062 40898 184094 41134
rect 183474 40814 184094 40898
rect 183474 40578 183506 40814
rect 183742 40578 183826 40814
rect 184062 40578 184094 40814
rect 183474 5134 184094 40578
rect 183474 4898 183506 5134
rect 183742 4898 183826 5134
rect 184062 4898 184094 5134
rect 183474 4814 184094 4898
rect 183474 4578 183506 4814
rect 183742 4578 183826 4814
rect 184062 4578 184094 4814
rect 183474 -2266 184094 4578
rect 183474 -2502 183506 -2266
rect 183742 -2502 183826 -2266
rect 184062 -2502 184094 -2266
rect 183474 -2586 184094 -2502
rect 183474 -2822 183506 -2586
rect 183742 -2822 183826 -2586
rect 184062 -2822 184094 -2586
rect 183474 -7654 184094 -2822
rect 184714 707718 185334 711590
rect 184714 707482 184746 707718
rect 184982 707482 185066 707718
rect 185302 707482 185334 707718
rect 184714 707398 185334 707482
rect 184714 707162 184746 707398
rect 184982 707162 185066 707398
rect 185302 707162 185334 707398
rect 184714 690374 185334 707162
rect 184714 690138 184746 690374
rect 184982 690138 185066 690374
rect 185302 690138 185334 690374
rect 184714 690054 185334 690138
rect 184714 689818 184746 690054
rect 184982 689818 185066 690054
rect 185302 689818 185334 690054
rect 184714 654374 185334 689818
rect 184714 654138 184746 654374
rect 184982 654138 185066 654374
rect 185302 654138 185334 654374
rect 184714 654054 185334 654138
rect 184714 653818 184746 654054
rect 184982 653818 185066 654054
rect 185302 653818 185334 654054
rect 184714 618374 185334 653818
rect 184714 618138 184746 618374
rect 184982 618138 185066 618374
rect 185302 618138 185334 618374
rect 184714 618054 185334 618138
rect 184714 617818 184746 618054
rect 184982 617818 185066 618054
rect 185302 617818 185334 618054
rect 184714 582374 185334 617818
rect 184714 582138 184746 582374
rect 184982 582138 185066 582374
rect 185302 582138 185334 582374
rect 184714 582054 185334 582138
rect 184714 581818 184746 582054
rect 184982 581818 185066 582054
rect 185302 581818 185334 582054
rect 184714 546374 185334 581818
rect 184714 546138 184746 546374
rect 184982 546138 185066 546374
rect 185302 546138 185334 546374
rect 184714 546054 185334 546138
rect 184714 545818 184746 546054
rect 184982 545818 185066 546054
rect 185302 545818 185334 546054
rect 184714 510374 185334 545818
rect 184714 510138 184746 510374
rect 184982 510138 185066 510374
rect 185302 510138 185334 510374
rect 184714 510054 185334 510138
rect 184714 509818 184746 510054
rect 184982 509818 185066 510054
rect 185302 509818 185334 510054
rect 184714 474374 185334 509818
rect 184714 474138 184746 474374
rect 184982 474138 185066 474374
rect 185302 474138 185334 474374
rect 184714 474054 185334 474138
rect 184714 473818 184746 474054
rect 184982 473818 185066 474054
rect 185302 473818 185334 474054
rect 184714 438374 185334 473818
rect 184714 438138 184746 438374
rect 184982 438138 185066 438374
rect 185302 438138 185334 438374
rect 184714 438054 185334 438138
rect 184714 437818 184746 438054
rect 184982 437818 185066 438054
rect 185302 437818 185334 438054
rect 184714 402374 185334 437818
rect 184714 402138 184746 402374
rect 184982 402138 185066 402374
rect 185302 402138 185334 402374
rect 184714 402054 185334 402138
rect 184714 401818 184746 402054
rect 184982 401818 185066 402054
rect 185302 401818 185334 402054
rect 184714 366374 185334 401818
rect 184714 366138 184746 366374
rect 184982 366138 185066 366374
rect 185302 366138 185334 366374
rect 184714 366054 185334 366138
rect 184714 365818 184746 366054
rect 184982 365818 185066 366054
rect 185302 365818 185334 366054
rect 184714 330374 185334 365818
rect 184714 330138 184746 330374
rect 184982 330138 185066 330374
rect 185302 330138 185334 330374
rect 184714 330054 185334 330138
rect 184714 329818 184746 330054
rect 184982 329818 185066 330054
rect 185302 329818 185334 330054
rect 184714 294374 185334 329818
rect 184714 294138 184746 294374
rect 184982 294138 185066 294374
rect 185302 294138 185334 294374
rect 184714 294054 185334 294138
rect 184714 293818 184746 294054
rect 184982 293818 185066 294054
rect 185302 293818 185334 294054
rect 184714 258374 185334 293818
rect 184714 258138 184746 258374
rect 184982 258138 185066 258374
rect 185302 258138 185334 258374
rect 184714 258054 185334 258138
rect 184714 257818 184746 258054
rect 184982 257818 185066 258054
rect 185302 257818 185334 258054
rect 184714 222374 185334 257818
rect 184714 222138 184746 222374
rect 184982 222138 185066 222374
rect 185302 222138 185334 222374
rect 184714 222054 185334 222138
rect 184714 221818 184746 222054
rect 184982 221818 185066 222054
rect 185302 221818 185334 222054
rect 184714 186374 185334 221818
rect 184714 186138 184746 186374
rect 184982 186138 185066 186374
rect 185302 186138 185334 186374
rect 184714 186054 185334 186138
rect 184714 185818 184746 186054
rect 184982 185818 185066 186054
rect 185302 185818 185334 186054
rect 184714 150374 185334 185818
rect 184714 150138 184746 150374
rect 184982 150138 185066 150374
rect 185302 150138 185334 150374
rect 184714 150054 185334 150138
rect 184714 149818 184746 150054
rect 184982 149818 185066 150054
rect 185302 149818 185334 150054
rect 184714 114374 185334 149818
rect 184714 114138 184746 114374
rect 184982 114138 185066 114374
rect 185302 114138 185334 114374
rect 184714 114054 185334 114138
rect 184714 113818 184746 114054
rect 184982 113818 185066 114054
rect 185302 113818 185334 114054
rect 184714 78374 185334 113818
rect 184714 78138 184746 78374
rect 184982 78138 185066 78374
rect 185302 78138 185334 78374
rect 184714 78054 185334 78138
rect 184714 77818 184746 78054
rect 184982 77818 185066 78054
rect 185302 77818 185334 78054
rect 184714 42374 185334 77818
rect 184714 42138 184746 42374
rect 184982 42138 185066 42374
rect 185302 42138 185334 42374
rect 184714 42054 185334 42138
rect 184714 41818 184746 42054
rect 184982 41818 185066 42054
rect 185302 41818 185334 42054
rect 184714 6374 185334 41818
rect 184714 6138 184746 6374
rect 184982 6138 185066 6374
rect 185302 6138 185334 6374
rect 184714 6054 185334 6138
rect 184714 5818 184746 6054
rect 184982 5818 185066 6054
rect 185302 5818 185334 6054
rect 184714 -3226 185334 5818
rect 184714 -3462 184746 -3226
rect 184982 -3462 185066 -3226
rect 185302 -3462 185334 -3226
rect 184714 -3546 185334 -3462
rect 184714 -3782 184746 -3546
rect 184982 -3782 185066 -3546
rect 185302 -3782 185334 -3546
rect 184714 -7654 185334 -3782
rect 185954 708678 186574 711590
rect 185954 708442 185986 708678
rect 186222 708442 186306 708678
rect 186542 708442 186574 708678
rect 185954 708358 186574 708442
rect 185954 708122 185986 708358
rect 186222 708122 186306 708358
rect 186542 708122 186574 708358
rect 185954 691614 186574 708122
rect 185954 691378 185986 691614
rect 186222 691378 186306 691614
rect 186542 691378 186574 691614
rect 185954 691294 186574 691378
rect 185954 691058 185986 691294
rect 186222 691058 186306 691294
rect 186542 691058 186574 691294
rect 185954 655614 186574 691058
rect 185954 655378 185986 655614
rect 186222 655378 186306 655614
rect 186542 655378 186574 655614
rect 185954 655294 186574 655378
rect 185954 655058 185986 655294
rect 186222 655058 186306 655294
rect 186542 655058 186574 655294
rect 185954 619614 186574 655058
rect 185954 619378 185986 619614
rect 186222 619378 186306 619614
rect 186542 619378 186574 619614
rect 185954 619294 186574 619378
rect 185954 619058 185986 619294
rect 186222 619058 186306 619294
rect 186542 619058 186574 619294
rect 185954 583614 186574 619058
rect 185954 583378 185986 583614
rect 186222 583378 186306 583614
rect 186542 583378 186574 583614
rect 185954 583294 186574 583378
rect 185954 583058 185986 583294
rect 186222 583058 186306 583294
rect 186542 583058 186574 583294
rect 185954 547614 186574 583058
rect 185954 547378 185986 547614
rect 186222 547378 186306 547614
rect 186542 547378 186574 547614
rect 185954 547294 186574 547378
rect 185954 547058 185986 547294
rect 186222 547058 186306 547294
rect 186542 547058 186574 547294
rect 185954 511614 186574 547058
rect 185954 511378 185986 511614
rect 186222 511378 186306 511614
rect 186542 511378 186574 511614
rect 185954 511294 186574 511378
rect 185954 511058 185986 511294
rect 186222 511058 186306 511294
rect 186542 511058 186574 511294
rect 185954 475614 186574 511058
rect 185954 475378 185986 475614
rect 186222 475378 186306 475614
rect 186542 475378 186574 475614
rect 185954 475294 186574 475378
rect 185954 475058 185986 475294
rect 186222 475058 186306 475294
rect 186542 475058 186574 475294
rect 185954 439614 186574 475058
rect 185954 439378 185986 439614
rect 186222 439378 186306 439614
rect 186542 439378 186574 439614
rect 185954 439294 186574 439378
rect 185954 439058 185986 439294
rect 186222 439058 186306 439294
rect 186542 439058 186574 439294
rect 185954 403614 186574 439058
rect 185954 403378 185986 403614
rect 186222 403378 186306 403614
rect 186542 403378 186574 403614
rect 185954 403294 186574 403378
rect 185954 403058 185986 403294
rect 186222 403058 186306 403294
rect 186542 403058 186574 403294
rect 185954 367614 186574 403058
rect 185954 367378 185986 367614
rect 186222 367378 186306 367614
rect 186542 367378 186574 367614
rect 185954 367294 186574 367378
rect 185954 367058 185986 367294
rect 186222 367058 186306 367294
rect 186542 367058 186574 367294
rect 185954 331614 186574 367058
rect 185954 331378 185986 331614
rect 186222 331378 186306 331614
rect 186542 331378 186574 331614
rect 185954 331294 186574 331378
rect 185954 331058 185986 331294
rect 186222 331058 186306 331294
rect 186542 331058 186574 331294
rect 185954 295614 186574 331058
rect 185954 295378 185986 295614
rect 186222 295378 186306 295614
rect 186542 295378 186574 295614
rect 185954 295294 186574 295378
rect 185954 295058 185986 295294
rect 186222 295058 186306 295294
rect 186542 295058 186574 295294
rect 185954 259614 186574 295058
rect 185954 259378 185986 259614
rect 186222 259378 186306 259614
rect 186542 259378 186574 259614
rect 185954 259294 186574 259378
rect 185954 259058 185986 259294
rect 186222 259058 186306 259294
rect 186542 259058 186574 259294
rect 185954 223614 186574 259058
rect 185954 223378 185986 223614
rect 186222 223378 186306 223614
rect 186542 223378 186574 223614
rect 185954 223294 186574 223378
rect 185954 223058 185986 223294
rect 186222 223058 186306 223294
rect 186542 223058 186574 223294
rect 185954 187614 186574 223058
rect 185954 187378 185986 187614
rect 186222 187378 186306 187614
rect 186542 187378 186574 187614
rect 185954 187294 186574 187378
rect 185954 187058 185986 187294
rect 186222 187058 186306 187294
rect 186542 187058 186574 187294
rect 185954 151614 186574 187058
rect 185954 151378 185986 151614
rect 186222 151378 186306 151614
rect 186542 151378 186574 151614
rect 185954 151294 186574 151378
rect 185954 151058 185986 151294
rect 186222 151058 186306 151294
rect 186542 151058 186574 151294
rect 185954 115614 186574 151058
rect 185954 115378 185986 115614
rect 186222 115378 186306 115614
rect 186542 115378 186574 115614
rect 185954 115294 186574 115378
rect 185954 115058 185986 115294
rect 186222 115058 186306 115294
rect 186542 115058 186574 115294
rect 185954 79614 186574 115058
rect 185954 79378 185986 79614
rect 186222 79378 186306 79614
rect 186542 79378 186574 79614
rect 185954 79294 186574 79378
rect 185954 79058 185986 79294
rect 186222 79058 186306 79294
rect 186542 79058 186574 79294
rect 185954 43614 186574 79058
rect 185954 43378 185986 43614
rect 186222 43378 186306 43614
rect 186542 43378 186574 43614
rect 185954 43294 186574 43378
rect 185954 43058 185986 43294
rect 186222 43058 186306 43294
rect 186542 43058 186574 43294
rect 185954 7614 186574 43058
rect 185954 7378 185986 7614
rect 186222 7378 186306 7614
rect 186542 7378 186574 7614
rect 185954 7294 186574 7378
rect 185954 7058 185986 7294
rect 186222 7058 186306 7294
rect 186542 7058 186574 7294
rect 185954 -4186 186574 7058
rect 185954 -4422 185986 -4186
rect 186222 -4422 186306 -4186
rect 186542 -4422 186574 -4186
rect 185954 -4506 186574 -4422
rect 185954 -4742 185986 -4506
rect 186222 -4742 186306 -4506
rect 186542 -4742 186574 -4506
rect 185954 -7654 186574 -4742
rect 187194 709638 187814 711590
rect 187194 709402 187226 709638
rect 187462 709402 187546 709638
rect 187782 709402 187814 709638
rect 187194 709318 187814 709402
rect 187194 709082 187226 709318
rect 187462 709082 187546 709318
rect 187782 709082 187814 709318
rect 187194 692854 187814 709082
rect 187194 692618 187226 692854
rect 187462 692618 187546 692854
rect 187782 692618 187814 692854
rect 187194 692534 187814 692618
rect 187194 692298 187226 692534
rect 187462 692298 187546 692534
rect 187782 692298 187814 692534
rect 187194 656854 187814 692298
rect 187194 656618 187226 656854
rect 187462 656618 187546 656854
rect 187782 656618 187814 656854
rect 187194 656534 187814 656618
rect 187194 656298 187226 656534
rect 187462 656298 187546 656534
rect 187782 656298 187814 656534
rect 187194 620854 187814 656298
rect 187194 620618 187226 620854
rect 187462 620618 187546 620854
rect 187782 620618 187814 620854
rect 187194 620534 187814 620618
rect 187194 620298 187226 620534
rect 187462 620298 187546 620534
rect 187782 620298 187814 620534
rect 187194 584854 187814 620298
rect 187194 584618 187226 584854
rect 187462 584618 187546 584854
rect 187782 584618 187814 584854
rect 187194 584534 187814 584618
rect 187194 584298 187226 584534
rect 187462 584298 187546 584534
rect 187782 584298 187814 584534
rect 187194 548854 187814 584298
rect 187194 548618 187226 548854
rect 187462 548618 187546 548854
rect 187782 548618 187814 548854
rect 187194 548534 187814 548618
rect 187194 548298 187226 548534
rect 187462 548298 187546 548534
rect 187782 548298 187814 548534
rect 187194 512854 187814 548298
rect 187194 512618 187226 512854
rect 187462 512618 187546 512854
rect 187782 512618 187814 512854
rect 187194 512534 187814 512618
rect 187194 512298 187226 512534
rect 187462 512298 187546 512534
rect 187782 512298 187814 512534
rect 187194 476854 187814 512298
rect 187194 476618 187226 476854
rect 187462 476618 187546 476854
rect 187782 476618 187814 476854
rect 187194 476534 187814 476618
rect 187194 476298 187226 476534
rect 187462 476298 187546 476534
rect 187782 476298 187814 476534
rect 187194 440854 187814 476298
rect 187194 440618 187226 440854
rect 187462 440618 187546 440854
rect 187782 440618 187814 440854
rect 187194 440534 187814 440618
rect 187194 440298 187226 440534
rect 187462 440298 187546 440534
rect 187782 440298 187814 440534
rect 187194 404854 187814 440298
rect 187194 404618 187226 404854
rect 187462 404618 187546 404854
rect 187782 404618 187814 404854
rect 187194 404534 187814 404618
rect 187194 404298 187226 404534
rect 187462 404298 187546 404534
rect 187782 404298 187814 404534
rect 187194 368854 187814 404298
rect 187194 368618 187226 368854
rect 187462 368618 187546 368854
rect 187782 368618 187814 368854
rect 187194 368534 187814 368618
rect 187194 368298 187226 368534
rect 187462 368298 187546 368534
rect 187782 368298 187814 368534
rect 187194 332854 187814 368298
rect 187194 332618 187226 332854
rect 187462 332618 187546 332854
rect 187782 332618 187814 332854
rect 187194 332534 187814 332618
rect 187194 332298 187226 332534
rect 187462 332298 187546 332534
rect 187782 332298 187814 332534
rect 187194 296854 187814 332298
rect 187194 296618 187226 296854
rect 187462 296618 187546 296854
rect 187782 296618 187814 296854
rect 187194 296534 187814 296618
rect 187194 296298 187226 296534
rect 187462 296298 187546 296534
rect 187782 296298 187814 296534
rect 187194 260854 187814 296298
rect 187194 260618 187226 260854
rect 187462 260618 187546 260854
rect 187782 260618 187814 260854
rect 187194 260534 187814 260618
rect 187194 260298 187226 260534
rect 187462 260298 187546 260534
rect 187782 260298 187814 260534
rect 187194 224854 187814 260298
rect 187194 224618 187226 224854
rect 187462 224618 187546 224854
rect 187782 224618 187814 224854
rect 187194 224534 187814 224618
rect 187194 224298 187226 224534
rect 187462 224298 187546 224534
rect 187782 224298 187814 224534
rect 187194 188854 187814 224298
rect 187194 188618 187226 188854
rect 187462 188618 187546 188854
rect 187782 188618 187814 188854
rect 187194 188534 187814 188618
rect 187194 188298 187226 188534
rect 187462 188298 187546 188534
rect 187782 188298 187814 188534
rect 187194 152854 187814 188298
rect 187194 152618 187226 152854
rect 187462 152618 187546 152854
rect 187782 152618 187814 152854
rect 187194 152534 187814 152618
rect 187194 152298 187226 152534
rect 187462 152298 187546 152534
rect 187782 152298 187814 152534
rect 187194 116854 187814 152298
rect 187194 116618 187226 116854
rect 187462 116618 187546 116854
rect 187782 116618 187814 116854
rect 187194 116534 187814 116618
rect 187194 116298 187226 116534
rect 187462 116298 187546 116534
rect 187782 116298 187814 116534
rect 187194 80854 187814 116298
rect 187194 80618 187226 80854
rect 187462 80618 187546 80854
rect 187782 80618 187814 80854
rect 187194 80534 187814 80618
rect 187194 80298 187226 80534
rect 187462 80298 187546 80534
rect 187782 80298 187814 80534
rect 187194 44854 187814 80298
rect 187194 44618 187226 44854
rect 187462 44618 187546 44854
rect 187782 44618 187814 44854
rect 187194 44534 187814 44618
rect 187194 44298 187226 44534
rect 187462 44298 187546 44534
rect 187782 44298 187814 44534
rect 187194 8854 187814 44298
rect 187194 8618 187226 8854
rect 187462 8618 187546 8854
rect 187782 8618 187814 8854
rect 187194 8534 187814 8618
rect 187194 8298 187226 8534
rect 187462 8298 187546 8534
rect 187782 8298 187814 8534
rect 187194 -5146 187814 8298
rect 187194 -5382 187226 -5146
rect 187462 -5382 187546 -5146
rect 187782 -5382 187814 -5146
rect 187194 -5466 187814 -5382
rect 187194 -5702 187226 -5466
rect 187462 -5702 187546 -5466
rect 187782 -5702 187814 -5466
rect 187194 -7654 187814 -5702
rect 188434 710598 189054 711590
rect 188434 710362 188466 710598
rect 188702 710362 188786 710598
rect 189022 710362 189054 710598
rect 188434 710278 189054 710362
rect 188434 710042 188466 710278
rect 188702 710042 188786 710278
rect 189022 710042 189054 710278
rect 188434 694094 189054 710042
rect 188434 693858 188466 694094
rect 188702 693858 188786 694094
rect 189022 693858 189054 694094
rect 188434 693774 189054 693858
rect 188434 693538 188466 693774
rect 188702 693538 188786 693774
rect 189022 693538 189054 693774
rect 188434 658094 189054 693538
rect 188434 657858 188466 658094
rect 188702 657858 188786 658094
rect 189022 657858 189054 658094
rect 188434 657774 189054 657858
rect 188434 657538 188466 657774
rect 188702 657538 188786 657774
rect 189022 657538 189054 657774
rect 188434 622094 189054 657538
rect 188434 621858 188466 622094
rect 188702 621858 188786 622094
rect 189022 621858 189054 622094
rect 188434 621774 189054 621858
rect 188434 621538 188466 621774
rect 188702 621538 188786 621774
rect 189022 621538 189054 621774
rect 188434 586094 189054 621538
rect 188434 585858 188466 586094
rect 188702 585858 188786 586094
rect 189022 585858 189054 586094
rect 188434 585774 189054 585858
rect 188434 585538 188466 585774
rect 188702 585538 188786 585774
rect 189022 585538 189054 585774
rect 188434 550094 189054 585538
rect 188434 549858 188466 550094
rect 188702 549858 188786 550094
rect 189022 549858 189054 550094
rect 188434 549774 189054 549858
rect 188434 549538 188466 549774
rect 188702 549538 188786 549774
rect 189022 549538 189054 549774
rect 188434 514094 189054 549538
rect 188434 513858 188466 514094
rect 188702 513858 188786 514094
rect 189022 513858 189054 514094
rect 188434 513774 189054 513858
rect 188434 513538 188466 513774
rect 188702 513538 188786 513774
rect 189022 513538 189054 513774
rect 188434 478094 189054 513538
rect 188434 477858 188466 478094
rect 188702 477858 188786 478094
rect 189022 477858 189054 478094
rect 188434 477774 189054 477858
rect 188434 477538 188466 477774
rect 188702 477538 188786 477774
rect 189022 477538 189054 477774
rect 188434 442094 189054 477538
rect 188434 441858 188466 442094
rect 188702 441858 188786 442094
rect 189022 441858 189054 442094
rect 188434 441774 189054 441858
rect 188434 441538 188466 441774
rect 188702 441538 188786 441774
rect 189022 441538 189054 441774
rect 188434 406094 189054 441538
rect 188434 405858 188466 406094
rect 188702 405858 188786 406094
rect 189022 405858 189054 406094
rect 188434 405774 189054 405858
rect 188434 405538 188466 405774
rect 188702 405538 188786 405774
rect 189022 405538 189054 405774
rect 188434 370094 189054 405538
rect 188434 369858 188466 370094
rect 188702 369858 188786 370094
rect 189022 369858 189054 370094
rect 188434 369774 189054 369858
rect 188434 369538 188466 369774
rect 188702 369538 188786 369774
rect 189022 369538 189054 369774
rect 188434 334094 189054 369538
rect 188434 333858 188466 334094
rect 188702 333858 188786 334094
rect 189022 333858 189054 334094
rect 188434 333774 189054 333858
rect 188434 333538 188466 333774
rect 188702 333538 188786 333774
rect 189022 333538 189054 333774
rect 188434 298094 189054 333538
rect 188434 297858 188466 298094
rect 188702 297858 188786 298094
rect 189022 297858 189054 298094
rect 188434 297774 189054 297858
rect 188434 297538 188466 297774
rect 188702 297538 188786 297774
rect 189022 297538 189054 297774
rect 188434 262094 189054 297538
rect 188434 261858 188466 262094
rect 188702 261858 188786 262094
rect 189022 261858 189054 262094
rect 188434 261774 189054 261858
rect 188434 261538 188466 261774
rect 188702 261538 188786 261774
rect 189022 261538 189054 261774
rect 188434 226094 189054 261538
rect 188434 225858 188466 226094
rect 188702 225858 188786 226094
rect 189022 225858 189054 226094
rect 188434 225774 189054 225858
rect 188434 225538 188466 225774
rect 188702 225538 188786 225774
rect 189022 225538 189054 225774
rect 188434 190094 189054 225538
rect 188434 189858 188466 190094
rect 188702 189858 188786 190094
rect 189022 189858 189054 190094
rect 188434 189774 189054 189858
rect 188434 189538 188466 189774
rect 188702 189538 188786 189774
rect 189022 189538 189054 189774
rect 188434 154094 189054 189538
rect 188434 153858 188466 154094
rect 188702 153858 188786 154094
rect 189022 153858 189054 154094
rect 188434 153774 189054 153858
rect 188434 153538 188466 153774
rect 188702 153538 188786 153774
rect 189022 153538 189054 153774
rect 188434 118094 189054 153538
rect 188434 117858 188466 118094
rect 188702 117858 188786 118094
rect 189022 117858 189054 118094
rect 188434 117774 189054 117858
rect 188434 117538 188466 117774
rect 188702 117538 188786 117774
rect 189022 117538 189054 117774
rect 188434 82094 189054 117538
rect 188434 81858 188466 82094
rect 188702 81858 188786 82094
rect 189022 81858 189054 82094
rect 188434 81774 189054 81858
rect 188434 81538 188466 81774
rect 188702 81538 188786 81774
rect 189022 81538 189054 81774
rect 188434 46094 189054 81538
rect 188434 45858 188466 46094
rect 188702 45858 188786 46094
rect 189022 45858 189054 46094
rect 188434 45774 189054 45858
rect 188434 45538 188466 45774
rect 188702 45538 188786 45774
rect 189022 45538 189054 45774
rect 188434 10094 189054 45538
rect 188434 9858 188466 10094
rect 188702 9858 188786 10094
rect 189022 9858 189054 10094
rect 188434 9774 189054 9858
rect 188434 9538 188466 9774
rect 188702 9538 188786 9774
rect 189022 9538 189054 9774
rect 188434 -6106 189054 9538
rect 188434 -6342 188466 -6106
rect 188702 -6342 188786 -6106
rect 189022 -6342 189054 -6106
rect 188434 -6426 189054 -6342
rect 188434 -6662 188466 -6426
rect 188702 -6662 188786 -6426
rect 189022 -6662 189054 -6426
rect 188434 -7654 189054 -6662
rect 189674 711558 190294 711590
rect 189674 711322 189706 711558
rect 189942 711322 190026 711558
rect 190262 711322 190294 711558
rect 189674 711238 190294 711322
rect 189674 711002 189706 711238
rect 189942 711002 190026 711238
rect 190262 711002 190294 711238
rect 189674 695334 190294 711002
rect 189674 695098 189706 695334
rect 189942 695098 190026 695334
rect 190262 695098 190294 695334
rect 189674 695014 190294 695098
rect 189674 694778 189706 695014
rect 189942 694778 190026 695014
rect 190262 694778 190294 695014
rect 189674 659334 190294 694778
rect 189674 659098 189706 659334
rect 189942 659098 190026 659334
rect 190262 659098 190294 659334
rect 189674 659014 190294 659098
rect 189674 658778 189706 659014
rect 189942 658778 190026 659014
rect 190262 658778 190294 659014
rect 189674 623334 190294 658778
rect 189674 623098 189706 623334
rect 189942 623098 190026 623334
rect 190262 623098 190294 623334
rect 189674 623014 190294 623098
rect 189674 622778 189706 623014
rect 189942 622778 190026 623014
rect 190262 622778 190294 623014
rect 189674 587334 190294 622778
rect 189674 587098 189706 587334
rect 189942 587098 190026 587334
rect 190262 587098 190294 587334
rect 189674 587014 190294 587098
rect 189674 586778 189706 587014
rect 189942 586778 190026 587014
rect 190262 586778 190294 587014
rect 189674 551334 190294 586778
rect 189674 551098 189706 551334
rect 189942 551098 190026 551334
rect 190262 551098 190294 551334
rect 189674 551014 190294 551098
rect 189674 550778 189706 551014
rect 189942 550778 190026 551014
rect 190262 550778 190294 551014
rect 189674 515334 190294 550778
rect 189674 515098 189706 515334
rect 189942 515098 190026 515334
rect 190262 515098 190294 515334
rect 189674 515014 190294 515098
rect 189674 514778 189706 515014
rect 189942 514778 190026 515014
rect 190262 514778 190294 515014
rect 189674 479334 190294 514778
rect 189674 479098 189706 479334
rect 189942 479098 190026 479334
rect 190262 479098 190294 479334
rect 189674 479014 190294 479098
rect 189674 478778 189706 479014
rect 189942 478778 190026 479014
rect 190262 478778 190294 479014
rect 189674 443334 190294 478778
rect 189674 443098 189706 443334
rect 189942 443098 190026 443334
rect 190262 443098 190294 443334
rect 189674 443014 190294 443098
rect 189674 442778 189706 443014
rect 189942 442778 190026 443014
rect 190262 442778 190294 443014
rect 189674 407334 190294 442778
rect 189674 407098 189706 407334
rect 189942 407098 190026 407334
rect 190262 407098 190294 407334
rect 189674 407014 190294 407098
rect 189674 406778 189706 407014
rect 189942 406778 190026 407014
rect 190262 406778 190294 407014
rect 189674 371334 190294 406778
rect 189674 371098 189706 371334
rect 189942 371098 190026 371334
rect 190262 371098 190294 371334
rect 189674 371014 190294 371098
rect 189674 370778 189706 371014
rect 189942 370778 190026 371014
rect 190262 370778 190294 371014
rect 189674 335334 190294 370778
rect 189674 335098 189706 335334
rect 189942 335098 190026 335334
rect 190262 335098 190294 335334
rect 189674 335014 190294 335098
rect 189674 334778 189706 335014
rect 189942 334778 190026 335014
rect 190262 334778 190294 335014
rect 189674 299334 190294 334778
rect 189674 299098 189706 299334
rect 189942 299098 190026 299334
rect 190262 299098 190294 299334
rect 189674 299014 190294 299098
rect 189674 298778 189706 299014
rect 189942 298778 190026 299014
rect 190262 298778 190294 299014
rect 189674 263334 190294 298778
rect 189674 263098 189706 263334
rect 189942 263098 190026 263334
rect 190262 263098 190294 263334
rect 189674 263014 190294 263098
rect 189674 262778 189706 263014
rect 189942 262778 190026 263014
rect 190262 262778 190294 263014
rect 189674 227334 190294 262778
rect 189674 227098 189706 227334
rect 189942 227098 190026 227334
rect 190262 227098 190294 227334
rect 189674 227014 190294 227098
rect 189674 226778 189706 227014
rect 189942 226778 190026 227014
rect 190262 226778 190294 227014
rect 189674 191334 190294 226778
rect 189674 191098 189706 191334
rect 189942 191098 190026 191334
rect 190262 191098 190294 191334
rect 189674 191014 190294 191098
rect 189674 190778 189706 191014
rect 189942 190778 190026 191014
rect 190262 190778 190294 191014
rect 189674 155334 190294 190778
rect 189674 155098 189706 155334
rect 189942 155098 190026 155334
rect 190262 155098 190294 155334
rect 189674 155014 190294 155098
rect 189674 154778 189706 155014
rect 189942 154778 190026 155014
rect 190262 154778 190294 155014
rect 189674 119334 190294 154778
rect 189674 119098 189706 119334
rect 189942 119098 190026 119334
rect 190262 119098 190294 119334
rect 189674 119014 190294 119098
rect 189674 118778 189706 119014
rect 189942 118778 190026 119014
rect 190262 118778 190294 119014
rect 189674 83334 190294 118778
rect 189674 83098 189706 83334
rect 189942 83098 190026 83334
rect 190262 83098 190294 83334
rect 189674 83014 190294 83098
rect 189674 82778 189706 83014
rect 189942 82778 190026 83014
rect 190262 82778 190294 83014
rect 189674 47334 190294 82778
rect 189674 47098 189706 47334
rect 189942 47098 190026 47334
rect 190262 47098 190294 47334
rect 189674 47014 190294 47098
rect 189674 46778 189706 47014
rect 189942 46778 190026 47014
rect 190262 46778 190294 47014
rect 189674 11334 190294 46778
rect 189674 11098 189706 11334
rect 189942 11098 190026 11334
rect 190262 11098 190294 11334
rect 189674 11014 190294 11098
rect 189674 10778 189706 11014
rect 189942 10778 190026 11014
rect 190262 10778 190294 11014
rect 189674 -7066 190294 10778
rect 189674 -7302 189706 -7066
rect 189942 -7302 190026 -7066
rect 190262 -7302 190294 -7066
rect 189674 -7386 190294 -7302
rect 189674 -7622 189706 -7386
rect 189942 -7622 190026 -7386
rect 190262 -7622 190294 -7386
rect 189674 -7654 190294 -7622
rect 216994 704838 217614 711590
rect 216994 704602 217026 704838
rect 217262 704602 217346 704838
rect 217582 704602 217614 704838
rect 216994 704518 217614 704602
rect 216994 704282 217026 704518
rect 217262 704282 217346 704518
rect 217582 704282 217614 704518
rect 216994 686654 217614 704282
rect 216994 686418 217026 686654
rect 217262 686418 217346 686654
rect 217582 686418 217614 686654
rect 216994 686334 217614 686418
rect 216994 686098 217026 686334
rect 217262 686098 217346 686334
rect 217582 686098 217614 686334
rect 216994 650654 217614 686098
rect 216994 650418 217026 650654
rect 217262 650418 217346 650654
rect 217582 650418 217614 650654
rect 216994 650334 217614 650418
rect 216994 650098 217026 650334
rect 217262 650098 217346 650334
rect 217582 650098 217614 650334
rect 216994 614654 217614 650098
rect 216994 614418 217026 614654
rect 217262 614418 217346 614654
rect 217582 614418 217614 614654
rect 216994 614334 217614 614418
rect 216994 614098 217026 614334
rect 217262 614098 217346 614334
rect 217582 614098 217614 614334
rect 216994 578654 217614 614098
rect 216994 578418 217026 578654
rect 217262 578418 217346 578654
rect 217582 578418 217614 578654
rect 216994 578334 217614 578418
rect 216994 578098 217026 578334
rect 217262 578098 217346 578334
rect 217582 578098 217614 578334
rect 216994 542654 217614 578098
rect 216994 542418 217026 542654
rect 217262 542418 217346 542654
rect 217582 542418 217614 542654
rect 216994 542334 217614 542418
rect 216994 542098 217026 542334
rect 217262 542098 217346 542334
rect 217582 542098 217614 542334
rect 216994 506654 217614 542098
rect 216994 506418 217026 506654
rect 217262 506418 217346 506654
rect 217582 506418 217614 506654
rect 216994 506334 217614 506418
rect 216994 506098 217026 506334
rect 217262 506098 217346 506334
rect 217582 506098 217614 506334
rect 216994 470654 217614 506098
rect 216994 470418 217026 470654
rect 217262 470418 217346 470654
rect 217582 470418 217614 470654
rect 216994 470334 217614 470418
rect 216994 470098 217026 470334
rect 217262 470098 217346 470334
rect 217582 470098 217614 470334
rect 216994 434654 217614 470098
rect 216994 434418 217026 434654
rect 217262 434418 217346 434654
rect 217582 434418 217614 434654
rect 216994 434334 217614 434418
rect 216994 434098 217026 434334
rect 217262 434098 217346 434334
rect 217582 434098 217614 434334
rect 216994 398654 217614 434098
rect 216994 398418 217026 398654
rect 217262 398418 217346 398654
rect 217582 398418 217614 398654
rect 216994 398334 217614 398418
rect 216994 398098 217026 398334
rect 217262 398098 217346 398334
rect 217582 398098 217614 398334
rect 216994 362654 217614 398098
rect 216994 362418 217026 362654
rect 217262 362418 217346 362654
rect 217582 362418 217614 362654
rect 216994 362334 217614 362418
rect 216994 362098 217026 362334
rect 217262 362098 217346 362334
rect 217582 362098 217614 362334
rect 216994 326654 217614 362098
rect 216994 326418 217026 326654
rect 217262 326418 217346 326654
rect 217582 326418 217614 326654
rect 216994 326334 217614 326418
rect 216994 326098 217026 326334
rect 217262 326098 217346 326334
rect 217582 326098 217614 326334
rect 216994 290654 217614 326098
rect 216994 290418 217026 290654
rect 217262 290418 217346 290654
rect 217582 290418 217614 290654
rect 216994 290334 217614 290418
rect 216994 290098 217026 290334
rect 217262 290098 217346 290334
rect 217582 290098 217614 290334
rect 216994 254654 217614 290098
rect 216994 254418 217026 254654
rect 217262 254418 217346 254654
rect 217582 254418 217614 254654
rect 216994 254334 217614 254418
rect 216994 254098 217026 254334
rect 217262 254098 217346 254334
rect 217582 254098 217614 254334
rect 216994 218654 217614 254098
rect 216994 218418 217026 218654
rect 217262 218418 217346 218654
rect 217582 218418 217614 218654
rect 216994 218334 217614 218418
rect 216994 218098 217026 218334
rect 217262 218098 217346 218334
rect 217582 218098 217614 218334
rect 216994 182654 217614 218098
rect 216994 182418 217026 182654
rect 217262 182418 217346 182654
rect 217582 182418 217614 182654
rect 216994 182334 217614 182418
rect 216994 182098 217026 182334
rect 217262 182098 217346 182334
rect 217582 182098 217614 182334
rect 216994 146654 217614 182098
rect 216994 146418 217026 146654
rect 217262 146418 217346 146654
rect 217582 146418 217614 146654
rect 216994 146334 217614 146418
rect 216994 146098 217026 146334
rect 217262 146098 217346 146334
rect 217582 146098 217614 146334
rect 216994 110654 217614 146098
rect 216994 110418 217026 110654
rect 217262 110418 217346 110654
rect 217582 110418 217614 110654
rect 216994 110334 217614 110418
rect 216994 110098 217026 110334
rect 217262 110098 217346 110334
rect 217582 110098 217614 110334
rect 216994 74654 217614 110098
rect 216994 74418 217026 74654
rect 217262 74418 217346 74654
rect 217582 74418 217614 74654
rect 216994 74334 217614 74418
rect 216994 74098 217026 74334
rect 217262 74098 217346 74334
rect 217582 74098 217614 74334
rect 216994 38654 217614 74098
rect 216994 38418 217026 38654
rect 217262 38418 217346 38654
rect 217582 38418 217614 38654
rect 216994 38334 217614 38418
rect 216994 38098 217026 38334
rect 217262 38098 217346 38334
rect 217582 38098 217614 38334
rect 216994 2654 217614 38098
rect 216994 2418 217026 2654
rect 217262 2418 217346 2654
rect 217582 2418 217614 2654
rect 216994 2334 217614 2418
rect 216994 2098 217026 2334
rect 217262 2098 217346 2334
rect 217582 2098 217614 2334
rect 216994 -346 217614 2098
rect 216994 -582 217026 -346
rect 217262 -582 217346 -346
rect 217582 -582 217614 -346
rect 216994 -666 217614 -582
rect 216994 -902 217026 -666
rect 217262 -902 217346 -666
rect 217582 -902 217614 -666
rect 216994 -7654 217614 -902
rect 218234 705798 218854 711590
rect 218234 705562 218266 705798
rect 218502 705562 218586 705798
rect 218822 705562 218854 705798
rect 218234 705478 218854 705562
rect 218234 705242 218266 705478
rect 218502 705242 218586 705478
rect 218822 705242 218854 705478
rect 218234 687894 218854 705242
rect 218234 687658 218266 687894
rect 218502 687658 218586 687894
rect 218822 687658 218854 687894
rect 218234 687574 218854 687658
rect 218234 687338 218266 687574
rect 218502 687338 218586 687574
rect 218822 687338 218854 687574
rect 218234 651894 218854 687338
rect 218234 651658 218266 651894
rect 218502 651658 218586 651894
rect 218822 651658 218854 651894
rect 218234 651574 218854 651658
rect 218234 651338 218266 651574
rect 218502 651338 218586 651574
rect 218822 651338 218854 651574
rect 218234 615894 218854 651338
rect 218234 615658 218266 615894
rect 218502 615658 218586 615894
rect 218822 615658 218854 615894
rect 218234 615574 218854 615658
rect 218234 615338 218266 615574
rect 218502 615338 218586 615574
rect 218822 615338 218854 615574
rect 218234 579894 218854 615338
rect 218234 579658 218266 579894
rect 218502 579658 218586 579894
rect 218822 579658 218854 579894
rect 218234 579574 218854 579658
rect 218234 579338 218266 579574
rect 218502 579338 218586 579574
rect 218822 579338 218854 579574
rect 218234 543894 218854 579338
rect 218234 543658 218266 543894
rect 218502 543658 218586 543894
rect 218822 543658 218854 543894
rect 218234 543574 218854 543658
rect 218234 543338 218266 543574
rect 218502 543338 218586 543574
rect 218822 543338 218854 543574
rect 218234 507894 218854 543338
rect 218234 507658 218266 507894
rect 218502 507658 218586 507894
rect 218822 507658 218854 507894
rect 218234 507574 218854 507658
rect 218234 507338 218266 507574
rect 218502 507338 218586 507574
rect 218822 507338 218854 507574
rect 218234 471894 218854 507338
rect 218234 471658 218266 471894
rect 218502 471658 218586 471894
rect 218822 471658 218854 471894
rect 218234 471574 218854 471658
rect 218234 471338 218266 471574
rect 218502 471338 218586 471574
rect 218822 471338 218854 471574
rect 218234 435894 218854 471338
rect 218234 435658 218266 435894
rect 218502 435658 218586 435894
rect 218822 435658 218854 435894
rect 218234 435574 218854 435658
rect 218234 435338 218266 435574
rect 218502 435338 218586 435574
rect 218822 435338 218854 435574
rect 218234 399894 218854 435338
rect 218234 399658 218266 399894
rect 218502 399658 218586 399894
rect 218822 399658 218854 399894
rect 218234 399574 218854 399658
rect 218234 399338 218266 399574
rect 218502 399338 218586 399574
rect 218822 399338 218854 399574
rect 218234 363894 218854 399338
rect 218234 363658 218266 363894
rect 218502 363658 218586 363894
rect 218822 363658 218854 363894
rect 218234 363574 218854 363658
rect 218234 363338 218266 363574
rect 218502 363338 218586 363574
rect 218822 363338 218854 363574
rect 218234 327894 218854 363338
rect 218234 327658 218266 327894
rect 218502 327658 218586 327894
rect 218822 327658 218854 327894
rect 218234 327574 218854 327658
rect 218234 327338 218266 327574
rect 218502 327338 218586 327574
rect 218822 327338 218854 327574
rect 218234 291894 218854 327338
rect 218234 291658 218266 291894
rect 218502 291658 218586 291894
rect 218822 291658 218854 291894
rect 218234 291574 218854 291658
rect 218234 291338 218266 291574
rect 218502 291338 218586 291574
rect 218822 291338 218854 291574
rect 218234 255894 218854 291338
rect 218234 255658 218266 255894
rect 218502 255658 218586 255894
rect 218822 255658 218854 255894
rect 218234 255574 218854 255658
rect 218234 255338 218266 255574
rect 218502 255338 218586 255574
rect 218822 255338 218854 255574
rect 218234 219894 218854 255338
rect 218234 219658 218266 219894
rect 218502 219658 218586 219894
rect 218822 219658 218854 219894
rect 218234 219574 218854 219658
rect 218234 219338 218266 219574
rect 218502 219338 218586 219574
rect 218822 219338 218854 219574
rect 218234 183894 218854 219338
rect 218234 183658 218266 183894
rect 218502 183658 218586 183894
rect 218822 183658 218854 183894
rect 218234 183574 218854 183658
rect 218234 183338 218266 183574
rect 218502 183338 218586 183574
rect 218822 183338 218854 183574
rect 218234 147894 218854 183338
rect 218234 147658 218266 147894
rect 218502 147658 218586 147894
rect 218822 147658 218854 147894
rect 218234 147574 218854 147658
rect 218234 147338 218266 147574
rect 218502 147338 218586 147574
rect 218822 147338 218854 147574
rect 218234 111894 218854 147338
rect 218234 111658 218266 111894
rect 218502 111658 218586 111894
rect 218822 111658 218854 111894
rect 218234 111574 218854 111658
rect 218234 111338 218266 111574
rect 218502 111338 218586 111574
rect 218822 111338 218854 111574
rect 218234 75894 218854 111338
rect 218234 75658 218266 75894
rect 218502 75658 218586 75894
rect 218822 75658 218854 75894
rect 218234 75574 218854 75658
rect 218234 75338 218266 75574
rect 218502 75338 218586 75574
rect 218822 75338 218854 75574
rect 218234 39894 218854 75338
rect 218234 39658 218266 39894
rect 218502 39658 218586 39894
rect 218822 39658 218854 39894
rect 218234 39574 218854 39658
rect 218234 39338 218266 39574
rect 218502 39338 218586 39574
rect 218822 39338 218854 39574
rect 218234 3894 218854 39338
rect 218234 3658 218266 3894
rect 218502 3658 218586 3894
rect 218822 3658 218854 3894
rect 218234 3574 218854 3658
rect 218234 3338 218266 3574
rect 218502 3338 218586 3574
rect 218822 3338 218854 3574
rect 218234 -1306 218854 3338
rect 218234 -1542 218266 -1306
rect 218502 -1542 218586 -1306
rect 218822 -1542 218854 -1306
rect 218234 -1626 218854 -1542
rect 218234 -1862 218266 -1626
rect 218502 -1862 218586 -1626
rect 218822 -1862 218854 -1626
rect 218234 -7654 218854 -1862
rect 219474 706758 220094 711590
rect 219474 706522 219506 706758
rect 219742 706522 219826 706758
rect 220062 706522 220094 706758
rect 219474 706438 220094 706522
rect 219474 706202 219506 706438
rect 219742 706202 219826 706438
rect 220062 706202 220094 706438
rect 219474 689134 220094 706202
rect 219474 688898 219506 689134
rect 219742 688898 219826 689134
rect 220062 688898 220094 689134
rect 219474 688814 220094 688898
rect 219474 688578 219506 688814
rect 219742 688578 219826 688814
rect 220062 688578 220094 688814
rect 219474 653134 220094 688578
rect 219474 652898 219506 653134
rect 219742 652898 219826 653134
rect 220062 652898 220094 653134
rect 219474 652814 220094 652898
rect 219474 652578 219506 652814
rect 219742 652578 219826 652814
rect 220062 652578 220094 652814
rect 219474 617134 220094 652578
rect 219474 616898 219506 617134
rect 219742 616898 219826 617134
rect 220062 616898 220094 617134
rect 219474 616814 220094 616898
rect 219474 616578 219506 616814
rect 219742 616578 219826 616814
rect 220062 616578 220094 616814
rect 219474 581134 220094 616578
rect 219474 580898 219506 581134
rect 219742 580898 219826 581134
rect 220062 580898 220094 581134
rect 219474 580814 220094 580898
rect 219474 580578 219506 580814
rect 219742 580578 219826 580814
rect 220062 580578 220094 580814
rect 219474 545134 220094 580578
rect 219474 544898 219506 545134
rect 219742 544898 219826 545134
rect 220062 544898 220094 545134
rect 219474 544814 220094 544898
rect 219474 544578 219506 544814
rect 219742 544578 219826 544814
rect 220062 544578 220094 544814
rect 219474 509134 220094 544578
rect 219474 508898 219506 509134
rect 219742 508898 219826 509134
rect 220062 508898 220094 509134
rect 219474 508814 220094 508898
rect 219474 508578 219506 508814
rect 219742 508578 219826 508814
rect 220062 508578 220094 508814
rect 219474 473134 220094 508578
rect 219474 472898 219506 473134
rect 219742 472898 219826 473134
rect 220062 472898 220094 473134
rect 219474 472814 220094 472898
rect 219474 472578 219506 472814
rect 219742 472578 219826 472814
rect 220062 472578 220094 472814
rect 219474 437134 220094 472578
rect 219474 436898 219506 437134
rect 219742 436898 219826 437134
rect 220062 436898 220094 437134
rect 219474 436814 220094 436898
rect 219474 436578 219506 436814
rect 219742 436578 219826 436814
rect 220062 436578 220094 436814
rect 219474 401134 220094 436578
rect 219474 400898 219506 401134
rect 219742 400898 219826 401134
rect 220062 400898 220094 401134
rect 219474 400814 220094 400898
rect 219474 400578 219506 400814
rect 219742 400578 219826 400814
rect 220062 400578 220094 400814
rect 219474 365134 220094 400578
rect 219474 364898 219506 365134
rect 219742 364898 219826 365134
rect 220062 364898 220094 365134
rect 219474 364814 220094 364898
rect 219474 364578 219506 364814
rect 219742 364578 219826 364814
rect 220062 364578 220094 364814
rect 219474 329134 220094 364578
rect 219474 328898 219506 329134
rect 219742 328898 219826 329134
rect 220062 328898 220094 329134
rect 219474 328814 220094 328898
rect 219474 328578 219506 328814
rect 219742 328578 219826 328814
rect 220062 328578 220094 328814
rect 219474 293134 220094 328578
rect 219474 292898 219506 293134
rect 219742 292898 219826 293134
rect 220062 292898 220094 293134
rect 219474 292814 220094 292898
rect 219474 292578 219506 292814
rect 219742 292578 219826 292814
rect 220062 292578 220094 292814
rect 219474 257134 220094 292578
rect 219474 256898 219506 257134
rect 219742 256898 219826 257134
rect 220062 256898 220094 257134
rect 219474 256814 220094 256898
rect 219474 256578 219506 256814
rect 219742 256578 219826 256814
rect 220062 256578 220094 256814
rect 219474 221134 220094 256578
rect 219474 220898 219506 221134
rect 219742 220898 219826 221134
rect 220062 220898 220094 221134
rect 219474 220814 220094 220898
rect 219474 220578 219506 220814
rect 219742 220578 219826 220814
rect 220062 220578 220094 220814
rect 219474 185134 220094 220578
rect 219474 184898 219506 185134
rect 219742 184898 219826 185134
rect 220062 184898 220094 185134
rect 219474 184814 220094 184898
rect 219474 184578 219506 184814
rect 219742 184578 219826 184814
rect 220062 184578 220094 184814
rect 219474 149134 220094 184578
rect 219474 148898 219506 149134
rect 219742 148898 219826 149134
rect 220062 148898 220094 149134
rect 219474 148814 220094 148898
rect 219474 148578 219506 148814
rect 219742 148578 219826 148814
rect 220062 148578 220094 148814
rect 219474 113134 220094 148578
rect 219474 112898 219506 113134
rect 219742 112898 219826 113134
rect 220062 112898 220094 113134
rect 219474 112814 220094 112898
rect 219474 112578 219506 112814
rect 219742 112578 219826 112814
rect 220062 112578 220094 112814
rect 219474 77134 220094 112578
rect 219474 76898 219506 77134
rect 219742 76898 219826 77134
rect 220062 76898 220094 77134
rect 219474 76814 220094 76898
rect 219474 76578 219506 76814
rect 219742 76578 219826 76814
rect 220062 76578 220094 76814
rect 219474 41134 220094 76578
rect 219474 40898 219506 41134
rect 219742 40898 219826 41134
rect 220062 40898 220094 41134
rect 219474 40814 220094 40898
rect 219474 40578 219506 40814
rect 219742 40578 219826 40814
rect 220062 40578 220094 40814
rect 219474 5134 220094 40578
rect 219474 4898 219506 5134
rect 219742 4898 219826 5134
rect 220062 4898 220094 5134
rect 219474 4814 220094 4898
rect 219474 4578 219506 4814
rect 219742 4578 219826 4814
rect 220062 4578 220094 4814
rect 219474 -2266 220094 4578
rect 219474 -2502 219506 -2266
rect 219742 -2502 219826 -2266
rect 220062 -2502 220094 -2266
rect 219474 -2586 220094 -2502
rect 219474 -2822 219506 -2586
rect 219742 -2822 219826 -2586
rect 220062 -2822 220094 -2586
rect 219474 -7654 220094 -2822
rect 220714 707718 221334 711590
rect 220714 707482 220746 707718
rect 220982 707482 221066 707718
rect 221302 707482 221334 707718
rect 220714 707398 221334 707482
rect 220714 707162 220746 707398
rect 220982 707162 221066 707398
rect 221302 707162 221334 707398
rect 220714 690374 221334 707162
rect 220714 690138 220746 690374
rect 220982 690138 221066 690374
rect 221302 690138 221334 690374
rect 220714 690054 221334 690138
rect 220714 689818 220746 690054
rect 220982 689818 221066 690054
rect 221302 689818 221334 690054
rect 220714 654374 221334 689818
rect 220714 654138 220746 654374
rect 220982 654138 221066 654374
rect 221302 654138 221334 654374
rect 220714 654054 221334 654138
rect 220714 653818 220746 654054
rect 220982 653818 221066 654054
rect 221302 653818 221334 654054
rect 220714 618374 221334 653818
rect 220714 618138 220746 618374
rect 220982 618138 221066 618374
rect 221302 618138 221334 618374
rect 220714 618054 221334 618138
rect 220714 617818 220746 618054
rect 220982 617818 221066 618054
rect 221302 617818 221334 618054
rect 220714 582374 221334 617818
rect 220714 582138 220746 582374
rect 220982 582138 221066 582374
rect 221302 582138 221334 582374
rect 220714 582054 221334 582138
rect 220714 581818 220746 582054
rect 220982 581818 221066 582054
rect 221302 581818 221334 582054
rect 220714 546374 221334 581818
rect 220714 546138 220746 546374
rect 220982 546138 221066 546374
rect 221302 546138 221334 546374
rect 220714 546054 221334 546138
rect 220714 545818 220746 546054
rect 220982 545818 221066 546054
rect 221302 545818 221334 546054
rect 220714 510374 221334 545818
rect 220714 510138 220746 510374
rect 220982 510138 221066 510374
rect 221302 510138 221334 510374
rect 220714 510054 221334 510138
rect 220714 509818 220746 510054
rect 220982 509818 221066 510054
rect 221302 509818 221334 510054
rect 220714 474374 221334 509818
rect 220714 474138 220746 474374
rect 220982 474138 221066 474374
rect 221302 474138 221334 474374
rect 220714 474054 221334 474138
rect 220714 473818 220746 474054
rect 220982 473818 221066 474054
rect 221302 473818 221334 474054
rect 220714 438374 221334 473818
rect 220714 438138 220746 438374
rect 220982 438138 221066 438374
rect 221302 438138 221334 438374
rect 220714 438054 221334 438138
rect 220714 437818 220746 438054
rect 220982 437818 221066 438054
rect 221302 437818 221334 438054
rect 220714 402374 221334 437818
rect 220714 402138 220746 402374
rect 220982 402138 221066 402374
rect 221302 402138 221334 402374
rect 220714 402054 221334 402138
rect 220714 401818 220746 402054
rect 220982 401818 221066 402054
rect 221302 401818 221334 402054
rect 220714 366374 221334 401818
rect 220714 366138 220746 366374
rect 220982 366138 221066 366374
rect 221302 366138 221334 366374
rect 220714 366054 221334 366138
rect 220714 365818 220746 366054
rect 220982 365818 221066 366054
rect 221302 365818 221334 366054
rect 220714 330374 221334 365818
rect 220714 330138 220746 330374
rect 220982 330138 221066 330374
rect 221302 330138 221334 330374
rect 220714 330054 221334 330138
rect 220714 329818 220746 330054
rect 220982 329818 221066 330054
rect 221302 329818 221334 330054
rect 220714 294374 221334 329818
rect 220714 294138 220746 294374
rect 220982 294138 221066 294374
rect 221302 294138 221334 294374
rect 220714 294054 221334 294138
rect 220714 293818 220746 294054
rect 220982 293818 221066 294054
rect 221302 293818 221334 294054
rect 220714 258374 221334 293818
rect 220714 258138 220746 258374
rect 220982 258138 221066 258374
rect 221302 258138 221334 258374
rect 220714 258054 221334 258138
rect 220714 257818 220746 258054
rect 220982 257818 221066 258054
rect 221302 257818 221334 258054
rect 220714 222374 221334 257818
rect 220714 222138 220746 222374
rect 220982 222138 221066 222374
rect 221302 222138 221334 222374
rect 220714 222054 221334 222138
rect 220714 221818 220746 222054
rect 220982 221818 221066 222054
rect 221302 221818 221334 222054
rect 220714 186374 221334 221818
rect 220714 186138 220746 186374
rect 220982 186138 221066 186374
rect 221302 186138 221334 186374
rect 220714 186054 221334 186138
rect 220714 185818 220746 186054
rect 220982 185818 221066 186054
rect 221302 185818 221334 186054
rect 220714 150374 221334 185818
rect 220714 150138 220746 150374
rect 220982 150138 221066 150374
rect 221302 150138 221334 150374
rect 220714 150054 221334 150138
rect 220714 149818 220746 150054
rect 220982 149818 221066 150054
rect 221302 149818 221334 150054
rect 220714 114374 221334 149818
rect 220714 114138 220746 114374
rect 220982 114138 221066 114374
rect 221302 114138 221334 114374
rect 220714 114054 221334 114138
rect 220714 113818 220746 114054
rect 220982 113818 221066 114054
rect 221302 113818 221334 114054
rect 220714 78374 221334 113818
rect 220714 78138 220746 78374
rect 220982 78138 221066 78374
rect 221302 78138 221334 78374
rect 220714 78054 221334 78138
rect 220714 77818 220746 78054
rect 220982 77818 221066 78054
rect 221302 77818 221334 78054
rect 220714 42374 221334 77818
rect 220714 42138 220746 42374
rect 220982 42138 221066 42374
rect 221302 42138 221334 42374
rect 220714 42054 221334 42138
rect 220714 41818 220746 42054
rect 220982 41818 221066 42054
rect 221302 41818 221334 42054
rect 220714 6374 221334 41818
rect 220714 6138 220746 6374
rect 220982 6138 221066 6374
rect 221302 6138 221334 6374
rect 220714 6054 221334 6138
rect 220714 5818 220746 6054
rect 220982 5818 221066 6054
rect 221302 5818 221334 6054
rect 220714 -3226 221334 5818
rect 220714 -3462 220746 -3226
rect 220982 -3462 221066 -3226
rect 221302 -3462 221334 -3226
rect 220714 -3546 221334 -3462
rect 220714 -3782 220746 -3546
rect 220982 -3782 221066 -3546
rect 221302 -3782 221334 -3546
rect 220714 -7654 221334 -3782
rect 221954 708678 222574 711590
rect 221954 708442 221986 708678
rect 222222 708442 222306 708678
rect 222542 708442 222574 708678
rect 221954 708358 222574 708442
rect 221954 708122 221986 708358
rect 222222 708122 222306 708358
rect 222542 708122 222574 708358
rect 221954 691614 222574 708122
rect 221954 691378 221986 691614
rect 222222 691378 222306 691614
rect 222542 691378 222574 691614
rect 221954 691294 222574 691378
rect 221954 691058 221986 691294
rect 222222 691058 222306 691294
rect 222542 691058 222574 691294
rect 221954 655614 222574 691058
rect 221954 655378 221986 655614
rect 222222 655378 222306 655614
rect 222542 655378 222574 655614
rect 221954 655294 222574 655378
rect 221954 655058 221986 655294
rect 222222 655058 222306 655294
rect 222542 655058 222574 655294
rect 221954 619614 222574 655058
rect 221954 619378 221986 619614
rect 222222 619378 222306 619614
rect 222542 619378 222574 619614
rect 221954 619294 222574 619378
rect 221954 619058 221986 619294
rect 222222 619058 222306 619294
rect 222542 619058 222574 619294
rect 221954 583614 222574 619058
rect 221954 583378 221986 583614
rect 222222 583378 222306 583614
rect 222542 583378 222574 583614
rect 221954 583294 222574 583378
rect 221954 583058 221986 583294
rect 222222 583058 222306 583294
rect 222542 583058 222574 583294
rect 221954 547614 222574 583058
rect 221954 547378 221986 547614
rect 222222 547378 222306 547614
rect 222542 547378 222574 547614
rect 221954 547294 222574 547378
rect 221954 547058 221986 547294
rect 222222 547058 222306 547294
rect 222542 547058 222574 547294
rect 221954 511614 222574 547058
rect 221954 511378 221986 511614
rect 222222 511378 222306 511614
rect 222542 511378 222574 511614
rect 221954 511294 222574 511378
rect 221954 511058 221986 511294
rect 222222 511058 222306 511294
rect 222542 511058 222574 511294
rect 221954 475614 222574 511058
rect 221954 475378 221986 475614
rect 222222 475378 222306 475614
rect 222542 475378 222574 475614
rect 221954 475294 222574 475378
rect 221954 475058 221986 475294
rect 222222 475058 222306 475294
rect 222542 475058 222574 475294
rect 221954 439614 222574 475058
rect 221954 439378 221986 439614
rect 222222 439378 222306 439614
rect 222542 439378 222574 439614
rect 221954 439294 222574 439378
rect 221954 439058 221986 439294
rect 222222 439058 222306 439294
rect 222542 439058 222574 439294
rect 221954 403614 222574 439058
rect 221954 403378 221986 403614
rect 222222 403378 222306 403614
rect 222542 403378 222574 403614
rect 221954 403294 222574 403378
rect 221954 403058 221986 403294
rect 222222 403058 222306 403294
rect 222542 403058 222574 403294
rect 221954 367614 222574 403058
rect 221954 367378 221986 367614
rect 222222 367378 222306 367614
rect 222542 367378 222574 367614
rect 221954 367294 222574 367378
rect 221954 367058 221986 367294
rect 222222 367058 222306 367294
rect 222542 367058 222574 367294
rect 221954 331614 222574 367058
rect 221954 331378 221986 331614
rect 222222 331378 222306 331614
rect 222542 331378 222574 331614
rect 221954 331294 222574 331378
rect 221954 331058 221986 331294
rect 222222 331058 222306 331294
rect 222542 331058 222574 331294
rect 221954 295614 222574 331058
rect 221954 295378 221986 295614
rect 222222 295378 222306 295614
rect 222542 295378 222574 295614
rect 221954 295294 222574 295378
rect 221954 295058 221986 295294
rect 222222 295058 222306 295294
rect 222542 295058 222574 295294
rect 221954 259614 222574 295058
rect 221954 259378 221986 259614
rect 222222 259378 222306 259614
rect 222542 259378 222574 259614
rect 221954 259294 222574 259378
rect 221954 259058 221986 259294
rect 222222 259058 222306 259294
rect 222542 259058 222574 259294
rect 221954 223614 222574 259058
rect 221954 223378 221986 223614
rect 222222 223378 222306 223614
rect 222542 223378 222574 223614
rect 221954 223294 222574 223378
rect 221954 223058 221986 223294
rect 222222 223058 222306 223294
rect 222542 223058 222574 223294
rect 221954 187614 222574 223058
rect 221954 187378 221986 187614
rect 222222 187378 222306 187614
rect 222542 187378 222574 187614
rect 221954 187294 222574 187378
rect 221954 187058 221986 187294
rect 222222 187058 222306 187294
rect 222542 187058 222574 187294
rect 221954 151614 222574 187058
rect 221954 151378 221986 151614
rect 222222 151378 222306 151614
rect 222542 151378 222574 151614
rect 221954 151294 222574 151378
rect 221954 151058 221986 151294
rect 222222 151058 222306 151294
rect 222542 151058 222574 151294
rect 221954 115614 222574 151058
rect 221954 115378 221986 115614
rect 222222 115378 222306 115614
rect 222542 115378 222574 115614
rect 221954 115294 222574 115378
rect 221954 115058 221986 115294
rect 222222 115058 222306 115294
rect 222542 115058 222574 115294
rect 221954 79614 222574 115058
rect 221954 79378 221986 79614
rect 222222 79378 222306 79614
rect 222542 79378 222574 79614
rect 221954 79294 222574 79378
rect 221954 79058 221986 79294
rect 222222 79058 222306 79294
rect 222542 79058 222574 79294
rect 221954 43614 222574 79058
rect 221954 43378 221986 43614
rect 222222 43378 222306 43614
rect 222542 43378 222574 43614
rect 221954 43294 222574 43378
rect 221954 43058 221986 43294
rect 222222 43058 222306 43294
rect 222542 43058 222574 43294
rect 221954 7614 222574 43058
rect 221954 7378 221986 7614
rect 222222 7378 222306 7614
rect 222542 7378 222574 7614
rect 221954 7294 222574 7378
rect 221954 7058 221986 7294
rect 222222 7058 222306 7294
rect 222542 7058 222574 7294
rect 221954 -4186 222574 7058
rect 221954 -4422 221986 -4186
rect 222222 -4422 222306 -4186
rect 222542 -4422 222574 -4186
rect 221954 -4506 222574 -4422
rect 221954 -4742 221986 -4506
rect 222222 -4742 222306 -4506
rect 222542 -4742 222574 -4506
rect 221954 -7654 222574 -4742
rect 223194 709638 223814 711590
rect 223194 709402 223226 709638
rect 223462 709402 223546 709638
rect 223782 709402 223814 709638
rect 223194 709318 223814 709402
rect 223194 709082 223226 709318
rect 223462 709082 223546 709318
rect 223782 709082 223814 709318
rect 223194 692854 223814 709082
rect 223194 692618 223226 692854
rect 223462 692618 223546 692854
rect 223782 692618 223814 692854
rect 223194 692534 223814 692618
rect 223194 692298 223226 692534
rect 223462 692298 223546 692534
rect 223782 692298 223814 692534
rect 223194 656854 223814 692298
rect 223194 656618 223226 656854
rect 223462 656618 223546 656854
rect 223782 656618 223814 656854
rect 223194 656534 223814 656618
rect 223194 656298 223226 656534
rect 223462 656298 223546 656534
rect 223782 656298 223814 656534
rect 223194 620854 223814 656298
rect 223194 620618 223226 620854
rect 223462 620618 223546 620854
rect 223782 620618 223814 620854
rect 223194 620534 223814 620618
rect 223194 620298 223226 620534
rect 223462 620298 223546 620534
rect 223782 620298 223814 620534
rect 223194 584854 223814 620298
rect 223194 584618 223226 584854
rect 223462 584618 223546 584854
rect 223782 584618 223814 584854
rect 223194 584534 223814 584618
rect 223194 584298 223226 584534
rect 223462 584298 223546 584534
rect 223782 584298 223814 584534
rect 223194 548854 223814 584298
rect 223194 548618 223226 548854
rect 223462 548618 223546 548854
rect 223782 548618 223814 548854
rect 223194 548534 223814 548618
rect 223194 548298 223226 548534
rect 223462 548298 223546 548534
rect 223782 548298 223814 548534
rect 223194 512854 223814 548298
rect 223194 512618 223226 512854
rect 223462 512618 223546 512854
rect 223782 512618 223814 512854
rect 223194 512534 223814 512618
rect 223194 512298 223226 512534
rect 223462 512298 223546 512534
rect 223782 512298 223814 512534
rect 223194 476854 223814 512298
rect 223194 476618 223226 476854
rect 223462 476618 223546 476854
rect 223782 476618 223814 476854
rect 223194 476534 223814 476618
rect 223194 476298 223226 476534
rect 223462 476298 223546 476534
rect 223782 476298 223814 476534
rect 223194 440854 223814 476298
rect 223194 440618 223226 440854
rect 223462 440618 223546 440854
rect 223782 440618 223814 440854
rect 223194 440534 223814 440618
rect 223194 440298 223226 440534
rect 223462 440298 223546 440534
rect 223782 440298 223814 440534
rect 223194 404854 223814 440298
rect 223194 404618 223226 404854
rect 223462 404618 223546 404854
rect 223782 404618 223814 404854
rect 223194 404534 223814 404618
rect 223194 404298 223226 404534
rect 223462 404298 223546 404534
rect 223782 404298 223814 404534
rect 223194 368854 223814 404298
rect 223194 368618 223226 368854
rect 223462 368618 223546 368854
rect 223782 368618 223814 368854
rect 223194 368534 223814 368618
rect 223194 368298 223226 368534
rect 223462 368298 223546 368534
rect 223782 368298 223814 368534
rect 223194 332854 223814 368298
rect 223194 332618 223226 332854
rect 223462 332618 223546 332854
rect 223782 332618 223814 332854
rect 223194 332534 223814 332618
rect 223194 332298 223226 332534
rect 223462 332298 223546 332534
rect 223782 332298 223814 332534
rect 223194 296854 223814 332298
rect 223194 296618 223226 296854
rect 223462 296618 223546 296854
rect 223782 296618 223814 296854
rect 223194 296534 223814 296618
rect 223194 296298 223226 296534
rect 223462 296298 223546 296534
rect 223782 296298 223814 296534
rect 223194 260854 223814 296298
rect 223194 260618 223226 260854
rect 223462 260618 223546 260854
rect 223782 260618 223814 260854
rect 223194 260534 223814 260618
rect 223194 260298 223226 260534
rect 223462 260298 223546 260534
rect 223782 260298 223814 260534
rect 223194 224854 223814 260298
rect 223194 224618 223226 224854
rect 223462 224618 223546 224854
rect 223782 224618 223814 224854
rect 223194 224534 223814 224618
rect 223194 224298 223226 224534
rect 223462 224298 223546 224534
rect 223782 224298 223814 224534
rect 223194 188854 223814 224298
rect 223194 188618 223226 188854
rect 223462 188618 223546 188854
rect 223782 188618 223814 188854
rect 223194 188534 223814 188618
rect 223194 188298 223226 188534
rect 223462 188298 223546 188534
rect 223782 188298 223814 188534
rect 223194 152854 223814 188298
rect 223194 152618 223226 152854
rect 223462 152618 223546 152854
rect 223782 152618 223814 152854
rect 223194 152534 223814 152618
rect 223194 152298 223226 152534
rect 223462 152298 223546 152534
rect 223782 152298 223814 152534
rect 223194 116854 223814 152298
rect 223194 116618 223226 116854
rect 223462 116618 223546 116854
rect 223782 116618 223814 116854
rect 223194 116534 223814 116618
rect 223194 116298 223226 116534
rect 223462 116298 223546 116534
rect 223782 116298 223814 116534
rect 223194 80854 223814 116298
rect 223194 80618 223226 80854
rect 223462 80618 223546 80854
rect 223782 80618 223814 80854
rect 223194 80534 223814 80618
rect 223194 80298 223226 80534
rect 223462 80298 223546 80534
rect 223782 80298 223814 80534
rect 223194 44854 223814 80298
rect 223194 44618 223226 44854
rect 223462 44618 223546 44854
rect 223782 44618 223814 44854
rect 223194 44534 223814 44618
rect 223194 44298 223226 44534
rect 223462 44298 223546 44534
rect 223782 44298 223814 44534
rect 223194 8854 223814 44298
rect 223194 8618 223226 8854
rect 223462 8618 223546 8854
rect 223782 8618 223814 8854
rect 223194 8534 223814 8618
rect 223194 8298 223226 8534
rect 223462 8298 223546 8534
rect 223782 8298 223814 8534
rect 223194 -5146 223814 8298
rect 223194 -5382 223226 -5146
rect 223462 -5382 223546 -5146
rect 223782 -5382 223814 -5146
rect 223194 -5466 223814 -5382
rect 223194 -5702 223226 -5466
rect 223462 -5702 223546 -5466
rect 223782 -5702 223814 -5466
rect 223194 -7654 223814 -5702
rect 224434 710598 225054 711590
rect 224434 710362 224466 710598
rect 224702 710362 224786 710598
rect 225022 710362 225054 710598
rect 224434 710278 225054 710362
rect 224434 710042 224466 710278
rect 224702 710042 224786 710278
rect 225022 710042 225054 710278
rect 224434 694094 225054 710042
rect 224434 693858 224466 694094
rect 224702 693858 224786 694094
rect 225022 693858 225054 694094
rect 224434 693774 225054 693858
rect 224434 693538 224466 693774
rect 224702 693538 224786 693774
rect 225022 693538 225054 693774
rect 224434 658094 225054 693538
rect 224434 657858 224466 658094
rect 224702 657858 224786 658094
rect 225022 657858 225054 658094
rect 224434 657774 225054 657858
rect 224434 657538 224466 657774
rect 224702 657538 224786 657774
rect 225022 657538 225054 657774
rect 224434 622094 225054 657538
rect 224434 621858 224466 622094
rect 224702 621858 224786 622094
rect 225022 621858 225054 622094
rect 224434 621774 225054 621858
rect 224434 621538 224466 621774
rect 224702 621538 224786 621774
rect 225022 621538 225054 621774
rect 224434 586094 225054 621538
rect 224434 585858 224466 586094
rect 224702 585858 224786 586094
rect 225022 585858 225054 586094
rect 224434 585774 225054 585858
rect 224434 585538 224466 585774
rect 224702 585538 224786 585774
rect 225022 585538 225054 585774
rect 224434 550094 225054 585538
rect 224434 549858 224466 550094
rect 224702 549858 224786 550094
rect 225022 549858 225054 550094
rect 224434 549774 225054 549858
rect 224434 549538 224466 549774
rect 224702 549538 224786 549774
rect 225022 549538 225054 549774
rect 224434 514094 225054 549538
rect 224434 513858 224466 514094
rect 224702 513858 224786 514094
rect 225022 513858 225054 514094
rect 224434 513774 225054 513858
rect 224434 513538 224466 513774
rect 224702 513538 224786 513774
rect 225022 513538 225054 513774
rect 224434 478094 225054 513538
rect 224434 477858 224466 478094
rect 224702 477858 224786 478094
rect 225022 477858 225054 478094
rect 224434 477774 225054 477858
rect 224434 477538 224466 477774
rect 224702 477538 224786 477774
rect 225022 477538 225054 477774
rect 224434 442094 225054 477538
rect 224434 441858 224466 442094
rect 224702 441858 224786 442094
rect 225022 441858 225054 442094
rect 224434 441774 225054 441858
rect 224434 441538 224466 441774
rect 224702 441538 224786 441774
rect 225022 441538 225054 441774
rect 224434 406094 225054 441538
rect 224434 405858 224466 406094
rect 224702 405858 224786 406094
rect 225022 405858 225054 406094
rect 224434 405774 225054 405858
rect 224434 405538 224466 405774
rect 224702 405538 224786 405774
rect 225022 405538 225054 405774
rect 224434 370094 225054 405538
rect 224434 369858 224466 370094
rect 224702 369858 224786 370094
rect 225022 369858 225054 370094
rect 224434 369774 225054 369858
rect 224434 369538 224466 369774
rect 224702 369538 224786 369774
rect 225022 369538 225054 369774
rect 224434 334094 225054 369538
rect 224434 333858 224466 334094
rect 224702 333858 224786 334094
rect 225022 333858 225054 334094
rect 224434 333774 225054 333858
rect 224434 333538 224466 333774
rect 224702 333538 224786 333774
rect 225022 333538 225054 333774
rect 224434 298094 225054 333538
rect 224434 297858 224466 298094
rect 224702 297858 224786 298094
rect 225022 297858 225054 298094
rect 224434 297774 225054 297858
rect 224434 297538 224466 297774
rect 224702 297538 224786 297774
rect 225022 297538 225054 297774
rect 224434 262094 225054 297538
rect 224434 261858 224466 262094
rect 224702 261858 224786 262094
rect 225022 261858 225054 262094
rect 224434 261774 225054 261858
rect 224434 261538 224466 261774
rect 224702 261538 224786 261774
rect 225022 261538 225054 261774
rect 224434 226094 225054 261538
rect 224434 225858 224466 226094
rect 224702 225858 224786 226094
rect 225022 225858 225054 226094
rect 224434 225774 225054 225858
rect 224434 225538 224466 225774
rect 224702 225538 224786 225774
rect 225022 225538 225054 225774
rect 224434 190094 225054 225538
rect 224434 189858 224466 190094
rect 224702 189858 224786 190094
rect 225022 189858 225054 190094
rect 224434 189774 225054 189858
rect 224434 189538 224466 189774
rect 224702 189538 224786 189774
rect 225022 189538 225054 189774
rect 224434 154094 225054 189538
rect 224434 153858 224466 154094
rect 224702 153858 224786 154094
rect 225022 153858 225054 154094
rect 224434 153774 225054 153858
rect 224434 153538 224466 153774
rect 224702 153538 224786 153774
rect 225022 153538 225054 153774
rect 224434 118094 225054 153538
rect 224434 117858 224466 118094
rect 224702 117858 224786 118094
rect 225022 117858 225054 118094
rect 224434 117774 225054 117858
rect 224434 117538 224466 117774
rect 224702 117538 224786 117774
rect 225022 117538 225054 117774
rect 224434 82094 225054 117538
rect 224434 81858 224466 82094
rect 224702 81858 224786 82094
rect 225022 81858 225054 82094
rect 224434 81774 225054 81858
rect 224434 81538 224466 81774
rect 224702 81538 224786 81774
rect 225022 81538 225054 81774
rect 224434 46094 225054 81538
rect 224434 45858 224466 46094
rect 224702 45858 224786 46094
rect 225022 45858 225054 46094
rect 224434 45774 225054 45858
rect 224434 45538 224466 45774
rect 224702 45538 224786 45774
rect 225022 45538 225054 45774
rect 224434 10094 225054 45538
rect 224434 9858 224466 10094
rect 224702 9858 224786 10094
rect 225022 9858 225054 10094
rect 224434 9774 225054 9858
rect 224434 9538 224466 9774
rect 224702 9538 224786 9774
rect 225022 9538 225054 9774
rect 224434 -6106 225054 9538
rect 224434 -6342 224466 -6106
rect 224702 -6342 224786 -6106
rect 225022 -6342 225054 -6106
rect 224434 -6426 225054 -6342
rect 224434 -6662 224466 -6426
rect 224702 -6662 224786 -6426
rect 225022 -6662 225054 -6426
rect 224434 -7654 225054 -6662
rect 225674 711558 226294 711590
rect 225674 711322 225706 711558
rect 225942 711322 226026 711558
rect 226262 711322 226294 711558
rect 225674 711238 226294 711322
rect 225674 711002 225706 711238
rect 225942 711002 226026 711238
rect 226262 711002 226294 711238
rect 225674 695334 226294 711002
rect 225674 695098 225706 695334
rect 225942 695098 226026 695334
rect 226262 695098 226294 695334
rect 225674 695014 226294 695098
rect 225674 694778 225706 695014
rect 225942 694778 226026 695014
rect 226262 694778 226294 695014
rect 225674 659334 226294 694778
rect 225674 659098 225706 659334
rect 225942 659098 226026 659334
rect 226262 659098 226294 659334
rect 225674 659014 226294 659098
rect 225674 658778 225706 659014
rect 225942 658778 226026 659014
rect 226262 658778 226294 659014
rect 225674 623334 226294 658778
rect 225674 623098 225706 623334
rect 225942 623098 226026 623334
rect 226262 623098 226294 623334
rect 225674 623014 226294 623098
rect 225674 622778 225706 623014
rect 225942 622778 226026 623014
rect 226262 622778 226294 623014
rect 225674 587334 226294 622778
rect 225674 587098 225706 587334
rect 225942 587098 226026 587334
rect 226262 587098 226294 587334
rect 225674 587014 226294 587098
rect 225674 586778 225706 587014
rect 225942 586778 226026 587014
rect 226262 586778 226294 587014
rect 225674 551334 226294 586778
rect 225674 551098 225706 551334
rect 225942 551098 226026 551334
rect 226262 551098 226294 551334
rect 225674 551014 226294 551098
rect 225674 550778 225706 551014
rect 225942 550778 226026 551014
rect 226262 550778 226294 551014
rect 225674 515334 226294 550778
rect 225674 515098 225706 515334
rect 225942 515098 226026 515334
rect 226262 515098 226294 515334
rect 225674 515014 226294 515098
rect 225674 514778 225706 515014
rect 225942 514778 226026 515014
rect 226262 514778 226294 515014
rect 225674 479334 226294 514778
rect 225674 479098 225706 479334
rect 225942 479098 226026 479334
rect 226262 479098 226294 479334
rect 225674 479014 226294 479098
rect 225674 478778 225706 479014
rect 225942 478778 226026 479014
rect 226262 478778 226294 479014
rect 225674 443334 226294 478778
rect 225674 443098 225706 443334
rect 225942 443098 226026 443334
rect 226262 443098 226294 443334
rect 225674 443014 226294 443098
rect 225674 442778 225706 443014
rect 225942 442778 226026 443014
rect 226262 442778 226294 443014
rect 225674 407334 226294 442778
rect 225674 407098 225706 407334
rect 225942 407098 226026 407334
rect 226262 407098 226294 407334
rect 225674 407014 226294 407098
rect 225674 406778 225706 407014
rect 225942 406778 226026 407014
rect 226262 406778 226294 407014
rect 225674 371334 226294 406778
rect 225674 371098 225706 371334
rect 225942 371098 226026 371334
rect 226262 371098 226294 371334
rect 225674 371014 226294 371098
rect 225674 370778 225706 371014
rect 225942 370778 226026 371014
rect 226262 370778 226294 371014
rect 225674 335334 226294 370778
rect 225674 335098 225706 335334
rect 225942 335098 226026 335334
rect 226262 335098 226294 335334
rect 225674 335014 226294 335098
rect 225674 334778 225706 335014
rect 225942 334778 226026 335014
rect 226262 334778 226294 335014
rect 225674 299334 226294 334778
rect 225674 299098 225706 299334
rect 225942 299098 226026 299334
rect 226262 299098 226294 299334
rect 225674 299014 226294 299098
rect 225674 298778 225706 299014
rect 225942 298778 226026 299014
rect 226262 298778 226294 299014
rect 225674 263334 226294 298778
rect 225674 263098 225706 263334
rect 225942 263098 226026 263334
rect 226262 263098 226294 263334
rect 225674 263014 226294 263098
rect 225674 262778 225706 263014
rect 225942 262778 226026 263014
rect 226262 262778 226294 263014
rect 225674 227334 226294 262778
rect 225674 227098 225706 227334
rect 225942 227098 226026 227334
rect 226262 227098 226294 227334
rect 225674 227014 226294 227098
rect 225674 226778 225706 227014
rect 225942 226778 226026 227014
rect 226262 226778 226294 227014
rect 225674 191334 226294 226778
rect 225674 191098 225706 191334
rect 225942 191098 226026 191334
rect 226262 191098 226294 191334
rect 225674 191014 226294 191098
rect 225674 190778 225706 191014
rect 225942 190778 226026 191014
rect 226262 190778 226294 191014
rect 225674 155334 226294 190778
rect 225674 155098 225706 155334
rect 225942 155098 226026 155334
rect 226262 155098 226294 155334
rect 225674 155014 226294 155098
rect 225674 154778 225706 155014
rect 225942 154778 226026 155014
rect 226262 154778 226294 155014
rect 225674 119334 226294 154778
rect 225674 119098 225706 119334
rect 225942 119098 226026 119334
rect 226262 119098 226294 119334
rect 225674 119014 226294 119098
rect 225674 118778 225706 119014
rect 225942 118778 226026 119014
rect 226262 118778 226294 119014
rect 225674 83334 226294 118778
rect 225674 83098 225706 83334
rect 225942 83098 226026 83334
rect 226262 83098 226294 83334
rect 225674 83014 226294 83098
rect 225674 82778 225706 83014
rect 225942 82778 226026 83014
rect 226262 82778 226294 83014
rect 225674 47334 226294 82778
rect 225674 47098 225706 47334
rect 225942 47098 226026 47334
rect 226262 47098 226294 47334
rect 225674 47014 226294 47098
rect 225674 46778 225706 47014
rect 225942 46778 226026 47014
rect 226262 46778 226294 47014
rect 225674 11334 226294 46778
rect 225674 11098 225706 11334
rect 225942 11098 226026 11334
rect 226262 11098 226294 11334
rect 225674 11014 226294 11098
rect 225674 10778 225706 11014
rect 225942 10778 226026 11014
rect 226262 10778 226294 11014
rect 225674 -7066 226294 10778
rect 225674 -7302 225706 -7066
rect 225942 -7302 226026 -7066
rect 226262 -7302 226294 -7066
rect 225674 -7386 226294 -7302
rect 225674 -7622 225706 -7386
rect 225942 -7622 226026 -7386
rect 226262 -7622 226294 -7386
rect 225674 -7654 226294 -7622
rect 252994 704838 253614 711590
rect 252994 704602 253026 704838
rect 253262 704602 253346 704838
rect 253582 704602 253614 704838
rect 252994 704518 253614 704602
rect 252994 704282 253026 704518
rect 253262 704282 253346 704518
rect 253582 704282 253614 704518
rect 252994 686654 253614 704282
rect 252994 686418 253026 686654
rect 253262 686418 253346 686654
rect 253582 686418 253614 686654
rect 252994 686334 253614 686418
rect 252994 686098 253026 686334
rect 253262 686098 253346 686334
rect 253582 686098 253614 686334
rect 252994 650654 253614 686098
rect 252994 650418 253026 650654
rect 253262 650418 253346 650654
rect 253582 650418 253614 650654
rect 252994 650334 253614 650418
rect 252994 650098 253026 650334
rect 253262 650098 253346 650334
rect 253582 650098 253614 650334
rect 252994 614654 253614 650098
rect 252994 614418 253026 614654
rect 253262 614418 253346 614654
rect 253582 614418 253614 614654
rect 252994 614334 253614 614418
rect 252994 614098 253026 614334
rect 253262 614098 253346 614334
rect 253582 614098 253614 614334
rect 252994 578654 253614 614098
rect 252994 578418 253026 578654
rect 253262 578418 253346 578654
rect 253582 578418 253614 578654
rect 252994 578334 253614 578418
rect 252994 578098 253026 578334
rect 253262 578098 253346 578334
rect 253582 578098 253614 578334
rect 252994 542654 253614 578098
rect 252994 542418 253026 542654
rect 253262 542418 253346 542654
rect 253582 542418 253614 542654
rect 252994 542334 253614 542418
rect 252994 542098 253026 542334
rect 253262 542098 253346 542334
rect 253582 542098 253614 542334
rect 252994 506654 253614 542098
rect 252994 506418 253026 506654
rect 253262 506418 253346 506654
rect 253582 506418 253614 506654
rect 252994 506334 253614 506418
rect 252994 506098 253026 506334
rect 253262 506098 253346 506334
rect 253582 506098 253614 506334
rect 252994 470654 253614 506098
rect 252994 470418 253026 470654
rect 253262 470418 253346 470654
rect 253582 470418 253614 470654
rect 252994 470334 253614 470418
rect 252994 470098 253026 470334
rect 253262 470098 253346 470334
rect 253582 470098 253614 470334
rect 252994 434654 253614 470098
rect 252994 434418 253026 434654
rect 253262 434418 253346 434654
rect 253582 434418 253614 434654
rect 252994 434334 253614 434418
rect 252994 434098 253026 434334
rect 253262 434098 253346 434334
rect 253582 434098 253614 434334
rect 252994 398654 253614 434098
rect 252994 398418 253026 398654
rect 253262 398418 253346 398654
rect 253582 398418 253614 398654
rect 252994 398334 253614 398418
rect 252994 398098 253026 398334
rect 253262 398098 253346 398334
rect 253582 398098 253614 398334
rect 252994 362654 253614 398098
rect 252994 362418 253026 362654
rect 253262 362418 253346 362654
rect 253582 362418 253614 362654
rect 252994 362334 253614 362418
rect 252994 362098 253026 362334
rect 253262 362098 253346 362334
rect 253582 362098 253614 362334
rect 252994 326654 253614 362098
rect 252994 326418 253026 326654
rect 253262 326418 253346 326654
rect 253582 326418 253614 326654
rect 252994 326334 253614 326418
rect 252994 326098 253026 326334
rect 253262 326098 253346 326334
rect 253582 326098 253614 326334
rect 252994 290654 253614 326098
rect 252994 290418 253026 290654
rect 253262 290418 253346 290654
rect 253582 290418 253614 290654
rect 252994 290334 253614 290418
rect 252994 290098 253026 290334
rect 253262 290098 253346 290334
rect 253582 290098 253614 290334
rect 252994 254654 253614 290098
rect 252994 254418 253026 254654
rect 253262 254418 253346 254654
rect 253582 254418 253614 254654
rect 252994 254334 253614 254418
rect 252994 254098 253026 254334
rect 253262 254098 253346 254334
rect 253582 254098 253614 254334
rect 252994 218654 253614 254098
rect 252994 218418 253026 218654
rect 253262 218418 253346 218654
rect 253582 218418 253614 218654
rect 252994 218334 253614 218418
rect 252994 218098 253026 218334
rect 253262 218098 253346 218334
rect 253582 218098 253614 218334
rect 252994 182654 253614 218098
rect 252994 182418 253026 182654
rect 253262 182418 253346 182654
rect 253582 182418 253614 182654
rect 252994 182334 253614 182418
rect 252994 182098 253026 182334
rect 253262 182098 253346 182334
rect 253582 182098 253614 182334
rect 252994 146654 253614 182098
rect 252994 146418 253026 146654
rect 253262 146418 253346 146654
rect 253582 146418 253614 146654
rect 252994 146334 253614 146418
rect 252994 146098 253026 146334
rect 253262 146098 253346 146334
rect 253582 146098 253614 146334
rect 252994 110654 253614 146098
rect 252994 110418 253026 110654
rect 253262 110418 253346 110654
rect 253582 110418 253614 110654
rect 252994 110334 253614 110418
rect 252994 110098 253026 110334
rect 253262 110098 253346 110334
rect 253582 110098 253614 110334
rect 252994 74654 253614 110098
rect 252994 74418 253026 74654
rect 253262 74418 253346 74654
rect 253582 74418 253614 74654
rect 252994 74334 253614 74418
rect 252994 74098 253026 74334
rect 253262 74098 253346 74334
rect 253582 74098 253614 74334
rect 252994 38654 253614 74098
rect 252994 38418 253026 38654
rect 253262 38418 253346 38654
rect 253582 38418 253614 38654
rect 252994 38334 253614 38418
rect 252994 38098 253026 38334
rect 253262 38098 253346 38334
rect 253582 38098 253614 38334
rect 252994 2654 253614 38098
rect 252994 2418 253026 2654
rect 253262 2418 253346 2654
rect 253582 2418 253614 2654
rect 252994 2334 253614 2418
rect 252994 2098 253026 2334
rect 253262 2098 253346 2334
rect 253582 2098 253614 2334
rect 252994 -346 253614 2098
rect 252994 -582 253026 -346
rect 253262 -582 253346 -346
rect 253582 -582 253614 -346
rect 252994 -666 253614 -582
rect 252994 -902 253026 -666
rect 253262 -902 253346 -666
rect 253582 -902 253614 -666
rect 252994 -7654 253614 -902
rect 254234 705798 254854 711590
rect 254234 705562 254266 705798
rect 254502 705562 254586 705798
rect 254822 705562 254854 705798
rect 254234 705478 254854 705562
rect 254234 705242 254266 705478
rect 254502 705242 254586 705478
rect 254822 705242 254854 705478
rect 254234 687894 254854 705242
rect 254234 687658 254266 687894
rect 254502 687658 254586 687894
rect 254822 687658 254854 687894
rect 254234 687574 254854 687658
rect 254234 687338 254266 687574
rect 254502 687338 254586 687574
rect 254822 687338 254854 687574
rect 254234 651894 254854 687338
rect 254234 651658 254266 651894
rect 254502 651658 254586 651894
rect 254822 651658 254854 651894
rect 254234 651574 254854 651658
rect 254234 651338 254266 651574
rect 254502 651338 254586 651574
rect 254822 651338 254854 651574
rect 254234 615894 254854 651338
rect 254234 615658 254266 615894
rect 254502 615658 254586 615894
rect 254822 615658 254854 615894
rect 254234 615574 254854 615658
rect 254234 615338 254266 615574
rect 254502 615338 254586 615574
rect 254822 615338 254854 615574
rect 254234 579894 254854 615338
rect 254234 579658 254266 579894
rect 254502 579658 254586 579894
rect 254822 579658 254854 579894
rect 254234 579574 254854 579658
rect 254234 579338 254266 579574
rect 254502 579338 254586 579574
rect 254822 579338 254854 579574
rect 254234 543894 254854 579338
rect 254234 543658 254266 543894
rect 254502 543658 254586 543894
rect 254822 543658 254854 543894
rect 254234 543574 254854 543658
rect 254234 543338 254266 543574
rect 254502 543338 254586 543574
rect 254822 543338 254854 543574
rect 254234 507894 254854 543338
rect 254234 507658 254266 507894
rect 254502 507658 254586 507894
rect 254822 507658 254854 507894
rect 254234 507574 254854 507658
rect 254234 507338 254266 507574
rect 254502 507338 254586 507574
rect 254822 507338 254854 507574
rect 254234 471894 254854 507338
rect 254234 471658 254266 471894
rect 254502 471658 254586 471894
rect 254822 471658 254854 471894
rect 254234 471574 254854 471658
rect 254234 471338 254266 471574
rect 254502 471338 254586 471574
rect 254822 471338 254854 471574
rect 254234 435894 254854 471338
rect 254234 435658 254266 435894
rect 254502 435658 254586 435894
rect 254822 435658 254854 435894
rect 254234 435574 254854 435658
rect 254234 435338 254266 435574
rect 254502 435338 254586 435574
rect 254822 435338 254854 435574
rect 254234 399894 254854 435338
rect 254234 399658 254266 399894
rect 254502 399658 254586 399894
rect 254822 399658 254854 399894
rect 254234 399574 254854 399658
rect 254234 399338 254266 399574
rect 254502 399338 254586 399574
rect 254822 399338 254854 399574
rect 254234 363894 254854 399338
rect 254234 363658 254266 363894
rect 254502 363658 254586 363894
rect 254822 363658 254854 363894
rect 254234 363574 254854 363658
rect 254234 363338 254266 363574
rect 254502 363338 254586 363574
rect 254822 363338 254854 363574
rect 254234 327894 254854 363338
rect 254234 327658 254266 327894
rect 254502 327658 254586 327894
rect 254822 327658 254854 327894
rect 254234 327574 254854 327658
rect 254234 327338 254266 327574
rect 254502 327338 254586 327574
rect 254822 327338 254854 327574
rect 254234 291894 254854 327338
rect 254234 291658 254266 291894
rect 254502 291658 254586 291894
rect 254822 291658 254854 291894
rect 254234 291574 254854 291658
rect 254234 291338 254266 291574
rect 254502 291338 254586 291574
rect 254822 291338 254854 291574
rect 254234 255894 254854 291338
rect 254234 255658 254266 255894
rect 254502 255658 254586 255894
rect 254822 255658 254854 255894
rect 254234 255574 254854 255658
rect 254234 255338 254266 255574
rect 254502 255338 254586 255574
rect 254822 255338 254854 255574
rect 254234 219894 254854 255338
rect 254234 219658 254266 219894
rect 254502 219658 254586 219894
rect 254822 219658 254854 219894
rect 254234 219574 254854 219658
rect 254234 219338 254266 219574
rect 254502 219338 254586 219574
rect 254822 219338 254854 219574
rect 254234 183894 254854 219338
rect 254234 183658 254266 183894
rect 254502 183658 254586 183894
rect 254822 183658 254854 183894
rect 254234 183574 254854 183658
rect 254234 183338 254266 183574
rect 254502 183338 254586 183574
rect 254822 183338 254854 183574
rect 254234 147894 254854 183338
rect 254234 147658 254266 147894
rect 254502 147658 254586 147894
rect 254822 147658 254854 147894
rect 254234 147574 254854 147658
rect 254234 147338 254266 147574
rect 254502 147338 254586 147574
rect 254822 147338 254854 147574
rect 254234 111894 254854 147338
rect 254234 111658 254266 111894
rect 254502 111658 254586 111894
rect 254822 111658 254854 111894
rect 254234 111574 254854 111658
rect 254234 111338 254266 111574
rect 254502 111338 254586 111574
rect 254822 111338 254854 111574
rect 254234 75894 254854 111338
rect 254234 75658 254266 75894
rect 254502 75658 254586 75894
rect 254822 75658 254854 75894
rect 254234 75574 254854 75658
rect 254234 75338 254266 75574
rect 254502 75338 254586 75574
rect 254822 75338 254854 75574
rect 254234 39894 254854 75338
rect 254234 39658 254266 39894
rect 254502 39658 254586 39894
rect 254822 39658 254854 39894
rect 254234 39574 254854 39658
rect 254234 39338 254266 39574
rect 254502 39338 254586 39574
rect 254822 39338 254854 39574
rect 254234 3894 254854 39338
rect 254234 3658 254266 3894
rect 254502 3658 254586 3894
rect 254822 3658 254854 3894
rect 254234 3574 254854 3658
rect 254234 3338 254266 3574
rect 254502 3338 254586 3574
rect 254822 3338 254854 3574
rect 254234 -1306 254854 3338
rect 254234 -1542 254266 -1306
rect 254502 -1542 254586 -1306
rect 254822 -1542 254854 -1306
rect 254234 -1626 254854 -1542
rect 254234 -1862 254266 -1626
rect 254502 -1862 254586 -1626
rect 254822 -1862 254854 -1626
rect 254234 -7654 254854 -1862
rect 255474 706758 256094 711590
rect 255474 706522 255506 706758
rect 255742 706522 255826 706758
rect 256062 706522 256094 706758
rect 255474 706438 256094 706522
rect 255474 706202 255506 706438
rect 255742 706202 255826 706438
rect 256062 706202 256094 706438
rect 255474 689134 256094 706202
rect 255474 688898 255506 689134
rect 255742 688898 255826 689134
rect 256062 688898 256094 689134
rect 255474 688814 256094 688898
rect 255474 688578 255506 688814
rect 255742 688578 255826 688814
rect 256062 688578 256094 688814
rect 255474 653134 256094 688578
rect 255474 652898 255506 653134
rect 255742 652898 255826 653134
rect 256062 652898 256094 653134
rect 255474 652814 256094 652898
rect 255474 652578 255506 652814
rect 255742 652578 255826 652814
rect 256062 652578 256094 652814
rect 255474 617134 256094 652578
rect 255474 616898 255506 617134
rect 255742 616898 255826 617134
rect 256062 616898 256094 617134
rect 255474 616814 256094 616898
rect 255474 616578 255506 616814
rect 255742 616578 255826 616814
rect 256062 616578 256094 616814
rect 255474 581134 256094 616578
rect 255474 580898 255506 581134
rect 255742 580898 255826 581134
rect 256062 580898 256094 581134
rect 255474 580814 256094 580898
rect 255474 580578 255506 580814
rect 255742 580578 255826 580814
rect 256062 580578 256094 580814
rect 255474 545134 256094 580578
rect 255474 544898 255506 545134
rect 255742 544898 255826 545134
rect 256062 544898 256094 545134
rect 255474 544814 256094 544898
rect 255474 544578 255506 544814
rect 255742 544578 255826 544814
rect 256062 544578 256094 544814
rect 255474 509134 256094 544578
rect 255474 508898 255506 509134
rect 255742 508898 255826 509134
rect 256062 508898 256094 509134
rect 255474 508814 256094 508898
rect 255474 508578 255506 508814
rect 255742 508578 255826 508814
rect 256062 508578 256094 508814
rect 255474 473134 256094 508578
rect 255474 472898 255506 473134
rect 255742 472898 255826 473134
rect 256062 472898 256094 473134
rect 255474 472814 256094 472898
rect 255474 472578 255506 472814
rect 255742 472578 255826 472814
rect 256062 472578 256094 472814
rect 255474 437134 256094 472578
rect 255474 436898 255506 437134
rect 255742 436898 255826 437134
rect 256062 436898 256094 437134
rect 255474 436814 256094 436898
rect 255474 436578 255506 436814
rect 255742 436578 255826 436814
rect 256062 436578 256094 436814
rect 255474 401134 256094 436578
rect 255474 400898 255506 401134
rect 255742 400898 255826 401134
rect 256062 400898 256094 401134
rect 255474 400814 256094 400898
rect 255474 400578 255506 400814
rect 255742 400578 255826 400814
rect 256062 400578 256094 400814
rect 255474 365134 256094 400578
rect 255474 364898 255506 365134
rect 255742 364898 255826 365134
rect 256062 364898 256094 365134
rect 255474 364814 256094 364898
rect 255474 364578 255506 364814
rect 255742 364578 255826 364814
rect 256062 364578 256094 364814
rect 255474 329134 256094 364578
rect 255474 328898 255506 329134
rect 255742 328898 255826 329134
rect 256062 328898 256094 329134
rect 255474 328814 256094 328898
rect 255474 328578 255506 328814
rect 255742 328578 255826 328814
rect 256062 328578 256094 328814
rect 255474 293134 256094 328578
rect 255474 292898 255506 293134
rect 255742 292898 255826 293134
rect 256062 292898 256094 293134
rect 255474 292814 256094 292898
rect 255474 292578 255506 292814
rect 255742 292578 255826 292814
rect 256062 292578 256094 292814
rect 255474 257134 256094 292578
rect 255474 256898 255506 257134
rect 255742 256898 255826 257134
rect 256062 256898 256094 257134
rect 255474 256814 256094 256898
rect 255474 256578 255506 256814
rect 255742 256578 255826 256814
rect 256062 256578 256094 256814
rect 255474 221134 256094 256578
rect 255474 220898 255506 221134
rect 255742 220898 255826 221134
rect 256062 220898 256094 221134
rect 255474 220814 256094 220898
rect 255474 220578 255506 220814
rect 255742 220578 255826 220814
rect 256062 220578 256094 220814
rect 255474 185134 256094 220578
rect 255474 184898 255506 185134
rect 255742 184898 255826 185134
rect 256062 184898 256094 185134
rect 255474 184814 256094 184898
rect 255474 184578 255506 184814
rect 255742 184578 255826 184814
rect 256062 184578 256094 184814
rect 255474 149134 256094 184578
rect 255474 148898 255506 149134
rect 255742 148898 255826 149134
rect 256062 148898 256094 149134
rect 255474 148814 256094 148898
rect 255474 148578 255506 148814
rect 255742 148578 255826 148814
rect 256062 148578 256094 148814
rect 255474 113134 256094 148578
rect 255474 112898 255506 113134
rect 255742 112898 255826 113134
rect 256062 112898 256094 113134
rect 255474 112814 256094 112898
rect 255474 112578 255506 112814
rect 255742 112578 255826 112814
rect 256062 112578 256094 112814
rect 255474 77134 256094 112578
rect 255474 76898 255506 77134
rect 255742 76898 255826 77134
rect 256062 76898 256094 77134
rect 255474 76814 256094 76898
rect 255474 76578 255506 76814
rect 255742 76578 255826 76814
rect 256062 76578 256094 76814
rect 255474 41134 256094 76578
rect 255474 40898 255506 41134
rect 255742 40898 255826 41134
rect 256062 40898 256094 41134
rect 255474 40814 256094 40898
rect 255474 40578 255506 40814
rect 255742 40578 255826 40814
rect 256062 40578 256094 40814
rect 255474 5134 256094 40578
rect 255474 4898 255506 5134
rect 255742 4898 255826 5134
rect 256062 4898 256094 5134
rect 255474 4814 256094 4898
rect 255474 4578 255506 4814
rect 255742 4578 255826 4814
rect 256062 4578 256094 4814
rect 255474 -2266 256094 4578
rect 255474 -2502 255506 -2266
rect 255742 -2502 255826 -2266
rect 256062 -2502 256094 -2266
rect 255474 -2586 256094 -2502
rect 255474 -2822 255506 -2586
rect 255742 -2822 255826 -2586
rect 256062 -2822 256094 -2586
rect 255474 -7654 256094 -2822
rect 256714 707718 257334 711590
rect 256714 707482 256746 707718
rect 256982 707482 257066 707718
rect 257302 707482 257334 707718
rect 256714 707398 257334 707482
rect 256714 707162 256746 707398
rect 256982 707162 257066 707398
rect 257302 707162 257334 707398
rect 256714 690374 257334 707162
rect 256714 690138 256746 690374
rect 256982 690138 257066 690374
rect 257302 690138 257334 690374
rect 256714 690054 257334 690138
rect 256714 689818 256746 690054
rect 256982 689818 257066 690054
rect 257302 689818 257334 690054
rect 256714 654374 257334 689818
rect 256714 654138 256746 654374
rect 256982 654138 257066 654374
rect 257302 654138 257334 654374
rect 256714 654054 257334 654138
rect 256714 653818 256746 654054
rect 256982 653818 257066 654054
rect 257302 653818 257334 654054
rect 256714 618374 257334 653818
rect 256714 618138 256746 618374
rect 256982 618138 257066 618374
rect 257302 618138 257334 618374
rect 256714 618054 257334 618138
rect 256714 617818 256746 618054
rect 256982 617818 257066 618054
rect 257302 617818 257334 618054
rect 256714 582374 257334 617818
rect 256714 582138 256746 582374
rect 256982 582138 257066 582374
rect 257302 582138 257334 582374
rect 256714 582054 257334 582138
rect 256714 581818 256746 582054
rect 256982 581818 257066 582054
rect 257302 581818 257334 582054
rect 256714 546374 257334 581818
rect 256714 546138 256746 546374
rect 256982 546138 257066 546374
rect 257302 546138 257334 546374
rect 256714 546054 257334 546138
rect 256714 545818 256746 546054
rect 256982 545818 257066 546054
rect 257302 545818 257334 546054
rect 256714 510374 257334 545818
rect 256714 510138 256746 510374
rect 256982 510138 257066 510374
rect 257302 510138 257334 510374
rect 256714 510054 257334 510138
rect 256714 509818 256746 510054
rect 256982 509818 257066 510054
rect 257302 509818 257334 510054
rect 256714 474374 257334 509818
rect 256714 474138 256746 474374
rect 256982 474138 257066 474374
rect 257302 474138 257334 474374
rect 256714 474054 257334 474138
rect 256714 473818 256746 474054
rect 256982 473818 257066 474054
rect 257302 473818 257334 474054
rect 256714 438374 257334 473818
rect 256714 438138 256746 438374
rect 256982 438138 257066 438374
rect 257302 438138 257334 438374
rect 256714 438054 257334 438138
rect 256714 437818 256746 438054
rect 256982 437818 257066 438054
rect 257302 437818 257334 438054
rect 256714 402374 257334 437818
rect 256714 402138 256746 402374
rect 256982 402138 257066 402374
rect 257302 402138 257334 402374
rect 256714 402054 257334 402138
rect 256714 401818 256746 402054
rect 256982 401818 257066 402054
rect 257302 401818 257334 402054
rect 256714 366374 257334 401818
rect 256714 366138 256746 366374
rect 256982 366138 257066 366374
rect 257302 366138 257334 366374
rect 256714 366054 257334 366138
rect 256714 365818 256746 366054
rect 256982 365818 257066 366054
rect 257302 365818 257334 366054
rect 256714 330374 257334 365818
rect 256714 330138 256746 330374
rect 256982 330138 257066 330374
rect 257302 330138 257334 330374
rect 256714 330054 257334 330138
rect 256714 329818 256746 330054
rect 256982 329818 257066 330054
rect 257302 329818 257334 330054
rect 256714 294374 257334 329818
rect 256714 294138 256746 294374
rect 256982 294138 257066 294374
rect 257302 294138 257334 294374
rect 256714 294054 257334 294138
rect 256714 293818 256746 294054
rect 256982 293818 257066 294054
rect 257302 293818 257334 294054
rect 256714 258374 257334 293818
rect 256714 258138 256746 258374
rect 256982 258138 257066 258374
rect 257302 258138 257334 258374
rect 256714 258054 257334 258138
rect 256714 257818 256746 258054
rect 256982 257818 257066 258054
rect 257302 257818 257334 258054
rect 256714 222374 257334 257818
rect 256714 222138 256746 222374
rect 256982 222138 257066 222374
rect 257302 222138 257334 222374
rect 256714 222054 257334 222138
rect 256714 221818 256746 222054
rect 256982 221818 257066 222054
rect 257302 221818 257334 222054
rect 256714 186374 257334 221818
rect 256714 186138 256746 186374
rect 256982 186138 257066 186374
rect 257302 186138 257334 186374
rect 256714 186054 257334 186138
rect 256714 185818 256746 186054
rect 256982 185818 257066 186054
rect 257302 185818 257334 186054
rect 256714 150374 257334 185818
rect 256714 150138 256746 150374
rect 256982 150138 257066 150374
rect 257302 150138 257334 150374
rect 256714 150054 257334 150138
rect 256714 149818 256746 150054
rect 256982 149818 257066 150054
rect 257302 149818 257334 150054
rect 256714 114374 257334 149818
rect 256714 114138 256746 114374
rect 256982 114138 257066 114374
rect 257302 114138 257334 114374
rect 256714 114054 257334 114138
rect 256714 113818 256746 114054
rect 256982 113818 257066 114054
rect 257302 113818 257334 114054
rect 256714 78374 257334 113818
rect 256714 78138 256746 78374
rect 256982 78138 257066 78374
rect 257302 78138 257334 78374
rect 256714 78054 257334 78138
rect 256714 77818 256746 78054
rect 256982 77818 257066 78054
rect 257302 77818 257334 78054
rect 256714 42374 257334 77818
rect 256714 42138 256746 42374
rect 256982 42138 257066 42374
rect 257302 42138 257334 42374
rect 256714 42054 257334 42138
rect 256714 41818 256746 42054
rect 256982 41818 257066 42054
rect 257302 41818 257334 42054
rect 256714 6374 257334 41818
rect 256714 6138 256746 6374
rect 256982 6138 257066 6374
rect 257302 6138 257334 6374
rect 256714 6054 257334 6138
rect 256714 5818 256746 6054
rect 256982 5818 257066 6054
rect 257302 5818 257334 6054
rect 256714 -3226 257334 5818
rect 256714 -3462 256746 -3226
rect 256982 -3462 257066 -3226
rect 257302 -3462 257334 -3226
rect 256714 -3546 257334 -3462
rect 256714 -3782 256746 -3546
rect 256982 -3782 257066 -3546
rect 257302 -3782 257334 -3546
rect 256714 -7654 257334 -3782
rect 257954 708678 258574 711590
rect 257954 708442 257986 708678
rect 258222 708442 258306 708678
rect 258542 708442 258574 708678
rect 257954 708358 258574 708442
rect 257954 708122 257986 708358
rect 258222 708122 258306 708358
rect 258542 708122 258574 708358
rect 257954 691614 258574 708122
rect 257954 691378 257986 691614
rect 258222 691378 258306 691614
rect 258542 691378 258574 691614
rect 257954 691294 258574 691378
rect 257954 691058 257986 691294
rect 258222 691058 258306 691294
rect 258542 691058 258574 691294
rect 257954 655614 258574 691058
rect 257954 655378 257986 655614
rect 258222 655378 258306 655614
rect 258542 655378 258574 655614
rect 257954 655294 258574 655378
rect 257954 655058 257986 655294
rect 258222 655058 258306 655294
rect 258542 655058 258574 655294
rect 257954 619614 258574 655058
rect 257954 619378 257986 619614
rect 258222 619378 258306 619614
rect 258542 619378 258574 619614
rect 257954 619294 258574 619378
rect 257954 619058 257986 619294
rect 258222 619058 258306 619294
rect 258542 619058 258574 619294
rect 257954 583614 258574 619058
rect 257954 583378 257986 583614
rect 258222 583378 258306 583614
rect 258542 583378 258574 583614
rect 257954 583294 258574 583378
rect 257954 583058 257986 583294
rect 258222 583058 258306 583294
rect 258542 583058 258574 583294
rect 257954 547614 258574 583058
rect 257954 547378 257986 547614
rect 258222 547378 258306 547614
rect 258542 547378 258574 547614
rect 257954 547294 258574 547378
rect 257954 547058 257986 547294
rect 258222 547058 258306 547294
rect 258542 547058 258574 547294
rect 257954 511614 258574 547058
rect 257954 511378 257986 511614
rect 258222 511378 258306 511614
rect 258542 511378 258574 511614
rect 257954 511294 258574 511378
rect 257954 511058 257986 511294
rect 258222 511058 258306 511294
rect 258542 511058 258574 511294
rect 257954 475614 258574 511058
rect 257954 475378 257986 475614
rect 258222 475378 258306 475614
rect 258542 475378 258574 475614
rect 257954 475294 258574 475378
rect 257954 475058 257986 475294
rect 258222 475058 258306 475294
rect 258542 475058 258574 475294
rect 257954 439614 258574 475058
rect 257954 439378 257986 439614
rect 258222 439378 258306 439614
rect 258542 439378 258574 439614
rect 257954 439294 258574 439378
rect 257954 439058 257986 439294
rect 258222 439058 258306 439294
rect 258542 439058 258574 439294
rect 257954 403614 258574 439058
rect 257954 403378 257986 403614
rect 258222 403378 258306 403614
rect 258542 403378 258574 403614
rect 257954 403294 258574 403378
rect 257954 403058 257986 403294
rect 258222 403058 258306 403294
rect 258542 403058 258574 403294
rect 257954 367614 258574 403058
rect 257954 367378 257986 367614
rect 258222 367378 258306 367614
rect 258542 367378 258574 367614
rect 257954 367294 258574 367378
rect 257954 367058 257986 367294
rect 258222 367058 258306 367294
rect 258542 367058 258574 367294
rect 257954 331614 258574 367058
rect 257954 331378 257986 331614
rect 258222 331378 258306 331614
rect 258542 331378 258574 331614
rect 257954 331294 258574 331378
rect 257954 331058 257986 331294
rect 258222 331058 258306 331294
rect 258542 331058 258574 331294
rect 257954 295614 258574 331058
rect 257954 295378 257986 295614
rect 258222 295378 258306 295614
rect 258542 295378 258574 295614
rect 257954 295294 258574 295378
rect 257954 295058 257986 295294
rect 258222 295058 258306 295294
rect 258542 295058 258574 295294
rect 257954 259614 258574 295058
rect 257954 259378 257986 259614
rect 258222 259378 258306 259614
rect 258542 259378 258574 259614
rect 257954 259294 258574 259378
rect 257954 259058 257986 259294
rect 258222 259058 258306 259294
rect 258542 259058 258574 259294
rect 257954 223614 258574 259058
rect 257954 223378 257986 223614
rect 258222 223378 258306 223614
rect 258542 223378 258574 223614
rect 257954 223294 258574 223378
rect 257954 223058 257986 223294
rect 258222 223058 258306 223294
rect 258542 223058 258574 223294
rect 257954 187614 258574 223058
rect 257954 187378 257986 187614
rect 258222 187378 258306 187614
rect 258542 187378 258574 187614
rect 257954 187294 258574 187378
rect 257954 187058 257986 187294
rect 258222 187058 258306 187294
rect 258542 187058 258574 187294
rect 257954 151614 258574 187058
rect 257954 151378 257986 151614
rect 258222 151378 258306 151614
rect 258542 151378 258574 151614
rect 257954 151294 258574 151378
rect 257954 151058 257986 151294
rect 258222 151058 258306 151294
rect 258542 151058 258574 151294
rect 257954 115614 258574 151058
rect 257954 115378 257986 115614
rect 258222 115378 258306 115614
rect 258542 115378 258574 115614
rect 257954 115294 258574 115378
rect 257954 115058 257986 115294
rect 258222 115058 258306 115294
rect 258542 115058 258574 115294
rect 257954 79614 258574 115058
rect 257954 79378 257986 79614
rect 258222 79378 258306 79614
rect 258542 79378 258574 79614
rect 257954 79294 258574 79378
rect 257954 79058 257986 79294
rect 258222 79058 258306 79294
rect 258542 79058 258574 79294
rect 257954 43614 258574 79058
rect 257954 43378 257986 43614
rect 258222 43378 258306 43614
rect 258542 43378 258574 43614
rect 257954 43294 258574 43378
rect 257954 43058 257986 43294
rect 258222 43058 258306 43294
rect 258542 43058 258574 43294
rect 257954 7614 258574 43058
rect 257954 7378 257986 7614
rect 258222 7378 258306 7614
rect 258542 7378 258574 7614
rect 257954 7294 258574 7378
rect 257954 7058 257986 7294
rect 258222 7058 258306 7294
rect 258542 7058 258574 7294
rect 257954 -4186 258574 7058
rect 257954 -4422 257986 -4186
rect 258222 -4422 258306 -4186
rect 258542 -4422 258574 -4186
rect 257954 -4506 258574 -4422
rect 257954 -4742 257986 -4506
rect 258222 -4742 258306 -4506
rect 258542 -4742 258574 -4506
rect 257954 -7654 258574 -4742
rect 259194 709638 259814 711590
rect 259194 709402 259226 709638
rect 259462 709402 259546 709638
rect 259782 709402 259814 709638
rect 259194 709318 259814 709402
rect 259194 709082 259226 709318
rect 259462 709082 259546 709318
rect 259782 709082 259814 709318
rect 259194 692854 259814 709082
rect 259194 692618 259226 692854
rect 259462 692618 259546 692854
rect 259782 692618 259814 692854
rect 259194 692534 259814 692618
rect 259194 692298 259226 692534
rect 259462 692298 259546 692534
rect 259782 692298 259814 692534
rect 259194 656854 259814 692298
rect 259194 656618 259226 656854
rect 259462 656618 259546 656854
rect 259782 656618 259814 656854
rect 259194 656534 259814 656618
rect 259194 656298 259226 656534
rect 259462 656298 259546 656534
rect 259782 656298 259814 656534
rect 259194 620854 259814 656298
rect 259194 620618 259226 620854
rect 259462 620618 259546 620854
rect 259782 620618 259814 620854
rect 259194 620534 259814 620618
rect 259194 620298 259226 620534
rect 259462 620298 259546 620534
rect 259782 620298 259814 620534
rect 259194 584854 259814 620298
rect 259194 584618 259226 584854
rect 259462 584618 259546 584854
rect 259782 584618 259814 584854
rect 259194 584534 259814 584618
rect 259194 584298 259226 584534
rect 259462 584298 259546 584534
rect 259782 584298 259814 584534
rect 259194 548854 259814 584298
rect 259194 548618 259226 548854
rect 259462 548618 259546 548854
rect 259782 548618 259814 548854
rect 259194 548534 259814 548618
rect 259194 548298 259226 548534
rect 259462 548298 259546 548534
rect 259782 548298 259814 548534
rect 259194 512854 259814 548298
rect 259194 512618 259226 512854
rect 259462 512618 259546 512854
rect 259782 512618 259814 512854
rect 259194 512534 259814 512618
rect 259194 512298 259226 512534
rect 259462 512298 259546 512534
rect 259782 512298 259814 512534
rect 259194 476854 259814 512298
rect 259194 476618 259226 476854
rect 259462 476618 259546 476854
rect 259782 476618 259814 476854
rect 259194 476534 259814 476618
rect 259194 476298 259226 476534
rect 259462 476298 259546 476534
rect 259782 476298 259814 476534
rect 259194 440854 259814 476298
rect 259194 440618 259226 440854
rect 259462 440618 259546 440854
rect 259782 440618 259814 440854
rect 259194 440534 259814 440618
rect 259194 440298 259226 440534
rect 259462 440298 259546 440534
rect 259782 440298 259814 440534
rect 259194 404854 259814 440298
rect 259194 404618 259226 404854
rect 259462 404618 259546 404854
rect 259782 404618 259814 404854
rect 259194 404534 259814 404618
rect 259194 404298 259226 404534
rect 259462 404298 259546 404534
rect 259782 404298 259814 404534
rect 259194 368854 259814 404298
rect 259194 368618 259226 368854
rect 259462 368618 259546 368854
rect 259782 368618 259814 368854
rect 259194 368534 259814 368618
rect 259194 368298 259226 368534
rect 259462 368298 259546 368534
rect 259782 368298 259814 368534
rect 259194 332854 259814 368298
rect 259194 332618 259226 332854
rect 259462 332618 259546 332854
rect 259782 332618 259814 332854
rect 259194 332534 259814 332618
rect 259194 332298 259226 332534
rect 259462 332298 259546 332534
rect 259782 332298 259814 332534
rect 259194 296854 259814 332298
rect 259194 296618 259226 296854
rect 259462 296618 259546 296854
rect 259782 296618 259814 296854
rect 259194 296534 259814 296618
rect 259194 296298 259226 296534
rect 259462 296298 259546 296534
rect 259782 296298 259814 296534
rect 259194 260854 259814 296298
rect 259194 260618 259226 260854
rect 259462 260618 259546 260854
rect 259782 260618 259814 260854
rect 259194 260534 259814 260618
rect 259194 260298 259226 260534
rect 259462 260298 259546 260534
rect 259782 260298 259814 260534
rect 259194 224854 259814 260298
rect 259194 224618 259226 224854
rect 259462 224618 259546 224854
rect 259782 224618 259814 224854
rect 259194 224534 259814 224618
rect 259194 224298 259226 224534
rect 259462 224298 259546 224534
rect 259782 224298 259814 224534
rect 259194 188854 259814 224298
rect 259194 188618 259226 188854
rect 259462 188618 259546 188854
rect 259782 188618 259814 188854
rect 259194 188534 259814 188618
rect 259194 188298 259226 188534
rect 259462 188298 259546 188534
rect 259782 188298 259814 188534
rect 259194 152854 259814 188298
rect 259194 152618 259226 152854
rect 259462 152618 259546 152854
rect 259782 152618 259814 152854
rect 259194 152534 259814 152618
rect 259194 152298 259226 152534
rect 259462 152298 259546 152534
rect 259782 152298 259814 152534
rect 259194 116854 259814 152298
rect 259194 116618 259226 116854
rect 259462 116618 259546 116854
rect 259782 116618 259814 116854
rect 259194 116534 259814 116618
rect 259194 116298 259226 116534
rect 259462 116298 259546 116534
rect 259782 116298 259814 116534
rect 259194 80854 259814 116298
rect 259194 80618 259226 80854
rect 259462 80618 259546 80854
rect 259782 80618 259814 80854
rect 259194 80534 259814 80618
rect 259194 80298 259226 80534
rect 259462 80298 259546 80534
rect 259782 80298 259814 80534
rect 259194 44854 259814 80298
rect 259194 44618 259226 44854
rect 259462 44618 259546 44854
rect 259782 44618 259814 44854
rect 259194 44534 259814 44618
rect 259194 44298 259226 44534
rect 259462 44298 259546 44534
rect 259782 44298 259814 44534
rect 259194 8854 259814 44298
rect 259194 8618 259226 8854
rect 259462 8618 259546 8854
rect 259782 8618 259814 8854
rect 259194 8534 259814 8618
rect 259194 8298 259226 8534
rect 259462 8298 259546 8534
rect 259782 8298 259814 8534
rect 259194 -5146 259814 8298
rect 259194 -5382 259226 -5146
rect 259462 -5382 259546 -5146
rect 259782 -5382 259814 -5146
rect 259194 -5466 259814 -5382
rect 259194 -5702 259226 -5466
rect 259462 -5702 259546 -5466
rect 259782 -5702 259814 -5466
rect 259194 -7654 259814 -5702
rect 260434 710598 261054 711590
rect 260434 710362 260466 710598
rect 260702 710362 260786 710598
rect 261022 710362 261054 710598
rect 260434 710278 261054 710362
rect 260434 710042 260466 710278
rect 260702 710042 260786 710278
rect 261022 710042 261054 710278
rect 260434 694094 261054 710042
rect 260434 693858 260466 694094
rect 260702 693858 260786 694094
rect 261022 693858 261054 694094
rect 260434 693774 261054 693858
rect 260434 693538 260466 693774
rect 260702 693538 260786 693774
rect 261022 693538 261054 693774
rect 260434 658094 261054 693538
rect 260434 657858 260466 658094
rect 260702 657858 260786 658094
rect 261022 657858 261054 658094
rect 260434 657774 261054 657858
rect 260434 657538 260466 657774
rect 260702 657538 260786 657774
rect 261022 657538 261054 657774
rect 260434 622094 261054 657538
rect 260434 621858 260466 622094
rect 260702 621858 260786 622094
rect 261022 621858 261054 622094
rect 260434 621774 261054 621858
rect 260434 621538 260466 621774
rect 260702 621538 260786 621774
rect 261022 621538 261054 621774
rect 260434 586094 261054 621538
rect 260434 585858 260466 586094
rect 260702 585858 260786 586094
rect 261022 585858 261054 586094
rect 260434 585774 261054 585858
rect 260434 585538 260466 585774
rect 260702 585538 260786 585774
rect 261022 585538 261054 585774
rect 260434 550094 261054 585538
rect 260434 549858 260466 550094
rect 260702 549858 260786 550094
rect 261022 549858 261054 550094
rect 260434 549774 261054 549858
rect 260434 549538 260466 549774
rect 260702 549538 260786 549774
rect 261022 549538 261054 549774
rect 260434 514094 261054 549538
rect 260434 513858 260466 514094
rect 260702 513858 260786 514094
rect 261022 513858 261054 514094
rect 260434 513774 261054 513858
rect 260434 513538 260466 513774
rect 260702 513538 260786 513774
rect 261022 513538 261054 513774
rect 260434 478094 261054 513538
rect 260434 477858 260466 478094
rect 260702 477858 260786 478094
rect 261022 477858 261054 478094
rect 260434 477774 261054 477858
rect 260434 477538 260466 477774
rect 260702 477538 260786 477774
rect 261022 477538 261054 477774
rect 260434 442094 261054 477538
rect 260434 441858 260466 442094
rect 260702 441858 260786 442094
rect 261022 441858 261054 442094
rect 260434 441774 261054 441858
rect 260434 441538 260466 441774
rect 260702 441538 260786 441774
rect 261022 441538 261054 441774
rect 260434 406094 261054 441538
rect 260434 405858 260466 406094
rect 260702 405858 260786 406094
rect 261022 405858 261054 406094
rect 260434 405774 261054 405858
rect 260434 405538 260466 405774
rect 260702 405538 260786 405774
rect 261022 405538 261054 405774
rect 260434 370094 261054 405538
rect 260434 369858 260466 370094
rect 260702 369858 260786 370094
rect 261022 369858 261054 370094
rect 260434 369774 261054 369858
rect 260434 369538 260466 369774
rect 260702 369538 260786 369774
rect 261022 369538 261054 369774
rect 260434 334094 261054 369538
rect 260434 333858 260466 334094
rect 260702 333858 260786 334094
rect 261022 333858 261054 334094
rect 260434 333774 261054 333858
rect 260434 333538 260466 333774
rect 260702 333538 260786 333774
rect 261022 333538 261054 333774
rect 260434 298094 261054 333538
rect 260434 297858 260466 298094
rect 260702 297858 260786 298094
rect 261022 297858 261054 298094
rect 260434 297774 261054 297858
rect 260434 297538 260466 297774
rect 260702 297538 260786 297774
rect 261022 297538 261054 297774
rect 260434 262094 261054 297538
rect 260434 261858 260466 262094
rect 260702 261858 260786 262094
rect 261022 261858 261054 262094
rect 260434 261774 261054 261858
rect 260434 261538 260466 261774
rect 260702 261538 260786 261774
rect 261022 261538 261054 261774
rect 260434 226094 261054 261538
rect 260434 225858 260466 226094
rect 260702 225858 260786 226094
rect 261022 225858 261054 226094
rect 260434 225774 261054 225858
rect 260434 225538 260466 225774
rect 260702 225538 260786 225774
rect 261022 225538 261054 225774
rect 260434 190094 261054 225538
rect 260434 189858 260466 190094
rect 260702 189858 260786 190094
rect 261022 189858 261054 190094
rect 260434 189774 261054 189858
rect 260434 189538 260466 189774
rect 260702 189538 260786 189774
rect 261022 189538 261054 189774
rect 260434 154094 261054 189538
rect 260434 153858 260466 154094
rect 260702 153858 260786 154094
rect 261022 153858 261054 154094
rect 260434 153774 261054 153858
rect 260434 153538 260466 153774
rect 260702 153538 260786 153774
rect 261022 153538 261054 153774
rect 260434 118094 261054 153538
rect 260434 117858 260466 118094
rect 260702 117858 260786 118094
rect 261022 117858 261054 118094
rect 260434 117774 261054 117858
rect 260434 117538 260466 117774
rect 260702 117538 260786 117774
rect 261022 117538 261054 117774
rect 260434 82094 261054 117538
rect 260434 81858 260466 82094
rect 260702 81858 260786 82094
rect 261022 81858 261054 82094
rect 260434 81774 261054 81858
rect 260434 81538 260466 81774
rect 260702 81538 260786 81774
rect 261022 81538 261054 81774
rect 260434 46094 261054 81538
rect 260434 45858 260466 46094
rect 260702 45858 260786 46094
rect 261022 45858 261054 46094
rect 260434 45774 261054 45858
rect 260434 45538 260466 45774
rect 260702 45538 260786 45774
rect 261022 45538 261054 45774
rect 260434 10094 261054 45538
rect 260434 9858 260466 10094
rect 260702 9858 260786 10094
rect 261022 9858 261054 10094
rect 260434 9774 261054 9858
rect 260434 9538 260466 9774
rect 260702 9538 260786 9774
rect 261022 9538 261054 9774
rect 260434 -6106 261054 9538
rect 260434 -6342 260466 -6106
rect 260702 -6342 260786 -6106
rect 261022 -6342 261054 -6106
rect 260434 -6426 261054 -6342
rect 260434 -6662 260466 -6426
rect 260702 -6662 260786 -6426
rect 261022 -6662 261054 -6426
rect 260434 -7654 261054 -6662
rect 261674 711558 262294 711590
rect 261674 711322 261706 711558
rect 261942 711322 262026 711558
rect 262262 711322 262294 711558
rect 261674 711238 262294 711322
rect 261674 711002 261706 711238
rect 261942 711002 262026 711238
rect 262262 711002 262294 711238
rect 261674 695334 262294 711002
rect 261674 695098 261706 695334
rect 261942 695098 262026 695334
rect 262262 695098 262294 695334
rect 261674 695014 262294 695098
rect 261674 694778 261706 695014
rect 261942 694778 262026 695014
rect 262262 694778 262294 695014
rect 261674 659334 262294 694778
rect 261674 659098 261706 659334
rect 261942 659098 262026 659334
rect 262262 659098 262294 659334
rect 261674 659014 262294 659098
rect 261674 658778 261706 659014
rect 261942 658778 262026 659014
rect 262262 658778 262294 659014
rect 261674 623334 262294 658778
rect 261674 623098 261706 623334
rect 261942 623098 262026 623334
rect 262262 623098 262294 623334
rect 261674 623014 262294 623098
rect 261674 622778 261706 623014
rect 261942 622778 262026 623014
rect 262262 622778 262294 623014
rect 261674 587334 262294 622778
rect 261674 587098 261706 587334
rect 261942 587098 262026 587334
rect 262262 587098 262294 587334
rect 261674 587014 262294 587098
rect 261674 586778 261706 587014
rect 261942 586778 262026 587014
rect 262262 586778 262294 587014
rect 261674 551334 262294 586778
rect 261674 551098 261706 551334
rect 261942 551098 262026 551334
rect 262262 551098 262294 551334
rect 261674 551014 262294 551098
rect 261674 550778 261706 551014
rect 261942 550778 262026 551014
rect 262262 550778 262294 551014
rect 261674 515334 262294 550778
rect 261674 515098 261706 515334
rect 261942 515098 262026 515334
rect 262262 515098 262294 515334
rect 261674 515014 262294 515098
rect 261674 514778 261706 515014
rect 261942 514778 262026 515014
rect 262262 514778 262294 515014
rect 261674 479334 262294 514778
rect 261674 479098 261706 479334
rect 261942 479098 262026 479334
rect 262262 479098 262294 479334
rect 261674 479014 262294 479098
rect 261674 478778 261706 479014
rect 261942 478778 262026 479014
rect 262262 478778 262294 479014
rect 261674 443334 262294 478778
rect 261674 443098 261706 443334
rect 261942 443098 262026 443334
rect 262262 443098 262294 443334
rect 261674 443014 262294 443098
rect 261674 442778 261706 443014
rect 261942 442778 262026 443014
rect 262262 442778 262294 443014
rect 261674 407334 262294 442778
rect 261674 407098 261706 407334
rect 261942 407098 262026 407334
rect 262262 407098 262294 407334
rect 261674 407014 262294 407098
rect 261674 406778 261706 407014
rect 261942 406778 262026 407014
rect 262262 406778 262294 407014
rect 261674 371334 262294 406778
rect 261674 371098 261706 371334
rect 261942 371098 262026 371334
rect 262262 371098 262294 371334
rect 261674 371014 262294 371098
rect 261674 370778 261706 371014
rect 261942 370778 262026 371014
rect 262262 370778 262294 371014
rect 261674 335334 262294 370778
rect 261674 335098 261706 335334
rect 261942 335098 262026 335334
rect 262262 335098 262294 335334
rect 261674 335014 262294 335098
rect 261674 334778 261706 335014
rect 261942 334778 262026 335014
rect 262262 334778 262294 335014
rect 261674 299334 262294 334778
rect 261674 299098 261706 299334
rect 261942 299098 262026 299334
rect 262262 299098 262294 299334
rect 261674 299014 262294 299098
rect 261674 298778 261706 299014
rect 261942 298778 262026 299014
rect 262262 298778 262294 299014
rect 261674 263334 262294 298778
rect 261674 263098 261706 263334
rect 261942 263098 262026 263334
rect 262262 263098 262294 263334
rect 261674 263014 262294 263098
rect 261674 262778 261706 263014
rect 261942 262778 262026 263014
rect 262262 262778 262294 263014
rect 261674 227334 262294 262778
rect 261674 227098 261706 227334
rect 261942 227098 262026 227334
rect 262262 227098 262294 227334
rect 261674 227014 262294 227098
rect 261674 226778 261706 227014
rect 261942 226778 262026 227014
rect 262262 226778 262294 227014
rect 261674 191334 262294 226778
rect 261674 191098 261706 191334
rect 261942 191098 262026 191334
rect 262262 191098 262294 191334
rect 261674 191014 262294 191098
rect 261674 190778 261706 191014
rect 261942 190778 262026 191014
rect 262262 190778 262294 191014
rect 261674 155334 262294 190778
rect 261674 155098 261706 155334
rect 261942 155098 262026 155334
rect 262262 155098 262294 155334
rect 261674 155014 262294 155098
rect 261674 154778 261706 155014
rect 261942 154778 262026 155014
rect 262262 154778 262294 155014
rect 261674 119334 262294 154778
rect 261674 119098 261706 119334
rect 261942 119098 262026 119334
rect 262262 119098 262294 119334
rect 261674 119014 262294 119098
rect 261674 118778 261706 119014
rect 261942 118778 262026 119014
rect 262262 118778 262294 119014
rect 261674 83334 262294 118778
rect 261674 83098 261706 83334
rect 261942 83098 262026 83334
rect 262262 83098 262294 83334
rect 261674 83014 262294 83098
rect 261674 82778 261706 83014
rect 261942 82778 262026 83014
rect 262262 82778 262294 83014
rect 261674 47334 262294 82778
rect 261674 47098 261706 47334
rect 261942 47098 262026 47334
rect 262262 47098 262294 47334
rect 261674 47014 262294 47098
rect 261674 46778 261706 47014
rect 261942 46778 262026 47014
rect 262262 46778 262294 47014
rect 261674 11334 262294 46778
rect 261674 11098 261706 11334
rect 261942 11098 262026 11334
rect 262262 11098 262294 11334
rect 261674 11014 262294 11098
rect 261674 10778 261706 11014
rect 261942 10778 262026 11014
rect 262262 10778 262294 11014
rect 261674 -7066 262294 10778
rect 261674 -7302 261706 -7066
rect 261942 -7302 262026 -7066
rect 262262 -7302 262294 -7066
rect 261674 -7386 262294 -7302
rect 261674 -7622 261706 -7386
rect 261942 -7622 262026 -7386
rect 262262 -7622 262294 -7386
rect 261674 -7654 262294 -7622
rect 288994 704838 289614 711590
rect 288994 704602 289026 704838
rect 289262 704602 289346 704838
rect 289582 704602 289614 704838
rect 288994 704518 289614 704602
rect 288994 704282 289026 704518
rect 289262 704282 289346 704518
rect 289582 704282 289614 704518
rect 288994 686654 289614 704282
rect 288994 686418 289026 686654
rect 289262 686418 289346 686654
rect 289582 686418 289614 686654
rect 288994 686334 289614 686418
rect 288994 686098 289026 686334
rect 289262 686098 289346 686334
rect 289582 686098 289614 686334
rect 288994 650654 289614 686098
rect 288994 650418 289026 650654
rect 289262 650418 289346 650654
rect 289582 650418 289614 650654
rect 288994 650334 289614 650418
rect 288994 650098 289026 650334
rect 289262 650098 289346 650334
rect 289582 650098 289614 650334
rect 288994 614654 289614 650098
rect 288994 614418 289026 614654
rect 289262 614418 289346 614654
rect 289582 614418 289614 614654
rect 288994 614334 289614 614418
rect 288994 614098 289026 614334
rect 289262 614098 289346 614334
rect 289582 614098 289614 614334
rect 288994 578654 289614 614098
rect 288994 578418 289026 578654
rect 289262 578418 289346 578654
rect 289582 578418 289614 578654
rect 288994 578334 289614 578418
rect 288994 578098 289026 578334
rect 289262 578098 289346 578334
rect 289582 578098 289614 578334
rect 288994 542654 289614 578098
rect 288994 542418 289026 542654
rect 289262 542418 289346 542654
rect 289582 542418 289614 542654
rect 288994 542334 289614 542418
rect 288994 542098 289026 542334
rect 289262 542098 289346 542334
rect 289582 542098 289614 542334
rect 288994 506654 289614 542098
rect 288994 506418 289026 506654
rect 289262 506418 289346 506654
rect 289582 506418 289614 506654
rect 288994 506334 289614 506418
rect 288994 506098 289026 506334
rect 289262 506098 289346 506334
rect 289582 506098 289614 506334
rect 288994 470654 289614 506098
rect 288994 470418 289026 470654
rect 289262 470418 289346 470654
rect 289582 470418 289614 470654
rect 288994 470334 289614 470418
rect 288994 470098 289026 470334
rect 289262 470098 289346 470334
rect 289582 470098 289614 470334
rect 288994 434654 289614 470098
rect 288994 434418 289026 434654
rect 289262 434418 289346 434654
rect 289582 434418 289614 434654
rect 288994 434334 289614 434418
rect 288994 434098 289026 434334
rect 289262 434098 289346 434334
rect 289582 434098 289614 434334
rect 288994 398654 289614 434098
rect 288994 398418 289026 398654
rect 289262 398418 289346 398654
rect 289582 398418 289614 398654
rect 288994 398334 289614 398418
rect 288994 398098 289026 398334
rect 289262 398098 289346 398334
rect 289582 398098 289614 398334
rect 288994 362654 289614 398098
rect 288994 362418 289026 362654
rect 289262 362418 289346 362654
rect 289582 362418 289614 362654
rect 288994 362334 289614 362418
rect 288994 362098 289026 362334
rect 289262 362098 289346 362334
rect 289582 362098 289614 362334
rect 288994 326654 289614 362098
rect 288994 326418 289026 326654
rect 289262 326418 289346 326654
rect 289582 326418 289614 326654
rect 288994 326334 289614 326418
rect 288994 326098 289026 326334
rect 289262 326098 289346 326334
rect 289582 326098 289614 326334
rect 288994 290654 289614 326098
rect 288994 290418 289026 290654
rect 289262 290418 289346 290654
rect 289582 290418 289614 290654
rect 288994 290334 289614 290418
rect 288994 290098 289026 290334
rect 289262 290098 289346 290334
rect 289582 290098 289614 290334
rect 288994 254654 289614 290098
rect 288994 254418 289026 254654
rect 289262 254418 289346 254654
rect 289582 254418 289614 254654
rect 288994 254334 289614 254418
rect 288994 254098 289026 254334
rect 289262 254098 289346 254334
rect 289582 254098 289614 254334
rect 288994 218654 289614 254098
rect 288994 218418 289026 218654
rect 289262 218418 289346 218654
rect 289582 218418 289614 218654
rect 288994 218334 289614 218418
rect 288994 218098 289026 218334
rect 289262 218098 289346 218334
rect 289582 218098 289614 218334
rect 288994 182654 289614 218098
rect 288994 182418 289026 182654
rect 289262 182418 289346 182654
rect 289582 182418 289614 182654
rect 288994 182334 289614 182418
rect 288994 182098 289026 182334
rect 289262 182098 289346 182334
rect 289582 182098 289614 182334
rect 288994 146654 289614 182098
rect 288994 146418 289026 146654
rect 289262 146418 289346 146654
rect 289582 146418 289614 146654
rect 288994 146334 289614 146418
rect 288994 146098 289026 146334
rect 289262 146098 289346 146334
rect 289582 146098 289614 146334
rect 288994 110654 289614 146098
rect 288994 110418 289026 110654
rect 289262 110418 289346 110654
rect 289582 110418 289614 110654
rect 288994 110334 289614 110418
rect 288994 110098 289026 110334
rect 289262 110098 289346 110334
rect 289582 110098 289614 110334
rect 288994 74654 289614 110098
rect 288994 74418 289026 74654
rect 289262 74418 289346 74654
rect 289582 74418 289614 74654
rect 288994 74334 289614 74418
rect 288994 74098 289026 74334
rect 289262 74098 289346 74334
rect 289582 74098 289614 74334
rect 288994 38654 289614 74098
rect 288994 38418 289026 38654
rect 289262 38418 289346 38654
rect 289582 38418 289614 38654
rect 288994 38334 289614 38418
rect 288994 38098 289026 38334
rect 289262 38098 289346 38334
rect 289582 38098 289614 38334
rect 288994 2654 289614 38098
rect 288994 2418 289026 2654
rect 289262 2418 289346 2654
rect 289582 2418 289614 2654
rect 288994 2334 289614 2418
rect 288994 2098 289026 2334
rect 289262 2098 289346 2334
rect 289582 2098 289614 2334
rect 288994 -346 289614 2098
rect 288994 -582 289026 -346
rect 289262 -582 289346 -346
rect 289582 -582 289614 -346
rect 288994 -666 289614 -582
rect 288994 -902 289026 -666
rect 289262 -902 289346 -666
rect 289582 -902 289614 -666
rect 288994 -7654 289614 -902
rect 290234 705798 290854 711590
rect 290234 705562 290266 705798
rect 290502 705562 290586 705798
rect 290822 705562 290854 705798
rect 290234 705478 290854 705562
rect 290234 705242 290266 705478
rect 290502 705242 290586 705478
rect 290822 705242 290854 705478
rect 290234 687894 290854 705242
rect 290234 687658 290266 687894
rect 290502 687658 290586 687894
rect 290822 687658 290854 687894
rect 290234 687574 290854 687658
rect 290234 687338 290266 687574
rect 290502 687338 290586 687574
rect 290822 687338 290854 687574
rect 290234 651894 290854 687338
rect 290234 651658 290266 651894
rect 290502 651658 290586 651894
rect 290822 651658 290854 651894
rect 290234 651574 290854 651658
rect 290234 651338 290266 651574
rect 290502 651338 290586 651574
rect 290822 651338 290854 651574
rect 290234 615894 290854 651338
rect 290234 615658 290266 615894
rect 290502 615658 290586 615894
rect 290822 615658 290854 615894
rect 290234 615574 290854 615658
rect 290234 615338 290266 615574
rect 290502 615338 290586 615574
rect 290822 615338 290854 615574
rect 290234 579894 290854 615338
rect 290234 579658 290266 579894
rect 290502 579658 290586 579894
rect 290822 579658 290854 579894
rect 290234 579574 290854 579658
rect 290234 579338 290266 579574
rect 290502 579338 290586 579574
rect 290822 579338 290854 579574
rect 290234 543894 290854 579338
rect 290234 543658 290266 543894
rect 290502 543658 290586 543894
rect 290822 543658 290854 543894
rect 290234 543574 290854 543658
rect 290234 543338 290266 543574
rect 290502 543338 290586 543574
rect 290822 543338 290854 543574
rect 290234 507894 290854 543338
rect 290234 507658 290266 507894
rect 290502 507658 290586 507894
rect 290822 507658 290854 507894
rect 290234 507574 290854 507658
rect 290234 507338 290266 507574
rect 290502 507338 290586 507574
rect 290822 507338 290854 507574
rect 290234 471894 290854 507338
rect 290234 471658 290266 471894
rect 290502 471658 290586 471894
rect 290822 471658 290854 471894
rect 290234 471574 290854 471658
rect 290234 471338 290266 471574
rect 290502 471338 290586 471574
rect 290822 471338 290854 471574
rect 290234 435894 290854 471338
rect 290234 435658 290266 435894
rect 290502 435658 290586 435894
rect 290822 435658 290854 435894
rect 290234 435574 290854 435658
rect 290234 435338 290266 435574
rect 290502 435338 290586 435574
rect 290822 435338 290854 435574
rect 290234 399894 290854 435338
rect 290234 399658 290266 399894
rect 290502 399658 290586 399894
rect 290822 399658 290854 399894
rect 290234 399574 290854 399658
rect 290234 399338 290266 399574
rect 290502 399338 290586 399574
rect 290822 399338 290854 399574
rect 290234 363894 290854 399338
rect 290234 363658 290266 363894
rect 290502 363658 290586 363894
rect 290822 363658 290854 363894
rect 290234 363574 290854 363658
rect 290234 363338 290266 363574
rect 290502 363338 290586 363574
rect 290822 363338 290854 363574
rect 290234 327894 290854 363338
rect 290234 327658 290266 327894
rect 290502 327658 290586 327894
rect 290822 327658 290854 327894
rect 290234 327574 290854 327658
rect 290234 327338 290266 327574
rect 290502 327338 290586 327574
rect 290822 327338 290854 327574
rect 290234 291894 290854 327338
rect 290234 291658 290266 291894
rect 290502 291658 290586 291894
rect 290822 291658 290854 291894
rect 290234 291574 290854 291658
rect 290234 291338 290266 291574
rect 290502 291338 290586 291574
rect 290822 291338 290854 291574
rect 290234 255894 290854 291338
rect 290234 255658 290266 255894
rect 290502 255658 290586 255894
rect 290822 255658 290854 255894
rect 290234 255574 290854 255658
rect 290234 255338 290266 255574
rect 290502 255338 290586 255574
rect 290822 255338 290854 255574
rect 290234 219894 290854 255338
rect 290234 219658 290266 219894
rect 290502 219658 290586 219894
rect 290822 219658 290854 219894
rect 290234 219574 290854 219658
rect 290234 219338 290266 219574
rect 290502 219338 290586 219574
rect 290822 219338 290854 219574
rect 290234 183894 290854 219338
rect 290234 183658 290266 183894
rect 290502 183658 290586 183894
rect 290822 183658 290854 183894
rect 290234 183574 290854 183658
rect 290234 183338 290266 183574
rect 290502 183338 290586 183574
rect 290822 183338 290854 183574
rect 290234 147894 290854 183338
rect 290234 147658 290266 147894
rect 290502 147658 290586 147894
rect 290822 147658 290854 147894
rect 290234 147574 290854 147658
rect 290234 147338 290266 147574
rect 290502 147338 290586 147574
rect 290822 147338 290854 147574
rect 290234 111894 290854 147338
rect 290234 111658 290266 111894
rect 290502 111658 290586 111894
rect 290822 111658 290854 111894
rect 290234 111574 290854 111658
rect 290234 111338 290266 111574
rect 290502 111338 290586 111574
rect 290822 111338 290854 111574
rect 290234 75894 290854 111338
rect 290234 75658 290266 75894
rect 290502 75658 290586 75894
rect 290822 75658 290854 75894
rect 290234 75574 290854 75658
rect 290234 75338 290266 75574
rect 290502 75338 290586 75574
rect 290822 75338 290854 75574
rect 290234 39894 290854 75338
rect 290234 39658 290266 39894
rect 290502 39658 290586 39894
rect 290822 39658 290854 39894
rect 290234 39574 290854 39658
rect 290234 39338 290266 39574
rect 290502 39338 290586 39574
rect 290822 39338 290854 39574
rect 290234 3894 290854 39338
rect 290234 3658 290266 3894
rect 290502 3658 290586 3894
rect 290822 3658 290854 3894
rect 290234 3574 290854 3658
rect 290234 3338 290266 3574
rect 290502 3338 290586 3574
rect 290822 3338 290854 3574
rect 290234 -1306 290854 3338
rect 290234 -1542 290266 -1306
rect 290502 -1542 290586 -1306
rect 290822 -1542 290854 -1306
rect 290234 -1626 290854 -1542
rect 290234 -1862 290266 -1626
rect 290502 -1862 290586 -1626
rect 290822 -1862 290854 -1626
rect 290234 -7654 290854 -1862
rect 291474 706758 292094 711590
rect 291474 706522 291506 706758
rect 291742 706522 291826 706758
rect 292062 706522 292094 706758
rect 291474 706438 292094 706522
rect 291474 706202 291506 706438
rect 291742 706202 291826 706438
rect 292062 706202 292094 706438
rect 291474 689134 292094 706202
rect 291474 688898 291506 689134
rect 291742 688898 291826 689134
rect 292062 688898 292094 689134
rect 291474 688814 292094 688898
rect 291474 688578 291506 688814
rect 291742 688578 291826 688814
rect 292062 688578 292094 688814
rect 291474 653134 292094 688578
rect 291474 652898 291506 653134
rect 291742 652898 291826 653134
rect 292062 652898 292094 653134
rect 291474 652814 292094 652898
rect 291474 652578 291506 652814
rect 291742 652578 291826 652814
rect 292062 652578 292094 652814
rect 291474 617134 292094 652578
rect 291474 616898 291506 617134
rect 291742 616898 291826 617134
rect 292062 616898 292094 617134
rect 291474 616814 292094 616898
rect 291474 616578 291506 616814
rect 291742 616578 291826 616814
rect 292062 616578 292094 616814
rect 291474 581134 292094 616578
rect 291474 580898 291506 581134
rect 291742 580898 291826 581134
rect 292062 580898 292094 581134
rect 291474 580814 292094 580898
rect 291474 580578 291506 580814
rect 291742 580578 291826 580814
rect 292062 580578 292094 580814
rect 291474 545134 292094 580578
rect 291474 544898 291506 545134
rect 291742 544898 291826 545134
rect 292062 544898 292094 545134
rect 291474 544814 292094 544898
rect 291474 544578 291506 544814
rect 291742 544578 291826 544814
rect 292062 544578 292094 544814
rect 291474 509134 292094 544578
rect 291474 508898 291506 509134
rect 291742 508898 291826 509134
rect 292062 508898 292094 509134
rect 291474 508814 292094 508898
rect 291474 508578 291506 508814
rect 291742 508578 291826 508814
rect 292062 508578 292094 508814
rect 291474 473134 292094 508578
rect 291474 472898 291506 473134
rect 291742 472898 291826 473134
rect 292062 472898 292094 473134
rect 291474 472814 292094 472898
rect 291474 472578 291506 472814
rect 291742 472578 291826 472814
rect 292062 472578 292094 472814
rect 291474 437134 292094 472578
rect 291474 436898 291506 437134
rect 291742 436898 291826 437134
rect 292062 436898 292094 437134
rect 291474 436814 292094 436898
rect 291474 436578 291506 436814
rect 291742 436578 291826 436814
rect 292062 436578 292094 436814
rect 291474 401134 292094 436578
rect 291474 400898 291506 401134
rect 291742 400898 291826 401134
rect 292062 400898 292094 401134
rect 291474 400814 292094 400898
rect 291474 400578 291506 400814
rect 291742 400578 291826 400814
rect 292062 400578 292094 400814
rect 291474 365134 292094 400578
rect 291474 364898 291506 365134
rect 291742 364898 291826 365134
rect 292062 364898 292094 365134
rect 291474 364814 292094 364898
rect 291474 364578 291506 364814
rect 291742 364578 291826 364814
rect 292062 364578 292094 364814
rect 291474 329134 292094 364578
rect 291474 328898 291506 329134
rect 291742 328898 291826 329134
rect 292062 328898 292094 329134
rect 291474 328814 292094 328898
rect 291474 328578 291506 328814
rect 291742 328578 291826 328814
rect 292062 328578 292094 328814
rect 291474 293134 292094 328578
rect 291474 292898 291506 293134
rect 291742 292898 291826 293134
rect 292062 292898 292094 293134
rect 291474 292814 292094 292898
rect 291474 292578 291506 292814
rect 291742 292578 291826 292814
rect 292062 292578 292094 292814
rect 291474 257134 292094 292578
rect 291474 256898 291506 257134
rect 291742 256898 291826 257134
rect 292062 256898 292094 257134
rect 291474 256814 292094 256898
rect 291474 256578 291506 256814
rect 291742 256578 291826 256814
rect 292062 256578 292094 256814
rect 291474 221134 292094 256578
rect 291474 220898 291506 221134
rect 291742 220898 291826 221134
rect 292062 220898 292094 221134
rect 291474 220814 292094 220898
rect 291474 220578 291506 220814
rect 291742 220578 291826 220814
rect 292062 220578 292094 220814
rect 291474 185134 292094 220578
rect 291474 184898 291506 185134
rect 291742 184898 291826 185134
rect 292062 184898 292094 185134
rect 291474 184814 292094 184898
rect 291474 184578 291506 184814
rect 291742 184578 291826 184814
rect 292062 184578 292094 184814
rect 291474 149134 292094 184578
rect 291474 148898 291506 149134
rect 291742 148898 291826 149134
rect 292062 148898 292094 149134
rect 291474 148814 292094 148898
rect 291474 148578 291506 148814
rect 291742 148578 291826 148814
rect 292062 148578 292094 148814
rect 291474 113134 292094 148578
rect 291474 112898 291506 113134
rect 291742 112898 291826 113134
rect 292062 112898 292094 113134
rect 291474 112814 292094 112898
rect 291474 112578 291506 112814
rect 291742 112578 291826 112814
rect 292062 112578 292094 112814
rect 291474 77134 292094 112578
rect 291474 76898 291506 77134
rect 291742 76898 291826 77134
rect 292062 76898 292094 77134
rect 291474 76814 292094 76898
rect 291474 76578 291506 76814
rect 291742 76578 291826 76814
rect 292062 76578 292094 76814
rect 291474 41134 292094 76578
rect 291474 40898 291506 41134
rect 291742 40898 291826 41134
rect 292062 40898 292094 41134
rect 291474 40814 292094 40898
rect 291474 40578 291506 40814
rect 291742 40578 291826 40814
rect 292062 40578 292094 40814
rect 291474 5134 292094 40578
rect 291474 4898 291506 5134
rect 291742 4898 291826 5134
rect 292062 4898 292094 5134
rect 291474 4814 292094 4898
rect 291474 4578 291506 4814
rect 291742 4578 291826 4814
rect 292062 4578 292094 4814
rect 291474 -2266 292094 4578
rect 291474 -2502 291506 -2266
rect 291742 -2502 291826 -2266
rect 292062 -2502 292094 -2266
rect 291474 -2586 292094 -2502
rect 291474 -2822 291506 -2586
rect 291742 -2822 291826 -2586
rect 292062 -2822 292094 -2586
rect 291474 -7654 292094 -2822
rect 292714 707718 293334 711590
rect 292714 707482 292746 707718
rect 292982 707482 293066 707718
rect 293302 707482 293334 707718
rect 292714 707398 293334 707482
rect 292714 707162 292746 707398
rect 292982 707162 293066 707398
rect 293302 707162 293334 707398
rect 292714 690374 293334 707162
rect 292714 690138 292746 690374
rect 292982 690138 293066 690374
rect 293302 690138 293334 690374
rect 292714 690054 293334 690138
rect 292714 689818 292746 690054
rect 292982 689818 293066 690054
rect 293302 689818 293334 690054
rect 292714 654374 293334 689818
rect 292714 654138 292746 654374
rect 292982 654138 293066 654374
rect 293302 654138 293334 654374
rect 292714 654054 293334 654138
rect 292714 653818 292746 654054
rect 292982 653818 293066 654054
rect 293302 653818 293334 654054
rect 292714 618374 293334 653818
rect 292714 618138 292746 618374
rect 292982 618138 293066 618374
rect 293302 618138 293334 618374
rect 292714 618054 293334 618138
rect 292714 617818 292746 618054
rect 292982 617818 293066 618054
rect 293302 617818 293334 618054
rect 292714 582374 293334 617818
rect 292714 582138 292746 582374
rect 292982 582138 293066 582374
rect 293302 582138 293334 582374
rect 292714 582054 293334 582138
rect 292714 581818 292746 582054
rect 292982 581818 293066 582054
rect 293302 581818 293334 582054
rect 292714 546374 293334 581818
rect 292714 546138 292746 546374
rect 292982 546138 293066 546374
rect 293302 546138 293334 546374
rect 292714 546054 293334 546138
rect 292714 545818 292746 546054
rect 292982 545818 293066 546054
rect 293302 545818 293334 546054
rect 292714 510374 293334 545818
rect 292714 510138 292746 510374
rect 292982 510138 293066 510374
rect 293302 510138 293334 510374
rect 292714 510054 293334 510138
rect 292714 509818 292746 510054
rect 292982 509818 293066 510054
rect 293302 509818 293334 510054
rect 292714 474374 293334 509818
rect 292714 474138 292746 474374
rect 292982 474138 293066 474374
rect 293302 474138 293334 474374
rect 292714 474054 293334 474138
rect 292714 473818 292746 474054
rect 292982 473818 293066 474054
rect 293302 473818 293334 474054
rect 292714 438374 293334 473818
rect 292714 438138 292746 438374
rect 292982 438138 293066 438374
rect 293302 438138 293334 438374
rect 292714 438054 293334 438138
rect 292714 437818 292746 438054
rect 292982 437818 293066 438054
rect 293302 437818 293334 438054
rect 292714 402374 293334 437818
rect 292714 402138 292746 402374
rect 292982 402138 293066 402374
rect 293302 402138 293334 402374
rect 292714 402054 293334 402138
rect 292714 401818 292746 402054
rect 292982 401818 293066 402054
rect 293302 401818 293334 402054
rect 292714 366374 293334 401818
rect 292714 366138 292746 366374
rect 292982 366138 293066 366374
rect 293302 366138 293334 366374
rect 292714 366054 293334 366138
rect 292714 365818 292746 366054
rect 292982 365818 293066 366054
rect 293302 365818 293334 366054
rect 292714 330374 293334 365818
rect 292714 330138 292746 330374
rect 292982 330138 293066 330374
rect 293302 330138 293334 330374
rect 292714 330054 293334 330138
rect 292714 329818 292746 330054
rect 292982 329818 293066 330054
rect 293302 329818 293334 330054
rect 292714 294374 293334 329818
rect 292714 294138 292746 294374
rect 292982 294138 293066 294374
rect 293302 294138 293334 294374
rect 292714 294054 293334 294138
rect 292714 293818 292746 294054
rect 292982 293818 293066 294054
rect 293302 293818 293334 294054
rect 292714 258374 293334 293818
rect 292714 258138 292746 258374
rect 292982 258138 293066 258374
rect 293302 258138 293334 258374
rect 292714 258054 293334 258138
rect 292714 257818 292746 258054
rect 292982 257818 293066 258054
rect 293302 257818 293334 258054
rect 292714 222374 293334 257818
rect 292714 222138 292746 222374
rect 292982 222138 293066 222374
rect 293302 222138 293334 222374
rect 292714 222054 293334 222138
rect 292714 221818 292746 222054
rect 292982 221818 293066 222054
rect 293302 221818 293334 222054
rect 292714 186374 293334 221818
rect 292714 186138 292746 186374
rect 292982 186138 293066 186374
rect 293302 186138 293334 186374
rect 292714 186054 293334 186138
rect 292714 185818 292746 186054
rect 292982 185818 293066 186054
rect 293302 185818 293334 186054
rect 292714 150374 293334 185818
rect 292714 150138 292746 150374
rect 292982 150138 293066 150374
rect 293302 150138 293334 150374
rect 292714 150054 293334 150138
rect 292714 149818 292746 150054
rect 292982 149818 293066 150054
rect 293302 149818 293334 150054
rect 292714 114374 293334 149818
rect 292714 114138 292746 114374
rect 292982 114138 293066 114374
rect 293302 114138 293334 114374
rect 292714 114054 293334 114138
rect 292714 113818 292746 114054
rect 292982 113818 293066 114054
rect 293302 113818 293334 114054
rect 292714 78374 293334 113818
rect 292714 78138 292746 78374
rect 292982 78138 293066 78374
rect 293302 78138 293334 78374
rect 292714 78054 293334 78138
rect 292714 77818 292746 78054
rect 292982 77818 293066 78054
rect 293302 77818 293334 78054
rect 292714 42374 293334 77818
rect 292714 42138 292746 42374
rect 292982 42138 293066 42374
rect 293302 42138 293334 42374
rect 292714 42054 293334 42138
rect 292714 41818 292746 42054
rect 292982 41818 293066 42054
rect 293302 41818 293334 42054
rect 292714 6374 293334 41818
rect 292714 6138 292746 6374
rect 292982 6138 293066 6374
rect 293302 6138 293334 6374
rect 292714 6054 293334 6138
rect 292714 5818 292746 6054
rect 292982 5818 293066 6054
rect 293302 5818 293334 6054
rect 292714 -3226 293334 5818
rect 292714 -3462 292746 -3226
rect 292982 -3462 293066 -3226
rect 293302 -3462 293334 -3226
rect 292714 -3546 293334 -3462
rect 292714 -3782 292746 -3546
rect 292982 -3782 293066 -3546
rect 293302 -3782 293334 -3546
rect 292714 -7654 293334 -3782
rect 293954 708678 294574 711590
rect 293954 708442 293986 708678
rect 294222 708442 294306 708678
rect 294542 708442 294574 708678
rect 293954 708358 294574 708442
rect 293954 708122 293986 708358
rect 294222 708122 294306 708358
rect 294542 708122 294574 708358
rect 293954 691614 294574 708122
rect 293954 691378 293986 691614
rect 294222 691378 294306 691614
rect 294542 691378 294574 691614
rect 293954 691294 294574 691378
rect 293954 691058 293986 691294
rect 294222 691058 294306 691294
rect 294542 691058 294574 691294
rect 293954 655614 294574 691058
rect 293954 655378 293986 655614
rect 294222 655378 294306 655614
rect 294542 655378 294574 655614
rect 293954 655294 294574 655378
rect 293954 655058 293986 655294
rect 294222 655058 294306 655294
rect 294542 655058 294574 655294
rect 293954 619614 294574 655058
rect 293954 619378 293986 619614
rect 294222 619378 294306 619614
rect 294542 619378 294574 619614
rect 293954 619294 294574 619378
rect 293954 619058 293986 619294
rect 294222 619058 294306 619294
rect 294542 619058 294574 619294
rect 293954 583614 294574 619058
rect 293954 583378 293986 583614
rect 294222 583378 294306 583614
rect 294542 583378 294574 583614
rect 293954 583294 294574 583378
rect 293954 583058 293986 583294
rect 294222 583058 294306 583294
rect 294542 583058 294574 583294
rect 293954 547614 294574 583058
rect 293954 547378 293986 547614
rect 294222 547378 294306 547614
rect 294542 547378 294574 547614
rect 293954 547294 294574 547378
rect 293954 547058 293986 547294
rect 294222 547058 294306 547294
rect 294542 547058 294574 547294
rect 293954 511614 294574 547058
rect 293954 511378 293986 511614
rect 294222 511378 294306 511614
rect 294542 511378 294574 511614
rect 293954 511294 294574 511378
rect 293954 511058 293986 511294
rect 294222 511058 294306 511294
rect 294542 511058 294574 511294
rect 293954 475614 294574 511058
rect 293954 475378 293986 475614
rect 294222 475378 294306 475614
rect 294542 475378 294574 475614
rect 293954 475294 294574 475378
rect 293954 475058 293986 475294
rect 294222 475058 294306 475294
rect 294542 475058 294574 475294
rect 293954 439614 294574 475058
rect 293954 439378 293986 439614
rect 294222 439378 294306 439614
rect 294542 439378 294574 439614
rect 293954 439294 294574 439378
rect 293954 439058 293986 439294
rect 294222 439058 294306 439294
rect 294542 439058 294574 439294
rect 293954 403614 294574 439058
rect 293954 403378 293986 403614
rect 294222 403378 294306 403614
rect 294542 403378 294574 403614
rect 293954 403294 294574 403378
rect 293954 403058 293986 403294
rect 294222 403058 294306 403294
rect 294542 403058 294574 403294
rect 293954 367614 294574 403058
rect 293954 367378 293986 367614
rect 294222 367378 294306 367614
rect 294542 367378 294574 367614
rect 293954 367294 294574 367378
rect 293954 367058 293986 367294
rect 294222 367058 294306 367294
rect 294542 367058 294574 367294
rect 293954 331614 294574 367058
rect 293954 331378 293986 331614
rect 294222 331378 294306 331614
rect 294542 331378 294574 331614
rect 293954 331294 294574 331378
rect 293954 331058 293986 331294
rect 294222 331058 294306 331294
rect 294542 331058 294574 331294
rect 293954 295614 294574 331058
rect 293954 295378 293986 295614
rect 294222 295378 294306 295614
rect 294542 295378 294574 295614
rect 293954 295294 294574 295378
rect 293954 295058 293986 295294
rect 294222 295058 294306 295294
rect 294542 295058 294574 295294
rect 293954 259614 294574 295058
rect 293954 259378 293986 259614
rect 294222 259378 294306 259614
rect 294542 259378 294574 259614
rect 293954 259294 294574 259378
rect 293954 259058 293986 259294
rect 294222 259058 294306 259294
rect 294542 259058 294574 259294
rect 293954 223614 294574 259058
rect 293954 223378 293986 223614
rect 294222 223378 294306 223614
rect 294542 223378 294574 223614
rect 293954 223294 294574 223378
rect 293954 223058 293986 223294
rect 294222 223058 294306 223294
rect 294542 223058 294574 223294
rect 293954 187614 294574 223058
rect 293954 187378 293986 187614
rect 294222 187378 294306 187614
rect 294542 187378 294574 187614
rect 293954 187294 294574 187378
rect 293954 187058 293986 187294
rect 294222 187058 294306 187294
rect 294542 187058 294574 187294
rect 293954 151614 294574 187058
rect 293954 151378 293986 151614
rect 294222 151378 294306 151614
rect 294542 151378 294574 151614
rect 293954 151294 294574 151378
rect 293954 151058 293986 151294
rect 294222 151058 294306 151294
rect 294542 151058 294574 151294
rect 293954 115614 294574 151058
rect 293954 115378 293986 115614
rect 294222 115378 294306 115614
rect 294542 115378 294574 115614
rect 293954 115294 294574 115378
rect 293954 115058 293986 115294
rect 294222 115058 294306 115294
rect 294542 115058 294574 115294
rect 293954 79614 294574 115058
rect 293954 79378 293986 79614
rect 294222 79378 294306 79614
rect 294542 79378 294574 79614
rect 293954 79294 294574 79378
rect 293954 79058 293986 79294
rect 294222 79058 294306 79294
rect 294542 79058 294574 79294
rect 293954 43614 294574 79058
rect 293954 43378 293986 43614
rect 294222 43378 294306 43614
rect 294542 43378 294574 43614
rect 293954 43294 294574 43378
rect 293954 43058 293986 43294
rect 294222 43058 294306 43294
rect 294542 43058 294574 43294
rect 293954 7614 294574 43058
rect 293954 7378 293986 7614
rect 294222 7378 294306 7614
rect 294542 7378 294574 7614
rect 293954 7294 294574 7378
rect 293954 7058 293986 7294
rect 294222 7058 294306 7294
rect 294542 7058 294574 7294
rect 293954 -4186 294574 7058
rect 293954 -4422 293986 -4186
rect 294222 -4422 294306 -4186
rect 294542 -4422 294574 -4186
rect 293954 -4506 294574 -4422
rect 293954 -4742 293986 -4506
rect 294222 -4742 294306 -4506
rect 294542 -4742 294574 -4506
rect 293954 -7654 294574 -4742
rect 295194 709638 295814 711590
rect 295194 709402 295226 709638
rect 295462 709402 295546 709638
rect 295782 709402 295814 709638
rect 295194 709318 295814 709402
rect 295194 709082 295226 709318
rect 295462 709082 295546 709318
rect 295782 709082 295814 709318
rect 295194 692854 295814 709082
rect 295194 692618 295226 692854
rect 295462 692618 295546 692854
rect 295782 692618 295814 692854
rect 295194 692534 295814 692618
rect 295194 692298 295226 692534
rect 295462 692298 295546 692534
rect 295782 692298 295814 692534
rect 295194 656854 295814 692298
rect 295194 656618 295226 656854
rect 295462 656618 295546 656854
rect 295782 656618 295814 656854
rect 295194 656534 295814 656618
rect 295194 656298 295226 656534
rect 295462 656298 295546 656534
rect 295782 656298 295814 656534
rect 295194 620854 295814 656298
rect 295194 620618 295226 620854
rect 295462 620618 295546 620854
rect 295782 620618 295814 620854
rect 295194 620534 295814 620618
rect 295194 620298 295226 620534
rect 295462 620298 295546 620534
rect 295782 620298 295814 620534
rect 295194 584854 295814 620298
rect 295194 584618 295226 584854
rect 295462 584618 295546 584854
rect 295782 584618 295814 584854
rect 295194 584534 295814 584618
rect 295194 584298 295226 584534
rect 295462 584298 295546 584534
rect 295782 584298 295814 584534
rect 295194 548854 295814 584298
rect 295194 548618 295226 548854
rect 295462 548618 295546 548854
rect 295782 548618 295814 548854
rect 295194 548534 295814 548618
rect 295194 548298 295226 548534
rect 295462 548298 295546 548534
rect 295782 548298 295814 548534
rect 295194 512854 295814 548298
rect 295194 512618 295226 512854
rect 295462 512618 295546 512854
rect 295782 512618 295814 512854
rect 295194 512534 295814 512618
rect 295194 512298 295226 512534
rect 295462 512298 295546 512534
rect 295782 512298 295814 512534
rect 295194 476854 295814 512298
rect 295194 476618 295226 476854
rect 295462 476618 295546 476854
rect 295782 476618 295814 476854
rect 295194 476534 295814 476618
rect 295194 476298 295226 476534
rect 295462 476298 295546 476534
rect 295782 476298 295814 476534
rect 295194 440854 295814 476298
rect 295194 440618 295226 440854
rect 295462 440618 295546 440854
rect 295782 440618 295814 440854
rect 295194 440534 295814 440618
rect 295194 440298 295226 440534
rect 295462 440298 295546 440534
rect 295782 440298 295814 440534
rect 295194 404854 295814 440298
rect 295194 404618 295226 404854
rect 295462 404618 295546 404854
rect 295782 404618 295814 404854
rect 295194 404534 295814 404618
rect 295194 404298 295226 404534
rect 295462 404298 295546 404534
rect 295782 404298 295814 404534
rect 295194 368854 295814 404298
rect 295194 368618 295226 368854
rect 295462 368618 295546 368854
rect 295782 368618 295814 368854
rect 295194 368534 295814 368618
rect 295194 368298 295226 368534
rect 295462 368298 295546 368534
rect 295782 368298 295814 368534
rect 295194 332854 295814 368298
rect 295194 332618 295226 332854
rect 295462 332618 295546 332854
rect 295782 332618 295814 332854
rect 295194 332534 295814 332618
rect 295194 332298 295226 332534
rect 295462 332298 295546 332534
rect 295782 332298 295814 332534
rect 295194 296854 295814 332298
rect 295194 296618 295226 296854
rect 295462 296618 295546 296854
rect 295782 296618 295814 296854
rect 295194 296534 295814 296618
rect 295194 296298 295226 296534
rect 295462 296298 295546 296534
rect 295782 296298 295814 296534
rect 295194 260854 295814 296298
rect 295194 260618 295226 260854
rect 295462 260618 295546 260854
rect 295782 260618 295814 260854
rect 295194 260534 295814 260618
rect 295194 260298 295226 260534
rect 295462 260298 295546 260534
rect 295782 260298 295814 260534
rect 295194 224854 295814 260298
rect 295194 224618 295226 224854
rect 295462 224618 295546 224854
rect 295782 224618 295814 224854
rect 295194 224534 295814 224618
rect 295194 224298 295226 224534
rect 295462 224298 295546 224534
rect 295782 224298 295814 224534
rect 295194 188854 295814 224298
rect 295194 188618 295226 188854
rect 295462 188618 295546 188854
rect 295782 188618 295814 188854
rect 295194 188534 295814 188618
rect 295194 188298 295226 188534
rect 295462 188298 295546 188534
rect 295782 188298 295814 188534
rect 295194 152854 295814 188298
rect 295194 152618 295226 152854
rect 295462 152618 295546 152854
rect 295782 152618 295814 152854
rect 295194 152534 295814 152618
rect 295194 152298 295226 152534
rect 295462 152298 295546 152534
rect 295782 152298 295814 152534
rect 295194 116854 295814 152298
rect 295194 116618 295226 116854
rect 295462 116618 295546 116854
rect 295782 116618 295814 116854
rect 295194 116534 295814 116618
rect 295194 116298 295226 116534
rect 295462 116298 295546 116534
rect 295782 116298 295814 116534
rect 295194 80854 295814 116298
rect 295194 80618 295226 80854
rect 295462 80618 295546 80854
rect 295782 80618 295814 80854
rect 295194 80534 295814 80618
rect 295194 80298 295226 80534
rect 295462 80298 295546 80534
rect 295782 80298 295814 80534
rect 295194 44854 295814 80298
rect 295194 44618 295226 44854
rect 295462 44618 295546 44854
rect 295782 44618 295814 44854
rect 295194 44534 295814 44618
rect 295194 44298 295226 44534
rect 295462 44298 295546 44534
rect 295782 44298 295814 44534
rect 295194 8854 295814 44298
rect 295194 8618 295226 8854
rect 295462 8618 295546 8854
rect 295782 8618 295814 8854
rect 295194 8534 295814 8618
rect 295194 8298 295226 8534
rect 295462 8298 295546 8534
rect 295782 8298 295814 8534
rect 295194 -5146 295814 8298
rect 295194 -5382 295226 -5146
rect 295462 -5382 295546 -5146
rect 295782 -5382 295814 -5146
rect 295194 -5466 295814 -5382
rect 295194 -5702 295226 -5466
rect 295462 -5702 295546 -5466
rect 295782 -5702 295814 -5466
rect 295194 -7654 295814 -5702
rect 296434 710598 297054 711590
rect 296434 710362 296466 710598
rect 296702 710362 296786 710598
rect 297022 710362 297054 710598
rect 296434 710278 297054 710362
rect 296434 710042 296466 710278
rect 296702 710042 296786 710278
rect 297022 710042 297054 710278
rect 296434 694094 297054 710042
rect 296434 693858 296466 694094
rect 296702 693858 296786 694094
rect 297022 693858 297054 694094
rect 296434 693774 297054 693858
rect 296434 693538 296466 693774
rect 296702 693538 296786 693774
rect 297022 693538 297054 693774
rect 296434 658094 297054 693538
rect 296434 657858 296466 658094
rect 296702 657858 296786 658094
rect 297022 657858 297054 658094
rect 296434 657774 297054 657858
rect 296434 657538 296466 657774
rect 296702 657538 296786 657774
rect 297022 657538 297054 657774
rect 296434 622094 297054 657538
rect 296434 621858 296466 622094
rect 296702 621858 296786 622094
rect 297022 621858 297054 622094
rect 296434 621774 297054 621858
rect 296434 621538 296466 621774
rect 296702 621538 296786 621774
rect 297022 621538 297054 621774
rect 296434 586094 297054 621538
rect 296434 585858 296466 586094
rect 296702 585858 296786 586094
rect 297022 585858 297054 586094
rect 296434 585774 297054 585858
rect 296434 585538 296466 585774
rect 296702 585538 296786 585774
rect 297022 585538 297054 585774
rect 296434 550094 297054 585538
rect 296434 549858 296466 550094
rect 296702 549858 296786 550094
rect 297022 549858 297054 550094
rect 296434 549774 297054 549858
rect 296434 549538 296466 549774
rect 296702 549538 296786 549774
rect 297022 549538 297054 549774
rect 296434 514094 297054 549538
rect 296434 513858 296466 514094
rect 296702 513858 296786 514094
rect 297022 513858 297054 514094
rect 296434 513774 297054 513858
rect 296434 513538 296466 513774
rect 296702 513538 296786 513774
rect 297022 513538 297054 513774
rect 296434 478094 297054 513538
rect 296434 477858 296466 478094
rect 296702 477858 296786 478094
rect 297022 477858 297054 478094
rect 296434 477774 297054 477858
rect 296434 477538 296466 477774
rect 296702 477538 296786 477774
rect 297022 477538 297054 477774
rect 296434 442094 297054 477538
rect 296434 441858 296466 442094
rect 296702 441858 296786 442094
rect 297022 441858 297054 442094
rect 296434 441774 297054 441858
rect 296434 441538 296466 441774
rect 296702 441538 296786 441774
rect 297022 441538 297054 441774
rect 296434 406094 297054 441538
rect 296434 405858 296466 406094
rect 296702 405858 296786 406094
rect 297022 405858 297054 406094
rect 296434 405774 297054 405858
rect 296434 405538 296466 405774
rect 296702 405538 296786 405774
rect 297022 405538 297054 405774
rect 296434 370094 297054 405538
rect 296434 369858 296466 370094
rect 296702 369858 296786 370094
rect 297022 369858 297054 370094
rect 296434 369774 297054 369858
rect 296434 369538 296466 369774
rect 296702 369538 296786 369774
rect 297022 369538 297054 369774
rect 296434 334094 297054 369538
rect 296434 333858 296466 334094
rect 296702 333858 296786 334094
rect 297022 333858 297054 334094
rect 296434 333774 297054 333858
rect 296434 333538 296466 333774
rect 296702 333538 296786 333774
rect 297022 333538 297054 333774
rect 296434 298094 297054 333538
rect 296434 297858 296466 298094
rect 296702 297858 296786 298094
rect 297022 297858 297054 298094
rect 296434 297774 297054 297858
rect 296434 297538 296466 297774
rect 296702 297538 296786 297774
rect 297022 297538 297054 297774
rect 296434 262094 297054 297538
rect 296434 261858 296466 262094
rect 296702 261858 296786 262094
rect 297022 261858 297054 262094
rect 296434 261774 297054 261858
rect 296434 261538 296466 261774
rect 296702 261538 296786 261774
rect 297022 261538 297054 261774
rect 296434 226094 297054 261538
rect 296434 225858 296466 226094
rect 296702 225858 296786 226094
rect 297022 225858 297054 226094
rect 296434 225774 297054 225858
rect 296434 225538 296466 225774
rect 296702 225538 296786 225774
rect 297022 225538 297054 225774
rect 296434 190094 297054 225538
rect 296434 189858 296466 190094
rect 296702 189858 296786 190094
rect 297022 189858 297054 190094
rect 296434 189774 297054 189858
rect 296434 189538 296466 189774
rect 296702 189538 296786 189774
rect 297022 189538 297054 189774
rect 296434 154094 297054 189538
rect 296434 153858 296466 154094
rect 296702 153858 296786 154094
rect 297022 153858 297054 154094
rect 296434 153774 297054 153858
rect 296434 153538 296466 153774
rect 296702 153538 296786 153774
rect 297022 153538 297054 153774
rect 296434 118094 297054 153538
rect 296434 117858 296466 118094
rect 296702 117858 296786 118094
rect 297022 117858 297054 118094
rect 296434 117774 297054 117858
rect 296434 117538 296466 117774
rect 296702 117538 296786 117774
rect 297022 117538 297054 117774
rect 296434 82094 297054 117538
rect 296434 81858 296466 82094
rect 296702 81858 296786 82094
rect 297022 81858 297054 82094
rect 296434 81774 297054 81858
rect 296434 81538 296466 81774
rect 296702 81538 296786 81774
rect 297022 81538 297054 81774
rect 296434 46094 297054 81538
rect 296434 45858 296466 46094
rect 296702 45858 296786 46094
rect 297022 45858 297054 46094
rect 296434 45774 297054 45858
rect 296434 45538 296466 45774
rect 296702 45538 296786 45774
rect 297022 45538 297054 45774
rect 296434 10094 297054 45538
rect 296434 9858 296466 10094
rect 296702 9858 296786 10094
rect 297022 9858 297054 10094
rect 296434 9774 297054 9858
rect 296434 9538 296466 9774
rect 296702 9538 296786 9774
rect 297022 9538 297054 9774
rect 296434 -6106 297054 9538
rect 296434 -6342 296466 -6106
rect 296702 -6342 296786 -6106
rect 297022 -6342 297054 -6106
rect 296434 -6426 297054 -6342
rect 296434 -6662 296466 -6426
rect 296702 -6662 296786 -6426
rect 297022 -6662 297054 -6426
rect 296434 -7654 297054 -6662
rect 297674 711558 298294 711590
rect 297674 711322 297706 711558
rect 297942 711322 298026 711558
rect 298262 711322 298294 711558
rect 297674 711238 298294 711322
rect 297674 711002 297706 711238
rect 297942 711002 298026 711238
rect 298262 711002 298294 711238
rect 297674 695334 298294 711002
rect 297674 695098 297706 695334
rect 297942 695098 298026 695334
rect 298262 695098 298294 695334
rect 297674 695014 298294 695098
rect 297674 694778 297706 695014
rect 297942 694778 298026 695014
rect 298262 694778 298294 695014
rect 297674 659334 298294 694778
rect 297674 659098 297706 659334
rect 297942 659098 298026 659334
rect 298262 659098 298294 659334
rect 297674 659014 298294 659098
rect 297674 658778 297706 659014
rect 297942 658778 298026 659014
rect 298262 658778 298294 659014
rect 297674 623334 298294 658778
rect 297674 623098 297706 623334
rect 297942 623098 298026 623334
rect 298262 623098 298294 623334
rect 297674 623014 298294 623098
rect 297674 622778 297706 623014
rect 297942 622778 298026 623014
rect 298262 622778 298294 623014
rect 297674 587334 298294 622778
rect 297674 587098 297706 587334
rect 297942 587098 298026 587334
rect 298262 587098 298294 587334
rect 297674 587014 298294 587098
rect 297674 586778 297706 587014
rect 297942 586778 298026 587014
rect 298262 586778 298294 587014
rect 297674 551334 298294 586778
rect 297674 551098 297706 551334
rect 297942 551098 298026 551334
rect 298262 551098 298294 551334
rect 297674 551014 298294 551098
rect 297674 550778 297706 551014
rect 297942 550778 298026 551014
rect 298262 550778 298294 551014
rect 297674 515334 298294 550778
rect 297674 515098 297706 515334
rect 297942 515098 298026 515334
rect 298262 515098 298294 515334
rect 297674 515014 298294 515098
rect 297674 514778 297706 515014
rect 297942 514778 298026 515014
rect 298262 514778 298294 515014
rect 297674 479334 298294 514778
rect 297674 479098 297706 479334
rect 297942 479098 298026 479334
rect 298262 479098 298294 479334
rect 297674 479014 298294 479098
rect 297674 478778 297706 479014
rect 297942 478778 298026 479014
rect 298262 478778 298294 479014
rect 297674 443334 298294 478778
rect 297674 443098 297706 443334
rect 297942 443098 298026 443334
rect 298262 443098 298294 443334
rect 297674 443014 298294 443098
rect 297674 442778 297706 443014
rect 297942 442778 298026 443014
rect 298262 442778 298294 443014
rect 297674 407334 298294 442778
rect 297674 407098 297706 407334
rect 297942 407098 298026 407334
rect 298262 407098 298294 407334
rect 297674 407014 298294 407098
rect 297674 406778 297706 407014
rect 297942 406778 298026 407014
rect 298262 406778 298294 407014
rect 297674 371334 298294 406778
rect 297674 371098 297706 371334
rect 297942 371098 298026 371334
rect 298262 371098 298294 371334
rect 297674 371014 298294 371098
rect 297674 370778 297706 371014
rect 297942 370778 298026 371014
rect 298262 370778 298294 371014
rect 297674 335334 298294 370778
rect 297674 335098 297706 335334
rect 297942 335098 298026 335334
rect 298262 335098 298294 335334
rect 297674 335014 298294 335098
rect 297674 334778 297706 335014
rect 297942 334778 298026 335014
rect 298262 334778 298294 335014
rect 297674 299334 298294 334778
rect 297674 299098 297706 299334
rect 297942 299098 298026 299334
rect 298262 299098 298294 299334
rect 297674 299014 298294 299098
rect 297674 298778 297706 299014
rect 297942 298778 298026 299014
rect 298262 298778 298294 299014
rect 297674 263334 298294 298778
rect 297674 263098 297706 263334
rect 297942 263098 298026 263334
rect 298262 263098 298294 263334
rect 297674 263014 298294 263098
rect 297674 262778 297706 263014
rect 297942 262778 298026 263014
rect 298262 262778 298294 263014
rect 297674 227334 298294 262778
rect 297674 227098 297706 227334
rect 297942 227098 298026 227334
rect 298262 227098 298294 227334
rect 297674 227014 298294 227098
rect 297674 226778 297706 227014
rect 297942 226778 298026 227014
rect 298262 226778 298294 227014
rect 297674 191334 298294 226778
rect 297674 191098 297706 191334
rect 297942 191098 298026 191334
rect 298262 191098 298294 191334
rect 297674 191014 298294 191098
rect 297674 190778 297706 191014
rect 297942 190778 298026 191014
rect 298262 190778 298294 191014
rect 297674 155334 298294 190778
rect 297674 155098 297706 155334
rect 297942 155098 298026 155334
rect 298262 155098 298294 155334
rect 297674 155014 298294 155098
rect 297674 154778 297706 155014
rect 297942 154778 298026 155014
rect 298262 154778 298294 155014
rect 297674 119334 298294 154778
rect 297674 119098 297706 119334
rect 297942 119098 298026 119334
rect 298262 119098 298294 119334
rect 297674 119014 298294 119098
rect 297674 118778 297706 119014
rect 297942 118778 298026 119014
rect 298262 118778 298294 119014
rect 297674 83334 298294 118778
rect 297674 83098 297706 83334
rect 297942 83098 298026 83334
rect 298262 83098 298294 83334
rect 297674 83014 298294 83098
rect 297674 82778 297706 83014
rect 297942 82778 298026 83014
rect 298262 82778 298294 83014
rect 297674 47334 298294 82778
rect 297674 47098 297706 47334
rect 297942 47098 298026 47334
rect 298262 47098 298294 47334
rect 297674 47014 298294 47098
rect 297674 46778 297706 47014
rect 297942 46778 298026 47014
rect 298262 46778 298294 47014
rect 297674 11334 298294 46778
rect 297674 11098 297706 11334
rect 297942 11098 298026 11334
rect 298262 11098 298294 11334
rect 297674 11014 298294 11098
rect 297674 10778 297706 11014
rect 297942 10778 298026 11014
rect 298262 10778 298294 11014
rect 297674 -7066 298294 10778
rect 297674 -7302 297706 -7066
rect 297942 -7302 298026 -7066
rect 298262 -7302 298294 -7066
rect 297674 -7386 298294 -7302
rect 297674 -7622 297706 -7386
rect 297942 -7622 298026 -7386
rect 298262 -7622 298294 -7386
rect 297674 -7654 298294 -7622
rect 324994 704838 325614 711590
rect 324994 704602 325026 704838
rect 325262 704602 325346 704838
rect 325582 704602 325614 704838
rect 324994 704518 325614 704602
rect 324994 704282 325026 704518
rect 325262 704282 325346 704518
rect 325582 704282 325614 704518
rect 324994 686654 325614 704282
rect 324994 686418 325026 686654
rect 325262 686418 325346 686654
rect 325582 686418 325614 686654
rect 324994 686334 325614 686418
rect 324994 686098 325026 686334
rect 325262 686098 325346 686334
rect 325582 686098 325614 686334
rect 324994 650654 325614 686098
rect 324994 650418 325026 650654
rect 325262 650418 325346 650654
rect 325582 650418 325614 650654
rect 324994 650334 325614 650418
rect 324994 650098 325026 650334
rect 325262 650098 325346 650334
rect 325582 650098 325614 650334
rect 324994 614654 325614 650098
rect 324994 614418 325026 614654
rect 325262 614418 325346 614654
rect 325582 614418 325614 614654
rect 324994 614334 325614 614418
rect 324994 614098 325026 614334
rect 325262 614098 325346 614334
rect 325582 614098 325614 614334
rect 324994 578654 325614 614098
rect 324994 578418 325026 578654
rect 325262 578418 325346 578654
rect 325582 578418 325614 578654
rect 324994 578334 325614 578418
rect 324994 578098 325026 578334
rect 325262 578098 325346 578334
rect 325582 578098 325614 578334
rect 324994 542654 325614 578098
rect 324994 542418 325026 542654
rect 325262 542418 325346 542654
rect 325582 542418 325614 542654
rect 324994 542334 325614 542418
rect 324994 542098 325026 542334
rect 325262 542098 325346 542334
rect 325582 542098 325614 542334
rect 324994 506654 325614 542098
rect 324994 506418 325026 506654
rect 325262 506418 325346 506654
rect 325582 506418 325614 506654
rect 324994 506334 325614 506418
rect 324994 506098 325026 506334
rect 325262 506098 325346 506334
rect 325582 506098 325614 506334
rect 324994 470654 325614 506098
rect 324994 470418 325026 470654
rect 325262 470418 325346 470654
rect 325582 470418 325614 470654
rect 324994 470334 325614 470418
rect 324994 470098 325026 470334
rect 325262 470098 325346 470334
rect 325582 470098 325614 470334
rect 324994 434654 325614 470098
rect 324994 434418 325026 434654
rect 325262 434418 325346 434654
rect 325582 434418 325614 434654
rect 324994 434334 325614 434418
rect 324994 434098 325026 434334
rect 325262 434098 325346 434334
rect 325582 434098 325614 434334
rect 324994 398654 325614 434098
rect 324994 398418 325026 398654
rect 325262 398418 325346 398654
rect 325582 398418 325614 398654
rect 324994 398334 325614 398418
rect 324994 398098 325026 398334
rect 325262 398098 325346 398334
rect 325582 398098 325614 398334
rect 324994 362654 325614 398098
rect 324994 362418 325026 362654
rect 325262 362418 325346 362654
rect 325582 362418 325614 362654
rect 324994 362334 325614 362418
rect 324994 362098 325026 362334
rect 325262 362098 325346 362334
rect 325582 362098 325614 362334
rect 324994 326654 325614 362098
rect 324994 326418 325026 326654
rect 325262 326418 325346 326654
rect 325582 326418 325614 326654
rect 324994 326334 325614 326418
rect 324994 326098 325026 326334
rect 325262 326098 325346 326334
rect 325582 326098 325614 326334
rect 324994 290654 325614 326098
rect 324994 290418 325026 290654
rect 325262 290418 325346 290654
rect 325582 290418 325614 290654
rect 324994 290334 325614 290418
rect 324994 290098 325026 290334
rect 325262 290098 325346 290334
rect 325582 290098 325614 290334
rect 324994 254654 325614 290098
rect 324994 254418 325026 254654
rect 325262 254418 325346 254654
rect 325582 254418 325614 254654
rect 324994 254334 325614 254418
rect 324994 254098 325026 254334
rect 325262 254098 325346 254334
rect 325582 254098 325614 254334
rect 324994 218654 325614 254098
rect 324994 218418 325026 218654
rect 325262 218418 325346 218654
rect 325582 218418 325614 218654
rect 324994 218334 325614 218418
rect 324994 218098 325026 218334
rect 325262 218098 325346 218334
rect 325582 218098 325614 218334
rect 324994 182654 325614 218098
rect 324994 182418 325026 182654
rect 325262 182418 325346 182654
rect 325582 182418 325614 182654
rect 324994 182334 325614 182418
rect 324994 182098 325026 182334
rect 325262 182098 325346 182334
rect 325582 182098 325614 182334
rect 324994 146654 325614 182098
rect 324994 146418 325026 146654
rect 325262 146418 325346 146654
rect 325582 146418 325614 146654
rect 324994 146334 325614 146418
rect 324994 146098 325026 146334
rect 325262 146098 325346 146334
rect 325582 146098 325614 146334
rect 324994 110654 325614 146098
rect 324994 110418 325026 110654
rect 325262 110418 325346 110654
rect 325582 110418 325614 110654
rect 324994 110334 325614 110418
rect 324994 110098 325026 110334
rect 325262 110098 325346 110334
rect 325582 110098 325614 110334
rect 324994 74654 325614 110098
rect 324994 74418 325026 74654
rect 325262 74418 325346 74654
rect 325582 74418 325614 74654
rect 324994 74334 325614 74418
rect 324994 74098 325026 74334
rect 325262 74098 325346 74334
rect 325582 74098 325614 74334
rect 324994 38654 325614 74098
rect 324994 38418 325026 38654
rect 325262 38418 325346 38654
rect 325582 38418 325614 38654
rect 324994 38334 325614 38418
rect 324994 38098 325026 38334
rect 325262 38098 325346 38334
rect 325582 38098 325614 38334
rect 324994 2654 325614 38098
rect 324994 2418 325026 2654
rect 325262 2418 325346 2654
rect 325582 2418 325614 2654
rect 324994 2334 325614 2418
rect 324994 2098 325026 2334
rect 325262 2098 325346 2334
rect 325582 2098 325614 2334
rect 324994 -346 325614 2098
rect 324994 -582 325026 -346
rect 325262 -582 325346 -346
rect 325582 -582 325614 -346
rect 324994 -666 325614 -582
rect 324994 -902 325026 -666
rect 325262 -902 325346 -666
rect 325582 -902 325614 -666
rect 324994 -7654 325614 -902
rect 326234 705798 326854 711590
rect 326234 705562 326266 705798
rect 326502 705562 326586 705798
rect 326822 705562 326854 705798
rect 326234 705478 326854 705562
rect 326234 705242 326266 705478
rect 326502 705242 326586 705478
rect 326822 705242 326854 705478
rect 326234 687894 326854 705242
rect 326234 687658 326266 687894
rect 326502 687658 326586 687894
rect 326822 687658 326854 687894
rect 326234 687574 326854 687658
rect 326234 687338 326266 687574
rect 326502 687338 326586 687574
rect 326822 687338 326854 687574
rect 326234 651894 326854 687338
rect 326234 651658 326266 651894
rect 326502 651658 326586 651894
rect 326822 651658 326854 651894
rect 326234 651574 326854 651658
rect 326234 651338 326266 651574
rect 326502 651338 326586 651574
rect 326822 651338 326854 651574
rect 326234 615894 326854 651338
rect 326234 615658 326266 615894
rect 326502 615658 326586 615894
rect 326822 615658 326854 615894
rect 326234 615574 326854 615658
rect 326234 615338 326266 615574
rect 326502 615338 326586 615574
rect 326822 615338 326854 615574
rect 326234 579894 326854 615338
rect 326234 579658 326266 579894
rect 326502 579658 326586 579894
rect 326822 579658 326854 579894
rect 326234 579574 326854 579658
rect 326234 579338 326266 579574
rect 326502 579338 326586 579574
rect 326822 579338 326854 579574
rect 326234 543894 326854 579338
rect 326234 543658 326266 543894
rect 326502 543658 326586 543894
rect 326822 543658 326854 543894
rect 326234 543574 326854 543658
rect 326234 543338 326266 543574
rect 326502 543338 326586 543574
rect 326822 543338 326854 543574
rect 326234 507894 326854 543338
rect 326234 507658 326266 507894
rect 326502 507658 326586 507894
rect 326822 507658 326854 507894
rect 326234 507574 326854 507658
rect 326234 507338 326266 507574
rect 326502 507338 326586 507574
rect 326822 507338 326854 507574
rect 326234 471894 326854 507338
rect 326234 471658 326266 471894
rect 326502 471658 326586 471894
rect 326822 471658 326854 471894
rect 326234 471574 326854 471658
rect 326234 471338 326266 471574
rect 326502 471338 326586 471574
rect 326822 471338 326854 471574
rect 326234 435894 326854 471338
rect 326234 435658 326266 435894
rect 326502 435658 326586 435894
rect 326822 435658 326854 435894
rect 326234 435574 326854 435658
rect 326234 435338 326266 435574
rect 326502 435338 326586 435574
rect 326822 435338 326854 435574
rect 326234 399894 326854 435338
rect 326234 399658 326266 399894
rect 326502 399658 326586 399894
rect 326822 399658 326854 399894
rect 326234 399574 326854 399658
rect 326234 399338 326266 399574
rect 326502 399338 326586 399574
rect 326822 399338 326854 399574
rect 326234 363894 326854 399338
rect 326234 363658 326266 363894
rect 326502 363658 326586 363894
rect 326822 363658 326854 363894
rect 326234 363574 326854 363658
rect 326234 363338 326266 363574
rect 326502 363338 326586 363574
rect 326822 363338 326854 363574
rect 326234 327894 326854 363338
rect 326234 327658 326266 327894
rect 326502 327658 326586 327894
rect 326822 327658 326854 327894
rect 326234 327574 326854 327658
rect 326234 327338 326266 327574
rect 326502 327338 326586 327574
rect 326822 327338 326854 327574
rect 326234 291894 326854 327338
rect 326234 291658 326266 291894
rect 326502 291658 326586 291894
rect 326822 291658 326854 291894
rect 326234 291574 326854 291658
rect 326234 291338 326266 291574
rect 326502 291338 326586 291574
rect 326822 291338 326854 291574
rect 326234 255894 326854 291338
rect 326234 255658 326266 255894
rect 326502 255658 326586 255894
rect 326822 255658 326854 255894
rect 326234 255574 326854 255658
rect 326234 255338 326266 255574
rect 326502 255338 326586 255574
rect 326822 255338 326854 255574
rect 326234 219894 326854 255338
rect 326234 219658 326266 219894
rect 326502 219658 326586 219894
rect 326822 219658 326854 219894
rect 326234 219574 326854 219658
rect 326234 219338 326266 219574
rect 326502 219338 326586 219574
rect 326822 219338 326854 219574
rect 326234 183894 326854 219338
rect 326234 183658 326266 183894
rect 326502 183658 326586 183894
rect 326822 183658 326854 183894
rect 326234 183574 326854 183658
rect 326234 183338 326266 183574
rect 326502 183338 326586 183574
rect 326822 183338 326854 183574
rect 326234 147894 326854 183338
rect 326234 147658 326266 147894
rect 326502 147658 326586 147894
rect 326822 147658 326854 147894
rect 326234 147574 326854 147658
rect 326234 147338 326266 147574
rect 326502 147338 326586 147574
rect 326822 147338 326854 147574
rect 326234 111894 326854 147338
rect 326234 111658 326266 111894
rect 326502 111658 326586 111894
rect 326822 111658 326854 111894
rect 326234 111574 326854 111658
rect 326234 111338 326266 111574
rect 326502 111338 326586 111574
rect 326822 111338 326854 111574
rect 326234 75894 326854 111338
rect 326234 75658 326266 75894
rect 326502 75658 326586 75894
rect 326822 75658 326854 75894
rect 326234 75574 326854 75658
rect 326234 75338 326266 75574
rect 326502 75338 326586 75574
rect 326822 75338 326854 75574
rect 326234 39894 326854 75338
rect 326234 39658 326266 39894
rect 326502 39658 326586 39894
rect 326822 39658 326854 39894
rect 326234 39574 326854 39658
rect 326234 39338 326266 39574
rect 326502 39338 326586 39574
rect 326822 39338 326854 39574
rect 326234 3894 326854 39338
rect 326234 3658 326266 3894
rect 326502 3658 326586 3894
rect 326822 3658 326854 3894
rect 326234 3574 326854 3658
rect 326234 3338 326266 3574
rect 326502 3338 326586 3574
rect 326822 3338 326854 3574
rect 326234 -1306 326854 3338
rect 326234 -1542 326266 -1306
rect 326502 -1542 326586 -1306
rect 326822 -1542 326854 -1306
rect 326234 -1626 326854 -1542
rect 326234 -1862 326266 -1626
rect 326502 -1862 326586 -1626
rect 326822 -1862 326854 -1626
rect 326234 -7654 326854 -1862
rect 327474 706758 328094 711590
rect 327474 706522 327506 706758
rect 327742 706522 327826 706758
rect 328062 706522 328094 706758
rect 327474 706438 328094 706522
rect 327474 706202 327506 706438
rect 327742 706202 327826 706438
rect 328062 706202 328094 706438
rect 327474 689134 328094 706202
rect 327474 688898 327506 689134
rect 327742 688898 327826 689134
rect 328062 688898 328094 689134
rect 327474 688814 328094 688898
rect 327474 688578 327506 688814
rect 327742 688578 327826 688814
rect 328062 688578 328094 688814
rect 327474 653134 328094 688578
rect 327474 652898 327506 653134
rect 327742 652898 327826 653134
rect 328062 652898 328094 653134
rect 327474 652814 328094 652898
rect 327474 652578 327506 652814
rect 327742 652578 327826 652814
rect 328062 652578 328094 652814
rect 327474 617134 328094 652578
rect 327474 616898 327506 617134
rect 327742 616898 327826 617134
rect 328062 616898 328094 617134
rect 327474 616814 328094 616898
rect 327474 616578 327506 616814
rect 327742 616578 327826 616814
rect 328062 616578 328094 616814
rect 327474 581134 328094 616578
rect 327474 580898 327506 581134
rect 327742 580898 327826 581134
rect 328062 580898 328094 581134
rect 327474 580814 328094 580898
rect 327474 580578 327506 580814
rect 327742 580578 327826 580814
rect 328062 580578 328094 580814
rect 327474 545134 328094 580578
rect 327474 544898 327506 545134
rect 327742 544898 327826 545134
rect 328062 544898 328094 545134
rect 327474 544814 328094 544898
rect 327474 544578 327506 544814
rect 327742 544578 327826 544814
rect 328062 544578 328094 544814
rect 327474 509134 328094 544578
rect 327474 508898 327506 509134
rect 327742 508898 327826 509134
rect 328062 508898 328094 509134
rect 327474 508814 328094 508898
rect 327474 508578 327506 508814
rect 327742 508578 327826 508814
rect 328062 508578 328094 508814
rect 327474 473134 328094 508578
rect 327474 472898 327506 473134
rect 327742 472898 327826 473134
rect 328062 472898 328094 473134
rect 327474 472814 328094 472898
rect 327474 472578 327506 472814
rect 327742 472578 327826 472814
rect 328062 472578 328094 472814
rect 327474 437134 328094 472578
rect 327474 436898 327506 437134
rect 327742 436898 327826 437134
rect 328062 436898 328094 437134
rect 327474 436814 328094 436898
rect 327474 436578 327506 436814
rect 327742 436578 327826 436814
rect 328062 436578 328094 436814
rect 327474 401134 328094 436578
rect 327474 400898 327506 401134
rect 327742 400898 327826 401134
rect 328062 400898 328094 401134
rect 327474 400814 328094 400898
rect 327474 400578 327506 400814
rect 327742 400578 327826 400814
rect 328062 400578 328094 400814
rect 327474 365134 328094 400578
rect 327474 364898 327506 365134
rect 327742 364898 327826 365134
rect 328062 364898 328094 365134
rect 327474 364814 328094 364898
rect 327474 364578 327506 364814
rect 327742 364578 327826 364814
rect 328062 364578 328094 364814
rect 327474 329134 328094 364578
rect 327474 328898 327506 329134
rect 327742 328898 327826 329134
rect 328062 328898 328094 329134
rect 327474 328814 328094 328898
rect 327474 328578 327506 328814
rect 327742 328578 327826 328814
rect 328062 328578 328094 328814
rect 327474 293134 328094 328578
rect 327474 292898 327506 293134
rect 327742 292898 327826 293134
rect 328062 292898 328094 293134
rect 327474 292814 328094 292898
rect 327474 292578 327506 292814
rect 327742 292578 327826 292814
rect 328062 292578 328094 292814
rect 327474 257134 328094 292578
rect 327474 256898 327506 257134
rect 327742 256898 327826 257134
rect 328062 256898 328094 257134
rect 327474 256814 328094 256898
rect 327474 256578 327506 256814
rect 327742 256578 327826 256814
rect 328062 256578 328094 256814
rect 327474 221134 328094 256578
rect 327474 220898 327506 221134
rect 327742 220898 327826 221134
rect 328062 220898 328094 221134
rect 327474 220814 328094 220898
rect 327474 220578 327506 220814
rect 327742 220578 327826 220814
rect 328062 220578 328094 220814
rect 327474 185134 328094 220578
rect 327474 184898 327506 185134
rect 327742 184898 327826 185134
rect 328062 184898 328094 185134
rect 327474 184814 328094 184898
rect 327474 184578 327506 184814
rect 327742 184578 327826 184814
rect 328062 184578 328094 184814
rect 327474 149134 328094 184578
rect 327474 148898 327506 149134
rect 327742 148898 327826 149134
rect 328062 148898 328094 149134
rect 327474 148814 328094 148898
rect 327474 148578 327506 148814
rect 327742 148578 327826 148814
rect 328062 148578 328094 148814
rect 327474 113134 328094 148578
rect 327474 112898 327506 113134
rect 327742 112898 327826 113134
rect 328062 112898 328094 113134
rect 327474 112814 328094 112898
rect 327474 112578 327506 112814
rect 327742 112578 327826 112814
rect 328062 112578 328094 112814
rect 327474 77134 328094 112578
rect 327474 76898 327506 77134
rect 327742 76898 327826 77134
rect 328062 76898 328094 77134
rect 327474 76814 328094 76898
rect 327474 76578 327506 76814
rect 327742 76578 327826 76814
rect 328062 76578 328094 76814
rect 327474 41134 328094 76578
rect 327474 40898 327506 41134
rect 327742 40898 327826 41134
rect 328062 40898 328094 41134
rect 327474 40814 328094 40898
rect 327474 40578 327506 40814
rect 327742 40578 327826 40814
rect 328062 40578 328094 40814
rect 327474 5134 328094 40578
rect 327474 4898 327506 5134
rect 327742 4898 327826 5134
rect 328062 4898 328094 5134
rect 327474 4814 328094 4898
rect 327474 4578 327506 4814
rect 327742 4578 327826 4814
rect 328062 4578 328094 4814
rect 327474 -2266 328094 4578
rect 327474 -2502 327506 -2266
rect 327742 -2502 327826 -2266
rect 328062 -2502 328094 -2266
rect 327474 -2586 328094 -2502
rect 327474 -2822 327506 -2586
rect 327742 -2822 327826 -2586
rect 328062 -2822 328094 -2586
rect 327474 -7654 328094 -2822
rect 328714 707718 329334 711590
rect 328714 707482 328746 707718
rect 328982 707482 329066 707718
rect 329302 707482 329334 707718
rect 328714 707398 329334 707482
rect 328714 707162 328746 707398
rect 328982 707162 329066 707398
rect 329302 707162 329334 707398
rect 328714 690374 329334 707162
rect 328714 690138 328746 690374
rect 328982 690138 329066 690374
rect 329302 690138 329334 690374
rect 328714 690054 329334 690138
rect 328714 689818 328746 690054
rect 328982 689818 329066 690054
rect 329302 689818 329334 690054
rect 328714 654374 329334 689818
rect 328714 654138 328746 654374
rect 328982 654138 329066 654374
rect 329302 654138 329334 654374
rect 328714 654054 329334 654138
rect 328714 653818 328746 654054
rect 328982 653818 329066 654054
rect 329302 653818 329334 654054
rect 328714 618374 329334 653818
rect 328714 618138 328746 618374
rect 328982 618138 329066 618374
rect 329302 618138 329334 618374
rect 328714 618054 329334 618138
rect 328714 617818 328746 618054
rect 328982 617818 329066 618054
rect 329302 617818 329334 618054
rect 328714 582374 329334 617818
rect 328714 582138 328746 582374
rect 328982 582138 329066 582374
rect 329302 582138 329334 582374
rect 328714 582054 329334 582138
rect 328714 581818 328746 582054
rect 328982 581818 329066 582054
rect 329302 581818 329334 582054
rect 328714 546374 329334 581818
rect 328714 546138 328746 546374
rect 328982 546138 329066 546374
rect 329302 546138 329334 546374
rect 328714 546054 329334 546138
rect 328714 545818 328746 546054
rect 328982 545818 329066 546054
rect 329302 545818 329334 546054
rect 328714 510374 329334 545818
rect 328714 510138 328746 510374
rect 328982 510138 329066 510374
rect 329302 510138 329334 510374
rect 328714 510054 329334 510138
rect 328714 509818 328746 510054
rect 328982 509818 329066 510054
rect 329302 509818 329334 510054
rect 328714 474374 329334 509818
rect 328714 474138 328746 474374
rect 328982 474138 329066 474374
rect 329302 474138 329334 474374
rect 328714 474054 329334 474138
rect 328714 473818 328746 474054
rect 328982 473818 329066 474054
rect 329302 473818 329334 474054
rect 328714 438374 329334 473818
rect 328714 438138 328746 438374
rect 328982 438138 329066 438374
rect 329302 438138 329334 438374
rect 328714 438054 329334 438138
rect 328714 437818 328746 438054
rect 328982 437818 329066 438054
rect 329302 437818 329334 438054
rect 328714 402374 329334 437818
rect 328714 402138 328746 402374
rect 328982 402138 329066 402374
rect 329302 402138 329334 402374
rect 328714 402054 329334 402138
rect 328714 401818 328746 402054
rect 328982 401818 329066 402054
rect 329302 401818 329334 402054
rect 328714 366374 329334 401818
rect 328714 366138 328746 366374
rect 328982 366138 329066 366374
rect 329302 366138 329334 366374
rect 328714 366054 329334 366138
rect 328714 365818 328746 366054
rect 328982 365818 329066 366054
rect 329302 365818 329334 366054
rect 328714 330374 329334 365818
rect 328714 330138 328746 330374
rect 328982 330138 329066 330374
rect 329302 330138 329334 330374
rect 328714 330054 329334 330138
rect 328714 329818 328746 330054
rect 328982 329818 329066 330054
rect 329302 329818 329334 330054
rect 328714 294374 329334 329818
rect 328714 294138 328746 294374
rect 328982 294138 329066 294374
rect 329302 294138 329334 294374
rect 328714 294054 329334 294138
rect 328714 293818 328746 294054
rect 328982 293818 329066 294054
rect 329302 293818 329334 294054
rect 328714 258374 329334 293818
rect 328714 258138 328746 258374
rect 328982 258138 329066 258374
rect 329302 258138 329334 258374
rect 328714 258054 329334 258138
rect 328714 257818 328746 258054
rect 328982 257818 329066 258054
rect 329302 257818 329334 258054
rect 328714 222374 329334 257818
rect 328714 222138 328746 222374
rect 328982 222138 329066 222374
rect 329302 222138 329334 222374
rect 328714 222054 329334 222138
rect 328714 221818 328746 222054
rect 328982 221818 329066 222054
rect 329302 221818 329334 222054
rect 328714 186374 329334 221818
rect 328714 186138 328746 186374
rect 328982 186138 329066 186374
rect 329302 186138 329334 186374
rect 328714 186054 329334 186138
rect 328714 185818 328746 186054
rect 328982 185818 329066 186054
rect 329302 185818 329334 186054
rect 328714 150374 329334 185818
rect 328714 150138 328746 150374
rect 328982 150138 329066 150374
rect 329302 150138 329334 150374
rect 328714 150054 329334 150138
rect 328714 149818 328746 150054
rect 328982 149818 329066 150054
rect 329302 149818 329334 150054
rect 328714 114374 329334 149818
rect 328714 114138 328746 114374
rect 328982 114138 329066 114374
rect 329302 114138 329334 114374
rect 328714 114054 329334 114138
rect 328714 113818 328746 114054
rect 328982 113818 329066 114054
rect 329302 113818 329334 114054
rect 328714 78374 329334 113818
rect 328714 78138 328746 78374
rect 328982 78138 329066 78374
rect 329302 78138 329334 78374
rect 328714 78054 329334 78138
rect 328714 77818 328746 78054
rect 328982 77818 329066 78054
rect 329302 77818 329334 78054
rect 328714 42374 329334 77818
rect 328714 42138 328746 42374
rect 328982 42138 329066 42374
rect 329302 42138 329334 42374
rect 328714 42054 329334 42138
rect 328714 41818 328746 42054
rect 328982 41818 329066 42054
rect 329302 41818 329334 42054
rect 328714 6374 329334 41818
rect 328714 6138 328746 6374
rect 328982 6138 329066 6374
rect 329302 6138 329334 6374
rect 328714 6054 329334 6138
rect 328714 5818 328746 6054
rect 328982 5818 329066 6054
rect 329302 5818 329334 6054
rect 328714 -3226 329334 5818
rect 328714 -3462 328746 -3226
rect 328982 -3462 329066 -3226
rect 329302 -3462 329334 -3226
rect 328714 -3546 329334 -3462
rect 328714 -3782 328746 -3546
rect 328982 -3782 329066 -3546
rect 329302 -3782 329334 -3546
rect 328714 -7654 329334 -3782
rect 329954 708678 330574 711590
rect 329954 708442 329986 708678
rect 330222 708442 330306 708678
rect 330542 708442 330574 708678
rect 329954 708358 330574 708442
rect 329954 708122 329986 708358
rect 330222 708122 330306 708358
rect 330542 708122 330574 708358
rect 329954 691614 330574 708122
rect 329954 691378 329986 691614
rect 330222 691378 330306 691614
rect 330542 691378 330574 691614
rect 329954 691294 330574 691378
rect 329954 691058 329986 691294
rect 330222 691058 330306 691294
rect 330542 691058 330574 691294
rect 329954 655614 330574 691058
rect 329954 655378 329986 655614
rect 330222 655378 330306 655614
rect 330542 655378 330574 655614
rect 329954 655294 330574 655378
rect 329954 655058 329986 655294
rect 330222 655058 330306 655294
rect 330542 655058 330574 655294
rect 329954 619614 330574 655058
rect 329954 619378 329986 619614
rect 330222 619378 330306 619614
rect 330542 619378 330574 619614
rect 329954 619294 330574 619378
rect 329954 619058 329986 619294
rect 330222 619058 330306 619294
rect 330542 619058 330574 619294
rect 329954 583614 330574 619058
rect 329954 583378 329986 583614
rect 330222 583378 330306 583614
rect 330542 583378 330574 583614
rect 329954 583294 330574 583378
rect 329954 583058 329986 583294
rect 330222 583058 330306 583294
rect 330542 583058 330574 583294
rect 329954 547614 330574 583058
rect 329954 547378 329986 547614
rect 330222 547378 330306 547614
rect 330542 547378 330574 547614
rect 329954 547294 330574 547378
rect 329954 547058 329986 547294
rect 330222 547058 330306 547294
rect 330542 547058 330574 547294
rect 329954 511614 330574 547058
rect 329954 511378 329986 511614
rect 330222 511378 330306 511614
rect 330542 511378 330574 511614
rect 329954 511294 330574 511378
rect 329954 511058 329986 511294
rect 330222 511058 330306 511294
rect 330542 511058 330574 511294
rect 329954 475614 330574 511058
rect 329954 475378 329986 475614
rect 330222 475378 330306 475614
rect 330542 475378 330574 475614
rect 329954 475294 330574 475378
rect 329954 475058 329986 475294
rect 330222 475058 330306 475294
rect 330542 475058 330574 475294
rect 329954 439614 330574 475058
rect 329954 439378 329986 439614
rect 330222 439378 330306 439614
rect 330542 439378 330574 439614
rect 329954 439294 330574 439378
rect 329954 439058 329986 439294
rect 330222 439058 330306 439294
rect 330542 439058 330574 439294
rect 329954 403614 330574 439058
rect 329954 403378 329986 403614
rect 330222 403378 330306 403614
rect 330542 403378 330574 403614
rect 329954 403294 330574 403378
rect 329954 403058 329986 403294
rect 330222 403058 330306 403294
rect 330542 403058 330574 403294
rect 329954 367614 330574 403058
rect 329954 367378 329986 367614
rect 330222 367378 330306 367614
rect 330542 367378 330574 367614
rect 329954 367294 330574 367378
rect 329954 367058 329986 367294
rect 330222 367058 330306 367294
rect 330542 367058 330574 367294
rect 329954 331614 330574 367058
rect 329954 331378 329986 331614
rect 330222 331378 330306 331614
rect 330542 331378 330574 331614
rect 329954 331294 330574 331378
rect 329954 331058 329986 331294
rect 330222 331058 330306 331294
rect 330542 331058 330574 331294
rect 329954 295614 330574 331058
rect 329954 295378 329986 295614
rect 330222 295378 330306 295614
rect 330542 295378 330574 295614
rect 329954 295294 330574 295378
rect 329954 295058 329986 295294
rect 330222 295058 330306 295294
rect 330542 295058 330574 295294
rect 329954 259614 330574 295058
rect 329954 259378 329986 259614
rect 330222 259378 330306 259614
rect 330542 259378 330574 259614
rect 329954 259294 330574 259378
rect 329954 259058 329986 259294
rect 330222 259058 330306 259294
rect 330542 259058 330574 259294
rect 329954 223614 330574 259058
rect 329954 223378 329986 223614
rect 330222 223378 330306 223614
rect 330542 223378 330574 223614
rect 329954 223294 330574 223378
rect 329954 223058 329986 223294
rect 330222 223058 330306 223294
rect 330542 223058 330574 223294
rect 329954 187614 330574 223058
rect 329954 187378 329986 187614
rect 330222 187378 330306 187614
rect 330542 187378 330574 187614
rect 329954 187294 330574 187378
rect 329954 187058 329986 187294
rect 330222 187058 330306 187294
rect 330542 187058 330574 187294
rect 329954 151614 330574 187058
rect 329954 151378 329986 151614
rect 330222 151378 330306 151614
rect 330542 151378 330574 151614
rect 329954 151294 330574 151378
rect 329954 151058 329986 151294
rect 330222 151058 330306 151294
rect 330542 151058 330574 151294
rect 329954 115614 330574 151058
rect 329954 115378 329986 115614
rect 330222 115378 330306 115614
rect 330542 115378 330574 115614
rect 329954 115294 330574 115378
rect 329954 115058 329986 115294
rect 330222 115058 330306 115294
rect 330542 115058 330574 115294
rect 329954 79614 330574 115058
rect 329954 79378 329986 79614
rect 330222 79378 330306 79614
rect 330542 79378 330574 79614
rect 329954 79294 330574 79378
rect 329954 79058 329986 79294
rect 330222 79058 330306 79294
rect 330542 79058 330574 79294
rect 329954 43614 330574 79058
rect 329954 43378 329986 43614
rect 330222 43378 330306 43614
rect 330542 43378 330574 43614
rect 329954 43294 330574 43378
rect 329954 43058 329986 43294
rect 330222 43058 330306 43294
rect 330542 43058 330574 43294
rect 329954 7614 330574 43058
rect 329954 7378 329986 7614
rect 330222 7378 330306 7614
rect 330542 7378 330574 7614
rect 329954 7294 330574 7378
rect 329954 7058 329986 7294
rect 330222 7058 330306 7294
rect 330542 7058 330574 7294
rect 329954 -4186 330574 7058
rect 329954 -4422 329986 -4186
rect 330222 -4422 330306 -4186
rect 330542 -4422 330574 -4186
rect 329954 -4506 330574 -4422
rect 329954 -4742 329986 -4506
rect 330222 -4742 330306 -4506
rect 330542 -4742 330574 -4506
rect 329954 -7654 330574 -4742
rect 331194 709638 331814 711590
rect 331194 709402 331226 709638
rect 331462 709402 331546 709638
rect 331782 709402 331814 709638
rect 331194 709318 331814 709402
rect 331194 709082 331226 709318
rect 331462 709082 331546 709318
rect 331782 709082 331814 709318
rect 331194 692854 331814 709082
rect 331194 692618 331226 692854
rect 331462 692618 331546 692854
rect 331782 692618 331814 692854
rect 331194 692534 331814 692618
rect 331194 692298 331226 692534
rect 331462 692298 331546 692534
rect 331782 692298 331814 692534
rect 331194 656854 331814 692298
rect 331194 656618 331226 656854
rect 331462 656618 331546 656854
rect 331782 656618 331814 656854
rect 331194 656534 331814 656618
rect 331194 656298 331226 656534
rect 331462 656298 331546 656534
rect 331782 656298 331814 656534
rect 331194 620854 331814 656298
rect 331194 620618 331226 620854
rect 331462 620618 331546 620854
rect 331782 620618 331814 620854
rect 331194 620534 331814 620618
rect 331194 620298 331226 620534
rect 331462 620298 331546 620534
rect 331782 620298 331814 620534
rect 331194 584854 331814 620298
rect 331194 584618 331226 584854
rect 331462 584618 331546 584854
rect 331782 584618 331814 584854
rect 331194 584534 331814 584618
rect 331194 584298 331226 584534
rect 331462 584298 331546 584534
rect 331782 584298 331814 584534
rect 331194 548854 331814 584298
rect 331194 548618 331226 548854
rect 331462 548618 331546 548854
rect 331782 548618 331814 548854
rect 331194 548534 331814 548618
rect 331194 548298 331226 548534
rect 331462 548298 331546 548534
rect 331782 548298 331814 548534
rect 331194 512854 331814 548298
rect 331194 512618 331226 512854
rect 331462 512618 331546 512854
rect 331782 512618 331814 512854
rect 331194 512534 331814 512618
rect 331194 512298 331226 512534
rect 331462 512298 331546 512534
rect 331782 512298 331814 512534
rect 331194 476854 331814 512298
rect 331194 476618 331226 476854
rect 331462 476618 331546 476854
rect 331782 476618 331814 476854
rect 331194 476534 331814 476618
rect 331194 476298 331226 476534
rect 331462 476298 331546 476534
rect 331782 476298 331814 476534
rect 331194 440854 331814 476298
rect 331194 440618 331226 440854
rect 331462 440618 331546 440854
rect 331782 440618 331814 440854
rect 331194 440534 331814 440618
rect 331194 440298 331226 440534
rect 331462 440298 331546 440534
rect 331782 440298 331814 440534
rect 331194 404854 331814 440298
rect 331194 404618 331226 404854
rect 331462 404618 331546 404854
rect 331782 404618 331814 404854
rect 331194 404534 331814 404618
rect 331194 404298 331226 404534
rect 331462 404298 331546 404534
rect 331782 404298 331814 404534
rect 331194 368854 331814 404298
rect 331194 368618 331226 368854
rect 331462 368618 331546 368854
rect 331782 368618 331814 368854
rect 331194 368534 331814 368618
rect 331194 368298 331226 368534
rect 331462 368298 331546 368534
rect 331782 368298 331814 368534
rect 331194 332854 331814 368298
rect 331194 332618 331226 332854
rect 331462 332618 331546 332854
rect 331782 332618 331814 332854
rect 331194 332534 331814 332618
rect 331194 332298 331226 332534
rect 331462 332298 331546 332534
rect 331782 332298 331814 332534
rect 331194 296854 331814 332298
rect 331194 296618 331226 296854
rect 331462 296618 331546 296854
rect 331782 296618 331814 296854
rect 331194 296534 331814 296618
rect 331194 296298 331226 296534
rect 331462 296298 331546 296534
rect 331782 296298 331814 296534
rect 331194 260854 331814 296298
rect 331194 260618 331226 260854
rect 331462 260618 331546 260854
rect 331782 260618 331814 260854
rect 331194 260534 331814 260618
rect 331194 260298 331226 260534
rect 331462 260298 331546 260534
rect 331782 260298 331814 260534
rect 331194 224854 331814 260298
rect 331194 224618 331226 224854
rect 331462 224618 331546 224854
rect 331782 224618 331814 224854
rect 331194 224534 331814 224618
rect 331194 224298 331226 224534
rect 331462 224298 331546 224534
rect 331782 224298 331814 224534
rect 331194 188854 331814 224298
rect 331194 188618 331226 188854
rect 331462 188618 331546 188854
rect 331782 188618 331814 188854
rect 331194 188534 331814 188618
rect 331194 188298 331226 188534
rect 331462 188298 331546 188534
rect 331782 188298 331814 188534
rect 331194 152854 331814 188298
rect 331194 152618 331226 152854
rect 331462 152618 331546 152854
rect 331782 152618 331814 152854
rect 331194 152534 331814 152618
rect 331194 152298 331226 152534
rect 331462 152298 331546 152534
rect 331782 152298 331814 152534
rect 331194 116854 331814 152298
rect 331194 116618 331226 116854
rect 331462 116618 331546 116854
rect 331782 116618 331814 116854
rect 331194 116534 331814 116618
rect 331194 116298 331226 116534
rect 331462 116298 331546 116534
rect 331782 116298 331814 116534
rect 331194 80854 331814 116298
rect 331194 80618 331226 80854
rect 331462 80618 331546 80854
rect 331782 80618 331814 80854
rect 331194 80534 331814 80618
rect 331194 80298 331226 80534
rect 331462 80298 331546 80534
rect 331782 80298 331814 80534
rect 331194 44854 331814 80298
rect 331194 44618 331226 44854
rect 331462 44618 331546 44854
rect 331782 44618 331814 44854
rect 331194 44534 331814 44618
rect 331194 44298 331226 44534
rect 331462 44298 331546 44534
rect 331782 44298 331814 44534
rect 331194 8854 331814 44298
rect 331194 8618 331226 8854
rect 331462 8618 331546 8854
rect 331782 8618 331814 8854
rect 331194 8534 331814 8618
rect 331194 8298 331226 8534
rect 331462 8298 331546 8534
rect 331782 8298 331814 8534
rect 331194 -5146 331814 8298
rect 331194 -5382 331226 -5146
rect 331462 -5382 331546 -5146
rect 331782 -5382 331814 -5146
rect 331194 -5466 331814 -5382
rect 331194 -5702 331226 -5466
rect 331462 -5702 331546 -5466
rect 331782 -5702 331814 -5466
rect 331194 -7654 331814 -5702
rect 332434 710598 333054 711590
rect 332434 710362 332466 710598
rect 332702 710362 332786 710598
rect 333022 710362 333054 710598
rect 332434 710278 333054 710362
rect 332434 710042 332466 710278
rect 332702 710042 332786 710278
rect 333022 710042 333054 710278
rect 332434 694094 333054 710042
rect 332434 693858 332466 694094
rect 332702 693858 332786 694094
rect 333022 693858 333054 694094
rect 332434 693774 333054 693858
rect 332434 693538 332466 693774
rect 332702 693538 332786 693774
rect 333022 693538 333054 693774
rect 332434 658094 333054 693538
rect 332434 657858 332466 658094
rect 332702 657858 332786 658094
rect 333022 657858 333054 658094
rect 332434 657774 333054 657858
rect 332434 657538 332466 657774
rect 332702 657538 332786 657774
rect 333022 657538 333054 657774
rect 332434 622094 333054 657538
rect 332434 621858 332466 622094
rect 332702 621858 332786 622094
rect 333022 621858 333054 622094
rect 332434 621774 333054 621858
rect 332434 621538 332466 621774
rect 332702 621538 332786 621774
rect 333022 621538 333054 621774
rect 332434 586094 333054 621538
rect 332434 585858 332466 586094
rect 332702 585858 332786 586094
rect 333022 585858 333054 586094
rect 332434 585774 333054 585858
rect 332434 585538 332466 585774
rect 332702 585538 332786 585774
rect 333022 585538 333054 585774
rect 332434 550094 333054 585538
rect 332434 549858 332466 550094
rect 332702 549858 332786 550094
rect 333022 549858 333054 550094
rect 332434 549774 333054 549858
rect 332434 549538 332466 549774
rect 332702 549538 332786 549774
rect 333022 549538 333054 549774
rect 332434 514094 333054 549538
rect 332434 513858 332466 514094
rect 332702 513858 332786 514094
rect 333022 513858 333054 514094
rect 332434 513774 333054 513858
rect 332434 513538 332466 513774
rect 332702 513538 332786 513774
rect 333022 513538 333054 513774
rect 332434 478094 333054 513538
rect 332434 477858 332466 478094
rect 332702 477858 332786 478094
rect 333022 477858 333054 478094
rect 332434 477774 333054 477858
rect 332434 477538 332466 477774
rect 332702 477538 332786 477774
rect 333022 477538 333054 477774
rect 332434 442094 333054 477538
rect 332434 441858 332466 442094
rect 332702 441858 332786 442094
rect 333022 441858 333054 442094
rect 332434 441774 333054 441858
rect 332434 441538 332466 441774
rect 332702 441538 332786 441774
rect 333022 441538 333054 441774
rect 332434 406094 333054 441538
rect 332434 405858 332466 406094
rect 332702 405858 332786 406094
rect 333022 405858 333054 406094
rect 332434 405774 333054 405858
rect 332434 405538 332466 405774
rect 332702 405538 332786 405774
rect 333022 405538 333054 405774
rect 332434 370094 333054 405538
rect 332434 369858 332466 370094
rect 332702 369858 332786 370094
rect 333022 369858 333054 370094
rect 332434 369774 333054 369858
rect 332434 369538 332466 369774
rect 332702 369538 332786 369774
rect 333022 369538 333054 369774
rect 332434 334094 333054 369538
rect 332434 333858 332466 334094
rect 332702 333858 332786 334094
rect 333022 333858 333054 334094
rect 332434 333774 333054 333858
rect 332434 333538 332466 333774
rect 332702 333538 332786 333774
rect 333022 333538 333054 333774
rect 332434 298094 333054 333538
rect 332434 297858 332466 298094
rect 332702 297858 332786 298094
rect 333022 297858 333054 298094
rect 332434 297774 333054 297858
rect 332434 297538 332466 297774
rect 332702 297538 332786 297774
rect 333022 297538 333054 297774
rect 332434 262094 333054 297538
rect 332434 261858 332466 262094
rect 332702 261858 332786 262094
rect 333022 261858 333054 262094
rect 332434 261774 333054 261858
rect 332434 261538 332466 261774
rect 332702 261538 332786 261774
rect 333022 261538 333054 261774
rect 332434 226094 333054 261538
rect 332434 225858 332466 226094
rect 332702 225858 332786 226094
rect 333022 225858 333054 226094
rect 332434 225774 333054 225858
rect 332434 225538 332466 225774
rect 332702 225538 332786 225774
rect 333022 225538 333054 225774
rect 332434 190094 333054 225538
rect 332434 189858 332466 190094
rect 332702 189858 332786 190094
rect 333022 189858 333054 190094
rect 332434 189774 333054 189858
rect 332434 189538 332466 189774
rect 332702 189538 332786 189774
rect 333022 189538 333054 189774
rect 332434 154094 333054 189538
rect 332434 153858 332466 154094
rect 332702 153858 332786 154094
rect 333022 153858 333054 154094
rect 332434 153774 333054 153858
rect 332434 153538 332466 153774
rect 332702 153538 332786 153774
rect 333022 153538 333054 153774
rect 332434 118094 333054 153538
rect 332434 117858 332466 118094
rect 332702 117858 332786 118094
rect 333022 117858 333054 118094
rect 332434 117774 333054 117858
rect 332434 117538 332466 117774
rect 332702 117538 332786 117774
rect 333022 117538 333054 117774
rect 332434 82094 333054 117538
rect 332434 81858 332466 82094
rect 332702 81858 332786 82094
rect 333022 81858 333054 82094
rect 332434 81774 333054 81858
rect 332434 81538 332466 81774
rect 332702 81538 332786 81774
rect 333022 81538 333054 81774
rect 332434 46094 333054 81538
rect 332434 45858 332466 46094
rect 332702 45858 332786 46094
rect 333022 45858 333054 46094
rect 332434 45774 333054 45858
rect 332434 45538 332466 45774
rect 332702 45538 332786 45774
rect 333022 45538 333054 45774
rect 332434 10094 333054 45538
rect 332434 9858 332466 10094
rect 332702 9858 332786 10094
rect 333022 9858 333054 10094
rect 332434 9774 333054 9858
rect 332434 9538 332466 9774
rect 332702 9538 332786 9774
rect 333022 9538 333054 9774
rect 332434 -6106 333054 9538
rect 332434 -6342 332466 -6106
rect 332702 -6342 332786 -6106
rect 333022 -6342 333054 -6106
rect 332434 -6426 333054 -6342
rect 332434 -6662 332466 -6426
rect 332702 -6662 332786 -6426
rect 333022 -6662 333054 -6426
rect 332434 -7654 333054 -6662
rect 333674 711558 334294 711590
rect 333674 711322 333706 711558
rect 333942 711322 334026 711558
rect 334262 711322 334294 711558
rect 333674 711238 334294 711322
rect 333674 711002 333706 711238
rect 333942 711002 334026 711238
rect 334262 711002 334294 711238
rect 333674 695334 334294 711002
rect 333674 695098 333706 695334
rect 333942 695098 334026 695334
rect 334262 695098 334294 695334
rect 333674 695014 334294 695098
rect 333674 694778 333706 695014
rect 333942 694778 334026 695014
rect 334262 694778 334294 695014
rect 333674 659334 334294 694778
rect 333674 659098 333706 659334
rect 333942 659098 334026 659334
rect 334262 659098 334294 659334
rect 333674 659014 334294 659098
rect 333674 658778 333706 659014
rect 333942 658778 334026 659014
rect 334262 658778 334294 659014
rect 333674 623334 334294 658778
rect 333674 623098 333706 623334
rect 333942 623098 334026 623334
rect 334262 623098 334294 623334
rect 333674 623014 334294 623098
rect 333674 622778 333706 623014
rect 333942 622778 334026 623014
rect 334262 622778 334294 623014
rect 333674 587334 334294 622778
rect 333674 587098 333706 587334
rect 333942 587098 334026 587334
rect 334262 587098 334294 587334
rect 333674 587014 334294 587098
rect 333674 586778 333706 587014
rect 333942 586778 334026 587014
rect 334262 586778 334294 587014
rect 333674 551334 334294 586778
rect 333674 551098 333706 551334
rect 333942 551098 334026 551334
rect 334262 551098 334294 551334
rect 333674 551014 334294 551098
rect 333674 550778 333706 551014
rect 333942 550778 334026 551014
rect 334262 550778 334294 551014
rect 333674 515334 334294 550778
rect 333674 515098 333706 515334
rect 333942 515098 334026 515334
rect 334262 515098 334294 515334
rect 333674 515014 334294 515098
rect 333674 514778 333706 515014
rect 333942 514778 334026 515014
rect 334262 514778 334294 515014
rect 333674 479334 334294 514778
rect 333674 479098 333706 479334
rect 333942 479098 334026 479334
rect 334262 479098 334294 479334
rect 333674 479014 334294 479098
rect 333674 478778 333706 479014
rect 333942 478778 334026 479014
rect 334262 478778 334294 479014
rect 333674 443334 334294 478778
rect 333674 443098 333706 443334
rect 333942 443098 334026 443334
rect 334262 443098 334294 443334
rect 333674 443014 334294 443098
rect 333674 442778 333706 443014
rect 333942 442778 334026 443014
rect 334262 442778 334294 443014
rect 333674 407334 334294 442778
rect 333674 407098 333706 407334
rect 333942 407098 334026 407334
rect 334262 407098 334294 407334
rect 333674 407014 334294 407098
rect 333674 406778 333706 407014
rect 333942 406778 334026 407014
rect 334262 406778 334294 407014
rect 333674 371334 334294 406778
rect 333674 371098 333706 371334
rect 333942 371098 334026 371334
rect 334262 371098 334294 371334
rect 333674 371014 334294 371098
rect 333674 370778 333706 371014
rect 333942 370778 334026 371014
rect 334262 370778 334294 371014
rect 333674 335334 334294 370778
rect 333674 335098 333706 335334
rect 333942 335098 334026 335334
rect 334262 335098 334294 335334
rect 333674 335014 334294 335098
rect 333674 334778 333706 335014
rect 333942 334778 334026 335014
rect 334262 334778 334294 335014
rect 333674 299334 334294 334778
rect 333674 299098 333706 299334
rect 333942 299098 334026 299334
rect 334262 299098 334294 299334
rect 333674 299014 334294 299098
rect 333674 298778 333706 299014
rect 333942 298778 334026 299014
rect 334262 298778 334294 299014
rect 333674 263334 334294 298778
rect 333674 263098 333706 263334
rect 333942 263098 334026 263334
rect 334262 263098 334294 263334
rect 333674 263014 334294 263098
rect 333674 262778 333706 263014
rect 333942 262778 334026 263014
rect 334262 262778 334294 263014
rect 333674 227334 334294 262778
rect 333674 227098 333706 227334
rect 333942 227098 334026 227334
rect 334262 227098 334294 227334
rect 333674 227014 334294 227098
rect 333674 226778 333706 227014
rect 333942 226778 334026 227014
rect 334262 226778 334294 227014
rect 333674 191334 334294 226778
rect 333674 191098 333706 191334
rect 333942 191098 334026 191334
rect 334262 191098 334294 191334
rect 333674 191014 334294 191098
rect 333674 190778 333706 191014
rect 333942 190778 334026 191014
rect 334262 190778 334294 191014
rect 333674 155334 334294 190778
rect 333674 155098 333706 155334
rect 333942 155098 334026 155334
rect 334262 155098 334294 155334
rect 333674 155014 334294 155098
rect 333674 154778 333706 155014
rect 333942 154778 334026 155014
rect 334262 154778 334294 155014
rect 333674 119334 334294 154778
rect 333674 119098 333706 119334
rect 333942 119098 334026 119334
rect 334262 119098 334294 119334
rect 333674 119014 334294 119098
rect 333674 118778 333706 119014
rect 333942 118778 334026 119014
rect 334262 118778 334294 119014
rect 333674 83334 334294 118778
rect 333674 83098 333706 83334
rect 333942 83098 334026 83334
rect 334262 83098 334294 83334
rect 333674 83014 334294 83098
rect 333674 82778 333706 83014
rect 333942 82778 334026 83014
rect 334262 82778 334294 83014
rect 333674 47334 334294 82778
rect 333674 47098 333706 47334
rect 333942 47098 334026 47334
rect 334262 47098 334294 47334
rect 333674 47014 334294 47098
rect 333674 46778 333706 47014
rect 333942 46778 334026 47014
rect 334262 46778 334294 47014
rect 333674 11334 334294 46778
rect 333674 11098 333706 11334
rect 333942 11098 334026 11334
rect 334262 11098 334294 11334
rect 333674 11014 334294 11098
rect 333674 10778 333706 11014
rect 333942 10778 334026 11014
rect 334262 10778 334294 11014
rect 333674 -7066 334294 10778
rect 333674 -7302 333706 -7066
rect 333942 -7302 334026 -7066
rect 334262 -7302 334294 -7066
rect 333674 -7386 334294 -7302
rect 333674 -7622 333706 -7386
rect 333942 -7622 334026 -7386
rect 334262 -7622 334294 -7386
rect 333674 -7654 334294 -7622
rect 360994 704838 361614 711590
rect 360994 704602 361026 704838
rect 361262 704602 361346 704838
rect 361582 704602 361614 704838
rect 360994 704518 361614 704602
rect 360994 704282 361026 704518
rect 361262 704282 361346 704518
rect 361582 704282 361614 704518
rect 360994 686654 361614 704282
rect 360994 686418 361026 686654
rect 361262 686418 361346 686654
rect 361582 686418 361614 686654
rect 360994 686334 361614 686418
rect 360994 686098 361026 686334
rect 361262 686098 361346 686334
rect 361582 686098 361614 686334
rect 360994 650654 361614 686098
rect 360994 650418 361026 650654
rect 361262 650418 361346 650654
rect 361582 650418 361614 650654
rect 360994 650334 361614 650418
rect 360994 650098 361026 650334
rect 361262 650098 361346 650334
rect 361582 650098 361614 650334
rect 360994 614654 361614 650098
rect 360994 614418 361026 614654
rect 361262 614418 361346 614654
rect 361582 614418 361614 614654
rect 360994 614334 361614 614418
rect 360994 614098 361026 614334
rect 361262 614098 361346 614334
rect 361582 614098 361614 614334
rect 360994 578654 361614 614098
rect 360994 578418 361026 578654
rect 361262 578418 361346 578654
rect 361582 578418 361614 578654
rect 360994 578334 361614 578418
rect 360994 578098 361026 578334
rect 361262 578098 361346 578334
rect 361582 578098 361614 578334
rect 360994 542654 361614 578098
rect 360994 542418 361026 542654
rect 361262 542418 361346 542654
rect 361582 542418 361614 542654
rect 360994 542334 361614 542418
rect 360994 542098 361026 542334
rect 361262 542098 361346 542334
rect 361582 542098 361614 542334
rect 360994 506654 361614 542098
rect 360994 506418 361026 506654
rect 361262 506418 361346 506654
rect 361582 506418 361614 506654
rect 360994 506334 361614 506418
rect 360994 506098 361026 506334
rect 361262 506098 361346 506334
rect 361582 506098 361614 506334
rect 360994 470654 361614 506098
rect 360994 470418 361026 470654
rect 361262 470418 361346 470654
rect 361582 470418 361614 470654
rect 360994 470334 361614 470418
rect 360994 470098 361026 470334
rect 361262 470098 361346 470334
rect 361582 470098 361614 470334
rect 360994 434654 361614 470098
rect 360994 434418 361026 434654
rect 361262 434418 361346 434654
rect 361582 434418 361614 434654
rect 360994 434334 361614 434418
rect 360994 434098 361026 434334
rect 361262 434098 361346 434334
rect 361582 434098 361614 434334
rect 360994 398654 361614 434098
rect 360994 398418 361026 398654
rect 361262 398418 361346 398654
rect 361582 398418 361614 398654
rect 360994 398334 361614 398418
rect 360994 398098 361026 398334
rect 361262 398098 361346 398334
rect 361582 398098 361614 398334
rect 360994 362654 361614 398098
rect 360994 362418 361026 362654
rect 361262 362418 361346 362654
rect 361582 362418 361614 362654
rect 360994 362334 361614 362418
rect 360994 362098 361026 362334
rect 361262 362098 361346 362334
rect 361582 362098 361614 362334
rect 360994 326654 361614 362098
rect 360994 326418 361026 326654
rect 361262 326418 361346 326654
rect 361582 326418 361614 326654
rect 360994 326334 361614 326418
rect 360994 326098 361026 326334
rect 361262 326098 361346 326334
rect 361582 326098 361614 326334
rect 360994 290654 361614 326098
rect 360994 290418 361026 290654
rect 361262 290418 361346 290654
rect 361582 290418 361614 290654
rect 360994 290334 361614 290418
rect 360994 290098 361026 290334
rect 361262 290098 361346 290334
rect 361582 290098 361614 290334
rect 360994 254654 361614 290098
rect 360994 254418 361026 254654
rect 361262 254418 361346 254654
rect 361582 254418 361614 254654
rect 360994 254334 361614 254418
rect 360994 254098 361026 254334
rect 361262 254098 361346 254334
rect 361582 254098 361614 254334
rect 360994 218654 361614 254098
rect 360994 218418 361026 218654
rect 361262 218418 361346 218654
rect 361582 218418 361614 218654
rect 360994 218334 361614 218418
rect 360994 218098 361026 218334
rect 361262 218098 361346 218334
rect 361582 218098 361614 218334
rect 360994 182654 361614 218098
rect 360994 182418 361026 182654
rect 361262 182418 361346 182654
rect 361582 182418 361614 182654
rect 360994 182334 361614 182418
rect 360994 182098 361026 182334
rect 361262 182098 361346 182334
rect 361582 182098 361614 182334
rect 360994 146654 361614 182098
rect 360994 146418 361026 146654
rect 361262 146418 361346 146654
rect 361582 146418 361614 146654
rect 360994 146334 361614 146418
rect 360994 146098 361026 146334
rect 361262 146098 361346 146334
rect 361582 146098 361614 146334
rect 360994 110654 361614 146098
rect 360994 110418 361026 110654
rect 361262 110418 361346 110654
rect 361582 110418 361614 110654
rect 360994 110334 361614 110418
rect 360994 110098 361026 110334
rect 361262 110098 361346 110334
rect 361582 110098 361614 110334
rect 360994 74654 361614 110098
rect 360994 74418 361026 74654
rect 361262 74418 361346 74654
rect 361582 74418 361614 74654
rect 360994 74334 361614 74418
rect 360994 74098 361026 74334
rect 361262 74098 361346 74334
rect 361582 74098 361614 74334
rect 360994 38654 361614 74098
rect 360994 38418 361026 38654
rect 361262 38418 361346 38654
rect 361582 38418 361614 38654
rect 360994 38334 361614 38418
rect 360994 38098 361026 38334
rect 361262 38098 361346 38334
rect 361582 38098 361614 38334
rect 360994 2654 361614 38098
rect 360994 2418 361026 2654
rect 361262 2418 361346 2654
rect 361582 2418 361614 2654
rect 360994 2334 361614 2418
rect 360994 2098 361026 2334
rect 361262 2098 361346 2334
rect 361582 2098 361614 2334
rect 360994 -346 361614 2098
rect 360994 -582 361026 -346
rect 361262 -582 361346 -346
rect 361582 -582 361614 -346
rect 360994 -666 361614 -582
rect 360994 -902 361026 -666
rect 361262 -902 361346 -666
rect 361582 -902 361614 -666
rect 360994 -7654 361614 -902
rect 362234 705798 362854 711590
rect 362234 705562 362266 705798
rect 362502 705562 362586 705798
rect 362822 705562 362854 705798
rect 362234 705478 362854 705562
rect 362234 705242 362266 705478
rect 362502 705242 362586 705478
rect 362822 705242 362854 705478
rect 362234 687894 362854 705242
rect 362234 687658 362266 687894
rect 362502 687658 362586 687894
rect 362822 687658 362854 687894
rect 362234 687574 362854 687658
rect 362234 687338 362266 687574
rect 362502 687338 362586 687574
rect 362822 687338 362854 687574
rect 362234 651894 362854 687338
rect 362234 651658 362266 651894
rect 362502 651658 362586 651894
rect 362822 651658 362854 651894
rect 362234 651574 362854 651658
rect 362234 651338 362266 651574
rect 362502 651338 362586 651574
rect 362822 651338 362854 651574
rect 362234 615894 362854 651338
rect 362234 615658 362266 615894
rect 362502 615658 362586 615894
rect 362822 615658 362854 615894
rect 362234 615574 362854 615658
rect 362234 615338 362266 615574
rect 362502 615338 362586 615574
rect 362822 615338 362854 615574
rect 362234 579894 362854 615338
rect 362234 579658 362266 579894
rect 362502 579658 362586 579894
rect 362822 579658 362854 579894
rect 362234 579574 362854 579658
rect 362234 579338 362266 579574
rect 362502 579338 362586 579574
rect 362822 579338 362854 579574
rect 362234 543894 362854 579338
rect 362234 543658 362266 543894
rect 362502 543658 362586 543894
rect 362822 543658 362854 543894
rect 362234 543574 362854 543658
rect 362234 543338 362266 543574
rect 362502 543338 362586 543574
rect 362822 543338 362854 543574
rect 362234 507894 362854 543338
rect 362234 507658 362266 507894
rect 362502 507658 362586 507894
rect 362822 507658 362854 507894
rect 362234 507574 362854 507658
rect 362234 507338 362266 507574
rect 362502 507338 362586 507574
rect 362822 507338 362854 507574
rect 362234 471894 362854 507338
rect 362234 471658 362266 471894
rect 362502 471658 362586 471894
rect 362822 471658 362854 471894
rect 362234 471574 362854 471658
rect 362234 471338 362266 471574
rect 362502 471338 362586 471574
rect 362822 471338 362854 471574
rect 362234 435894 362854 471338
rect 362234 435658 362266 435894
rect 362502 435658 362586 435894
rect 362822 435658 362854 435894
rect 362234 435574 362854 435658
rect 362234 435338 362266 435574
rect 362502 435338 362586 435574
rect 362822 435338 362854 435574
rect 362234 399894 362854 435338
rect 362234 399658 362266 399894
rect 362502 399658 362586 399894
rect 362822 399658 362854 399894
rect 362234 399574 362854 399658
rect 362234 399338 362266 399574
rect 362502 399338 362586 399574
rect 362822 399338 362854 399574
rect 362234 363894 362854 399338
rect 362234 363658 362266 363894
rect 362502 363658 362586 363894
rect 362822 363658 362854 363894
rect 362234 363574 362854 363658
rect 362234 363338 362266 363574
rect 362502 363338 362586 363574
rect 362822 363338 362854 363574
rect 362234 327894 362854 363338
rect 362234 327658 362266 327894
rect 362502 327658 362586 327894
rect 362822 327658 362854 327894
rect 362234 327574 362854 327658
rect 362234 327338 362266 327574
rect 362502 327338 362586 327574
rect 362822 327338 362854 327574
rect 362234 291894 362854 327338
rect 362234 291658 362266 291894
rect 362502 291658 362586 291894
rect 362822 291658 362854 291894
rect 362234 291574 362854 291658
rect 362234 291338 362266 291574
rect 362502 291338 362586 291574
rect 362822 291338 362854 291574
rect 362234 255894 362854 291338
rect 362234 255658 362266 255894
rect 362502 255658 362586 255894
rect 362822 255658 362854 255894
rect 362234 255574 362854 255658
rect 362234 255338 362266 255574
rect 362502 255338 362586 255574
rect 362822 255338 362854 255574
rect 362234 219894 362854 255338
rect 362234 219658 362266 219894
rect 362502 219658 362586 219894
rect 362822 219658 362854 219894
rect 362234 219574 362854 219658
rect 362234 219338 362266 219574
rect 362502 219338 362586 219574
rect 362822 219338 362854 219574
rect 362234 183894 362854 219338
rect 362234 183658 362266 183894
rect 362502 183658 362586 183894
rect 362822 183658 362854 183894
rect 362234 183574 362854 183658
rect 362234 183338 362266 183574
rect 362502 183338 362586 183574
rect 362822 183338 362854 183574
rect 362234 147894 362854 183338
rect 362234 147658 362266 147894
rect 362502 147658 362586 147894
rect 362822 147658 362854 147894
rect 362234 147574 362854 147658
rect 362234 147338 362266 147574
rect 362502 147338 362586 147574
rect 362822 147338 362854 147574
rect 362234 111894 362854 147338
rect 362234 111658 362266 111894
rect 362502 111658 362586 111894
rect 362822 111658 362854 111894
rect 362234 111574 362854 111658
rect 362234 111338 362266 111574
rect 362502 111338 362586 111574
rect 362822 111338 362854 111574
rect 362234 75894 362854 111338
rect 362234 75658 362266 75894
rect 362502 75658 362586 75894
rect 362822 75658 362854 75894
rect 362234 75574 362854 75658
rect 362234 75338 362266 75574
rect 362502 75338 362586 75574
rect 362822 75338 362854 75574
rect 362234 39894 362854 75338
rect 362234 39658 362266 39894
rect 362502 39658 362586 39894
rect 362822 39658 362854 39894
rect 362234 39574 362854 39658
rect 362234 39338 362266 39574
rect 362502 39338 362586 39574
rect 362822 39338 362854 39574
rect 362234 3894 362854 39338
rect 362234 3658 362266 3894
rect 362502 3658 362586 3894
rect 362822 3658 362854 3894
rect 362234 3574 362854 3658
rect 362234 3338 362266 3574
rect 362502 3338 362586 3574
rect 362822 3338 362854 3574
rect 362234 -1306 362854 3338
rect 362234 -1542 362266 -1306
rect 362502 -1542 362586 -1306
rect 362822 -1542 362854 -1306
rect 362234 -1626 362854 -1542
rect 362234 -1862 362266 -1626
rect 362502 -1862 362586 -1626
rect 362822 -1862 362854 -1626
rect 362234 -7654 362854 -1862
rect 363474 706758 364094 711590
rect 363474 706522 363506 706758
rect 363742 706522 363826 706758
rect 364062 706522 364094 706758
rect 363474 706438 364094 706522
rect 363474 706202 363506 706438
rect 363742 706202 363826 706438
rect 364062 706202 364094 706438
rect 363474 689134 364094 706202
rect 363474 688898 363506 689134
rect 363742 688898 363826 689134
rect 364062 688898 364094 689134
rect 363474 688814 364094 688898
rect 363474 688578 363506 688814
rect 363742 688578 363826 688814
rect 364062 688578 364094 688814
rect 363474 653134 364094 688578
rect 363474 652898 363506 653134
rect 363742 652898 363826 653134
rect 364062 652898 364094 653134
rect 363474 652814 364094 652898
rect 363474 652578 363506 652814
rect 363742 652578 363826 652814
rect 364062 652578 364094 652814
rect 363474 617134 364094 652578
rect 363474 616898 363506 617134
rect 363742 616898 363826 617134
rect 364062 616898 364094 617134
rect 363474 616814 364094 616898
rect 363474 616578 363506 616814
rect 363742 616578 363826 616814
rect 364062 616578 364094 616814
rect 363474 581134 364094 616578
rect 363474 580898 363506 581134
rect 363742 580898 363826 581134
rect 364062 580898 364094 581134
rect 363474 580814 364094 580898
rect 363474 580578 363506 580814
rect 363742 580578 363826 580814
rect 364062 580578 364094 580814
rect 363474 545134 364094 580578
rect 363474 544898 363506 545134
rect 363742 544898 363826 545134
rect 364062 544898 364094 545134
rect 363474 544814 364094 544898
rect 363474 544578 363506 544814
rect 363742 544578 363826 544814
rect 364062 544578 364094 544814
rect 363474 509134 364094 544578
rect 363474 508898 363506 509134
rect 363742 508898 363826 509134
rect 364062 508898 364094 509134
rect 363474 508814 364094 508898
rect 363474 508578 363506 508814
rect 363742 508578 363826 508814
rect 364062 508578 364094 508814
rect 363474 473134 364094 508578
rect 363474 472898 363506 473134
rect 363742 472898 363826 473134
rect 364062 472898 364094 473134
rect 363474 472814 364094 472898
rect 363474 472578 363506 472814
rect 363742 472578 363826 472814
rect 364062 472578 364094 472814
rect 363474 437134 364094 472578
rect 363474 436898 363506 437134
rect 363742 436898 363826 437134
rect 364062 436898 364094 437134
rect 363474 436814 364094 436898
rect 363474 436578 363506 436814
rect 363742 436578 363826 436814
rect 364062 436578 364094 436814
rect 363474 401134 364094 436578
rect 363474 400898 363506 401134
rect 363742 400898 363826 401134
rect 364062 400898 364094 401134
rect 363474 400814 364094 400898
rect 363474 400578 363506 400814
rect 363742 400578 363826 400814
rect 364062 400578 364094 400814
rect 363474 365134 364094 400578
rect 363474 364898 363506 365134
rect 363742 364898 363826 365134
rect 364062 364898 364094 365134
rect 363474 364814 364094 364898
rect 363474 364578 363506 364814
rect 363742 364578 363826 364814
rect 364062 364578 364094 364814
rect 363474 329134 364094 364578
rect 363474 328898 363506 329134
rect 363742 328898 363826 329134
rect 364062 328898 364094 329134
rect 363474 328814 364094 328898
rect 363474 328578 363506 328814
rect 363742 328578 363826 328814
rect 364062 328578 364094 328814
rect 363474 293134 364094 328578
rect 363474 292898 363506 293134
rect 363742 292898 363826 293134
rect 364062 292898 364094 293134
rect 363474 292814 364094 292898
rect 363474 292578 363506 292814
rect 363742 292578 363826 292814
rect 364062 292578 364094 292814
rect 363474 257134 364094 292578
rect 363474 256898 363506 257134
rect 363742 256898 363826 257134
rect 364062 256898 364094 257134
rect 363474 256814 364094 256898
rect 363474 256578 363506 256814
rect 363742 256578 363826 256814
rect 364062 256578 364094 256814
rect 363474 221134 364094 256578
rect 363474 220898 363506 221134
rect 363742 220898 363826 221134
rect 364062 220898 364094 221134
rect 363474 220814 364094 220898
rect 363474 220578 363506 220814
rect 363742 220578 363826 220814
rect 364062 220578 364094 220814
rect 363474 185134 364094 220578
rect 363474 184898 363506 185134
rect 363742 184898 363826 185134
rect 364062 184898 364094 185134
rect 363474 184814 364094 184898
rect 363474 184578 363506 184814
rect 363742 184578 363826 184814
rect 364062 184578 364094 184814
rect 363474 149134 364094 184578
rect 363474 148898 363506 149134
rect 363742 148898 363826 149134
rect 364062 148898 364094 149134
rect 363474 148814 364094 148898
rect 363474 148578 363506 148814
rect 363742 148578 363826 148814
rect 364062 148578 364094 148814
rect 363474 113134 364094 148578
rect 363474 112898 363506 113134
rect 363742 112898 363826 113134
rect 364062 112898 364094 113134
rect 363474 112814 364094 112898
rect 363474 112578 363506 112814
rect 363742 112578 363826 112814
rect 364062 112578 364094 112814
rect 363474 77134 364094 112578
rect 363474 76898 363506 77134
rect 363742 76898 363826 77134
rect 364062 76898 364094 77134
rect 363474 76814 364094 76898
rect 363474 76578 363506 76814
rect 363742 76578 363826 76814
rect 364062 76578 364094 76814
rect 363474 41134 364094 76578
rect 363474 40898 363506 41134
rect 363742 40898 363826 41134
rect 364062 40898 364094 41134
rect 363474 40814 364094 40898
rect 363474 40578 363506 40814
rect 363742 40578 363826 40814
rect 364062 40578 364094 40814
rect 363474 5134 364094 40578
rect 363474 4898 363506 5134
rect 363742 4898 363826 5134
rect 364062 4898 364094 5134
rect 363474 4814 364094 4898
rect 363474 4578 363506 4814
rect 363742 4578 363826 4814
rect 364062 4578 364094 4814
rect 363474 -2266 364094 4578
rect 363474 -2502 363506 -2266
rect 363742 -2502 363826 -2266
rect 364062 -2502 364094 -2266
rect 363474 -2586 364094 -2502
rect 363474 -2822 363506 -2586
rect 363742 -2822 363826 -2586
rect 364062 -2822 364094 -2586
rect 363474 -7654 364094 -2822
rect 364714 707718 365334 711590
rect 364714 707482 364746 707718
rect 364982 707482 365066 707718
rect 365302 707482 365334 707718
rect 364714 707398 365334 707482
rect 364714 707162 364746 707398
rect 364982 707162 365066 707398
rect 365302 707162 365334 707398
rect 364714 690374 365334 707162
rect 364714 690138 364746 690374
rect 364982 690138 365066 690374
rect 365302 690138 365334 690374
rect 364714 690054 365334 690138
rect 364714 689818 364746 690054
rect 364982 689818 365066 690054
rect 365302 689818 365334 690054
rect 364714 654374 365334 689818
rect 364714 654138 364746 654374
rect 364982 654138 365066 654374
rect 365302 654138 365334 654374
rect 364714 654054 365334 654138
rect 364714 653818 364746 654054
rect 364982 653818 365066 654054
rect 365302 653818 365334 654054
rect 364714 618374 365334 653818
rect 364714 618138 364746 618374
rect 364982 618138 365066 618374
rect 365302 618138 365334 618374
rect 364714 618054 365334 618138
rect 364714 617818 364746 618054
rect 364982 617818 365066 618054
rect 365302 617818 365334 618054
rect 364714 582374 365334 617818
rect 364714 582138 364746 582374
rect 364982 582138 365066 582374
rect 365302 582138 365334 582374
rect 364714 582054 365334 582138
rect 364714 581818 364746 582054
rect 364982 581818 365066 582054
rect 365302 581818 365334 582054
rect 364714 546374 365334 581818
rect 364714 546138 364746 546374
rect 364982 546138 365066 546374
rect 365302 546138 365334 546374
rect 364714 546054 365334 546138
rect 364714 545818 364746 546054
rect 364982 545818 365066 546054
rect 365302 545818 365334 546054
rect 364714 510374 365334 545818
rect 364714 510138 364746 510374
rect 364982 510138 365066 510374
rect 365302 510138 365334 510374
rect 364714 510054 365334 510138
rect 364714 509818 364746 510054
rect 364982 509818 365066 510054
rect 365302 509818 365334 510054
rect 364714 474374 365334 509818
rect 364714 474138 364746 474374
rect 364982 474138 365066 474374
rect 365302 474138 365334 474374
rect 364714 474054 365334 474138
rect 364714 473818 364746 474054
rect 364982 473818 365066 474054
rect 365302 473818 365334 474054
rect 364714 438374 365334 473818
rect 364714 438138 364746 438374
rect 364982 438138 365066 438374
rect 365302 438138 365334 438374
rect 364714 438054 365334 438138
rect 364714 437818 364746 438054
rect 364982 437818 365066 438054
rect 365302 437818 365334 438054
rect 364714 402374 365334 437818
rect 364714 402138 364746 402374
rect 364982 402138 365066 402374
rect 365302 402138 365334 402374
rect 364714 402054 365334 402138
rect 364714 401818 364746 402054
rect 364982 401818 365066 402054
rect 365302 401818 365334 402054
rect 364714 366374 365334 401818
rect 364714 366138 364746 366374
rect 364982 366138 365066 366374
rect 365302 366138 365334 366374
rect 364714 366054 365334 366138
rect 364714 365818 364746 366054
rect 364982 365818 365066 366054
rect 365302 365818 365334 366054
rect 364714 330374 365334 365818
rect 364714 330138 364746 330374
rect 364982 330138 365066 330374
rect 365302 330138 365334 330374
rect 364714 330054 365334 330138
rect 364714 329818 364746 330054
rect 364982 329818 365066 330054
rect 365302 329818 365334 330054
rect 364714 294374 365334 329818
rect 364714 294138 364746 294374
rect 364982 294138 365066 294374
rect 365302 294138 365334 294374
rect 364714 294054 365334 294138
rect 364714 293818 364746 294054
rect 364982 293818 365066 294054
rect 365302 293818 365334 294054
rect 364714 258374 365334 293818
rect 364714 258138 364746 258374
rect 364982 258138 365066 258374
rect 365302 258138 365334 258374
rect 364714 258054 365334 258138
rect 364714 257818 364746 258054
rect 364982 257818 365066 258054
rect 365302 257818 365334 258054
rect 364714 222374 365334 257818
rect 364714 222138 364746 222374
rect 364982 222138 365066 222374
rect 365302 222138 365334 222374
rect 364714 222054 365334 222138
rect 364714 221818 364746 222054
rect 364982 221818 365066 222054
rect 365302 221818 365334 222054
rect 364714 186374 365334 221818
rect 364714 186138 364746 186374
rect 364982 186138 365066 186374
rect 365302 186138 365334 186374
rect 364714 186054 365334 186138
rect 364714 185818 364746 186054
rect 364982 185818 365066 186054
rect 365302 185818 365334 186054
rect 364714 150374 365334 185818
rect 364714 150138 364746 150374
rect 364982 150138 365066 150374
rect 365302 150138 365334 150374
rect 364714 150054 365334 150138
rect 364714 149818 364746 150054
rect 364982 149818 365066 150054
rect 365302 149818 365334 150054
rect 364714 114374 365334 149818
rect 364714 114138 364746 114374
rect 364982 114138 365066 114374
rect 365302 114138 365334 114374
rect 364714 114054 365334 114138
rect 364714 113818 364746 114054
rect 364982 113818 365066 114054
rect 365302 113818 365334 114054
rect 364714 78374 365334 113818
rect 364714 78138 364746 78374
rect 364982 78138 365066 78374
rect 365302 78138 365334 78374
rect 364714 78054 365334 78138
rect 364714 77818 364746 78054
rect 364982 77818 365066 78054
rect 365302 77818 365334 78054
rect 364714 42374 365334 77818
rect 364714 42138 364746 42374
rect 364982 42138 365066 42374
rect 365302 42138 365334 42374
rect 364714 42054 365334 42138
rect 364714 41818 364746 42054
rect 364982 41818 365066 42054
rect 365302 41818 365334 42054
rect 364714 6374 365334 41818
rect 364714 6138 364746 6374
rect 364982 6138 365066 6374
rect 365302 6138 365334 6374
rect 364714 6054 365334 6138
rect 364714 5818 364746 6054
rect 364982 5818 365066 6054
rect 365302 5818 365334 6054
rect 364714 -3226 365334 5818
rect 364714 -3462 364746 -3226
rect 364982 -3462 365066 -3226
rect 365302 -3462 365334 -3226
rect 364714 -3546 365334 -3462
rect 364714 -3782 364746 -3546
rect 364982 -3782 365066 -3546
rect 365302 -3782 365334 -3546
rect 364714 -7654 365334 -3782
rect 365954 708678 366574 711590
rect 365954 708442 365986 708678
rect 366222 708442 366306 708678
rect 366542 708442 366574 708678
rect 365954 708358 366574 708442
rect 365954 708122 365986 708358
rect 366222 708122 366306 708358
rect 366542 708122 366574 708358
rect 365954 691614 366574 708122
rect 365954 691378 365986 691614
rect 366222 691378 366306 691614
rect 366542 691378 366574 691614
rect 365954 691294 366574 691378
rect 365954 691058 365986 691294
rect 366222 691058 366306 691294
rect 366542 691058 366574 691294
rect 365954 655614 366574 691058
rect 365954 655378 365986 655614
rect 366222 655378 366306 655614
rect 366542 655378 366574 655614
rect 365954 655294 366574 655378
rect 365954 655058 365986 655294
rect 366222 655058 366306 655294
rect 366542 655058 366574 655294
rect 365954 619614 366574 655058
rect 365954 619378 365986 619614
rect 366222 619378 366306 619614
rect 366542 619378 366574 619614
rect 365954 619294 366574 619378
rect 365954 619058 365986 619294
rect 366222 619058 366306 619294
rect 366542 619058 366574 619294
rect 365954 583614 366574 619058
rect 365954 583378 365986 583614
rect 366222 583378 366306 583614
rect 366542 583378 366574 583614
rect 365954 583294 366574 583378
rect 365954 583058 365986 583294
rect 366222 583058 366306 583294
rect 366542 583058 366574 583294
rect 365954 547614 366574 583058
rect 365954 547378 365986 547614
rect 366222 547378 366306 547614
rect 366542 547378 366574 547614
rect 365954 547294 366574 547378
rect 365954 547058 365986 547294
rect 366222 547058 366306 547294
rect 366542 547058 366574 547294
rect 365954 511614 366574 547058
rect 365954 511378 365986 511614
rect 366222 511378 366306 511614
rect 366542 511378 366574 511614
rect 365954 511294 366574 511378
rect 365954 511058 365986 511294
rect 366222 511058 366306 511294
rect 366542 511058 366574 511294
rect 365954 475614 366574 511058
rect 365954 475378 365986 475614
rect 366222 475378 366306 475614
rect 366542 475378 366574 475614
rect 365954 475294 366574 475378
rect 365954 475058 365986 475294
rect 366222 475058 366306 475294
rect 366542 475058 366574 475294
rect 365954 439614 366574 475058
rect 365954 439378 365986 439614
rect 366222 439378 366306 439614
rect 366542 439378 366574 439614
rect 365954 439294 366574 439378
rect 365954 439058 365986 439294
rect 366222 439058 366306 439294
rect 366542 439058 366574 439294
rect 365954 403614 366574 439058
rect 365954 403378 365986 403614
rect 366222 403378 366306 403614
rect 366542 403378 366574 403614
rect 365954 403294 366574 403378
rect 365954 403058 365986 403294
rect 366222 403058 366306 403294
rect 366542 403058 366574 403294
rect 365954 367614 366574 403058
rect 365954 367378 365986 367614
rect 366222 367378 366306 367614
rect 366542 367378 366574 367614
rect 365954 367294 366574 367378
rect 365954 367058 365986 367294
rect 366222 367058 366306 367294
rect 366542 367058 366574 367294
rect 365954 331614 366574 367058
rect 365954 331378 365986 331614
rect 366222 331378 366306 331614
rect 366542 331378 366574 331614
rect 365954 331294 366574 331378
rect 365954 331058 365986 331294
rect 366222 331058 366306 331294
rect 366542 331058 366574 331294
rect 365954 295614 366574 331058
rect 365954 295378 365986 295614
rect 366222 295378 366306 295614
rect 366542 295378 366574 295614
rect 365954 295294 366574 295378
rect 365954 295058 365986 295294
rect 366222 295058 366306 295294
rect 366542 295058 366574 295294
rect 365954 259614 366574 295058
rect 365954 259378 365986 259614
rect 366222 259378 366306 259614
rect 366542 259378 366574 259614
rect 365954 259294 366574 259378
rect 365954 259058 365986 259294
rect 366222 259058 366306 259294
rect 366542 259058 366574 259294
rect 365954 223614 366574 259058
rect 365954 223378 365986 223614
rect 366222 223378 366306 223614
rect 366542 223378 366574 223614
rect 365954 223294 366574 223378
rect 365954 223058 365986 223294
rect 366222 223058 366306 223294
rect 366542 223058 366574 223294
rect 365954 187614 366574 223058
rect 365954 187378 365986 187614
rect 366222 187378 366306 187614
rect 366542 187378 366574 187614
rect 365954 187294 366574 187378
rect 365954 187058 365986 187294
rect 366222 187058 366306 187294
rect 366542 187058 366574 187294
rect 365954 151614 366574 187058
rect 365954 151378 365986 151614
rect 366222 151378 366306 151614
rect 366542 151378 366574 151614
rect 365954 151294 366574 151378
rect 365954 151058 365986 151294
rect 366222 151058 366306 151294
rect 366542 151058 366574 151294
rect 365954 115614 366574 151058
rect 365954 115378 365986 115614
rect 366222 115378 366306 115614
rect 366542 115378 366574 115614
rect 365954 115294 366574 115378
rect 365954 115058 365986 115294
rect 366222 115058 366306 115294
rect 366542 115058 366574 115294
rect 365954 79614 366574 115058
rect 365954 79378 365986 79614
rect 366222 79378 366306 79614
rect 366542 79378 366574 79614
rect 365954 79294 366574 79378
rect 365954 79058 365986 79294
rect 366222 79058 366306 79294
rect 366542 79058 366574 79294
rect 365954 43614 366574 79058
rect 365954 43378 365986 43614
rect 366222 43378 366306 43614
rect 366542 43378 366574 43614
rect 365954 43294 366574 43378
rect 365954 43058 365986 43294
rect 366222 43058 366306 43294
rect 366542 43058 366574 43294
rect 365954 7614 366574 43058
rect 365954 7378 365986 7614
rect 366222 7378 366306 7614
rect 366542 7378 366574 7614
rect 365954 7294 366574 7378
rect 365954 7058 365986 7294
rect 366222 7058 366306 7294
rect 366542 7058 366574 7294
rect 365954 -4186 366574 7058
rect 365954 -4422 365986 -4186
rect 366222 -4422 366306 -4186
rect 366542 -4422 366574 -4186
rect 365954 -4506 366574 -4422
rect 365954 -4742 365986 -4506
rect 366222 -4742 366306 -4506
rect 366542 -4742 366574 -4506
rect 365954 -7654 366574 -4742
rect 367194 709638 367814 711590
rect 367194 709402 367226 709638
rect 367462 709402 367546 709638
rect 367782 709402 367814 709638
rect 367194 709318 367814 709402
rect 367194 709082 367226 709318
rect 367462 709082 367546 709318
rect 367782 709082 367814 709318
rect 367194 692854 367814 709082
rect 367194 692618 367226 692854
rect 367462 692618 367546 692854
rect 367782 692618 367814 692854
rect 367194 692534 367814 692618
rect 367194 692298 367226 692534
rect 367462 692298 367546 692534
rect 367782 692298 367814 692534
rect 367194 656854 367814 692298
rect 367194 656618 367226 656854
rect 367462 656618 367546 656854
rect 367782 656618 367814 656854
rect 367194 656534 367814 656618
rect 367194 656298 367226 656534
rect 367462 656298 367546 656534
rect 367782 656298 367814 656534
rect 367194 620854 367814 656298
rect 367194 620618 367226 620854
rect 367462 620618 367546 620854
rect 367782 620618 367814 620854
rect 367194 620534 367814 620618
rect 367194 620298 367226 620534
rect 367462 620298 367546 620534
rect 367782 620298 367814 620534
rect 367194 584854 367814 620298
rect 367194 584618 367226 584854
rect 367462 584618 367546 584854
rect 367782 584618 367814 584854
rect 367194 584534 367814 584618
rect 367194 584298 367226 584534
rect 367462 584298 367546 584534
rect 367782 584298 367814 584534
rect 367194 548854 367814 584298
rect 367194 548618 367226 548854
rect 367462 548618 367546 548854
rect 367782 548618 367814 548854
rect 367194 548534 367814 548618
rect 367194 548298 367226 548534
rect 367462 548298 367546 548534
rect 367782 548298 367814 548534
rect 367194 512854 367814 548298
rect 367194 512618 367226 512854
rect 367462 512618 367546 512854
rect 367782 512618 367814 512854
rect 367194 512534 367814 512618
rect 367194 512298 367226 512534
rect 367462 512298 367546 512534
rect 367782 512298 367814 512534
rect 367194 476854 367814 512298
rect 367194 476618 367226 476854
rect 367462 476618 367546 476854
rect 367782 476618 367814 476854
rect 367194 476534 367814 476618
rect 367194 476298 367226 476534
rect 367462 476298 367546 476534
rect 367782 476298 367814 476534
rect 367194 440854 367814 476298
rect 367194 440618 367226 440854
rect 367462 440618 367546 440854
rect 367782 440618 367814 440854
rect 367194 440534 367814 440618
rect 367194 440298 367226 440534
rect 367462 440298 367546 440534
rect 367782 440298 367814 440534
rect 367194 404854 367814 440298
rect 367194 404618 367226 404854
rect 367462 404618 367546 404854
rect 367782 404618 367814 404854
rect 367194 404534 367814 404618
rect 367194 404298 367226 404534
rect 367462 404298 367546 404534
rect 367782 404298 367814 404534
rect 367194 368854 367814 404298
rect 367194 368618 367226 368854
rect 367462 368618 367546 368854
rect 367782 368618 367814 368854
rect 367194 368534 367814 368618
rect 367194 368298 367226 368534
rect 367462 368298 367546 368534
rect 367782 368298 367814 368534
rect 367194 332854 367814 368298
rect 367194 332618 367226 332854
rect 367462 332618 367546 332854
rect 367782 332618 367814 332854
rect 367194 332534 367814 332618
rect 367194 332298 367226 332534
rect 367462 332298 367546 332534
rect 367782 332298 367814 332534
rect 367194 296854 367814 332298
rect 367194 296618 367226 296854
rect 367462 296618 367546 296854
rect 367782 296618 367814 296854
rect 367194 296534 367814 296618
rect 367194 296298 367226 296534
rect 367462 296298 367546 296534
rect 367782 296298 367814 296534
rect 367194 260854 367814 296298
rect 367194 260618 367226 260854
rect 367462 260618 367546 260854
rect 367782 260618 367814 260854
rect 367194 260534 367814 260618
rect 367194 260298 367226 260534
rect 367462 260298 367546 260534
rect 367782 260298 367814 260534
rect 367194 224854 367814 260298
rect 367194 224618 367226 224854
rect 367462 224618 367546 224854
rect 367782 224618 367814 224854
rect 367194 224534 367814 224618
rect 367194 224298 367226 224534
rect 367462 224298 367546 224534
rect 367782 224298 367814 224534
rect 367194 188854 367814 224298
rect 367194 188618 367226 188854
rect 367462 188618 367546 188854
rect 367782 188618 367814 188854
rect 367194 188534 367814 188618
rect 367194 188298 367226 188534
rect 367462 188298 367546 188534
rect 367782 188298 367814 188534
rect 367194 152854 367814 188298
rect 367194 152618 367226 152854
rect 367462 152618 367546 152854
rect 367782 152618 367814 152854
rect 367194 152534 367814 152618
rect 367194 152298 367226 152534
rect 367462 152298 367546 152534
rect 367782 152298 367814 152534
rect 367194 116854 367814 152298
rect 367194 116618 367226 116854
rect 367462 116618 367546 116854
rect 367782 116618 367814 116854
rect 367194 116534 367814 116618
rect 367194 116298 367226 116534
rect 367462 116298 367546 116534
rect 367782 116298 367814 116534
rect 367194 80854 367814 116298
rect 367194 80618 367226 80854
rect 367462 80618 367546 80854
rect 367782 80618 367814 80854
rect 367194 80534 367814 80618
rect 367194 80298 367226 80534
rect 367462 80298 367546 80534
rect 367782 80298 367814 80534
rect 367194 44854 367814 80298
rect 367194 44618 367226 44854
rect 367462 44618 367546 44854
rect 367782 44618 367814 44854
rect 367194 44534 367814 44618
rect 367194 44298 367226 44534
rect 367462 44298 367546 44534
rect 367782 44298 367814 44534
rect 367194 8854 367814 44298
rect 367194 8618 367226 8854
rect 367462 8618 367546 8854
rect 367782 8618 367814 8854
rect 367194 8534 367814 8618
rect 367194 8298 367226 8534
rect 367462 8298 367546 8534
rect 367782 8298 367814 8534
rect 367194 -5146 367814 8298
rect 367194 -5382 367226 -5146
rect 367462 -5382 367546 -5146
rect 367782 -5382 367814 -5146
rect 367194 -5466 367814 -5382
rect 367194 -5702 367226 -5466
rect 367462 -5702 367546 -5466
rect 367782 -5702 367814 -5466
rect 367194 -7654 367814 -5702
rect 368434 710598 369054 711590
rect 368434 710362 368466 710598
rect 368702 710362 368786 710598
rect 369022 710362 369054 710598
rect 368434 710278 369054 710362
rect 368434 710042 368466 710278
rect 368702 710042 368786 710278
rect 369022 710042 369054 710278
rect 368434 694094 369054 710042
rect 368434 693858 368466 694094
rect 368702 693858 368786 694094
rect 369022 693858 369054 694094
rect 368434 693774 369054 693858
rect 368434 693538 368466 693774
rect 368702 693538 368786 693774
rect 369022 693538 369054 693774
rect 368434 658094 369054 693538
rect 368434 657858 368466 658094
rect 368702 657858 368786 658094
rect 369022 657858 369054 658094
rect 368434 657774 369054 657858
rect 368434 657538 368466 657774
rect 368702 657538 368786 657774
rect 369022 657538 369054 657774
rect 368434 622094 369054 657538
rect 368434 621858 368466 622094
rect 368702 621858 368786 622094
rect 369022 621858 369054 622094
rect 368434 621774 369054 621858
rect 368434 621538 368466 621774
rect 368702 621538 368786 621774
rect 369022 621538 369054 621774
rect 368434 586094 369054 621538
rect 368434 585858 368466 586094
rect 368702 585858 368786 586094
rect 369022 585858 369054 586094
rect 368434 585774 369054 585858
rect 368434 585538 368466 585774
rect 368702 585538 368786 585774
rect 369022 585538 369054 585774
rect 368434 550094 369054 585538
rect 368434 549858 368466 550094
rect 368702 549858 368786 550094
rect 369022 549858 369054 550094
rect 368434 549774 369054 549858
rect 368434 549538 368466 549774
rect 368702 549538 368786 549774
rect 369022 549538 369054 549774
rect 368434 514094 369054 549538
rect 368434 513858 368466 514094
rect 368702 513858 368786 514094
rect 369022 513858 369054 514094
rect 368434 513774 369054 513858
rect 368434 513538 368466 513774
rect 368702 513538 368786 513774
rect 369022 513538 369054 513774
rect 368434 478094 369054 513538
rect 368434 477858 368466 478094
rect 368702 477858 368786 478094
rect 369022 477858 369054 478094
rect 368434 477774 369054 477858
rect 368434 477538 368466 477774
rect 368702 477538 368786 477774
rect 369022 477538 369054 477774
rect 368434 442094 369054 477538
rect 368434 441858 368466 442094
rect 368702 441858 368786 442094
rect 369022 441858 369054 442094
rect 368434 441774 369054 441858
rect 368434 441538 368466 441774
rect 368702 441538 368786 441774
rect 369022 441538 369054 441774
rect 368434 406094 369054 441538
rect 368434 405858 368466 406094
rect 368702 405858 368786 406094
rect 369022 405858 369054 406094
rect 368434 405774 369054 405858
rect 368434 405538 368466 405774
rect 368702 405538 368786 405774
rect 369022 405538 369054 405774
rect 368434 370094 369054 405538
rect 368434 369858 368466 370094
rect 368702 369858 368786 370094
rect 369022 369858 369054 370094
rect 368434 369774 369054 369858
rect 368434 369538 368466 369774
rect 368702 369538 368786 369774
rect 369022 369538 369054 369774
rect 368434 334094 369054 369538
rect 368434 333858 368466 334094
rect 368702 333858 368786 334094
rect 369022 333858 369054 334094
rect 368434 333774 369054 333858
rect 368434 333538 368466 333774
rect 368702 333538 368786 333774
rect 369022 333538 369054 333774
rect 368434 298094 369054 333538
rect 368434 297858 368466 298094
rect 368702 297858 368786 298094
rect 369022 297858 369054 298094
rect 368434 297774 369054 297858
rect 368434 297538 368466 297774
rect 368702 297538 368786 297774
rect 369022 297538 369054 297774
rect 368434 262094 369054 297538
rect 368434 261858 368466 262094
rect 368702 261858 368786 262094
rect 369022 261858 369054 262094
rect 368434 261774 369054 261858
rect 368434 261538 368466 261774
rect 368702 261538 368786 261774
rect 369022 261538 369054 261774
rect 368434 226094 369054 261538
rect 368434 225858 368466 226094
rect 368702 225858 368786 226094
rect 369022 225858 369054 226094
rect 368434 225774 369054 225858
rect 368434 225538 368466 225774
rect 368702 225538 368786 225774
rect 369022 225538 369054 225774
rect 368434 190094 369054 225538
rect 368434 189858 368466 190094
rect 368702 189858 368786 190094
rect 369022 189858 369054 190094
rect 368434 189774 369054 189858
rect 368434 189538 368466 189774
rect 368702 189538 368786 189774
rect 369022 189538 369054 189774
rect 368434 154094 369054 189538
rect 368434 153858 368466 154094
rect 368702 153858 368786 154094
rect 369022 153858 369054 154094
rect 368434 153774 369054 153858
rect 368434 153538 368466 153774
rect 368702 153538 368786 153774
rect 369022 153538 369054 153774
rect 368434 118094 369054 153538
rect 368434 117858 368466 118094
rect 368702 117858 368786 118094
rect 369022 117858 369054 118094
rect 368434 117774 369054 117858
rect 368434 117538 368466 117774
rect 368702 117538 368786 117774
rect 369022 117538 369054 117774
rect 368434 82094 369054 117538
rect 368434 81858 368466 82094
rect 368702 81858 368786 82094
rect 369022 81858 369054 82094
rect 368434 81774 369054 81858
rect 368434 81538 368466 81774
rect 368702 81538 368786 81774
rect 369022 81538 369054 81774
rect 368434 46094 369054 81538
rect 368434 45858 368466 46094
rect 368702 45858 368786 46094
rect 369022 45858 369054 46094
rect 368434 45774 369054 45858
rect 368434 45538 368466 45774
rect 368702 45538 368786 45774
rect 369022 45538 369054 45774
rect 368434 10094 369054 45538
rect 368434 9858 368466 10094
rect 368702 9858 368786 10094
rect 369022 9858 369054 10094
rect 368434 9774 369054 9858
rect 368434 9538 368466 9774
rect 368702 9538 368786 9774
rect 369022 9538 369054 9774
rect 368434 -6106 369054 9538
rect 368434 -6342 368466 -6106
rect 368702 -6342 368786 -6106
rect 369022 -6342 369054 -6106
rect 368434 -6426 369054 -6342
rect 368434 -6662 368466 -6426
rect 368702 -6662 368786 -6426
rect 369022 -6662 369054 -6426
rect 368434 -7654 369054 -6662
rect 369674 711558 370294 711590
rect 369674 711322 369706 711558
rect 369942 711322 370026 711558
rect 370262 711322 370294 711558
rect 369674 711238 370294 711322
rect 369674 711002 369706 711238
rect 369942 711002 370026 711238
rect 370262 711002 370294 711238
rect 369674 695334 370294 711002
rect 369674 695098 369706 695334
rect 369942 695098 370026 695334
rect 370262 695098 370294 695334
rect 369674 695014 370294 695098
rect 369674 694778 369706 695014
rect 369942 694778 370026 695014
rect 370262 694778 370294 695014
rect 369674 659334 370294 694778
rect 369674 659098 369706 659334
rect 369942 659098 370026 659334
rect 370262 659098 370294 659334
rect 369674 659014 370294 659098
rect 369674 658778 369706 659014
rect 369942 658778 370026 659014
rect 370262 658778 370294 659014
rect 369674 623334 370294 658778
rect 369674 623098 369706 623334
rect 369942 623098 370026 623334
rect 370262 623098 370294 623334
rect 369674 623014 370294 623098
rect 369674 622778 369706 623014
rect 369942 622778 370026 623014
rect 370262 622778 370294 623014
rect 369674 587334 370294 622778
rect 369674 587098 369706 587334
rect 369942 587098 370026 587334
rect 370262 587098 370294 587334
rect 369674 587014 370294 587098
rect 369674 586778 369706 587014
rect 369942 586778 370026 587014
rect 370262 586778 370294 587014
rect 369674 551334 370294 586778
rect 369674 551098 369706 551334
rect 369942 551098 370026 551334
rect 370262 551098 370294 551334
rect 369674 551014 370294 551098
rect 369674 550778 369706 551014
rect 369942 550778 370026 551014
rect 370262 550778 370294 551014
rect 369674 515334 370294 550778
rect 369674 515098 369706 515334
rect 369942 515098 370026 515334
rect 370262 515098 370294 515334
rect 369674 515014 370294 515098
rect 369674 514778 369706 515014
rect 369942 514778 370026 515014
rect 370262 514778 370294 515014
rect 369674 479334 370294 514778
rect 369674 479098 369706 479334
rect 369942 479098 370026 479334
rect 370262 479098 370294 479334
rect 369674 479014 370294 479098
rect 369674 478778 369706 479014
rect 369942 478778 370026 479014
rect 370262 478778 370294 479014
rect 369674 443334 370294 478778
rect 369674 443098 369706 443334
rect 369942 443098 370026 443334
rect 370262 443098 370294 443334
rect 369674 443014 370294 443098
rect 369674 442778 369706 443014
rect 369942 442778 370026 443014
rect 370262 442778 370294 443014
rect 369674 407334 370294 442778
rect 369674 407098 369706 407334
rect 369942 407098 370026 407334
rect 370262 407098 370294 407334
rect 369674 407014 370294 407098
rect 369674 406778 369706 407014
rect 369942 406778 370026 407014
rect 370262 406778 370294 407014
rect 369674 371334 370294 406778
rect 369674 371098 369706 371334
rect 369942 371098 370026 371334
rect 370262 371098 370294 371334
rect 369674 371014 370294 371098
rect 369674 370778 369706 371014
rect 369942 370778 370026 371014
rect 370262 370778 370294 371014
rect 369674 335334 370294 370778
rect 369674 335098 369706 335334
rect 369942 335098 370026 335334
rect 370262 335098 370294 335334
rect 369674 335014 370294 335098
rect 369674 334778 369706 335014
rect 369942 334778 370026 335014
rect 370262 334778 370294 335014
rect 369674 299334 370294 334778
rect 369674 299098 369706 299334
rect 369942 299098 370026 299334
rect 370262 299098 370294 299334
rect 369674 299014 370294 299098
rect 369674 298778 369706 299014
rect 369942 298778 370026 299014
rect 370262 298778 370294 299014
rect 369674 263334 370294 298778
rect 369674 263098 369706 263334
rect 369942 263098 370026 263334
rect 370262 263098 370294 263334
rect 369674 263014 370294 263098
rect 369674 262778 369706 263014
rect 369942 262778 370026 263014
rect 370262 262778 370294 263014
rect 369674 227334 370294 262778
rect 369674 227098 369706 227334
rect 369942 227098 370026 227334
rect 370262 227098 370294 227334
rect 369674 227014 370294 227098
rect 369674 226778 369706 227014
rect 369942 226778 370026 227014
rect 370262 226778 370294 227014
rect 369674 191334 370294 226778
rect 369674 191098 369706 191334
rect 369942 191098 370026 191334
rect 370262 191098 370294 191334
rect 369674 191014 370294 191098
rect 369674 190778 369706 191014
rect 369942 190778 370026 191014
rect 370262 190778 370294 191014
rect 369674 155334 370294 190778
rect 369674 155098 369706 155334
rect 369942 155098 370026 155334
rect 370262 155098 370294 155334
rect 369674 155014 370294 155098
rect 369674 154778 369706 155014
rect 369942 154778 370026 155014
rect 370262 154778 370294 155014
rect 369674 119334 370294 154778
rect 369674 119098 369706 119334
rect 369942 119098 370026 119334
rect 370262 119098 370294 119334
rect 369674 119014 370294 119098
rect 369674 118778 369706 119014
rect 369942 118778 370026 119014
rect 370262 118778 370294 119014
rect 369674 83334 370294 118778
rect 369674 83098 369706 83334
rect 369942 83098 370026 83334
rect 370262 83098 370294 83334
rect 369674 83014 370294 83098
rect 369674 82778 369706 83014
rect 369942 82778 370026 83014
rect 370262 82778 370294 83014
rect 369674 47334 370294 82778
rect 369674 47098 369706 47334
rect 369942 47098 370026 47334
rect 370262 47098 370294 47334
rect 369674 47014 370294 47098
rect 369674 46778 369706 47014
rect 369942 46778 370026 47014
rect 370262 46778 370294 47014
rect 369674 11334 370294 46778
rect 369674 11098 369706 11334
rect 369942 11098 370026 11334
rect 370262 11098 370294 11334
rect 369674 11014 370294 11098
rect 369674 10778 369706 11014
rect 369942 10778 370026 11014
rect 370262 10778 370294 11014
rect 369674 -7066 370294 10778
rect 369674 -7302 369706 -7066
rect 369942 -7302 370026 -7066
rect 370262 -7302 370294 -7066
rect 369674 -7386 370294 -7302
rect 369674 -7622 369706 -7386
rect 369942 -7622 370026 -7386
rect 370262 -7622 370294 -7386
rect 369674 -7654 370294 -7622
rect 396994 704838 397614 711590
rect 396994 704602 397026 704838
rect 397262 704602 397346 704838
rect 397582 704602 397614 704838
rect 396994 704518 397614 704602
rect 396994 704282 397026 704518
rect 397262 704282 397346 704518
rect 397582 704282 397614 704518
rect 396994 686654 397614 704282
rect 396994 686418 397026 686654
rect 397262 686418 397346 686654
rect 397582 686418 397614 686654
rect 396994 686334 397614 686418
rect 396994 686098 397026 686334
rect 397262 686098 397346 686334
rect 397582 686098 397614 686334
rect 396994 650654 397614 686098
rect 396994 650418 397026 650654
rect 397262 650418 397346 650654
rect 397582 650418 397614 650654
rect 396994 650334 397614 650418
rect 396994 650098 397026 650334
rect 397262 650098 397346 650334
rect 397582 650098 397614 650334
rect 396994 614654 397614 650098
rect 396994 614418 397026 614654
rect 397262 614418 397346 614654
rect 397582 614418 397614 614654
rect 396994 614334 397614 614418
rect 396994 614098 397026 614334
rect 397262 614098 397346 614334
rect 397582 614098 397614 614334
rect 396994 578654 397614 614098
rect 396994 578418 397026 578654
rect 397262 578418 397346 578654
rect 397582 578418 397614 578654
rect 396994 578334 397614 578418
rect 396994 578098 397026 578334
rect 397262 578098 397346 578334
rect 397582 578098 397614 578334
rect 396994 542654 397614 578098
rect 396994 542418 397026 542654
rect 397262 542418 397346 542654
rect 397582 542418 397614 542654
rect 396994 542334 397614 542418
rect 396994 542098 397026 542334
rect 397262 542098 397346 542334
rect 397582 542098 397614 542334
rect 396994 506654 397614 542098
rect 396994 506418 397026 506654
rect 397262 506418 397346 506654
rect 397582 506418 397614 506654
rect 396994 506334 397614 506418
rect 396994 506098 397026 506334
rect 397262 506098 397346 506334
rect 397582 506098 397614 506334
rect 396994 470654 397614 506098
rect 396994 470418 397026 470654
rect 397262 470418 397346 470654
rect 397582 470418 397614 470654
rect 396994 470334 397614 470418
rect 396994 470098 397026 470334
rect 397262 470098 397346 470334
rect 397582 470098 397614 470334
rect 396994 434654 397614 470098
rect 396994 434418 397026 434654
rect 397262 434418 397346 434654
rect 397582 434418 397614 434654
rect 396994 434334 397614 434418
rect 396994 434098 397026 434334
rect 397262 434098 397346 434334
rect 397582 434098 397614 434334
rect 396994 398654 397614 434098
rect 396994 398418 397026 398654
rect 397262 398418 397346 398654
rect 397582 398418 397614 398654
rect 396994 398334 397614 398418
rect 396994 398098 397026 398334
rect 397262 398098 397346 398334
rect 397582 398098 397614 398334
rect 396994 362654 397614 398098
rect 396994 362418 397026 362654
rect 397262 362418 397346 362654
rect 397582 362418 397614 362654
rect 396994 362334 397614 362418
rect 396994 362098 397026 362334
rect 397262 362098 397346 362334
rect 397582 362098 397614 362334
rect 396994 326654 397614 362098
rect 396994 326418 397026 326654
rect 397262 326418 397346 326654
rect 397582 326418 397614 326654
rect 396994 326334 397614 326418
rect 396994 326098 397026 326334
rect 397262 326098 397346 326334
rect 397582 326098 397614 326334
rect 396994 290654 397614 326098
rect 396994 290418 397026 290654
rect 397262 290418 397346 290654
rect 397582 290418 397614 290654
rect 396994 290334 397614 290418
rect 396994 290098 397026 290334
rect 397262 290098 397346 290334
rect 397582 290098 397614 290334
rect 396994 254654 397614 290098
rect 396994 254418 397026 254654
rect 397262 254418 397346 254654
rect 397582 254418 397614 254654
rect 396994 254334 397614 254418
rect 396994 254098 397026 254334
rect 397262 254098 397346 254334
rect 397582 254098 397614 254334
rect 396994 218654 397614 254098
rect 396994 218418 397026 218654
rect 397262 218418 397346 218654
rect 397582 218418 397614 218654
rect 396994 218334 397614 218418
rect 396994 218098 397026 218334
rect 397262 218098 397346 218334
rect 397582 218098 397614 218334
rect 396994 182654 397614 218098
rect 396994 182418 397026 182654
rect 397262 182418 397346 182654
rect 397582 182418 397614 182654
rect 396994 182334 397614 182418
rect 396994 182098 397026 182334
rect 397262 182098 397346 182334
rect 397582 182098 397614 182334
rect 396994 146654 397614 182098
rect 396994 146418 397026 146654
rect 397262 146418 397346 146654
rect 397582 146418 397614 146654
rect 396994 146334 397614 146418
rect 396994 146098 397026 146334
rect 397262 146098 397346 146334
rect 397582 146098 397614 146334
rect 396994 110654 397614 146098
rect 396994 110418 397026 110654
rect 397262 110418 397346 110654
rect 397582 110418 397614 110654
rect 396994 110334 397614 110418
rect 396994 110098 397026 110334
rect 397262 110098 397346 110334
rect 397582 110098 397614 110334
rect 396994 74654 397614 110098
rect 396994 74418 397026 74654
rect 397262 74418 397346 74654
rect 397582 74418 397614 74654
rect 396994 74334 397614 74418
rect 396994 74098 397026 74334
rect 397262 74098 397346 74334
rect 397582 74098 397614 74334
rect 396994 38654 397614 74098
rect 396994 38418 397026 38654
rect 397262 38418 397346 38654
rect 397582 38418 397614 38654
rect 396994 38334 397614 38418
rect 396994 38098 397026 38334
rect 397262 38098 397346 38334
rect 397582 38098 397614 38334
rect 396994 2654 397614 38098
rect 396994 2418 397026 2654
rect 397262 2418 397346 2654
rect 397582 2418 397614 2654
rect 396994 2334 397614 2418
rect 396994 2098 397026 2334
rect 397262 2098 397346 2334
rect 397582 2098 397614 2334
rect 396994 -346 397614 2098
rect 396994 -582 397026 -346
rect 397262 -582 397346 -346
rect 397582 -582 397614 -346
rect 396994 -666 397614 -582
rect 396994 -902 397026 -666
rect 397262 -902 397346 -666
rect 397582 -902 397614 -666
rect 396994 -7654 397614 -902
rect 398234 705798 398854 711590
rect 398234 705562 398266 705798
rect 398502 705562 398586 705798
rect 398822 705562 398854 705798
rect 398234 705478 398854 705562
rect 398234 705242 398266 705478
rect 398502 705242 398586 705478
rect 398822 705242 398854 705478
rect 398234 687894 398854 705242
rect 398234 687658 398266 687894
rect 398502 687658 398586 687894
rect 398822 687658 398854 687894
rect 398234 687574 398854 687658
rect 398234 687338 398266 687574
rect 398502 687338 398586 687574
rect 398822 687338 398854 687574
rect 398234 651894 398854 687338
rect 398234 651658 398266 651894
rect 398502 651658 398586 651894
rect 398822 651658 398854 651894
rect 398234 651574 398854 651658
rect 398234 651338 398266 651574
rect 398502 651338 398586 651574
rect 398822 651338 398854 651574
rect 398234 615894 398854 651338
rect 398234 615658 398266 615894
rect 398502 615658 398586 615894
rect 398822 615658 398854 615894
rect 398234 615574 398854 615658
rect 398234 615338 398266 615574
rect 398502 615338 398586 615574
rect 398822 615338 398854 615574
rect 398234 579894 398854 615338
rect 398234 579658 398266 579894
rect 398502 579658 398586 579894
rect 398822 579658 398854 579894
rect 398234 579574 398854 579658
rect 398234 579338 398266 579574
rect 398502 579338 398586 579574
rect 398822 579338 398854 579574
rect 398234 543894 398854 579338
rect 398234 543658 398266 543894
rect 398502 543658 398586 543894
rect 398822 543658 398854 543894
rect 398234 543574 398854 543658
rect 398234 543338 398266 543574
rect 398502 543338 398586 543574
rect 398822 543338 398854 543574
rect 398234 507894 398854 543338
rect 398234 507658 398266 507894
rect 398502 507658 398586 507894
rect 398822 507658 398854 507894
rect 398234 507574 398854 507658
rect 398234 507338 398266 507574
rect 398502 507338 398586 507574
rect 398822 507338 398854 507574
rect 398234 471894 398854 507338
rect 398234 471658 398266 471894
rect 398502 471658 398586 471894
rect 398822 471658 398854 471894
rect 398234 471574 398854 471658
rect 398234 471338 398266 471574
rect 398502 471338 398586 471574
rect 398822 471338 398854 471574
rect 398234 435894 398854 471338
rect 398234 435658 398266 435894
rect 398502 435658 398586 435894
rect 398822 435658 398854 435894
rect 398234 435574 398854 435658
rect 398234 435338 398266 435574
rect 398502 435338 398586 435574
rect 398822 435338 398854 435574
rect 398234 399894 398854 435338
rect 398234 399658 398266 399894
rect 398502 399658 398586 399894
rect 398822 399658 398854 399894
rect 398234 399574 398854 399658
rect 398234 399338 398266 399574
rect 398502 399338 398586 399574
rect 398822 399338 398854 399574
rect 398234 363894 398854 399338
rect 398234 363658 398266 363894
rect 398502 363658 398586 363894
rect 398822 363658 398854 363894
rect 398234 363574 398854 363658
rect 398234 363338 398266 363574
rect 398502 363338 398586 363574
rect 398822 363338 398854 363574
rect 398234 327894 398854 363338
rect 398234 327658 398266 327894
rect 398502 327658 398586 327894
rect 398822 327658 398854 327894
rect 398234 327574 398854 327658
rect 398234 327338 398266 327574
rect 398502 327338 398586 327574
rect 398822 327338 398854 327574
rect 398234 291894 398854 327338
rect 398234 291658 398266 291894
rect 398502 291658 398586 291894
rect 398822 291658 398854 291894
rect 398234 291574 398854 291658
rect 398234 291338 398266 291574
rect 398502 291338 398586 291574
rect 398822 291338 398854 291574
rect 398234 255894 398854 291338
rect 398234 255658 398266 255894
rect 398502 255658 398586 255894
rect 398822 255658 398854 255894
rect 398234 255574 398854 255658
rect 398234 255338 398266 255574
rect 398502 255338 398586 255574
rect 398822 255338 398854 255574
rect 398234 219894 398854 255338
rect 398234 219658 398266 219894
rect 398502 219658 398586 219894
rect 398822 219658 398854 219894
rect 398234 219574 398854 219658
rect 398234 219338 398266 219574
rect 398502 219338 398586 219574
rect 398822 219338 398854 219574
rect 398234 183894 398854 219338
rect 398234 183658 398266 183894
rect 398502 183658 398586 183894
rect 398822 183658 398854 183894
rect 398234 183574 398854 183658
rect 398234 183338 398266 183574
rect 398502 183338 398586 183574
rect 398822 183338 398854 183574
rect 398234 147894 398854 183338
rect 398234 147658 398266 147894
rect 398502 147658 398586 147894
rect 398822 147658 398854 147894
rect 398234 147574 398854 147658
rect 398234 147338 398266 147574
rect 398502 147338 398586 147574
rect 398822 147338 398854 147574
rect 398234 111894 398854 147338
rect 398234 111658 398266 111894
rect 398502 111658 398586 111894
rect 398822 111658 398854 111894
rect 398234 111574 398854 111658
rect 398234 111338 398266 111574
rect 398502 111338 398586 111574
rect 398822 111338 398854 111574
rect 398234 75894 398854 111338
rect 398234 75658 398266 75894
rect 398502 75658 398586 75894
rect 398822 75658 398854 75894
rect 398234 75574 398854 75658
rect 398234 75338 398266 75574
rect 398502 75338 398586 75574
rect 398822 75338 398854 75574
rect 398234 39894 398854 75338
rect 398234 39658 398266 39894
rect 398502 39658 398586 39894
rect 398822 39658 398854 39894
rect 398234 39574 398854 39658
rect 398234 39338 398266 39574
rect 398502 39338 398586 39574
rect 398822 39338 398854 39574
rect 398234 3894 398854 39338
rect 398234 3658 398266 3894
rect 398502 3658 398586 3894
rect 398822 3658 398854 3894
rect 398234 3574 398854 3658
rect 398234 3338 398266 3574
rect 398502 3338 398586 3574
rect 398822 3338 398854 3574
rect 398234 -1306 398854 3338
rect 398234 -1542 398266 -1306
rect 398502 -1542 398586 -1306
rect 398822 -1542 398854 -1306
rect 398234 -1626 398854 -1542
rect 398234 -1862 398266 -1626
rect 398502 -1862 398586 -1626
rect 398822 -1862 398854 -1626
rect 398234 -7654 398854 -1862
rect 399474 706758 400094 711590
rect 399474 706522 399506 706758
rect 399742 706522 399826 706758
rect 400062 706522 400094 706758
rect 399474 706438 400094 706522
rect 399474 706202 399506 706438
rect 399742 706202 399826 706438
rect 400062 706202 400094 706438
rect 399474 689134 400094 706202
rect 399474 688898 399506 689134
rect 399742 688898 399826 689134
rect 400062 688898 400094 689134
rect 399474 688814 400094 688898
rect 399474 688578 399506 688814
rect 399742 688578 399826 688814
rect 400062 688578 400094 688814
rect 399474 653134 400094 688578
rect 399474 652898 399506 653134
rect 399742 652898 399826 653134
rect 400062 652898 400094 653134
rect 399474 652814 400094 652898
rect 399474 652578 399506 652814
rect 399742 652578 399826 652814
rect 400062 652578 400094 652814
rect 399474 617134 400094 652578
rect 399474 616898 399506 617134
rect 399742 616898 399826 617134
rect 400062 616898 400094 617134
rect 399474 616814 400094 616898
rect 399474 616578 399506 616814
rect 399742 616578 399826 616814
rect 400062 616578 400094 616814
rect 399474 581134 400094 616578
rect 399474 580898 399506 581134
rect 399742 580898 399826 581134
rect 400062 580898 400094 581134
rect 399474 580814 400094 580898
rect 399474 580578 399506 580814
rect 399742 580578 399826 580814
rect 400062 580578 400094 580814
rect 399474 545134 400094 580578
rect 399474 544898 399506 545134
rect 399742 544898 399826 545134
rect 400062 544898 400094 545134
rect 399474 544814 400094 544898
rect 399474 544578 399506 544814
rect 399742 544578 399826 544814
rect 400062 544578 400094 544814
rect 399474 509134 400094 544578
rect 399474 508898 399506 509134
rect 399742 508898 399826 509134
rect 400062 508898 400094 509134
rect 399474 508814 400094 508898
rect 399474 508578 399506 508814
rect 399742 508578 399826 508814
rect 400062 508578 400094 508814
rect 399474 473134 400094 508578
rect 399474 472898 399506 473134
rect 399742 472898 399826 473134
rect 400062 472898 400094 473134
rect 399474 472814 400094 472898
rect 399474 472578 399506 472814
rect 399742 472578 399826 472814
rect 400062 472578 400094 472814
rect 399474 437134 400094 472578
rect 399474 436898 399506 437134
rect 399742 436898 399826 437134
rect 400062 436898 400094 437134
rect 399474 436814 400094 436898
rect 399474 436578 399506 436814
rect 399742 436578 399826 436814
rect 400062 436578 400094 436814
rect 399474 401134 400094 436578
rect 399474 400898 399506 401134
rect 399742 400898 399826 401134
rect 400062 400898 400094 401134
rect 399474 400814 400094 400898
rect 399474 400578 399506 400814
rect 399742 400578 399826 400814
rect 400062 400578 400094 400814
rect 399474 365134 400094 400578
rect 399474 364898 399506 365134
rect 399742 364898 399826 365134
rect 400062 364898 400094 365134
rect 399474 364814 400094 364898
rect 399474 364578 399506 364814
rect 399742 364578 399826 364814
rect 400062 364578 400094 364814
rect 399474 329134 400094 364578
rect 399474 328898 399506 329134
rect 399742 328898 399826 329134
rect 400062 328898 400094 329134
rect 399474 328814 400094 328898
rect 399474 328578 399506 328814
rect 399742 328578 399826 328814
rect 400062 328578 400094 328814
rect 399474 293134 400094 328578
rect 399474 292898 399506 293134
rect 399742 292898 399826 293134
rect 400062 292898 400094 293134
rect 399474 292814 400094 292898
rect 399474 292578 399506 292814
rect 399742 292578 399826 292814
rect 400062 292578 400094 292814
rect 399474 257134 400094 292578
rect 399474 256898 399506 257134
rect 399742 256898 399826 257134
rect 400062 256898 400094 257134
rect 399474 256814 400094 256898
rect 399474 256578 399506 256814
rect 399742 256578 399826 256814
rect 400062 256578 400094 256814
rect 399474 221134 400094 256578
rect 399474 220898 399506 221134
rect 399742 220898 399826 221134
rect 400062 220898 400094 221134
rect 399474 220814 400094 220898
rect 399474 220578 399506 220814
rect 399742 220578 399826 220814
rect 400062 220578 400094 220814
rect 399474 185134 400094 220578
rect 399474 184898 399506 185134
rect 399742 184898 399826 185134
rect 400062 184898 400094 185134
rect 399474 184814 400094 184898
rect 399474 184578 399506 184814
rect 399742 184578 399826 184814
rect 400062 184578 400094 184814
rect 399474 149134 400094 184578
rect 399474 148898 399506 149134
rect 399742 148898 399826 149134
rect 400062 148898 400094 149134
rect 399474 148814 400094 148898
rect 399474 148578 399506 148814
rect 399742 148578 399826 148814
rect 400062 148578 400094 148814
rect 399474 113134 400094 148578
rect 399474 112898 399506 113134
rect 399742 112898 399826 113134
rect 400062 112898 400094 113134
rect 399474 112814 400094 112898
rect 399474 112578 399506 112814
rect 399742 112578 399826 112814
rect 400062 112578 400094 112814
rect 399474 77134 400094 112578
rect 399474 76898 399506 77134
rect 399742 76898 399826 77134
rect 400062 76898 400094 77134
rect 399474 76814 400094 76898
rect 399474 76578 399506 76814
rect 399742 76578 399826 76814
rect 400062 76578 400094 76814
rect 399474 41134 400094 76578
rect 399474 40898 399506 41134
rect 399742 40898 399826 41134
rect 400062 40898 400094 41134
rect 399474 40814 400094 40898
rect 399474 40578 399506 40814
rect 399742 40578 399826 40814
rect 400062 40578 400094 40814
rect 399474 5134 400094 40578
rect 399474 4898 399506 5134
rect 399742 4898 399826 5134
rect 400062 4898 400094 5134
rect 399474 4814 400094 4898
rect 399474 4578 399506 4814
rect 399742 4578 399826 4814
rect 400062 4578 400094 4814
rect 399474 -2266 400094 4578
rect 399474 -2502 399506 -2266
rect 399742 -2502 399826 -2266
rect 400062 -2502 400094 -2266
rect 399474 -2586 400094 -2502
rect 399474 -2822 399506 -2586
rect 399742 -2822 399826 -2586
rect 400062 -2822 400094 -2586
rect 399474 -7654 400094 -2822
rect 400714 707718 401334 711590
rect 400714 707482 400746 707718
rect 400982 707482 401066 707718
rect 401302 707482 401334 707718
rect 400714 707398 401334 707482
rect 400714 707162 400746 707398
rect 400982 707162 401066 707398
rect 401302 707162 401334 707398
rect 400714 690374 401334 707162
rect 400714 690138 400746 690374
rect 400982 690138 401066 690374
rect 401302 690138 401334 690374
rect 400714 690054 401334 690138
rect 400714 689818 400746 690054
rect 400982 689818 401066 690054
rect 401302 689818 401334 690054
rect 400714 654374 401334 689818
rect 400714 654138 400746 654374
rect 400982 654138 401066 654374
rect 401302 654138 401334 654374
rect 400714 654054 401334 654138
rect 400714 653818 400746 654054
rect 400982 653818 401066 654054
rect 401302 653818 401334 654054
rect 400714 618374 401334 653818
rect 400714 618138 400746 618374
rect 400982 618138 401066 618374
rect 401302 618138 401334 618374
rect 400714 618054 401334 618138
rect 400714 617818 400746 618054
rect 400982 617818 401066 618054
rect 401302 617818 401334 618054
rect 400714 582374 401334 617818
rect 400714 582138 400746 582374
rect 400982 582138 401066 582374
rect 401302 582138 401334 582374
rect 400714 582054 401334 582138
rect 400714 581818 400746 582054
rect 400982 581818 401066 582054
rect 401302 581818 401334 582054
rect 400714 546374 401334 581818
rect 400714 546138 400746 546374
rect 400982 546138 401066 546374
rect 401302 546138 401334 546374
rect 400714 546054 401334 546138
rect 400714 545818 400746 546054
rect 400982 545818 401066 546054
rect 401302 545818 401334 546054
rect 400714 510374 401334 545818
rect 400714 510138 400746 510374
rect 400982 510138 401066 510374
rect 401302 510138 401334 510374
rect 400714 510054 401334 510138
rect 400714 509818 400746 510054
rect 400982 509818 401066 510054
rect 401302 509818 401334 510054
rect 400714 474374 401334 509818
rect 400714 474138 400746 474374
rect 400982 474138 401066 474374
rect 401302 474138 401334 474374
rect 400714 474054 401334 474138
rect 400714 473818 400746 474054
rect 400982 473818 401066 474054
rect 401302 473818 401334 474054
rect 400714 438374 401334 473818
rect 400714 438138 400746 438374
rect 400982 438138 401066 438374
rect 401302 438138 401334 438374
rect 400714 438054 401334 438138
rect 400714 437818 400746 438054
rect 400982 437818 401066 438054
rect 401302 437818 401334 438054
rect 400714 402374 401334 437818
rect 400714 402138 400746 402374
rect 400982 402138 401066 402374
rect 401302 402138 401334 402374
rect 400714 402054 401334 402138
rect 400714 401818 400746 402054
rect 400982 401818 401066 402054
rect 401302 401818 401334 402054
rect 400714 366374 401334 401818
rect 400714 366138 400746 366374
rect 400982 366138 401066 366374
rect 401302 366138 401334 366374
rect 400714 366054 401334 366138
rect 400714 365818 400746 366054
rect 400982 365818 401066 366054
rect 401302 365818 401334 366054
rect 400714 330374 401334 365818
rect 400714 330138 400746 330374
rect 400982 330138 401066 330374
rect 401302 330138 401334 330374
rect 400714 330054 401334 330138
rect 400714 329818 400746 330054
rect 400982 329818 401066 330054
rect 401302 329818 401334 330054
rect 400714 294374 401334 329818
rect 400714 294138 400746 294374
rect 400982 294138 401066 294374
rect 401302 294138 401334 294374
rect 400714 294054 401334 294138
rect 400714 293818 400746 294054
rect 400982 293818 401066 294054
rect 401302 293818 401334 294054
rect 400714 258374 401334 293818
rect 400714 258138 400746 258374
rect 400982 258138 401066 258374
rect 401302 258138 401334 258374
rect 400714 258054 401334 258138
rect 400714 257818 400746 258054
rect 400982 257818 401066 258054
rect 401302 257818 401334 258054
rect 400714 222374 401334 257818
rect 400714 222138 400746 222374
rect 400982 222138 401066 222374
rect 401302 222138 401334 222374
rect 400714 222054 401334 222138
rect 400714 221818 400746 222054
rect 400982 221818 401066 222054
rect 401302 221818 401334 222054
rect 400714 186374 401334 221818
rect 400714 186138 400746 186374
rect 400982 186138 401066 186374
rect 401302 186138 401334 186374
rect 400714 186054 401334 186138
rect 400714 185818 400746 186054
rect 400982 185818 401066 186054
rect 401302 185818 401334 186054
rect 400714 150374 401334 185818
rect 400714 150138 400746 150374
rect 400982 150138 401066 150374
rect 401302 150138 401334 150374
rect 400714 150054 401334 150138
rect 400714 149818 400746 150054
rect 400982 149818 401066 150054
rect 401302 149818 401334 150054
rect 400714 114374 401334 149818
rect 400714 114138 400746 114374
rect 400982 114138 401066 114374
rect 401302 114138 401334 114374
rect 400714 114054 401334 114138
rect 400714 113818 400746 114054
rect 400982 113818 401066 114054
rect 401302 113818 401334 114054
rect 400714 78374 401334 113818
rect 400714 78138 400746 78374
rect 400982 78138 401066 78374
rect 401302 78138 401334 78374
rect 400714 78054 401334 78138
rect 400714 77818 400746 78054
rect 400982 77818 401066 78054
rect 401302 77818 401334 78054
rect 400714 42374 401334 77818
rect 400714 42138 400746 42374
rect 400982 42138 401066 42374
rect 401302 42138 401334 42374
rect 400714 42054 401334 42138
rect 400714 41818 400746 42054
rect 400982 41818 401066 42054
rect 401302 41818 401334 42054
rect 400714 6374 401334 41818
rect 400714 6138 400746 6374
rect 400982 6138 401066 6374
rect 401302 6138 401334 6374
rect 400714 6054 401334 6138
rect 400714 5818 400746 6054
rect 400982 5818 401066 6054
rect 401302 5818 401334 6054
rect 400714 -3226 401334 5818
rect 400714 -3462 400746 -3226
rect 400982 -3462 401066 -3226
rect 401302 -3462 401334 -3226
rect 400714 -3546 401334 -3462
rect 400714 -3782 400746 -3546
rect 400982 -3782 401066 -3546
rect 401302 -3782 401334 -3546
rect 400714 -7654 401334 -3782
rect 401954 708678 402574 711590
rect 401954 708442 401986 708678
rect 402222 708442 402306 708678
rect 402542 708442 402574 708678
rect 401954 708358 402574 708442
rect 401954 708122 401986 708358
rect 402222 708122 402306 708358
rect 402542 708122 402574 708358
rect 401954 691614 402574 708122
rect 401954 691378 401986 691614
rect 402222 691378 402306 691614
rect 402542 691378 402574 691614
rect 401954 691294 402574 691378
rect 401954 691058 401986 691294
rect 402222 691058 402306 691294
rect 402542 691058 402574 691294
rect 401954 655614 402574 691058
rect 401954 655378 401986 655614
rect 402222 655378 402306 655614
rect 402542 655378 402574 655614
rect 401954 655294 402574 655378
rect 401954 655058 401986 655294
rect 402222 655058 402306 655294
rect 402542 655058 402574 655294
rect 401954 619614 402574 655058
rect 401954 619378 401986 619614
rect 402222 619378 402306 619614
rect 402542 619378 402574 619614
rect 401954 619294 402574 619378
rect 401954 619058 401986 619294
rect 402222 619058 402306 619294
rect 402542 619058 402574 619294
rect 401954 583614 402574 619058
rect 401954 583378 401986 583614
rect 402222 583378 402306 583614
rect 402542 583378 402574 583614
rect 401954 583294 402574 583378
rect 401954 583058 401986 583294
rect 402222 583058 402306 583294
rect 402542 583058 402574 583294
rect 401954 547614 402574 583058
rect 401954 547378 401986 547614
rect 402222 547378 402306 547614
rect 402542 547378 402574 547614
rect 401954 547294 402574 547378
rect 401954 547058 401986 547294
rect 402222 547058 402306 547294
rect 402542 547058 402574 547294
rect 401954 511614 402574 547058
rect 401954 511378 401986 511614
rect 402222 511378 402306 511614
rect 402542 511378 402574 511614
rect 401954 511294 402574 511378
rect 401954 511058 401986 511294
rect 402222 511058 402306 511294
rect 402542 511058 402574 511294
rect 401954 475614 402574 511058
rect 401954 475378 401986 475614
rect 402222 475378 402306 475614
rect 402542 475378 402574 475614
rect 401954 475294 402574 475378
rect 401954 475058 401986 475294
rect 402222 475058 402306 475294
rect 402542 475058 402574 475294
rect 401954 439614 402574 475058
rect 401954 439378 401986 439614
rect 402222 439378 402306 439614
rect 402542 439378 402574 439614
rect 401954 439294 402574 439378
rect 401954 439058 401986 439294
rect 402222 439058 402306 439294
rect 402542 439058 402574 439294
rect 401954 403614 402574 439058
rect 401954 403378 401986 403614
rect 402222 403378 402306 403614
rect 402542 403378 402574 403614
rect 401954 403294 402574 403378
rect 401954 403058 401986 403294
rect 402222 403058 402306 403294
rect 402542 403058 402574 403294
rect 401954 367614 402574 403058
rect 401954 367378 401986 367614
rect 402222 367378 402306 367614
rect 402542 367378 402574 367614
rect 401954 367294 402574 367378
rect 401954 367058 401986 367294
rect 402222 367058 402306 367294
rect 402542 367058 402574 367294
rect 401954 331614 402574 367058
rect 401954 331378 401986 331614
rect 402222 331378 402306 331614
rect 402542 331378 402574 331614
rect 401954 331294 402574 331378
rect 401954 331058 401986 331294
rect 402222 331058 402306 331294
rect 402542 331058 402574 331294
rect 401954 295614 402574 331058
rect 401954 295378 401986 295614
rect 402222 295378 402306 295614
rect 402542 295378 402574 295614
rect 401954 295294 402574 295378
rect 401954 295058 401986 295294
rect 402222 295058 402306 295294
rect 402542 295058 402574 295294
rect 401954 259614 402574 295058
rect 401954 259378 401986 259614
rect 402222 259378 402306 259614
rect 402542 259378 402574 259614
rect 401954 259294 402574 259378
rect 401954 259058 401986 259294
rect 402222 259058 402306 259294
rect 402542 259058 402574 259294
rect 401954 223614 402574 259058
rect 401954 223378 401986 223614
rect 402222 223378 402306 223614
rect 402542 223378 402574 223614
rect 401954 223294 402574 223378
rect 401954 223058 401986 223294
rect 402222 223058 402306 223294
rect 402542 223058 402574 223294
rect 401954 187614 402574 223058
rect 401954 187378 401986 187614
rect 402222 187378 402306 187614
rect 402542 187378 402574 187614
rect 401954 187294 402574 187378
rect 401954 187058 401986 187294
rect 402222 187058 402306 187294
rect 402542 187058 402574 187294
rect 401954 151614 402574 187058
rect 401954 151378 401986 151614
rect 402222 151378 402306 151614
rect 402542 151378 402574 151614
rect 401954 151294 402574 151378
rect 401954 151058 401986 151294
rect 402222 151058 402306 151294
rect 402542 151058 402574 151294
rect 401954 115614 402574 151058
rect 401954 115378 401986 115614
rect 402222 115378 402306 115614
rect 402542 115378 402574 115614
rect 401954 115294 402574 115378
rect 401954 115058 401986 115294
rect 402222 115058 402306 115294
rect 402542 115058 402574 115294
rect 401954 79614 402574 115058
rect 401954 79378 401986 79614
rect 402222 79378 402306 79614
rect 402542 79378 402574 79614
rect 401954 79294 402574 79378
rect 401954 79058 401986 79294
rect 402222 79058 402306 79294
rect 402542 79058 402574 79294
rect 401954 43614 402574 79058
rect 401954 43378 401986 43614
rect 402222 43378 402306 43614
rect 402542 43378 402574 43614
rect 401954 43294 402574 43378
rect 401954 43058 401986 43294
rect 402222 43058 402306 43294
rect 402542 43058 402574 43294
rect 401954 7614 402574 43058
rect 401954 7378 401986 7614
rect 402222 7378 402306 7614
rect 402542 7378 402574 7614
rect 401954 7294 402574 7378
rect 401954 7058 401986 7294
rect 402222 7058 402306 7294
rect 402542 7058 402574 7294
rect 401954 -4186 402574 7058
rect 401954 -4422 401986 -4186
rect 402222 -4422 402306 -4186
rect 402542 -4422 402574 -4186
rect 401954 -4506 402574 -4422
rect 401954 -4742 401986 -4506
rect 402222 -4742 402306 -4506
rect 402542 -4742 402574 -4506
rect 401954 -7654 402574 -4742
rect 403194 709638 403814 711590
rect 403194 709402 403226 709638
rect 403462 709402 403546 709638
rect 403782 709402 403814 709638
rect 403194 709318 403814 709402
rect 403194 709082 403226 709318
rect 403462 709082 403546 709318
rect 403782 709082 403814 709318
rect 403194 692854 403814 709082
rect 403194 692618 403226 692854
rect 403462 692618 403546 692854
rect 403782 692618 403814 692854
rect 403194 692534 403814 692618
rect 403194 692298 403226 692534
rect 403462 692298 403546 692534
rect 403782 692298 403814 692534
rect 403194 656854 403814 692298
rect 403194 656618 403226 656854
rect 403462 656618 403546 656854
rect 403782 656618 403814 656854
rect 403194 656534 403814 656618
rect 403194 656298 403226 656534
rect 403462 656298 403546 656534
rect 403782 656298 403814 656534
rect 403194 620854 403814 656298
rect 403194 620618 403226 620854
rect 403462 620618 403546 620854
rect 403782 620618 403814 620854
rect 403194 620534 403814 620618
rect 403194 620298 403226 620534
rect 403462 620298 403546 620534
rect 403782 620298 403814 620534
rect 403194 584854 403814 620298
rect 403194 584618 403226 584854
rect 403462 584618 403546 584854
rect 403782 584618 403814 584854
rect 403194 584534 403814 584618
rect 403194 584298 403226 584534
rect 403462 584298 403546 584534
rect 403782 584298 403814 584534
rect 403194 548854 403814 584298
rect 403194 548618 403226 548854
rect 403462 548618 403546 548854
rect 403782 548618 403814 548854
rect 403194 548534 403814 548618
rect 403194 548298 403226 548534
rect 403462 548298 403546 548534
rect 403782 548298 403814 548534
rect 403194 512854 403814 548298
rect 403194 512618 403226 512854
rect 403462 512618 403546 512854
rect 403782 512618 403814 512854
rect 403194 512534 403814 512618
rect 403194 512298 403226 512534
rect 403462 512298 403546 512534
rect 403782 512298 403814 512534
rect 403194 476854 403814 512298
rect 403194 476618 403226 476854
rect 403462 476618 403546 476854
rect 403782 476618 403814 476854
rect 403194 476534 403814 476618
rect 403194 476298 403226 476534
rect 403462 476298 403546 476534
rect 403782 476298 403814 476534
rect 403194 440854 403814 476298
rect 403194 440618 403226 440854
rect 403462 440618 403546 440854
rect 403782 440618 403814 440854
rect 403194 440534 403814 440618
rect 403194 440298 403226 440534
rect 403462 440298 403546 440534
rect 403782 440298 403814 440534
rect 403194 404854 403814 440298
rect 403194 404618 403226 404854
rect 403462 404618 403546 404854
rect 403782 404618 403814 404854
rect 403194 404534 403814 404618
rect 403194 404298 403226 404534
rect 403462 404298 403546 404534
rect 403782 404298 403814 404534
rect 403194 368854 403814 404298
rect 403194 368618 403226 368854
rect 403462 368618 403546 368854
rect 403782 368618 403814 368854
rect 403194 368534 403814 368618
rect 403194 368298 403226 368534
rect 403462 368298 403546 368534
rect 403782 368298 403814 368534
rect 403194 332854 403814 368298
rect 403194 332618 403226 332854
rect 403462 332618 403546 332854
rect 403782 332618 403814 332854
rect 403194 332534 403814 332618
rect 403194 332298 403226 332534
rect 403462 332298 403546 332534
rect 403782 332298 403814 332534
rect 403194 296854 403814 332298
rect 403194 296618 403226 296854
rect 403462 296618 403546 296854
rect 403782 296618 403814 296854
rect 403194 296534 403814 296618
rect 403194 296298 403226 296534
rect 403462 296298 403546 296534
rect 403782 296298 403814 296534
rect 403194 260854 403814 296298
rect 403194 260618 403226 260854
rect 403462 260618 403546 260854
rect 403782 260618 403814 260854
rect 403194 260534 403814 260618
rect 403194 260298 403226 260534
rect 403462 260298 403546 260534
rect 403782 260298 403814 260534
rect 403194 224854 403814 260298
rect 403194 224618 403226 224854
rect 403462 224618 403546 224854
rect 403782 224618 403814 224854
rect 403194 224534 403814 224618
rect 403194 224298 403226 224534
rect 403462 224298 403546 224534
rect 403782 224298 403814 224534
rect 403194 188854 403814 224298
rect 403194 188618 403226 188854
rect 403462 188618 403546 188854
rect 403782 188618 403814 188854
rect 403194 188534 403814 188618
rect 403194 188298 403226 188534
rect 403462 188298 403546 188534
rect 403782 188298 403814 188534
rect 403194 152854 403814 188298
rect 403194 152618 403226 152854
rect 403462 152618 403546 152854
rect 403782 152618 403814 152854
rect 403194 152534 403814 152618
rect 403194 152298 403226 152534
rect 403462 152298 403546 152534
rect 403782 152298 403814 152534
rect 403194 116854 403814 152298
rect 403194 116618 403226 116854
rect 403462 116618 403546 116854
rect 403782 116618 403814 116854
rect 403194 116534 403814 116618
rect 403194 116298 403226 116534
rect 403462 116298 403546 116534
rect 403782 116298 403814 116534
rect 403194 80854 403814 116298
rect 403194 80618 403226 80854
rect 403462 80618 403546 80854
rect 403782 80618 403814 80854
rect 403194 80534 403814 80618
rect 403194 80298 403226 80534
rect 403462 80298 403546 80534
rect 403782 80298 403814 80534
rect 403194 44854 403814 80298
rect 403194 44618 403226 44854
rect 403462 44618 403546 44854
rect 403782 44618 403814 44854
rect 403194 44534 403814 44618
rect 403194 44298 403226 44534
rect 403462 44298 403546 44534
rect 403782 44298 403814 44534
rect 403194 8854 403814 44298
rect 403194 8618 403226 8854
rect 403462 8618 403546 8854
rect 403782 8618 403814 8854
rect 403194 8534 403814 8618
rect 403194 8298 403226 8534
rect 403462 8298 403546 8534
rect 403782 8298 403814 8534
rect 403194 -5146 403814 8298
rect 403194 -5382 403226 -5146
rect 403462 -5382 403546 -5146
rect 403782 -5382 403814 -5146
rect 403194 -5466 403814 -5382
rect 403194 -5702 403226 -5466
rect 403462 -5702 403546 -5466
rect 403782 -5702 403814 -5466
rect 403194 -7654 403814 -5702
rect 404434 710598 405054 711590
rect 404434 710362 404466 710598
rect 404702 710362 404786 710598
rect 405022 710362 405054 710598
rect 404434 710278 405054 710362
rect 404434 710042 404466 710278
rect 404702 710042 404786 710278
rect 405022 710042 405054 710278
rect 404434 694094 405054 710042
rect 404434 693858 404466 694094
rect 404702 693858 404786 694094
rect 405022 693858 405054 694094
rect 404434 693774 405054 693858
rect 404434 693538 404466 693774
rect 404702 693538 404786 693774
rect 405022 693538 405054 693774
rect 404434 658094 405054 693538
rect 404434 657858 404466 658094
rect 404702 657858 404786 658094
rect 405022 657858 405054 658094
rect 404434 657774 405054 657858
rect 404434 657538 404466 657774
rect 404702 657538 404786 657774
rect 405022 657538 405054 657774
rect 404434 622094 405054 657538
rect 404434 621858 404466 622094
rect 404702 621858 404786 622094
rect 405022 621858 405054 622094
rect 404434 621774 405054 621858
rect 404434 621538 404466 621774
rect 404702 621538 404786 621774
rect 405022 621538 405054 621774
rect 404434 586094 405054 621538
rect 404434 585858 404466 586094
rect 404702 585858 404786 586094
rect 405022 585858 405054 586094
rect 404434 585774 405054 585858
rect 404434 585538 404466 585774
rect 404702 585538 404786 585774
rect 405022 585538 405054 585774
rect 404434 550094 405054 585538
rect 404434 549858 404466 550094
rect 404702 549858 404786 550094
rect 405022 549858 405054 550094
rect 404434 549774 405054 549858
rect 404434 549538 404466 549774
rect 404702 549538 404786 549774
rect 405022 549538 405054 549774
rect 404434 514094 405054 549538
rect 404434 513858 404466 514094
rect 404702 513858 404786 514094
rect 405022 513858 405054 514094
rect 404434 513774 405054 513858
rect 404434 513538 404466 513774
rect 404702 513538 404786 513774
rect 405022 513538 405054 513774
rect 404434 478094 405054 513538
rect 404434 477858 404466 478094
rect 404702 477858 404786 478094
rect 405022 477858 405054 478094
rect 404434 477774 405054 477858
rect 404434 477538 404466 477774
rect 404702 477538 404786 477774
rect 405022 477538 405054 477774
rect 404434 442094 405054 477538
rect 404434 441858 404466 442094
rect 404702 441858 404786 442094
rect 405022 441858 405054 442094
rect 404434 441774 405054 441858
rect 404434 441538 404466 441774
rect 404702 441538 404786 441774
rect 405022 441538 405054 441774
rect 404434 406094 405054 441538
rect 404434 405858 404466 406094
rect 404702 405858 404786 406094
rect 405022 405858 405054 406094
rect 404434 405774 405054 405858
rect 404434 405538 404466 405774
rect 404702 405538 404786 405774
rect 405022 405538 405054 405774
rect 404434 370094 405054 405538
rect 404434 369858 404466 370094
rect 404702 369858 404786 370094
rect 405022 369858 405054 370094
rect 404434 369774 405054 369858
rect 404434 369538 404466 369774
rect 404702 369538 404786 369774
rect 405022 369538 405054 369774
rect 404434 334094 405054 369538
rect 404434 333858 404466 334094
rect 404702 333858 404786 334094
rect 405022 333858 405054 334094
rect 404434 333774 405054 333858
rect 404434 333538 404466 333774
rect 404702 333538 404786 333774
rect 405022 333538 405054 333774
rect 404434 298094 405054 333538
rect 404434 297858 404466 298094
rect 404702 297858 404786 298094
rect 405022 297858 405054 298094
rect 404434 297774 405054 297858
rect 404434 297538 404466 297774
rect 404702 297538 404786 297774
rect 405022 297538 405054 297774
rect 404434 262094 405054 297538
rect 404434 261858 404466 262094
rect 404702 261858 404786 262094
rect 405022 261858 405054 262094
rect 404434 261774 405054 261858
rect 404434 261538 404466 261774
rect 404702 261538 404786 261774
rect 405022 261538 405054 261774
rect 404434 226094 405054 261538
rect 404434 225858 404466 226094
rect 404702 225858 404786 226094
rect 405022 225858 405054 226094
rect 404434 225774 405054 225858
rect 404434 225538 404466 225774
rect 404702 225538 404786 225774
rect 405022 225538 405054 225774
rect 404434 190094 405054 225538
rect 404434 189858 404466 190094
rect 404702 189858 404786 190094
rect 405022 189858 405054 190094
rect 404434 189774 405054 189858
rect 404434 189538 404466 189774
rect 404702 189538 404786 189774
rect 405022 189538 405054 189774
rect 404434 154094 405054 189538
rect 404434 153858 404466 154094
rect 404702 153858 404786 154094
rect 405022 153858 405054 154094
rect 404434 153774 405054 153858
rect 404434 153538 404466 153774
rect 404702 153538 404786 153774
rect 405022 153538 405054 153774
rect 404434 118094 405054 153538
rect 404434 117858 404466 118094
rect 404702 117858 404786 118094
rect 405022 117858 405054 118094
rect 404434 117774 405054 117858
rect 404434 117538 404466 117774
rect 404702 117538 404786 117774
rect 405022 117538 405054 117774
rect 404434 82094 405054 117538
rect 404434 81858 404466 82094
rect 404702 81858 404786 82094
rect 405022 81858 405054 82094
rect 404434 81774 405054 81858
rect 404434 81538 404466 81774
rect 404702 81538 404786 81774
rect 405022 81538 405054 81774
rect 404434 46094 405054 81538
rect 404434 45858 404466 46094
rect 404702 45858 404786 46094
rect 405022 45858 405054 46094
rect 404434 45774 405054 45858
rect 404434 45538 404466 45774
rect 404702 45538 404786 45774
rect 405022 45538 405054 45774
rect 404434 10094 405054 45538
rect 404434 9858 404466 10094
rect 404702 9858 404786 10094
rect 405022 9858 405054 10094
rect 404434 9774 405054 9858
rect 404434 9538 404466 9774
rect 404702 9538 404786 9774
rect 405022 9538 405054 9774
rect 404434 -6106 405054 9538
rect 404434 -6342 404466 -6106
rect 404702 -6342 404786 -6106
rect 405022 -6342 405054 -6106
rect 404434 -6426 405054 -6342
rect 404434 -6662 404466 -6426
rect 404702 -6662 404786 -6426
rect 405022 -6662 405054 -6426
rect 404434 -7654 405054 -6662
rect 405674 711558 406294 711590
rect 405674 711322 405706 711558
rect 405942 711322 406026 711558
rect 406262 711322 406294 711558
rect 405674 711238 406294 711322
rect 405674 711002 405706 711238
rect 405942 711002 406026 711238
rect 406262 711002 406294 711238
rect 405674 695334 406294 711002
rect 405674 695098 405706 695334
rect 405942 695098 406026 695334
rect 406262 695098 406294 695334
rect 405674 695014 406294 695098
rect 405674 694778 405706 695014
rect 405942 694778 406026 695014
rect 406262 694778 406294 695014
rect 405674 659334 406294 694778
rect 405674 659098 405706 659334
rect 405942 659098 406026 659334
rect 406262 659098 406294 659334
rect 405674 659014 406294 659098
rect 405674 658778 405706 659014
rect 405942 658778 406026 659014
rect 406262 658778 406294 659014
rect 405674 623334 406294 658778
rect 405674 623098 405706 623334
rect 405942 623098 406026 623334
rect 406262 623098 406294 623334
rect 405674 623014 406294 623098
rect 405674 622778 405706 623014
rect 405942 622778 406026 623014
rect 406262 622778 406294 623014
rect 405674 587334 406294 622778
rect 405674 587098 405706 587334
rect 405942 587098 406026 587334
rect 406262 587098 406294 587334
rect 405674 587014 406294 587098
rect 405674 586778 405706 587014
rect 405942 586778 406026 587014
rect 406262 586778 406294 587014
rect 405674 551334 406294 586778
rect 405674 551098 405706 551334
rect 405942 551098 406026 551334
rect 406262 551098 406294 551334
rect 405674 551014 406294 551098
rect 405674 550778 405706 551014
rect 405942 550778 406026 551014
rect 406262 550778 406294 551014
rect 405674 515334 406294 550778
rect 405674 515098 405706 515334
rect 405942 515098 406026 515334
rect 406262 515098 406294 515334
rect 405674 515014 406294 515098
rect 405674 514778 405706 515014
rect 405942 514778 406026 515014
rect 406262 514778 406294 515014
rect 405674 479334 406294 514778
rect 405674 479098 405706 479334
rect 405942 479098 406026 479334
rect 406262 479098 406294 479334
rect 405674 479014 406294 479098
rect 405674 478778 405706 479014
rect 405942 478778 406026 479014
rect 406262 478778 406294 479014
rect 405674 443334 406294 478778
rect 405674 443098 405706 443334
rect 405942 443098 406026 443334
rect 406262 443098 406294 443334
rect 405674 443014 406294 443098
rect 405674 442778 405706 443014
rect 405942 442778 406026 443014
rect 406262 442778 406294 443014
rect 405674 407334 406294 442778
rect 405674 407098 405706 407334
rect 405942 407098 406026 407334
rect 406262 407098 406294 407334
rect 405674 407014 406294 407098
rect 405674 406778 405706 407014
rect 405942 406778 406026 407014
rect 406262 406778 406294 407014
rect 405674 371334 406294 406778
rect 405674 371098 405706 371334
rect 405942 371098 406026 371334
rect 406262 371098 406294 371334
rect 405674 371014 406294 371098
rect 405674 370778 405706 371014
rect 405942 370778 406026 371014
rect 406262 370778 406294 371014
rect 405674 335334 406294 370778
rect 405674 335098 405706 335334
rect 405942 335098 406026 335334
rect 406262 335098 406294 335334
rect 405674 335014 406294 335098
rect 405674 334778 405706 335014
rect 405942 334778 406026 335014
rect 406262 334778 406294 335014
rect 405674 299334 406294 334778
rect 405674 299098 405706 299334
rect 405942 299098 406026 299334
rect 406262 299098 406294 299334
rect 405674 299014 406294 299098
rect 405674 298778 405706 299014
rect 405942 298778 406026 299014
rect 406262 298778 406294 299014
rect 405674 263334 406294 298778
rect 405674 263098 405706 263334
rect 405942 263098 406026 263334
rect 406262 263098 406294 263334
rect 405674 263014 406294 263098
rect 405674 262778 405706 263014
rect 405942 262778 406026 263014
rect 406262 262778 406294 263014
rect 405674 227334 406294 262778
rect 405674 227098 405706 227334
rect 405942 227098 406026 227334
rect 406262 227098 406294 227334
rect 405674 227014 406294 227098
rect 405674 226778 405706 227014
rect 405942 226778 406026 227014
rect 406262 226778 406294 227014
rect 405674 191334 406294 226778
rect 405674 191098 405706 191334
rect 405942 191098 406026 191334
rect 406262 191098 406294 191334
rect 405674 191014 406294 191098
rect 405674 190778 405706 191014
rect 405942 190778 406026 191014
rect 406262 190778 406294 191014
rect 405674 155334 406294 190778
rect 405674 155098 405706 155334
rect 405942 155098 406026 155334
rect 406262 155098 406294 155334
rect 405674 155014 406294 155098
rect 405674 154778 405706 155014
rect 405942 154778 406026 155014
rect 406262 154778 406294 155014
rect 405674 119334 406294 154778
rect 405674 119098 405706 119334
rect 405942 119098 406026 119334
rect 406262 119098 406294 119334
rect 405674 119014 406294 119098
rect 405674 118778 405706 119014
rect 405942 118778 406026 119014
rect 406262 118778 406294 119014
rect 405674 83334 406294 118778
rect 405674 83098 405706 83334
rect 405942 83098 406026 83334
rect 406262 83098 406294 83334
rect 405674 83014 406294 83098
rect 405674 82778 405706 83014
rect 405942 82778 406026 83014
rect 406262 82778 406294 83014
rect 405674 47334 406294 82778
rect 405674 47098 405706 47334
rect 405942 47098 406026 47334
rect 406262 47098 406294 47334
rect 405674 47014 406294 47098
rect 405674 46778 405706 47014
rect 405942 46778 406026 47014
rect 406262 46778 406294 47014
rect 405674 11334 406294 46778
rect 405674 11098 405706 11334
rect 405942 11098 406026 11334
rect 406262 11098 406294 11334
rect 405674 11014 406294 11098
rect 405674 10778 405706 11014
rect 405942 10778 406026 11014
rect 406262 10778 406294 11014
rect 405674 -7066 406294 10778
rect 405674 -7302 405706 -7066
rect 405942 -7302 406026 -7066
rect 406262 -7302 406294 -7066
rect 405674 -7386 406294 -7302
rect 405674 -7622 405706 -7386
rect 405942 -7622 406026 -7386
rect 406262 -7622 406294 -7386
rect 405674 -7654 406294 -7622
rect 432994 704838 433614 711590
rect 432994 704602 433026 704838
rect 433262 704602 433346 704838
rect 433582 704602 433614 704838
rect 432994 704518 433614 704602
rect 432994 704282 433026 704518
rect 433262 704282 433346 704518
rect 433582 704282 433614 704518
rect 432994 686654 433614 704282
rect 432994 686418 433026 686654
rect 433262 686418 433346 686654
rect 433582 686418 433614 686654
rect 432994 686334 433614 686418
rect 432994 686098 433026 686334
rect 433262 686098 433346 686334
rect 433582 686098 433614 686334
rect 432994 650654 433614 686098
rect 432994 650418 433026 650654
rect 433262 650418 433346 650654
rect 433582 650418 433614 650654
rect 432994 650334 433614 650418
rect 432994 650098 433026 650334
rect 433262 650098 433346 650334
rect 433582 650098 433614 650334
rect 432994 614654 433614 650098
rect 432994 614418 433026 614654
rect 433262 614418 433346 614654
rect 433582 614418 433614 614654
rect 432994 614334 433614 614418
rect 432994 614098 433026 614334
rect 433262 614098 433346 614334
rect 433582 614098 433614 614334
rect 432994 578654 433614 614098
rect 432994 578418 433026 578654
rect 433262 578418 433346 578654
rect 433582 578418 433614 578654
rect 432994 578334 433614 578418
rect 432994 578098 433026 578334
rect 433262 578098 433346 578334
rect 433582 578098 433614 578334
rect 432994 542654 433614 578098
rect 432994 542418 433026 542654
rect 433262 542418 433346 542654
rect 433582 542418 433614 542654
rect 432994 542334 433614 542418
rect 432994 542098 433026 542334
rect 433262 542098 433346 542334
rect 433582 542098 433614 542334
rect 432994 506654 433614 542098
rect 432994 506418 433026 506654
rect 433262 506418 433346 506654
rect 433582 506418 433614 506654
rect 432994 506334 433614 506418
rect 432994 506098 433026 506334
rect 433262 506098 433346 506334
rect 433582 506098 433614 506334
rect 432994 470654 433614 506098
rect 432994 470418 433026 470654
rect 433262 470418 433346 470654
rect 433582 470418 433614 470654
rect 432994 470334 433614 470418
rect 432994 470098 433026 470334
rect 433262 470098 433346 470334
rect 433582 470098 433614 470334
rect 432994 434654 433614 470098
rect 432994 434418 433026 434654
rect 433262 434418 433346 434654
rect 433582 434418 433614 434654
rect 432994 434334 433614 434418
rect 432994 434098 433026 434334
rect 433262 434098 433346 434334
rect 433582 434098 433614 434334
rect 432994 398654 433614 434098
rect 432994 398418 433026 398654
rect 433262 398418 433346 398654
rect 433582 398418 433614 398654
rect 432994 398334 433614 398418
rect 432994 398098 433026 398334
rect 433262 398098 433346 398334
rect 433582 398098 433614 398334
rect 432994 362654 433614 398098
rect 432994 362418 433026 362654
rect 433262 362418 433346 362654
rect 433582 362418 433614 362654
rect 432994 362334 433614 362418
rect 432994 362098 433026 362334
rect 433262 362098 433346 362334
rect 433582 362098 433614 362334
rect 432994 326654 433614 362098
rect 432994 326418 433026 326654
rect 433262 326418 433346 326654
rect 433582 326418 433614 326654
rect 432994 326334 433614 326418
rect 432994 326098 433026 326334
rect 433262 326098 433346 326334
rect 433582 326098 433614 326334
rect 432994 290654 433614 326098
rect 432994 290418 433026 290654
rect 433262 290418 433346 290654
rect 433582 290418 433614 290654
rect 432994 290334 433614 290418
rect 432994 290098 433026 290334
rect 433262 290098 433346 290334
rect 433582 290098 433614 290334
rect 432994 254654 433614 290098
rect 432994 254418 433026 254654
rect 433262 254418 433346 254654
rect 433582 254418 433614 254654
rect 432994 254334 433614 254418
rect 432994 254098 433026 254334
rect 433262 254098 433346 254334
rect 433582 254098 433614 254334
rect 432994 218654 433614 254098
rect 432994 218418 433026 218654
rect 433262 218418 433346 218654
rect 433582 218418 433614 218654
rect 432994 218334 433614 218418
rect 432994 218098 433026 218334
rect 433262 218098 433346 218334
rect 433582 218098 433614 218334
rect 432994 182654 433614 218098
rect 432994 182418 433026 182654
rect 433262 182418 433346 182654
rect 433582 182418 433614 182654
rect 432994 182334 433614 182418
rect 432994 182098 433026 182334
rect 433262 182098 433346 182334
rect 433582 182098 433614 182334
rect 432994 146654 433614 182098
rect 432994 146418 433026 146654
rect 433262 146418 433346 146654
rect 433582 146418 433614 146654
rect 432994 146334 433614 146418
rect 432994 146098 433026 146334
rect 433262 146098 433346 146334
rect 433582 146098 433614 146334
rect 432994 110654 433614 146098
rect 432994 110418 433026 110654
rect 433262 110418 433346 110654
rect 433582 110418 433614 110654
rect 432994 110334 433614 110418
rect 432994 110098 433026 110334
rect 433262 110098 433346 110334
rect 433582 110098 433614 110334
rect 432994 74654 433614 110098
rect 432994 74418 433026 74654
rect 433262 74418 433346 74654
rect 433582 74418 433614 74654
rect 432994 74334 433614 74418
rect 432994 74098 433026 74334
rect 433262 74098 433346 74334
rect 433582 74098 433614 74334
rect 432994 38654 433614 74098
rect 432994 38418 433026 38654
rect 433262 38418 433346 38654
rect 433582 38418 433614 38654
rect 432994 38334 433614 38418
rect 432994 38098 433026 38334
rect 433262 38098 433346 38334
rect 433582 38098 433614 38334
rect 432994 2654 433614 38098
rect 432994 2418 433026 2654
rect 433262 2418 433346 2654
rect 433582 2418 433614 2654
rect 432994 2334 433614 2418
rect 432994 2098 433026 2334
rect 433262 2098 433346 2334
rect 433582 2098 433614 2334
rect 432994 -346 433614 2098
rect 432994 -582 433026 -346
rect 433262 -582 433346 -346
rect 433582 -582 433614 -346
rect 432994 -666 433614 -582
rect 432994 -902 433026 -666
rect 433262 -902 433346 -666
rect 433582 -902 433614 -666
rect 432994 -7654 433614 -902
rect 434234 705798 434854 711590
rect 434234 705562 434266 705798
rect 434502 705562 434586 705798
rect 434822 705562 434854 705798
rect 434234 705478 434854 705562
rect 434234 705242 434266 705478
rect 434502 705242 434586 705478
rect 434822 705242 434854 705478
rect 434234 687894 434854 705242
rect 434234 687658 434266 687894
rect 434502 687658 434586 687894
rect 434822 687658 434854 687894
rect 434234 687574 434854 687658
rect 434234 687338 434266 687574
rect 434502 687338 434586 687574
rect 434822 687338 434854 687574
rect 434234 651894 434854 687338
rect 434234 651658 434266 651894
rect 434502 651658 434586 651894
rect 434822 651658 434854 651894
rect 434234 651574 434854 651658
rect 434234 651338 434266 651574
rect 434502 651338 434586 651574
rect 434822 651338 434854 651574
rect 434234 615894 434854 651338
rect 434234 615658 434266 615894
rect 434502 615658 434586 615894
rect 434822 615658 434854 615894
rect 434234 615574 434854 615658
rect 434234 615338 434266 615574
rect 434502 615338 434586 615574
rect 434822 615338 434854 615574
rect 434234 579894 434854 615338
rect 434234 579658 434266 579894
rect 434502 579658 434586 579894
rect 434822 579658 434854 579894
rect 434234 579574 434854 579658
rect 434234 579338 434266 579574
rect 434502 579338 434586 579574
rect 434822 579338 434854 579574
rect 434234 543894 434854 579338
rect 434234 543658 434266 543894
rect 434502 543658 434586 543894
rect 434822 543658 434854 543894
rect 434234 543574 434854 543658
rect 434234 543338 434266 543574
rect 434502 543338 434586 543574
rect 434822 543338 434854 543574
rect 434234 507894 434854 543338
rect 434234 507658 434266 507894
rect 434502 507658 434586 507894
rect 434822 507658 434854 507894
rect 434234 507574 434854 507658
rect 434234 507338 434266 507574
rect 434502 507338 434586 507574
rect 434822 507338 434854 507574
rect 434234 471894 434854 507338
rect 434234 471658 434266 471894
rect 434502 471658 434586 471894
rect 434822 471658 434854 471894
rect 434234 471574 434854 471658
rect 434234 471338 434266 471574
rect 434502 471338 434586 471574
rect 434822 471338 434854 471574
rect 434234 435894 434854 471338
rect 434234 435658 434266 435894
rect 434502 435658 434586 435894
rect 434822 435658 434854 435894
rect 434234 435574 434854 435658
rect 434234 435338 434266 435574
rect 434502 435338 434586 435574
rect 434822 435338 434854 435574
rect 434234 399894 434854 435338
rect 434234 399658 434266 399894
rect 434502 399658 434586 399894
rect 434822 399658 434854 399894
rect 434234 399574 434854 399658
rect 434234 399338 434266 399574
rect 434502 399338 434586 399574
rect 434822 399338 434854 399574
rect 434234 363894 434854 399338
rect 434234 363658 434266 363894
rect 434502 363658 434586 363894
rect 434822 363658 434854 363894
rect 434234 363574 434854 363658
rect 434234 363338 434266 363574
rect 434502 363338 434586 363574
rect 434822 363338 434854 363574
rect 434234 327894 434854 363338
rect 434234 327658 434266 327894
rect 434502 327658 434586 327894
rect 434822 327658 434854 327894
rect 434234 327574 434854 327658
rect 434234 327338 434266 327574
rect 434502 327338 434586 327574
rect 434822 327338 434854 327574
rect 434234 291894 434854 327338
rect 434234 291658 434266 291894
rect 434502 291658 434586 291894
rect 434822 291658 434854 291894
rect 434234 291574 434854 291658
rect 434234 291338 434266 291574
rect 434502 291338 434586 291574
rect 434822 291338 434854 291574
rect 434234 255894 434854 291338
rect 434234 255658 434266 255894
rect 434502 255658 434586 255894
rect 434822 255658 434854 255894
rect 434234 255574 434854 255658
rect 434234 255338 434266 255574
rect 434502 255338 434586 255574
rect 434822 255338 434854 255574
rect 434234 219894 434854 255338
rect 434234 219658 434266 219894
rect 434502 219658 434586 219894
rect 434822 219658 434854 219894
rect 434234 219574 434854 219658
rect 434234 219338 434266 219574
rect 434502 219338 434586 219574
rect 434822 219338 434854 219574
rect 434234 183894 434854 219338
rect 434234 183658 434266 183894
rect 434502 183658 434586 183894
rect 434822 183658 434854 183894
rect 434234 183574 434854 183658
rect 434234 183338 434266 183574
rect 434502 183338 434586 183574
rect 434822 183338 434854 183574
rect 434234 147894 434854 183338
rect 434234 147658 434266 147894
rect 434502 147658 434586 147894
rect 434822 147658 434854 147894
rect 434234 147574 434854 147658
rect 434234 147338 434266 147574
rect 434502 147338 434586 147574
rect 434822 147338 434854 147574
rect 434234 111894 434854 147338
rect 434234 111658 434266 111894
rect 434502 111658 434586 111894
rect 434822 111658 434854 111894
rect 434234 111574 434854 111658
rect 434234 111338 434266 111574
rect 434502 111338 434586 111574
rect 434822 111338 434854 111574
rect 434234 75894 434854 111338
rect 434234 75658 434266 75894
rect 434502 75658 434586 75894
rect 434822 75658 434854 75894
rect 434234 75574 434854 75658
rect 434234 75338 434266 75574
rect 434502 75338 434586 75574
rect 434822 75338 434854 75574
rect 434234 39894 434854 75338
rect 434234 39658 434266 39894
rect 434502 39658 434586 39894
rect 434822 39658 434854 39894
rect 434234 39574 434854 39658
rect 434234 39338 434266 39574
rect 434502 39338 434586 39574
rect 434822 39338 434854 39574
rect 434234 3894 434854 39338
rect 434234 3658 434266 3894
rect 434502 3658 434586 3894
rect 434822 3658 434854 3894
rect 434234 3574 434854 3658
rect 434234 3338 434266 3574
rect 434502 3338 434586 3574
rect 434822 3338 434854 3574
rect 434234 -1306 434854 3338
rect 434234 -1542 434266 -1306
rect 434502 -1542 434586 -1306
rect 434822 -1542 434854 -1306
rect 434234 -1626 434854 -1542
rect 434234 -1862 434266 -1626
rect 434502 -1862 434586 -1626
rect 434822 -1862 434854 -1626
rect 434234 -7654 434854 -1862
rect 435474 706758 436094 711590
rect 435474 706522 435506 706758
rect 435742 706522 435826 706758
rect 436062 706522 436094 706758
rect 435474 706438 436094 706522
rect 435474 706202 435506 706438
rect 435742 706202 435826 706438
rect 436062 706202 436094 706438
rect 435474 689134 436094 706202
rect 435474 688898 435506 689134
rect 435742 688898 435826 689134
rect 436062 688898 436094 689134
rect 435474 688814 436094 688898
rect 435474 688578 435506 688814
rect 435742 688578 435826 688814
rect 436062 688578 436094 688814
rect 435474 653134 436094 688578
rect 435474 652898 435506 653134
rect 435742 652898 435826 653134
rect 436062 652898 436094 653134
rect 435474 652814 436094 652898
rect 435474 652578 435506 652814
rect 435742 652578 435826 652814
rect 436062 652578 436094 652814
rect 435474 617134 436094 652578
rect 435474 616898 435506 617134
rect 435742 616898 435826 617134
rect 436062 616898 436094 617134
rect 435474 616814 436094 616898
rect 435474 616578 435506 616814
rect 435742 616578 435826 616814
rect 436062 616578 436094 616814
rect 435474 581134 436094 616578
rect 435474 580898 435506 581134
rect 435742 580898 435826 581134
rect 436062 580898 436094 581134
rect 435474 580814 436094 580898
rect 435474 580578 435506 580814
rect 435742 580578 435826 580814
rect 436062 580578 436094 580814
rect 435474 545134 436094 580578
rect 435474 544898 435506 545134
rect 435742 544898 435826 545134
rect 436062 544898 436094 545134
rect 435474 544814 436094 544898
rect 435474 544578 435506 544814
rect 435742 544578 435826 544814
rect 436062 544578 436094 544814
rect 435474 509134 436094 544578
rect 435474 508898 435506 509134
rect 435742 508898 435826 509134
rect 436062 508898 436094 509134
rect 435474 508814 436094 508898
rect 435474 508578 435506 508814
rect 435742 508578 435826 508814
rect 436062 508578 436094 508814
rect 435474 473134 436094 508578
rect 435474 472898 435506 473134
rect 435742 472898 435826 473134
rect 436062 472898 436094 473134
rect 435474 472814 436094 472898
rect 435474 472578 435506 472814
rect 435742 472578 435826 472814
rect 436062 472578 436094 472814
rect 435474 437134 436094 472578
rect 435474 436898 435506 437134
rect 435742 436898 435826 437134
rect 436062 436898 436094 437134
rect 435474 436814 436094 436898
rect 435474 436578 435506 436814
rect 435742 436578 435826 436814
rect 436062 436578 436094 436814
rect 435474 401134 436094 436578
rect 435474 400898 435506 401134
rect 435742 400898 435826 401134
rect 436062 400898 436094 401134
rect 435474 400814 436094 400898
rect 435474 400578 435506 400814
rect 435742 400578 435826 400814
rect 436062 400578 436094 400814
rect 435474 365134 436094 400578
rect 435474 364898 435506 365134
rect 435742 364898 435826 365134
rect 436062 364898 436094 365134
rect 435474 364814 436094 364898
rect 435474 364578 435506 364814
rect 435742 364578 435826 364814
rect 436062 364578 436094 364814
rect 435474 329134 436094 364578
rect 435474 328898 435506 329134
rect 435742 328898 435826 329134
rect 436062 328898 436094 329134
rect 435474 328814 436094 328898
rect 435474 328578 435506 328814
rect 435742 328578 435826 328814
rect 436062 328578 436094 328814
rect 435474 293134 436094 328578
rect 435474 292898 435506 293134
rect 435742 292898 435826 293134
rect 436062 292898 436094 293134
rect 435474 292814 436094 292898
rect 435474 292578 435506 292814
rect 435742 292578 435826 292814
rect 436062 292578 436094 292814
rect 435474 257134 436094 292578
rect 435474 256898 435506 257134
rect 435742 256898 435826 257134
rect 436062 256898 436094 257134
rect 435474 256814 436094 256898
rect 435474 256578 435506 256814
rect 435742 256578 435826 256814
rect 436062 256578 436094 256814
rect 435474 221134 436094 256578
rect 435474 220898 435506 221134
rect 435742 220898 435826 221134
rect 436062 220898 436094 221134
rect 435474 220814 436094 220898
rect 435474 220578 435506 220814
rect 435742 220578 435826 220814
rect 436062 220578 436094 220814
rect 435474 185134 436094 220578
rect 435474 184898 435506 185134
rect 435742 184898 435826 185134
rect 436062 184898 436094 185134
rect 435474 184814 436094 184898
rect 435474 184578 435506 184814
rect 435742 184578 435826 184814
rect 436062 184578 436094 184814
rect 435474 149134 436094 184578
rect 435474 148898 435506 149134
rect 435742 148898 435826 149134
rect 436062 148898 436094 149134
rect 435474 148814 436094 148898
rect 435474 148578 435506 148814
rect 435742 148578 435826 148814
rect 436062 148578 436094 148814
rect 435474 113134 436094 148578
rect 435474 112898 435506 113134
rect 435742 112898 435826 113134
rect 436062 112898 436094 113134
rect 435474 112814 436094 112898
rect 435474 112578 435506 112814
rect 435742 112578 435826 112814
rect 436062 112578 436094 112814
rect 435474 77134 436094 112578
rect 435474 76898 435506 77134
rect 435742 76898 435826 77134
rect 436062 76898 436094 77134
rect 435474 76814 436094 76898
rect 435474 76578 435506 76814
rect 435742 76578 435826 76814
rect 436062 76578 436094 76814
rect 435474 41134 436094 76578
rect 435474 40898 435506 41134
rect 435742 40898 435826 41134
rect 436062 40898 436094 41134
rect 435474 40814 436094 40898
rect 435474 40578 435506 40814
rect 435742 40578 435826 40814
rect 436062 40578 436094 40814
rect 435474 5134 436094 40578
rect 435474 4898 435506 5134
rect 435742 4898 435826 5134
rect 436062 4898 436094 5134
rect 435474 4814 436094 4898
rect 435474 4578 435506 4814
rect 435742 4578 435826 4814
rect 436062 4578 436094 4814
rect 435474 -2266 436094 4578
rect 435474 -2502 435506 -2266
rect 435742 -2502 435826 -2266
rect 436062 -2502 436094 -2266
rect 435474 -2586 436094 -2502
rect 435474 -2822 435506 -2586
rect 435742 -2822 435826 -2586
rect 436062 -2822 436094 -2586
rect 435474 -7654 436094 -2822
rect 436714 707718 437334 711590
rect 436714 707482 436746 707718
rect 436982 707482 437066 707718
rect 437302 707482 437334 707718
rect 436714 707398 437334 707482
rect 436714 707162 436746 707398
rect 436982 707162 437066 707398
rect 437302 707162 437334 707398
rect 436714 690374 437334 707162
rect 436714 690138 436746 690374
rect 436982 690138 437066 690374
rect 437302 690138 437334 690374
rect 436714 690054 437334 690138
rect 436714 689818 436746 690054
rect 436982 689818 437066 690054
rect 437302 689818 437334 690054
rect 436714 654374 437334 689818
rect 436714 654138 436746 654374
rect 436982 654138 437066 654374
rect 437302 654138 437334 654374
rect 436714 654054 437334 654138
rect 436714 653818 436746 654054
rect 436982 653818 437066 654054
rect 437302 653818 437334 654054
rect 436714 618374 437334 653818
rect 436714 618138 436746 618374
rect 436982 618138 437066 618374
rect 437302 618138 437334 618374
rect 436714 618054 437334 618138
rect 436714 617818 436746 618054
rect 436982 617818 437066 618054
rect 437302 617818 437334 618054
rect 436714 582374 437334 617818
rect 436714 582138 436746 582374
rect 436982 582138 437066 582374
rect 437302 582138 437334 582374
rect 436714 582054 437334 582138
rect 436714 581818 436746 582054
rect 436982 581818 437066 582054
rect 437302 581818 437334 582054
rect 436714 546374 437334 581818
rect 436714 546138 436746 546374
rect 436982 546138 437066 546374
rect 437302 546138 437334 546374
rect 436714 546054 437334 546138
rect 436714 545818 436746 546054
rect 436982 545818 437066 546054
rect 437302 545818 437334 546054
rect 436714 510374 437334 545818
rect 436714 510138 436746 510374
rect 436982 510138 437066 510374
rect 437302 510138 437334 510374
rect 436714 510054 437334 510138
rect 436714 509818 436746 510054
rect 436982 509818 437066 510054
rect 437302 509818 437334 510054
rect 436714 474374 437334 509818
rect 436714 474138 436746 474374
rect 436982 474138 437066 474374
rect 437302 474138 437334 474374
rect 436714 474054 437334 474138
rect 436714 473818 436746 474054
rect 436982 473818 437066 474054
rect 437302 473818 437334 474054
rect 436714 438374 437334 473818
rect 436714 438138 436746 438374
rect 436982 438138 437066 438374
rect 437302 438138 437334 438374
rect 436714 438054 437334 438138
rect 436714 437818 436746 438054
rect 436982 437818 437066 438054
rect 437302 437818 437334 438054
rect 436714 402374 437334 437818
rect 436714 402138 436746 402374
rect 436982 402138 437066 402374
rect 437302 402138 437334 402374
rect 436714 402054 437334 402138
rect 436714 401818 436746 402054
rect 436982 401818 437066 402054
rect 437302 401818 437334 402054
rect 436714 366374 437334 401818
rect 436714 366138 436746 366374
rect 436982 366138 437066 366374
rect 437302 366138 437334 366374
rect 436714 366054 437334 366138
rect 436714 365818 436746 366054
rect 436982 365818 437066 366054
rect 437302 365818 437334 366054
rect 436714 330374 437334 365818
rect 436714 330138 436746 330374
rect 436982 330138 437066 330374
rect 437302 330138 437334 330374
rect 436714 330054 437334 330138
rect 436714 329818 436746 330054
rect 436982 329818 437066 330054
rect 437302 329818 437334 330054
rect 436714 294374 437334 329818
rect 436714 294138 436746 294374
rect 436982 294138 437066 294374
rect 437302 294138 437334 294374
rect 436714 294054 437334 294138
rect 436714 293818 436746 294054
rect 436982 293818 437066 294054
rect 437302 293818 437334 294054
rect 436714 258374 437334 293818
rect 436714 258138 436746 258374
rect 436982 258138 437066 258374
rect 437302 258138 437334 258374
rect 436714 258054 437334 258138
rect 436714 257818 436746 258054
rect 436982 257818 437066 258054
rect 437302 257818 437334 258054
rect 436714 222374 437334 257818
rect 436714 222138 436746 222374
rect 436982 222138 437066 222374
rect 437302 222138 437334 222374
rect 436714 222054 437334 222138
rect 436714 221818 436746 222054
rect 436982 221818 437066 222054
rect 437302 221818 437334 222054
rect 436714 186374 437334 221818
rect 436714 186138 436746 186374
rect 436982 186138 437066 186374
rect 437302 186138 437334 186374
rect 436714 186054 437334 186138
rect 436714 185818 436746 186054
rect 436982 185818 437066 186054
rect 437302 185818 437334 186054
rect 436714 150374 437334 185818
rect 436714 150138 436746 150374
rect 436982 150138 437066 150374
rect 437302 150138 437334 150374
rect 436714 150054 437334 150138
rect 436714 149818 436746 150054
rect 436982 149818 437066 150054
rect 437302 149818 437334 150054
rect 436714 114374 437334 149818
rect 436714 114138 436746 114374
rect 436982 114138 437066 114374
rect 437302 114138 437334 114374
rect 436714 114054 437334 114138
rect 436714 113818 436746 114054
rect 436982 113818 437066 114054
rect 437302 113818 437334 114054
rect 436714 78374 437334 113818
rect 436714 78138 436746 78374
rect 436982 78138 437066 78374
rect 437302 78138 437334 78374
rect 436714 78054 437334 78138
rect 436714 77818 436746 78054
rect 436982 77818 437066 78054
rect 437302 77818 437334 78054
rect 436714 42374 437334 77818
rect 436714 42138 436746 42374
rect 436982 42138 437066 42374
rect 437302 42138 437334 42374
rect 436714 42054 437334 42138
rect 436714 41818 436746 42054
rect 436982 41818 437066 42054
rect 437302 41818 437334 42054
rect 436714 6374 437334 41818
rect 436714 6138 436746 6374
rect 436982 6138 437066 6374
rect 437302 6138 437334 6374
rect 436714 6054 437334 6138
rect 436714 5818 436746 6054
rect 436982 5818 437066 6054
rect 437302 5818 437334 6054
rect 436714 -3226 437334 5818
rect 436714 -3462 436746 -3226
rect 436982 -3462 437066 -3226
rect 437302 -3462 437334 -3226
rect 436714 -3546 437334 -3462
rect 436714 -3782 436746 -3546
rect 436982 -3782 437066 -3546
rect 437302 -3782 437334 -3546
rect 436714 -7654 437334 -3782
rect 437954 708678 438574 711590
rect 437954 708442 437986 708678
rect 438222 708442 438306 708678
rect 438542 708442 438574 708678
rect 437954 708358 438574 708442
rect 437954 708122 437986 708358
rect 438222 708122 438306 708358
rect 438542 708122 438574 708358
rect 437954 691614 438574 708122
rect 437954 691378 437986 691614
rect 438222 691378 438306 691614
rect 438542 691378 438574 691614
rect 437954 691294 438574 691378
rect 437954 691058 437986 691294
rect 438222 691058 438306 691294
rect 438542 691058 438574 691294
rect 437954 655614 438574 691058
rect 437954 655378 437986 655614
rect 438222 655378 438306 655614
rect 438542 655378 438574 655614
rect 437954 655294 438574 655378
rect 437954 655058 437986 655294
rect 438222 655058 438306 655294
rect 438542 655058 438574 655294
rect 437954 619614 438574 655058
rect 437954 619378 437986 619614
rect 438222 619378 438306 619614
rect 438542 619378 438574 619614
rect 437954 619294 438574 619378
rect 437954 619058 437986 619294
rect 438222 619058 438306 619294
rect 438542 619058 438574 619294
rect 437954 583614 438574 619058
rect 437954 583378 437986 583614
rect 438222 583378 438306 583614
rect 438542 583378 438574 583614
rect 437954 583294 438574 583378
rect 437954 583058 437986 583294
rect 438222 583058 438306 583294
rect 438542 583058 438574 583294
rect 437954 547614 438574 583058
rect 437954 547378 437986 547614
rect 438222 547378 438306 547614
rect 438542 547378 438574 547614
rect 437954 547294 438574 547378
rect 437954 547058 437986 547294
rect 438222 547058 438306 547294
rect 438542 547058 438574 547294
rect 437954 511614 438574 547058
rect 437954 511378 437986 511614
rect 438222 511378 438306 511614
rect 438542 511378 438574 511614
rect 437954 511294 438574 511378
rect 437954 511058 437986 511294
rect 438222 511058 438306 511294
rect 438542 511058 438574 511294
rect 437954 475614 438574 511058
rect 437954 475378 437986 475614
rect 438222 475378 438306 475614
rect 438542 475378 438574 475614
rect 437954 475294 438574 475378
rect 437954 475058 437986 475294
rect 438222 475058 438306 475294
rect 438542 475058 438574 475294
rect 437954 439614 438574 475058
rect 437954 439378 437986 439614
rect 438222 439378 438306 439614
rect 438542 439378 438574 439614
rect 437954 439294 438574 439378
rect 437954 439058 437986 439294
rect 438222 439058 438306 439294
rect 438542 439058 438574 439294
rect 437954 403614 438574 439058
rect 437954 403378 437986 403614
rect 438222 403378 438306 403614
rect 438542 403378 438574 403614
rect 437954 403294 438574 403378
rect 437954 403058 437986 403294
rect 438222 403058 438306 403294
rect 438542 403058 438574 403294
rect 437954 367614 438574 403058
rect 437954 367378 437986 367614
rect 438222 367378 438306 367614
rect 438542 367378 438574 367614
rect 437954 367294 438574 367378
rect 437954 367058 437986 367294
rect 438222 367058 438306 367294
rect 438542 367058 438574 367294
rect 437954 331614 438574 367058
rect 437954 331378 437986 331614
rect 438222 331378 438306 331614
rect 438542 331378 438574 331614
rect 437954 331294 438574 331378
rect 437954 331058 437986 331294
rect 438222 331058 438306 331294
rect 438542 331058 438574 331294
rect 437954 295614 438574 331058
rect 437954 295378 437986 295614
rect 438222 295378 438306 295614
rect 438542 295378 438574 295614
rect 437954 295294 438574 295378
rect 437954 295058 437986 295294
rect 438222 295058 438306 295294
rect 438542 295058 438574 295294
rect 437954 259614 438574 295058
rect 437954 259378 437986 259614
rect 438222 259378 438306 259614
rect 438542 259378 438574 259614
rect 437954 259294 438574 259378
rect 437954 259058 437986 259294
rect 438222 259058 438306 259294
rect 438542 259058 438574 259294
rect 437954 223614 438574 259058
rect 437954 223378 437986 223614
rect 438222 223378 438306 223614
rect 438542 223378 438574 223614
rect 437954 223294 438574 223378
rect 437954 223058 437986 223294
rect 438222 223058 438306 223294
rect 438542 223058 438574 223294
rect 437954 187614 438574 223058
rect 437954 187378 437986 187614
rect 438222 187378 438306 187614
rect 438542 187378 438574 187614
rect 437954 187294 438574 187378
rect 437954 187058 437986 187294
rect 438222 187058 438306 187294
rect 438542 187058 438574 187294
rect 437954 151614 438574 187058
rect 437954 151378 437986 151614
rect 438222 151378 438306 151614
rect 438542 151378 438574 151614
rect 437954 151294 438574 151378
rect 437954 151058 437986 151294
rect 438222 151058 438306 151294
rect 438542 151058 438574 151294
rect 437954 115614 438574 151058
rect 437954 115378 437986 115614
rect 438222 115378 438306 115614
rect 438542 115378 438574 115614
rect 437954 115294 438574 115378
rect 437954 115058 437986 115294
rect 438222 115058 438306 115294
rect 438542 115058 438574 115294
rect 437954 79614 438574 115058
rect 437954 79378 437986 79614
rect 438222 79378 438306 79614
rect 438542 79378 438574 79614
rect 437954 79294 438574 79378
rect 437954 79058 437986 79294
rect 438222 79058 438306 79294
rect 438542 79058 438574 79294
rect 437954 43614 438574 79058
rect 437954 43378 437986 43614
rect 438222 43378 438306 43614
rect 438542 43378 438574 43614
rect 437954 43294 438574 43378
rect 437954 43058 437986 43294
rect 438222 43058 438306 43294
rect 438542 43058 438574 43294
rect 437954 7614 438574 43058
rect 437954 7378 437986 7614
rect 438222 7378 438306 7614
rect 438542 7378 438574 7614
rect 437954 7294 438574 7378
rect 437954 7058 437986 7294
rect 438222 7058 438306 7294
rect 438542 7058 438574 7294
rect 437954 -4186 438574 7058
rect 437954 -4422 437986 -4186
rect 438222 -4422 438306 -4186
rect 438542 -4422 438574 -4186
rect 437954 -4506 438574 -4422
rect 437954 -4742 437986 -4506
rect 438222 -4742 438306 -4506
rect 438542 -4742 438574 -4506
rect 437954 -7654 438574 -4742
rect 439194 709638 439814 711590
rect 439194 709402 439226 709638
rect 439462 709402 439546 709638
rect 439782 709402 439814 709638
rect 439194 709318 439814 709402
rect 439194 709082 439226 709318
rect 439462 709082 439546 709318
rect 439782 709082 439814 709318
rect 439194 692854 439814 709082
rect 439194 692618 439226 692854
rect 439462 692618 439546 692854
rect 439782 692618 439814 692854
rect 439194 692534 439814 692618
rect 439194 692298 439226 692534
rect 439462 692298 439546 692534
rect 439782 692298 439814 692534
rect 439194 656854 439814 692298
rect 439194 656618 439226 656854
rect 439462 656618 439546 656854
rect 439782 656618 439814 656854
rect 439194 656534 439814 656618
rect 439194 656298 439226 656534
rect 439462 656298 439546 656534
rect 439782 656298 439814 656534
rect 439194 620854 439814 656298
rect 439194 620618 439226 620854
rect 439462 620618 439546 620854
rect 439782 620618 439814 620854
rect 439194 620534 439814 620618
rect 439194 620298 439226 620534
rect 439462 620298 439546 620534
rect 439782 620298 439814 620534
rect 439194 584854 439814 620298
rect 439194 584618 439226 584854
rect 439462 584618 439546 584854
rect 439782 584618 439814 584854
rect 439194 584534 439814 584618
rect 439194 584298 439226 584534
rect 439462 584298 439546 584534
rect 439782 584298 439814 584534
rect 439194 548854 439814 584298
rect 439194 548618 439226 548854
rect 439462 548618 439546 548854
rect 439782 548618 439814 548854
rect 439194 548534 439814 548618
rect 439194 548298 439226 548534
rect 439462 548298 439546 548534
rect 439782 548298 439814 548534
rect 439194 512854 439814 548298
rect 439194 512618 439226 512854
rect 439462 512618 439546 512854
rect 439782 512618 439814 512854
rect 439194 512534 439814 512618
rect 439194 512298 439226 512534
rect 439462 512298 439546 512534
rect 439782 512298 439814 512534
rect 439194 476854 439814 512298
rect 439194 476618 439226 476854
rect 439462 476618 439546 476854
rect 439782 476618 439814 476854
rect 439194 476534 439814 476618
rect 439194 476298 439226 476534
rect 439462 476298 439546 476534
rect 439782 476298 439814 476534
rect 439194 440854 439814 476298
rect 439194 440618 439226 440854
rect 439462 440618 439546 440854
rect 439782 440618 439814 440854
rect 439194 440534 439814 440618
rect 439194 440298 439226 440534
rect 439462 440298 439546 440534
rect 439782 440298 439814 440534
rect 439194 404854 439814 440298
rect 439194 404618 439226 404854
rect 439462 404618 439546 404854
rect 439782 404618 439814 404854
rect 439194 404534 439814 404618
rect 439194 404298 439226 404534
rect 439462 404298 439546 404534
rect 439782 404298 439814 404534
rect 439194 368854 439814 404298
rect 439194 368618 439226 368854
rect 439462 368618 439546 368854
rect 439782 368618 439814 368854
rect 439194 368534 439814 368618
rect 439194 368298 439226 368534
rect 439462 368298 439546 368534
rect 439782 368298 439814 368534
rect 439194 332854 439814 368298
rect 439194 332618 439226 332854
rect 439462 332618 439546 332854
rect 439782 332618 439814 332854
rect 439194 332534 439814 332618
rect 439194 332298 439226 332534
rect 439462 332298 439546 332534
rect 439782 332298 439814 332534
rect 439194 296854 439814 332298
rect 439194 296618 439226 296854
rect 439462 296618 439546 296854
rect 439782 296618 439814 296854
rect 439194 296534 439814 296618
rect 439194 296298 439226 296534
rect 439462 296298 439546 296534
rect 439782 296298 439814 296534
rect 439194 260854 439814 296298
rect 439194 260618 439226 260854
rect 439462 260618 439546 260854
rect 439782 260618 439814 260854
rect 439194 260534 439814 260618
rect 439194 260298 439226 260534
rect 439462 260298 439546 260534
rect 439782 260298 439814 260534
rect 439194 224854 439814 260298
rect 439194 224618 439226 224854
rect 439462 224618 439546 224854
rect 439782 224618 439814 224854
rect 439194 224534 439814 224618
rect 439194 224298 439226 224534
rect 439462 224298 439546 224534
rect 439782 224298 439814 224534
rect 439194 188854 439814 224298
rect 439194 188618 439226 188854
rect 439462 188618 439546 188854
rect 439782 188618 439814 188854
rect 439194 188534 439814 188618
rect 439194 188298 439226 188534
rect 439462 188298 439546 188534
rect 439782 188298 439814 188534
rect 439194 152854 439814 188298
rect 439194 152618 439226 152854
rect 439462 152618 439546 152854
rect 439782 152618 439814 152854
rect 439194 152534 439814 152618
rect 439194 152298 439226 152534
rect 439462 152298 439546 152534
rect 439782 152298 439814 152534
rect 439194 116854 439814 152298
rect 439194 116618 439226 116854
rect 439462 116618 439546 116854
rect 439782 116618 439814 116854
rect 439194 116534 439814 116618
rect 439194 116298 439226 116534
rect 439462 116298 439546 116534
rect 439782 116298 439814 116534
rect 439194 80854 439814 116298
rect 439194 80618 439226 80854
rect 439462 80618 439546 80854
rect 439782 80618 439814 80854
rect 439194 80534 439814 80618
rect 439194 80298 439226 80534
rect 439462 80298 439546 80534
rect 439782 80298 439814 80534
rect 439194 44854 439814 80298
rect 439194 44618 439226 44854
rect 439462 44618 439546 44854
rect 439782 44618 439814 44854
rect 439194 44534 439814 44618
rect 439194 44298 439226 44534
rect 439462 44298 439546 44534
rect 439782 44298 439814 44534
rect 439194 8854 439814 44298
rect 439194 8618 439226 8854
rect 439462 8618 439546 8854
rect 439782 8618 439814 8854
rect 439194 8534 439814 8618
rect 439194 8298 439226 8534
rect 439462 8298 439546 8534
rect 439782 8298 439814 8534
rect 439194 -5146 439814 8298
rect 439194 -5382 439226 -5146
rect 439462 -5382 439546 -5146
rect 439782 -5382 439814 -5146
rect 439194 -5466 439814 -5382
rect 439194 -5702 439226 -5466
rect 439462 -5702 439546 -5466
rect 439782 -5702 439814 -5466
rect 439194 -7654 439814 -5702
rect 440434 710598 441054 711590
rect 440434 710362 440466 710598
rect 440702 710362 440786 710598
rect 441022 710362 441054 710598
rect 440434 710278 441054 710362
rect 440434 710042 440466 710278
rect 440702 710042 440786 710278
rect 441022 710042 441054 710278
rect 440434 694094 441054 710042
rect 440434 693858 440466 694094
rect 440702 693858 440786 694094
rect 441022 693858 441054 694094
rect 440434 693774 441054 693858
rect 440434 693538 440466 693774
rect 440702 693538 440786 693774
rect 441022 693538 441054 693774
rect 440434 658094 441054 693538
rect 440434 657858 440466 658094
rect 440702 657858 440786 658094
rect 441022 657858 441054 658094
rect 440434 657774 441054 657858
rect 440434 657538 440466 657774
rect 440702 657538 440786 657774
rect 441022 657538 441054 657774
rect 440434 622094 441054 657538
rect 440434 621858 440466 622094
rect 440702 621858 440786 622094
rect 441022 621858 441054 622094
rect 440434 621774 441054 621858
rect 440434 621538 440466 621774
rect 440702 621538 440786 621774
rect 441022 621538 441054 621774
rect 440434 586094 441054 621538
rect 440434 585858 440466 586094
rect 440702 585858 440786 586094
rect 441022 585858 441054 586094
rect 440434 585774 441054 585858
rect 440434 585538 440466 585774
rect 440702 585538 440786 585774
rect 441022 585538 441054 585774
rect 440434 550094 441054 585538
rect 440434 549858 440466 550094
rect 440702 549858 440786 550094
rect 441022 549858 441054 550094
rect 440434 549774 441054 549858
rect 440434 549538 440466 549774
rect 440702 549538 440786 549774
rect 441022 549538 441054 549774
rect 440434 514094 441054 549538
rect 440434 513858 440466 514094
rect 440702 513858 440786 514094
rect 441022 513858 441054 514094
rect 440434 513774 441054 513858
rect 440434 513538 440466 513774
rect 440702 513538 440786 513774
rect 441022 513538 441054 513774
rect 440434 478094 441054 513538
rect 440434 477858 440466 478094
rect 440702 477858 440786 478094
rect 441022 477858 441054 478094
rect 440434 477774 441054 477858
rect 440434 477538 440466 477774
rect 440702 477538 440786 477774
rect 441022 477538 441054 477774
rect 440434 442094 441054 477538
rect 440434 441858 440466 442094
rect 440702 441858 440786 442094
rect 441022 441858 441054 442094
rect 440434 441774 441054 441858
rect 440434 441538 440466 441774
rect 440702 441538 440786 441774
rect 441022 441538 441054 441774
rect 440434 406094 441054 441538
rect 440434 405858 440466 406094
rect 440702 405858 440786 406094
rect 441022 405858 441054 406094
rect 440434 405774 441054 405858
rect 440434 405538 440466 405774
rect 440702 405538 440786 405774
rect 441022 405538 441054 405774
rect 440434 370094 441054 405538
rect 440434 369858 440466 370094
rect 440702 369858 440786 370094
rect 441022 369858 441054 370094
rect 440434 369774 441054 369858
rect 440434 369538 440466 369774
rect 440702 369538 440786 369774
rect 441022 369538 441054 369774
rect 440434 334094 441054 369538
rect 440434 333858 440466 334094
rect 440702 333858 440786 334094
rect 441022 333858 441054 334094
rect 440434 333774 441054 333858
rect 440434 333538 440466 333774
rect 440702 333538 440786 333774
rect 441022 333538 441054 333774
rect 440434 298094 441054 333538
rect 440434 297858 440466 298094
rect 440702 297858 440786 298094
rect 441022 297858 441054 298094
rect 440434 297774 441054 297858
rect 440434 297538 440466 297774
rect 440702 297538 440786 297774
rect 441022 297538 441054 297774
rect 440434 262094 441054 297538
rect 440434 261858 440466 262094
rect 440702 261858 440786 262094
rect 441022 261858 441054 262094
rect 440434 261774 441054 261858
rect 440434 261538 440466 261774
rect 440702 261538 440786 261774
rect 441022 261538 441054 261774
rect 440434 226094 441054 261538
rect 440434 225858 440466 226094
rect 440702 225858 440786 226094
rect 441022 225858 441054 226094
rect 440434 225774 441054 225858
rect 440434 225538 440466 225774
rect 440702 225538 440786 225774
rect 441022 225538 441054 225774
rect 440434 190094 441054 225538
rect 440434 189858 440466 190094
rect 440702 189858 440786 190094
rect 441022 189858 441054 190094
rect 440434 189774 441054 189858
rect 440434 189538 440466 189774
rect 440702 189538 440786 189774
rect 441022 189538 441054 189774
rect 440434 154094 441054 189538
rect 440434 153858 440466 154094
rect 440702 153858 440786 154094
rect 441022 153858 441054 154094
rect 440434 153774 441054 153858
rect 440434 153538 440466 153774
rect 440702 153538 440786 153774
rect 441022 153538 441054 153774
rect 440434 118094 441054 153538
rect 440434 117858 440466 118094
rect 440702 117858 440786 118094
rect 441022 117858 441054 118094
rect 440434 117774 441054 117858
rect 440434 117538 440466 117774
rect 440702 117538 440786 117774
rect 441022 117538 441054 117774
rect 440434 82094 441054 117538
rect 440434 81858 440466 82094
rect 440702 81858 440786 82094
rect 441022 81858 441054 82094
rect 440434 81774 441054 81858
rect 440434 81538 440466 81774
rect 440702 81538 440786 81774
rect 441022 81538 441054 81774
rect 440434 46094 441054 81538
rect 440434 45858 440466 46094
rect 440702 45858 440786 46094
rect 441022 45858 441054 46094
rect 440434 45774 441054 45858
rect 440434 45538 440466 45774
rect 440702 45538 440786 45774
rect 441022 45538 441054 45774
rect 440434 10094 441054 45538
rect 440434 9858 440466 10094
rect 440702 9858 440786 10094
rect 441022 9858 441054 10094
rect 440434 9774 441054 9858
rect 440434 9538 440466 9774
rect 440702 9538 440786 9774
rect 441022 9538 441054 9774
rect 440434 -6106 441054 9538
rect 440434 -6342 440466 -6106
rect 440702 -6342 440786 -6106
rect 441022 -6342 441054 -6106
rect 440434 -6426 441054 -6342
rect 440434 -6662 440466 -6426
rect 440702 -6662 440786 -6426
rect 441022 -6662 441054 -6426
rect 440434 -7654 441054 -6662
rect 441674 711558 442294 711590
rect 441674 711322 441706 711558
rect 441942 711322 442026 711558
rect 442262 711322 442294 711558
rect 441674 711238 442294 711322
rect 441674 711002 441706 711238
rect 441942 711002 442026 711238
rect 442262 711002 442294 711238
rect 441674 695334 442294 711002
rect 441674 695098 441706 695334
rect 441942 695098 442026 695334
rect 442262 695098 442294 695334
rect 441674 695014 442294 695098
rect 441674 694778 441706 695014
rect 441942 694778 442026 695014
rect 442262 694778 442294 695014
rect 441674 659334 442294 694778
rect 441674 659098 441706 659334
rect 441942 659098 442026 659334
rect 442262 659098 442294 659334
rect 441674 659014 442294 659098
rect 441674 658778 441706 659014
rect 441942 658778 442026 659014
rect 442262 658778 442294 659014
rect 441674 623334 442294 658778
rect 441674 623098 441706 623334
rect 441942 623098 442026 623334
rect 442262 623098 442294 623334
rect 441674 623014 442294 623098
rect 441674 622778 441706 623014
rect 441942 622778 442026 623014
rect 442262 622778 442294 623014
rect 441674 587334 442294 622778
rect 441674 587098 441706 587334
rect 441942 587098 442026 587334
rect 442262 587098 442294 587334
rect 441674 587014 442294 587098
rect 441674 586778 441706 587014
rect 441942 586778 442026 587014
rect 442262 586778 442294 587014
rect 441674 551334 442294 586778
rect 441674 551098 441706 551334
rect 441942 551098 442026 551334
rect 442262 551098 442294 551334
rect 441674 551014 442294 551098
rect 441674 550778 441706 551014
rect 441942 550778 442026 551014
rect 442262 550778 442294 551014
rect 441674 515334 442294 550778
rect 441674 515098 441706 515334
rect 441942 515098 442026 515334
rect 442262 515098 442294 515334
rect 441674 515014 442294 515098
rect 441674 514778 441706 515014
rect 441942 514778 442026 515014
rect 442262 514778 442294 515014
rect 441674 479334 442294 514778
rect 441674 479098 441706 479334
rect 441942 479098 442026 479334
rect 442262 479098 442294 479334
rect 441674 479014 442294 479098
rect 441674 478778 441706 479014
rect 441942 478778 442026 479014
rect 442262 478778 442294 479014
rect 441674 443334 442294 478778
rect 441674 443098 441706 443334
rect 441942 443098 442026 443334
rect 442262 443098 442294 443334
rect 441674 443014 442294 443098
rect 441674 442778 441706 443014
rect 441942 442778 442026 443014
rect 442262 442778 442294 443014
rect 441674 407334 442294 442778
rect 441674 407098 441706 407334
rect 441942 407098 442026 407334
rect 442262 407098 442294 407334
rect 441674 407014 442294 407098
rect 441674 406778 441706 407014
rect 441942 406778 442026 407014
rect 442262 406778 442294 407014
rect 441674 371334 442294 406778
rect 441674 371098 441706 371334
rect 441942 371098 442026 371334
rect 442262 371098 442294 371334
rect 441674 371014 442294 371098
rect 441674 370778 441706 371014
rect 441942 370778 442026 371014
rect 442262 370778 442294 371014
rect 441674 335334 442294 370778
rect 441674 335098 441706 335334
rect 441942 335098 442026 335334
rect 442262 335098 442294 335334
rect 441674 335014 442294 335098
rect 441674 334778 441706 335014
rect 441942 334778 442026 335014
rect 442262 334778 442294 335014
rect 441674 299334 442294 334778
rect 441674 299098 441706 299334
rect 441942 299098 442026 299334
rect 442262 299098 442294 299334
rect 441674 299014 442294 299098
rect 441674 298778 441706 299014
rect 441942 298778 442026 299014
rect 442262 298778 442294 299014
rect 441674 263334 442294 298778
rect 441674 263098 441706 263334
rect 441942 263098 442026 263334
rect 442262 263098 442294 263334
rect 441674 263014 442294 263098
rect 441674 262778 441706 263014
rect 441942 262778 442026 263014
rect 442262 262778 442294 263014
rect 441674 227334 442294 262778
rect 441674 227098 441706 227334
rect 441942 227098 442026 227334
rect 442262 227098 442294 227334
rect 441674 227014 442294 227098
rect 441674 226778 441706 227014
rect 441942 226778 442026 227014
rect 442262 226778 442294 227014
rect 441674 191334 442294 226778
rect 441674 191098 441706 191334
rect 441942 191098 442026 191334
rect 442262 191098 442294 191334
rect 441674 191014 442294 191098
rect 441674 190778 441706 191014
rect 441942 190778 442026 191014
rect 442262 190778 442294 191014
rect 441674 155334 442294 190778
rect 441674 155098 441706 155334
rect 441942 155098 442026 155334
rect 442262 155098 442294 155334
rect 441674 155014 442294 155098
rect 441674 154778 441706 155014
rect 441942 154778 442026 155014
rect 442262 154778 442294 155014
rect 441674 119334 442294 154778
rect 441674 119098 441706 119334
rect 441942 119098 442026 119334
rect 442262 119098 442294 119334
rect 441674 119014 442294 119098
rect 441674 118778 441706 119014
rect 441942 118778 442026 119014
rect 442262 118778 442294 119014
rect 441674 83334 442294 118778
rect 441674 83098 441706 83334
rect 441942 83098 442026 83334
rect 442262 83098 442294 83334
rect 441674 83014 442294 83098
rect 441674 82778 441706 83014
rect 441942 82778 442026 83014
rect 442262 82778 442294 83014
rect 441674 47334 442294 82778
rect 441674 47098 441706 47334
rect 441942 47098 442026 47334
rect 442262 47098 442294 47334
rect 441674 47014 442294 47098
rect 441674 46778 441706 47014
rect 441942 46778 442026 47014
rect 442262 46778 442294 47014
rect 441674 11334 442294 46778
rect 441674 11098 441706 11334
rect 441942 11098 442026 11334
rect 442262 11098 442294 11334
rect 441674 11014 442294 11098
rect 441674 10778 441706 11014
rect 441942 10778 442026 11014
rect 442262 10778 442294 11014
rect 441674 -7066 442294 10778
rect 441674 -7302 441706 -7066
rect 441942 -7302 442026 -7066
rect 442262 -7302 442294 -7066
rect 441674 -7386 442294 -7302
rect 441674 -7622 441706 -7386
rect 441942 -7622 442026 -7386
rect 442262 -7622 442294 -7386
rect 441674 -7654 442294 -7622
rect 468994 704838 469614 711590
rect 468994 704602 469026 704838
rect 469262 704602 469346 704838
rect 469582 704602 469614 704838
rect 468994 704518 469614 704602
rect 468994 704282 469026 704518
rect 469262 704282 469346 704518
rect 469582 704282 469614 704518
rect 468994 686654 469614 704282
rect 468994 686418 469026 686654
rect 469262 686418 469346 686654
rect 469582 686418 469614 686654
rect 468994 686334 469614 686418
rect 468994 686098 469026 686334
rect 469262 686098 469346 686334
rect 469582 686098 469614 686334
rect 468994 650654 469614 686098
rect 468994 650418 469026 650654
rect 469262 650418 469346 650654
rect 469582 650418 469614 650654
rect 468994 650334 469614 650418
rect 468994 650098 469026 650334
rect 469262 650098 469346 650334
rect 469582 650098 469614 650334
rect 468994 614654 469614 650098
rect 468994 614418 469026 614654
rect 469262 614418 469346 614654
rect 469582 614418 469614 614654
rect 468994 614334 469614 614418
rect 468994 614098 469026 614334
rect 469262 614098 469346 614334
rect 469582 614098 469614 614334
rect 468994 578654 469614 614098
rect 468994 578418 469026 578654
rect 469262 578418 469346 578654
rect 469582 578418 469614 578654
rect 468994 578334 469614 578418
rect 468994 578098 469026 578334
rect 469262 578098 469346 578334
rect 469582 578098 469614 578334
rect 468994 542654 469614 578098
rect 468994 542418 469026 542654
rect 469262 542418 469346 542654
rect 469582 542418 469614 542654
rect 468994 542334 469614 542418
rect 468994 542098 469026 542334
rect 469262 542098 469346 542334
rect 469582 542098 469614 542334
rect 468994 506654 469614 542098
rect 468994 506418 469026 506654
rect 469262 506418 469346 506654
rect 469582 506418 469614 506654
rect 468994 506334 469614 506418
rect 468994 506098 469026 506334
rect 469262 506098 469346 506334
rect 469582 506098 469614 506334
rect 468994 470654 469614 506098
rect 468994 470418 469026 470654
rect 469262 470418 469346 470654
rect 469582 470418 469614 470654
rect 468994 470334 469614 470418
rect 468994 470098 469026 470334
rect 469262 470098 469346 470334
rect 469582 470098 469614 470334
rect 468994 450397 469614 470098
rect 468994 450333 469032 450397
rect 469096 450333 469112 450397
rect 469176 450333 469192 450397
rect 469256 450333 469272 450397
rect 469336 450333 469352 450397
rect 469416 450333 469432 450397
rect 469496 450333 469512 450397
rect 469576 450333 469614 450397
rect 468994 450317 469614 450333
rect 468994 450253 469032 450317
rect 469096 450253 469112 450317
rect 469176 450253 469192 450317
rect 469256 450253 469272 450317
rect 469336 450253 469352 450317
rect 469416 450253 469432 450317
rect 469496 450253 469512 450317
rect 469576 450253 469614 450317
rect 468994 450237 469614 450253
rect 468994 450173 469032 450237
rect 469096 450173 469112 450237
rect 469176 450173 469192 450237
rect 469256 450173 469272 450237
rect 469336 450173 469352 450237
rect 469416 450173 469432 450237
rect 469496 450173 469512 450237
rect 469576 450173 469614 450237
rect 468994 450157 469614 450173
rect 468994 450093 469032 450157
rect 469096 450093 469112 450157
rect 469176 450093 469192 450157
rect 469256 450093 469272 450157
rect 469336 450093 469352 450157
rect 469416 450093 469432 450157
rect 469496 450093 469512 450157
rect 469576 450093 469614 450157
rect 468994 434654 469614 450093
rect 468994 434418 469026 434654
rect 469262 434418 469346 434654
rect 469582 434418 469614 434654
rect 468994 434334 469614 434418
rect 468994 434098 469026 434334
rect 469262 434098 469346 434334
rect 469582 434098 469614 434334
rect 468994 431997 469614 434098
rect 468994 431933 469032 431997
rect 469096 431933 469112 431997
rect 469176 431933 469192 431997
rect 469256 431933 469272 431997
rect 469336 431933 469352 431997
rect 469416 431933 469432 431997
rect 469496 431933 469512 431997
rect 469576 431933 469614 431997
rect 468994 431917 469614 431933
rect 468994 431853 469032 431917
rect 469096 431853 469112 431917
rect 469176 431853 469192 431917
rect 469256 431853 469272 431917
rect 469336 431853 469352 431917
rect 469416 431853 469432 431917
rect 469496 431853 469512 431917
rect 469576 431853 469614 431917
rect 468994 431837 469614 431853
rect 468994 431773 469032 431837
rect 469096 431773 469112 431837
rect 469176 431773 469192 431837
rect 469256 431773 469272 431837
rect 469336 431773 469352 431837
rect 469416 431773 469432 431837
rect 469496 431773 469512 431837
rect 469576 431773 469614 431837
rect 468994 431757 469614 431773
rect 468994 431693 469032 431757
rect 469096 431693 469112 431757
rect 469176 431693 469192 431757
rect 469256 431693 469272 431757
rect 469336 431693 469352 431757
rect 469416 431693 469432 431757
rect 469496 431693 469512 431757
rect 469576 431693 469614 431757
rect 468994 410998 469614 431693
rect 468994 410934 469032 410998
rect 469096 410934 469112 410998
rect 469176 410934 469192 410998
rect 469256 410934 469272 410998
rect 469336 410934 469352 410998
rect 469416 410934 469432 410998
rect 469496 410934 469512 410998
rect 469576 410934 469614 410998
rect 468994 410918 469614 410934
rect 468994 410854 469032 410918
rect 469096 410854 469112 410918
rect 469176 410854 469192 410918
rect 469256 410854 469272 410918
rect 469336 410854 469352 410918
rect 469416 410854 469432 410918
rect 469496 410854 469512 410918
rect 469576 410854 469614 410918
rect 468994 410838 469614 410854
rect 468994 410774 469032 410838
rect 469096 410774 469112 410838
rect 469176 410774 469192 410838
rect 469256 410774 469272 410838
rect 469336 410774 469352 410838
rect 469416 410774 469432 410838
rect 469496 410774 469512 410838
rect 469576 410774 469614 410838
rect 468994 410758 469614 410774
rect 468994 410694 469032 410758
rect 469096 410694 469112 410758
rect 469176 410694 469192 410758
rect 469256 410694 469272 410758
rect 469336 410694 469352 410758
rect 469416 410694 469432 410758
rect 469496 410694 469512 410758
rect 469576 410694 469614 410758
rect 468994 398654 469614 410694
rect 468994 398418 469026 398654
rect 469262 398418 469346 398654
rect 469582 398418 469614 398654
rect 468994 398334 469614 398418
rect 468994 398098 469026 398334
rect 469262 398098 469346 398334
rect 469582 398098 469614 398334
rect 468994 390002 469614 398098
rect 468994 389938 469032 390002
rect 469096 389938 469112 390002
rect 469176 389938 469192 390002
rect 469256 389938 469272 390002
rect 469336 389938 469352 390002
rect 469416 389938 469432 390002
rect 469496 389938 469512 390002
rect 469576 389938 469614 390002
rect 468994 389922 469614 389938
rect 468994 389858 469032 389922
rect 469096 389858 469112 389922
rect 469176 389858 469192 389922
rect 469256 389858 469272 389922
rect 469336 389858 469352 389922
rect 469416 389858 469432 389922
rect 469496 389858 469512 389922
rect 469576 389858 469614 389922
rect 468994 389842 469614 389858
rect 468994 389778 469032 389842
rect 469096 389778 469112 389842
rect 469176 389778 469192 389842
rect 469256 389778 469272 389842
rect 469336 389778 469352 389842
rect 469416 389778 469432 389842
rect 469496 389778 469512 389842
rect 469576 389778 469614 389842
rect 468994 389762 469614 389778
rect 468994 389698 469032 389762
rect 469096 389698 469112 389762
rect 469176 389698 469192 389762
rect 469256 389698 469272 389762
rect 469336 389698 469352 389762
rect 469416 389698 469432 389762
rect 469496 389698 469512 389762
rect 469576 389698 469614 389762
rect 468994 362654 469614 389698
rect 468994 362418 469026 362654
rect 469262 362418 469346 362654
rect 469582 362418 469614 362654
rect 468994 362334 469614 362418
rect 468994 362098 469026 362334
rect 469262 362098 469346 362334
rect 469582 362098 469614 362334
rect 468994 357399 469614 362098
rect 468994 357335 469032 357399
rect 469096 357335 469112 357399
rect 469176 357335 469192 357399
rect 469256 357335 469272 357399
rect 469336 357335 469352 357399
rect 469416 357335 469432 357399
rect 469496 357335 469512 357399
rect 469576 357335 469614 357399
rect 468994 357319 469614 357335
rect 468994 357255 469032 357319
rect 469096 357255 469112 357319
rect 469176 357255 469192 357319
rect 469256 357255 469272 357319
rect 469336 357255 469352 357319
rect 469416 357255 469432 357319
rect 469496 357255 469512 357319
rect 469576 357255 469614 357319
rect 468994 357239 469614 357255
rect 468994 357175 469032 357239
rect 469096 357175 469112 357239
rect 469176 357175 469192 357239
rect 469256 357175 469272 357239
rect 469336 357175 469352 357239
rect 469416 357175 469432 357239
rect 469496 357175 469512 357239
rect 469576 357175 469614 357239
rect 468994 357159 469614 357175
rect 468994 357095 469032 357159
rect 469096 357095 469112 357159
rect 469176 357095 469192 357159
rect 469256 357095 469272 357159
rect 469336 357095 469352 357159
rect 469416 357095 469432 357159
rect 469496 357095 469512 357159
rect 469576 357095 469614 357159
rect 468994 341397 469614 357095
rect 468994 341333 469032 341397
rect 469096 341333 469112 341397
rect 469176 341333 469192 341397
rect 469256 341333 469272 341397
rect 469336 341333 469352 341397
rect 469416 341333 469432 341397
rect 469496 341333 469512 341397
rect 469576 341333 469614 341397
rect 468994 341317 469614 341333
rect 468994 341253 469032 341317
rect 469096 341253 469112 341317
rect 469176 341253 469192 341317
rect 469256 341253 469272 341317
rect 469336 341253 469352 341317
rect 469416 341253 469432 341317
rect 469496 341253 469512 341317
rect 469576 341253 469614 341317
rect 468994 341237 469614 341253
rect 468994 341173 469032 341237
rect 469096 341173 469112 341237
rect 469176 341173 469192 341237
rect 469256 341173 469272 341237
rect 469336 341173 469352 341237
rect 469416 341173 469432 341237
rect 469496 341173 469512 341237
rect 469576 341173 469614 341237
rect 468994 341157 469614 341173
rect 468994 341093 469032 341157
rect 469096 341093 469112 341157
rect 469176 341093 469192 341157
rect 469256 341093 469272 341157
rect 469336 341093 469352 341157
rect 469416 341093 469432 341157
rect 469496 341093 469512 341157
rect 469576 341093 469614 341157
rect 468994 326654 469614 341093
rect 468994 326418 469026 326654
rect 469262 326418 469346 326654
rect 469582 326418 469614 326654
rect 468994 326334 469614 326418
rect 468994 326098 469026 326334
rect 469262 326098 469346 326334
rect 469582 326098 469614 326334
rect 468994 321397 469614 326098
rect 468994 321333 469032 321397
rect 469096 321333 469112 321397
rect 469176 321333 469192 321397
rect 469256 321333 469272 321397
rect 469336 321333 469352 321397
rect 469416 321333 469432 321397
rect 469496 321333 469512 321397
rect 469576 321333 469614 321397
rect 468994 321317 469614 321333
rect 468994 321253 469032 321317
rect 469096 321253 469112 321317
rect 469176 321253 469192 321317
rect 469256 321253 469272 321317
rect 469336 321253 469352 321317
rect 469416 321253 469432 321317
rect 469496 321253 469512 321317
rect 469576 321253 469614 321317
rect 468994 321237 469614 321253
rect 468994 321173 469032 321237
rect 469096 321173 469112 321237
rect 469176 321173 469192 321237
rect 469256 321173 469272 321237
rect 469336 321173 469352 321237
rect 469416 321173 469432 321237
rect 469496 321173 469512 321237
rect 469576 321173 469614 321237
rect 468994 321157 469614 321173
rect 468994 321093 469032 321157
rect 469096 321093 469112 321157
rect 469176 321093 469192 321157
rect 469256 321093 469272 321157
rect 469336 321093 469352 321157
rect 469416 321093 469432 321157
rect 469496 321093 469512 321157
rect 469576 321093 469614 321157
rect 468994 305999 469614 321093
rect 468994 305935 469032 305999
rect 469096 305935 469112 305999
rect 469176 305935 469192 305999
rect 469256 305935 469272 305999
rect 469336 305935 469352 305999
rect 469416 305935 469432 305999
rect 469496 305935 469512 305999
rect 469576 305935 469614 305999
rect 468994 305919 469614 305935
rect 468994 305855 469032 305919
rect 469096 305855 469112 305919
rect 469176 305855 469192 305919
rect 469256 305855 469272 305919
rect 469336 305855 469352 305919
rect 469416 305855 469432 305919
rect 469496 305855 469512 305919
rect 469576 305855 469614 305919
rect 468994 305839 469614 305855
rect 468994 305775 469032 305839
rect 469096 305775 469112 305839
rect 469176 305775 469192 305839
rect 469256 305775 469272 305839
rect 469336 305775 469352 305839
rect 469416 305775 469432 305839
rect 469496 305775 469512 305839
rect 469576 305775 469614 305839
rect 468994 305759 469614 305775
rect 468994 305695 469032 305759
rect 469096 305695 469112 305759
rect 469176 305695 469192 305759
rect 469256 305695 469272 305759
rect 469336 305695 469352 305759
rect 469416 305695 469432 305759
rect 469496 305695 469512 305759
rect 469576 305695 469614 305759
rect 468994 290654 469614 305695
rect 468994 290418 469026 290654
rect 469262 290418 469346 290654
rect 469582 290418 469614 290654
rect 468994 290334 469614 290418
rect 468994 290098 469026 290334
rect 469262 290098 469346 290334
rect 469582 290098 469614 290334
rect 468994 286400 469614 290098
rect 468994 286336 469032 286400
rect 469096 286336 469112 286400
rect 469176 286336 469192 286400
rect 469256 286336 469272 286400
rect 469336 286336 469352 286400
rect 469416 286336 469432 286400
rect 469496 286336 469512 286400
rect 469576 286336 469614 286400
rect 468994 286320 469614 286336
rect 468994 286256 469032 286320
rect 469096 286256 469112 286320
rect 469176 286256 469192 286320
rect 469256 286256 469272 286320
rect 469336 286256 469352 286320
rect 469416 286256 469432 286320
rect 469496 286256 469512 286320
rect 469576 286256 469614 286320
rect 468994 286240 469614 286256
rect 468994 286176 469032 286240
rect 469096 286176 469112 286240
rect 469176 286176 469192 286240
rect 469256 286176 469272 286240
rect 469336 286176 469352 286240
rect 469416 286176 469432 286240
rect 469496 286176 469512 286240
rect 469576 286176 469614 286240
rect 468994 286160 469614 286176
rect 468994 286096 469032 286160
rect 469096 286096 469112 286160
rect 469176 286096 469192 286160
rect 469256 286096 469272 286160
rect 469336 286096 469352 286160
rect 469416 286096 469432 286160
rect 469496 286096 469512 286160
rect 469576 286096 469614 286160
rect 468994 266399 469614 286096
rect 468994 266335 469032 266399
rect 469096 266335 469112 266399
rect 469176 266335 469192 266399
rect 469256 266335 469272 266399
rect 469336 266335 469352 266399
rect 469416 266335 469432 266399
rect 469496 266335 469512 266399
rect 469576 266335 469614 266399
rect 468994 266319 469614 266335
rect 468994 266255 469032 266319
rect 469096 266255 469112 266319
rect 469176 266255 469192 266319
rect 469256 266255 469272 266319
rect 469336 266255 469352 266319
rect 469416 266255 469432 266319
rect 469496 266255 469512 266319
rect 469576 266255 469614 266319
rect 468994 266239 469614 266255
rect 468994 266175 469032 266239
rect 469096 266175 469112 266239
rect 469176 266175 469192 266239
rect 469256 266175 469272 266239
rect 469336 266175 469352 266239
rect 469416 266175 469432 266239
rect 469496 266175 469512 266239
rect 469576 266175 469614 266239
rect 468994 266159 469614 266175
rect 468994 266095 469032 266159
rect 469096 266095 469112 266159
rect 469176 266095 469192 266159
rect 469256 266095 469272 266159
rect 469336 266095 469352 266159
rect 469416 266095 469432 266159
rect 469496 266095 469512 266159
rect 469576 266095 469614 266159
rect 468994 254654 469614 266095
rect 468994 254418 469026 254654
rect 469262 254418 469346 254654
rect 469582 254418 469614 254654
rect 468994 254334 469614 254418
rect 468994 254098 469026 254334
rect 469262 254098 469346 254334
rect 469582 254098 469614 254334
rect 468994 218654 469614 254098
rect 468994 218418 469026 218654
rect 469262 218418 469346 218654
rect 469582 218418 469614 218654
rect 468994 218334 469614 218418
rect 468994 218098 469026 218334
rect 469262 218098 469346 218334
rect 469582 218098 469614 218334
rect 468994 182654 469614 218098
rect 468994 182418 469026 182654
rect 469262 182418 469346 182654
rect 469582 182418 469614 182654
rect 468994 182334 469614 182418
rect 468994 182098 469026 182334
rect 469262 182098 469346 182334
rect 469582 182098 469614 182334
rect 468994 146654 469614 182098
rect 468994 146418 469026 146654
rect 469262 146418 469346 146654
rect 469582 146418 469614 146654
rect 468994 146334 469614 146418
rect 468994 146098 469026 146334
rect 469262 146098 469346 146334
rect 469582 146098 469614 146334
rect 468994 110654 469614 146098
rect 468994 110418 469026 110654
rect 469262 110418 469346 110654
rect 469582 110418 469614 110654
rect 468994 110334 469614 110418
rect 468994 110098 469026 110334
rect 469262 110098 469346 110334
rect 469582 110098 469614 110334
rect 468994 74654 469614 110098
rect 468994 74418 469026 74654
rect 469262 74418 469346 74654
rect 469582 74418 469614 74654
rect 468994 74334 469614 74418
rect 468994 74098 469026 74334
rect 469262 74098 469346 74334
rect 469582 74098 469614 74334
rect 468994 38654 469614 74098
rect 468994 38418 469026 38654
rect 469262 38418 469346 38654
rect 469582 38418 469614 38654
rect 468994 38334 469614 38418
rect 468994 38098 469026 38334
rect 469262 38098 469346 38334
rect 469582 38098 469614 38334
rect 468994 2654 469614 38098
rect 468994 2418 469026 2654
rect 469262 2418 469346 2654
rect 469582 2418 469614 2654
rect 468994 2334 469614 2418
rect 468994 2098 469026 2334
rect 469262 2098 469346 2334
rect 469582 2098 469614 2334
rect 468994 -346 469614 2098
rect 468994 -582 469026 -346
rect 469262 -582 469346 -346
rect 469582 -582 469614 -346
rect 468994 -666 469614 -582
rect 468994 -902 469026 -666
rect 469262 -902 469346 -666
rect 469582 -902 469614 -666
rect 468994 -7654 469614 -902
rect 470234 705798 470854 711590
rect 470234 705562 470266 705798
rect 470502 705562 470586 705798
rect 470822 705562 470854 705798
rect 470234 705478 470854 705562
rect 470234 705242 470266 705478
rect 470502 705242 470586 705478
rect 470822 705242 470854 705478
rect 470234 687894 470854 705242
rect 470234 687658 470266 687894
rect 470502 687658 470586 687894
rect 470822 687658 470854 687894
rect 470234 687574 470854 687658
rect 470234 687338 470266 687574
rect 470502 687338 470586 687574
rect 470822 687338 470854 687574
rect 470234 651894 470854 687338
rect 470234 651658 470266 651894
rect 470502 651658 470586 651894
rect 470822 651658 470854 651894
rect 470234 651574 470854 651658
rect 470234 651338 470266 651574
rect 470502 651338 470586 651574
rect 470822 651338 470854 651574
rect 470234 615894 470854 651338
rect 470234 615658 470266 615894
rect 470502 615658 470586 615894
rect 470822 615658 470854 615894
rect 470234 615574 470854 615658
rect 470234 615338 470266 615574
rect 470502 615338 470586 615574
rect 470822 615338 470854 615574
rect 470234 579894 470854 615338
rect 470234 579658 470266 579894
rect 470502 579658 470586 579894
rect 470822 579658 470854 579894
rect 470234 579574 470854 579658
rect 470234 579338 470266 579574
rect 470502 579338 470586 579574
rect 470822 579338 470854 579574
rect 470234 543894 470854 579338
rect 470234 543658 470266 543894
rect 470502 543658 470586 543894
rect 470822 543658 470854 543894
rect 470234 543574 470854 543658
rect 470234 543338 470266 543574
rect 470502 543338 470586 543574
rect 470822 543338 470854 543574
rect 470234 507894 470854 543338
rect 470234 507658 470266 507894
rect 470502 507658 470586 507894
rect 470822 507658 470854 507894
rect 470234 507574 470854 507658
rect 470234 507338 470266 507574
rect 470502 507338 470586 507574
rect 470822 507338 470854 507574
rect 470234 471894 470854 507338
rect 470234 471658 470266 471894
rect 470502 471658 470586 471894
rect 470822 471658 470854 471894
rect 470234 471574 470854 471658
rect 470234 471338 470266 471574
rect 470502 471338 470586 471574
rect 470822 471338 470854 471574
rect 470234 451483 470854 471338
rect 470234 451419 470272 451483
rect 470336 451419 470352 451483
rect 470416 451419 470432 451483
rect 470496 451419 470512 451483
rect 470576 451419 470592 451483
rect 470656 451419 470672 451483
rect 470736 451419 470752 451483
rect 470816 451419 470854 451483
rect 470234 451403 470854 451419
rect 470234 451339 470272 451403
rect 470336 451339 470352 451403
rect 470416 451339 470432 451403
rect 470496 451339 470512 451403
rect 470576 451339 470592 451403
rect 470656 451339 470672 451403
rect 470736 451339 470752 451403
rect 470816 451339 470854 451403
rect 470234 451323 470854 451339
rect 470234 451259 470272 451323
rect 470336 451259 470352 451323
rect 470416 451259 470432 451323
rect 470496 451259 470512 451323
rect 470576 451259 470592 451323
rect 470656 451259 470672 451323
rect 470736 451259 470752 451323
rect 470816 451259 470854 451323
rect 470234 451243 470854 451259
rect 470234 451179 470272 451243
rect 470336 451179 470352 451243
rect 470416 451179 470432 451243
rect 470496 451179 470512 451243
rect 470576 451179 470592 451243
rect 470656 451179 470672 451243
rect 470736 451179 470752 451243
rect 470816 451179 470854 451243
rect 470234 449312 470854 451179
rect 470234 449248 470272 449312
rect 470336 449248 470352 449312
rect 470416 449248 470432 449312
rect 470496 449248 470512 449312
rect 470576 449248 470592 449312
rect 470656 449248 470672 449312
rect 470736 449248 470752 449312
rect 470816 449248 470854 449312
rect 470234 449232 470854 449248
rect 470234 449168 470272 449232
rect 470336 449168 470352 449232
rect 470416 449168 470432 449232
rect 470496 449168 470512 449232
rect 470576 449168 470592 449232
rect 470656 449168 470672 449232
rect 470736 449168 470752 449232
rect 470816 449168 470854 449232
rect 470234 449152 470854 449168
rect 470234 449088 470272 449152
rect 470336 449088 470352 449152
rect 470416 449088 470432 449152
rect 470496 449088 470512 449152
rect 470576 449088 470592 449152
rect 470656 449088 470672 449152
rect 470736 449088 470752 449152
rect 470816 449088 470854 449152
rect 470234 449072 470854 449088
rect 470234 449008 470272 449072
rect 470336 449008 470352 449072
rect 470416 449008 470432 449072
rect 470496 449008 470512 449072
rect 470576 449008 470592 449072
rect 470656 449008 470672 449072
rect 470736 449008 470752 449072
rect 470816 449008 470854 449072
rect 470234 435894 470854 449008
rect 470234 435658 470266 435894
rect 470502 435658 470586 435894
rect 470822 435658 470854 435894
rect 470234 435574 470854 435658
rect 470234 435338 470266 435574
rect 470502 435338 470586 435574
rect 470822 435338 470854 435574
rect 470234 433084 470854 435338
rect 470234 433020 470272 433084
rect 470336 433020 470352 433084
rect 470416 433020 470432 433084
rect 470496 433020 470512 433084
rect 470576 433020 470592 433084
rect 470656 433020 470672 433084
rect 470736 433020 470752 433084
rect 470816 433020 470854 433084
rect 470234 433004 470854 433020
rect 470234 432940 470272 433004
rect 470336 432940 470352 433004
rect 470416 432940 470432 433004
rect 470496 432940 470512 433004
rect 470576 432940 470592 433004
rect 470656 432940 470672 433004
rect 470736 432940 470752 433004
rect 470816 432940 470854 433004
rect 470234 432924 470854 432940
rect 470234 432860 470272 432924
rect 470336 432860 470352 432924
rect 470416 432860 470432 432924
rect 470496 432860 470512 432924
rect 470576 432860 470592 432924
rect 470656 432860 470672 432924
rect 470736 432860 470752 432924
rect 470816 432860 470854 432924
rect 470234 432844 470854 432860
rect 470234 432780 470272 432844
rect 470336 432780 470352 432844
rect 470416 432780 470432 432844
rect 470496 432780 470512 432844
rect 470576 432780 470592 432844
rect 470656 432780 470672 432844
rect 470736 432780 470752 432844
rect 470816 432780 470854 432844
rect 470234 430912 470854 432780
rect 470234 430848 470272 430912
rect 470336 430848 470352 430912
rect 470416 430848 470432 430912
rect 470496 430848 470512 430912
rect 470576 430848 470592 430912
rect 470656 430848 470672 430912
rect 470736 430848 470752 430912
rect 470816 430848 470854 430912
rect 470234 430832 470854 430848
rect 470234 430768 470272 430832
rect 470336 430768 470352 430832
rect 470416 430768 470432 430832
rect 470496 430768 470512 430832
rect 470576 430768 470592 430832
rect 470656 430768 470672 430832
rect 470736 430768 470752 430832
rect 470816 430768 470854 430832
rect 470234 430752 470854 430768
rect 470234 430688 470272 430752
rect 470336 430688 470352 430752
rect 470416 430688 470432 430752
rect 470496 430688 470512 430752
rect 470576 430688 470592 430752
rect 470656 430688 470672 430752
rect 470736 430688 470752 430752
rect 470816 430688 470854 430752
rect 470234 430672 470854 430688
rect 470234 430608 470272 430672
rect 470336 430608 470352 430672
rect 470416 430608 470432 430672
rect 470496 430608 470512 430672
rect 470576 430608 470592 430672
rect 470656 430608 470672 430672
rect 470736 430608 470752 430672
rect 470816 430608 470854 430672
rect 470234 412084 470854 430608
rect 470234 412020 470272 412084
rect 470336 412020 470352 412084
rect 470416 412020 470432 412084
rect 470496 412020 470512 412084
rect 470576 412020 470592 412084
rect 470656 412020 470672 412084
rect 470736 412020 470752 412084
rect 470816 412020 470854 412084
rect 470234 412004 470854 412020
rect 470234 411940 470272 412004
rect 470336 411940 470352 412004
rect 470416 411940 470432 412004
rect 470496 411940 470512 412004
rect 470576 411940 470592 412004
rect 470656 411940 470672 412004
rect 470736 411940 470752 412004
rect 470816 411940 470854 412004
rect 470234 411924 470854 411940
rect 470234 411860 470272 411924
rect 470336 411860 470352 411924
rect 470416 411860 470432 411924
rect 470496 411860 470512 411924
rect 470576 411860 470592 411924
rect 470656 411860 470672 411924
rect 470736 411860 470752 411924
rect 470816 411860 470854 411924
rect 470234 411844 470854 411860
rect 470234 411780 470272 411844
rect 470336 411780 470352 411844
rect 470416 411780 470432 411844
rect 470496 411780 470512 411844
rect 470576 411780 470592 411844
rect 470656 411780 470672 411844
rect 470736 411780 470752 411844
rect 470816 411780 470854 411844
rect 470234 409912 470854 411780
rect 470234 409848 470272 409912
rect 470336 409848 470352 409912
rect 470416 409848 470432 409912
rect 470496 409848 470512 409912
rect 470576 409848 470592 409912
rect 470656 409848 470672 409912
rect 470736 409848 470752 409912
rect 470816 409848 470854 409912
rect 470234 409832 470854 409848
rect 470234 409768 470272 409832
rect 470336 409768 470352 409832
rect 470416 409768 470432 409832
rect 470496 409768 470512 409832
rect 470576 409768 470592 409832
rect 470656 409768 470672 409832
rect 470736 409768 470752 409832
rect 470816 409768 470854 409832
rect 470234 409752 470854 409768
rect 470234 409688 470272 409752
rect 470336 409688 470352 409752
rect 470416 409688 470432 409752
rect 470496 409688 470512 409752
rect 470576 409688 470592 409752
rect 470656 409688 470672 409752
rect 470736 409688 470752 409752
rect 470816 409688 470854 409752
rect 470234 409672 470854 409688
rect 470234 409608 470272 409672
rect 470336 409608 470352 409672
rect 470416 409608 470432 409672
rect 470496 409608 470512 409672
rect 470576 409608 470592 409672
rect 470656 409608 470672 409672
rect 470736 409608 470752 409672
rect 470816 409608 470854 409672
rect 470234 399894 470854 409608
rect 470234 399658 470266 399894
rect 470502 399658 470586 399894
rect 470822 399658 470854 399894
rect 470234 399574 470854 399658
rect 470234 399338 470266 399574
rect 470502 399338 470586 399574
rect 470822 399338 470854 399574
rect 470234 391085 470854 399338
rect 470234 391021 470272 391085
rect 470336 391021 470352 391085
rect 470416 391021 470432 391085
rect 470496 391021 470512 391085
rect 470576 391021 470592 391085
rect 470656 391021 470672 391085
rect 470736 391021 470752 391085
rect 470816 391021 470854 391085
rect 470234 391005 470854 391021
rect 470234 390941 470272 391005
rect 470336 390941 470352 391005
rect 470416 390941 470432 391005
rect 470496 390941 470512 391005
rect 470576 390941 470592 391005
rect 470656 390941 470672 391005
rect 470736 390941 470752 391005
rect 470816 390941 470854 391005
rect 470234 390925 470854 390941
rect 470234 390861 470272 390925
rect 470336 390861 470352 390925
rect 470416 390861 470432 390925
rect 470496 390861 470512 390925
rect 470576 390861 470592 390925
rect 470656 390861 470672 390925
rect 470736 390861 470752 390925
rect 470816 390861 470854 390925
rect 470234 390845 470854 390861
rect 470234 390781 470272 390845
rect 470336 390781 470352 390845
rect 470416 390781 470432 390845
rect 470496 390781 470512 390845
rect 470576 390781 470592 390845
rect 470656 390781 470672 390845
rect 470736 390781 470752 390845
rect 470816 390781 470854 390845
rect 470234 388912 470854 390781
rect 470234 388848 470272 388912
rect 470336 388848 470352 388912
rect 470416 388848 470432 388912
rect 470496 388848 470512 388912
rect 470576 388848 470592 388912
rect 470656 388848 470672 388912
rect 470736 388848 470752 388912
rect 470816 388848 470854 388912
rect 470234 388832 470854 388848
rect 470234 388768 470272 388832
rect 470336 388768 470352 388832
rect 470416 388768 470432 388832
rect 470496 388768 470512 388832
rect 470576 388768 470592 388832
rect 470656 388768 470672 388832
rect 470736 388768 470752 388832
rect 470816 388768 470854 388832
rect 470234 388752 470854 388768
rect 470234 388688 470272 388752
rect 470336 388688 470352 388752
rect 470416 388688 470432 388752
rect 470496 388688 470512 388752
rect 470576 388688 470592 388752
rect 470656 388688 470672 388752
rect 470736 388688 470752 388752
rect 470816 388688 470854 388752
rect 470234 388672 470854 388688
rect 470234 388608 470272 388672
rect 470336 388608 470352 388672
rect 470416 388608 470432 388672
rect 470496 388608 470512 388672
rect 470576 388608 470592 388672
rect 470656 388608 470672 388672
rect 470736 388608 470752 388672
rect 470816 388608 470854 388672
rect 470234 363894 470854 388608
rect 470234 363658 470266 363894
rect 470502 363658 470586 363894
rect 470822 363658 470854 363894
rect 470234 363574 470854 363658
rect 470234 363338 470266 363574
rect 470502 363338 470586 363574
rect 470822 363338 470854 363574
rect 470234 358485 470854 363338
rect 470234 358421 470272 358485
rect 470336 358421 470352 358485
rect 470416 358421 470432 358485
rect 470496 358421 470512 358485
rect 470576 358421 470592 358485
rect 470656 358421 470672 358485
rect 470736 358421 470752 358485
rect 470816 358421 470854 358485
rect 470234 358405 470854 358421
rect 470234 358341 470272 358405
rect 470336 358341 470352 358405
rect 470416 358341 470432 358405
rect 470496 358341 470512 358405
rect 470576 358341 470592 358405
rect 470656 358341 470672 358405
rect 470736 358341 470752 358405
rect 470816 358341 470854 358405
rect 470234 358325 470854 358341
rect 470234 358261 470272 358325
rect 470336 358261 470352 358325
rect 470416 358261 470432 358325
rect 470496 358261 470512 358325
rect 470576 358261 470592 358325
rect 470656 358261 470672 358325
rect 470736 358261 470752 358325
rect 470816 358261 470854 358325
rect 470234 358245 470854 358261
rect 470234 358181 470272 358245
rect 470336 358181 470352 358245
rect 470416 358181 470432 358245
rect 470496 358181 470512 358245
rect 470576 358181 470592 358245
rect 470656 358181 470672 358245
rect 470736 358181 470752 358245
rect 470816 358181 470854 358245
rect 470234 356312 470854 358181
rect 470234 356248 470272 356312
rect 470336 356248 470352 356312
rect 470416 356248 470432 356312
rect 470496 356248 470512 356312
rect 470576 356248 470592 356312
rect 470656 356248 470672 356312
rect 470736 356248 470752 356312
rect 470816 356248 470854 356312
rect 470234 356232 470854 356248
rect 470234 356168 470272 356232
rect 470336 356168 470352 356232
rect 470416 356168 470432 356232
rect 470496 356168 470512 356232
rect 470576 356168 470592 356232
rect 470656 356168 470672 356232
rect 470736 356168 470752 356232
rect 470816 356168 470854 356232
rect 470234 356152 470854 356168
rect 470234 356088 470272 356152
rect 470336 356088 470352 356152
rect 470416 356088 470432 356152
rect 470496 356088 470512 356152
rect 470576 356088 470592 356152
rect 470656 356088 470672 356152
rect 470736 356088 470752 356152
rect 470816 356088 470854 356152
rect 470234 356072 470854 356088
rect 470234 356008 470272 356072
rect 470336 356008 470352 356072
rect 470416 356008 470432 356072
rect 470496 356008 470512 356072
rect 470576 356008 470592 356072
rect 470656 356008 470672 356072
rect 470736 356008 470752 356072
rect 470816 356008 470854 356072
rect 470234 342484 470854 356008
rect 470234 342420 470272 342484
rect 470336 342420 470352 342484
rect 470416 342420 470432 342484
rect 470496 342420 470512 342484
rect 470576 342420 470592 342484
rect 470656 342420 470672 342484
rect 470736 342420 470752 342484
rect 470816 342420 470854 342484
rect 470234 342404 470854 342420
rect 470234 342340 470272 342404
rect 470336 342340 470352 342404
rect 470416 342340 470432 342404
rect 470496 342340 470512 342404
rect 470576 342340 470592 342404
rect 470656 342340 470672 342404
rect 470736 342340 470752 342404
rect 470816 342340 470854 342404
rect 470234 342324 470854 342340
rect 470234 342260 470272 342324
rect 470336 342260 470352 342324
rect 470416 342260 470432 342324
rect 470496 342260 470512 342324
rect 470576 342260 470592 342324
rect 470656 342260 470672 342324
rect 470736 342260 470752 342324
rect 470816 342260 470854 342324
rect 470234 342244 470854 342260
rect 470234 342180 470272 342244
rect 470336 342180 470352 342244
rect 470416 342180 470432 342244
rect 470496 342180 470512 342244
rect 470576 342180 470592 342244
rect 470656 342180 470672 342244
rect 470736 342180 470752 342244
rect 470816 342180 470854 342244
rect 470234 340312 470854 342180
rect 470234 340248 470272 340312
rect 470336 340248 470352 340312
rect 470416 340248 470432 340312
rect 470496 340248 470512 340312
rect 470576 340248 470592 340312
rect 470656 340248 470672 340312
rect 470736 340248 470752 340312
rect 470816 340248 470854 340312
rect 470234 340232 470854 340248
rect 470234 340168 470272 340232
rect 470336 340168 470352 340232
rect 470416 340168 470432 340232
rect 470496 340168 470512 340232
rect 470576 340168 470592 340232
rect 470656 340168 470672 340232
rect 470736 340168 470752 340232
rect 470816 340168 470854 340232
rect 470234 340152 470854 340168
rect 470234 340088 470272 340152
rect 470336 340088 470352 340152
rect 470416 340088 470432 340152
rect 470496 340088 470512 340152
rect 470576 340088 470592 340152
rect 470656 340088 470672 340152
rect 470736 340088 470752 340152
rect 470816 340088 470854 340152
rect 470234 340072 470854 340088
rect 470234 340008 470272 340072
rect 470336 340008 470352 340072
rect 470416 340008 470432 340072
rect 470496 340008 470512 340072
rect 470576 340008 470592 340072
rect 470656 340008 470672 340072
rect 470736 340008 470752 340072
rect 470816 340008 470854 340072
rect 470234 327894 470854 340008
rect 470234 327658 470266 327894
rect 470502 327658 470586 327894
rect 470822 327658 470854 327894
rect 470234 327574 470854 327658
rect 470234 327338 470266 327574
rect 470502 327338 470586 327574
rect 470822 327338 470854 327574
rect 470234 322484 470854 327338
rect 470234 322420 470272 322484
rect 470336 322420 470352 322484
rect 470416 322420 470432 322484
rect 470496 322420 470512 322484
rect 470576 322420 470592 322484
rect 470656 322420 470672 322484
rect 470736 322420 470752 322484
rect 470816 322420 470854 322484
rect 470234 322404 470854 322420
rect 470234 322340 470272 322404
rect 470336 322340 470352 322404
rect 470416 322340 470432 322404
rect 470496 322340 470512 322404
rect 470576 322340 470592 322404
rect 470656 322340 470672 322404
rect 470736 322340 470752 322404
rect 470816 322340 470854 322404
rect 470234 322324 470854 322340
rect 470234 322260 470272 322324
rect 470336 322260 470352 322324
rect 470416 322260 470432 322324
rect 470496 322260 470512 322324
rect 470576 322260 470592 322324
rect 470656 322260 470672 322324
rect 470736 322260 470752 322324
rect 470816 322260 470854 322324
rect 470234 322244 470854 322260
rect 470234 322180 470272 322244
rect 470336 322180 470352 322244
rect 470416 322180 470432 322244
rect 470496 322180 470512 322244
rect 470576 322180 470592 322244
rect 470656 322180 470672 322244
rect 470736 322180 470752 322244
rect 470816 322180 470854 322244
rect 470234 320312 470854 322180
rect 470234 320248 470272 320312
rect 470336 320248 470352 320312
rect 470416 320248 470432 320312
rect 470496 320248 470512 320312
rect 470576 320248 470592 320312
rect 470656 320248 470672 320312
rect 470736 320248 470752 320312
rect 470816 320248 470854 320312
rect 470234 320232 470854 320248
rect 470234 320168 470272 320232
rect 470336 320168 470352 320232
rect 470416 320168 470432 320232
rect 470496 320168 470512 320232
rect 470576 320168 470592 320232
rect 470656 320168 470672 320232
rect 470736 320168 470752 320232
rect 470816 320168 470854 320232
rect 470234 320152 470854 320168
rect 470234 320088 470272 320152
rect 470336 320088 470352 320152
rect 470416 320088 470432 320152
rect 470496 320088 470512 320152
rect 470576 320088 470592 320152
rect 470656 320088 470672 320152
rect 470736 320088 470752 320152
rect 470816 320088 470854 320152
rect 470234 320072 470854 320088
rect 470234 320008 470272 320072
rect 470336 320008 470352 320072
rect 470416 320008 470432 320072
rect 470496 320008 470512 320072
rect 470576 320008 470592 320072
rect 470656 320008 470672 320072
rect 470736 320008 470752 320072
rect 470816 320008 470854 320072
rect 470234 307084 470854 320008
rect 470234 307020 470272 307084
rect 470336 307020 470352 307084
rect 470416 307020 470432 307084
rect 470496 307020 470512 307084
rect 470576 307020 470592 307084
rect 470656 307020 470672 307084
rect 470736 307020 470752 307084
rect 470816 307020 470854 307084
rect 470234 307004 470854 307020
rect 470234 306940 470272 307004
rect 470336 306940 470352 307004
rect 470416 306940 470432 307004
rect 470496 306940 470512 307004
rect 470576 306940 470592 307004
rect 470656 306940 470672 307004
rect 470736 306940 470752 307004
rect 470816 306940 470854 307004
rect 470234 306924 470854 306940
rect 470234 306860 470272 306924
rect 470336 306860 470352 306924
rect 470416 306860 470432 306924
rect 470496 306860 470512 306924
rect 470576 306860 470592 306924
rect 470656 306860 470672 306924
rect 470736 306860 470752 306924
rect 470816 306860 470854 306924
rect 470234 306844 470854 306860
rect 470234 306780 470272 306844
rect 470336 306780 470352 306844
rect 470416 306780 470432 306844
rect 470496 306780 470512 306844
rect 470576 306780 470592 306844
rect 470656 306780 470672 306844
rect 470736 306780 470752 306844
rect 470816 306780 470854 306844
rect 470234 304912 470854 306780
rect 470234 304848 470272 304912
rect 470336 304848 470352 304912
rect 470416 304848 470432 304912
rect 470496 304848 470512 304912
rect 470576 304848 470592 304912
rect 470656 304848 470672 304912
rect 470736 304848 470752 304912
rect 470816 304848 470854 304912
rect 470234 304832 470854 304848
rect 470234 304768 470272 304832
rect 470336 304768 470352 304832
rect 470416 304768 470432 304832
rect 470496 304768 470512 304832
rect 470576 304768 470592 304832
rect 470656 304768 470672 304832
rect 470736 304768 470752 304832
rect 470816 304768 470854 304832
rect 470234 304752 470854 304768
rect 470234 304688 470272 304752
rect 470336 304688 470352 304752
rect 470416 304688 470432 304752
rect 470496 304688 470512 304752
rect 470576 304688 470592 304752
rect 470656 304688 470672 304752
rect 470736 304688 470752 304752
rect 470816 304688 470854 304752
rect 470234 304672 470854 304688
rect 470234 304608 470272 304672
rect 470336 304608 470352 304672
rect 470416 304608 470432 304672
rect 470496 304608 470512 304672
rect 470576 304608 470592 304672
rect 470656 304608 470672 304672
rect 470736 304608 470752 304672
rect 470816 304608 470854 304672
rect 470234 291894 470854 304608
rect 470234 291658 470266 291894
rect 470502 291658 470586 291894
rect 470822 291658 470854 291894
rect 470234 291574 470854 291658
rect 470234 291338 470266 291574
rect 470502 291338 470586 291574
rect 470822 291338 470854 291574
rect 470234 287485 470854 291338
rect 470234 287421 470272 287485
rect 470336 287421 470352 287485
rect 470416 287421 470432 287485
rect 470496 287421 470512 287485
rect 470576 287421 470592 287485
rect 470656 287421 470672 287485
rect 470736 287421 470752 287485
rect 470816 287421 470854 287485
rect 470234 287405 470854 287421
rect 470234 287341 470272 287405
rect 470336 287341 470352 287405
rect 470416 287341 470432 287405
rect 470496 287341 470512 287405
rect 470576 287341 470592 287405
rect 470656 287341 470672 287405
rect 470736 287341 470752 287405
rect 470816 287341 470854 287405
rect 470234 287325 470854 287341
rect 470234 287261 470272 287325
rect 470336 287261 470352 287325
rect 470416 287261 470432 287325
rect 470496 287261 470512 287325
rect 470576 287261 470592 287325
rect 470656 287261 470672 287325
rect 470736 287261 470752 287325
rect 470816 287261 470854 287325
rect 470234 287245 470854 287261
rect 470234 287181 470272 287245
rect 470336 287181 470352 287245
rect 470416 287181 470432 287245
rect 470496 287181 470512 287245
rect 470576 287181 470592 287245
rect 470656 287181 470672 287245
rect 470736 287181 470752 287245
rect 470816 287181 470854 287245
rect 470234 285312 470854 287181
rect 470234 285248 470272 285312
rect 470336 285248 470352 285312
rect 470416 285248 470432 285312
rect 470496 285248 470512 285312
rect 470576 285248 470592 285312
rect 470656 285248 470672 285312
rect 470736 285248 470752 285312
rect 470816 285248 470854 285312
rect 470234 285232 470854 285248
rect 470234 285168 470272 285232
rect 470336 285168 470352 285232
rect 470416 285168 470432 285232
rect 470496 285168 470512 285232
rect 470576 285168 470592 285232
rect 470656 285168 470672 285232
rect 470736 285168 470752 285232
rect 470816 285168 470854 285232
rect 470234 285152 470854 285168
rect 470234 285088 470272 285152
rect 470336 285088 470352 285152
rect 470416 285088 470432 285152
rect 470496 285088 470512 285152
rect 470576 285088 470592 285152
rect 470656 285088 470672 285152
rect 470736 285088 470752 285152
rect 470816 285088 470854 285152
rect 470234 285072 470854 285088
rect 470234 285008 470272 285072
rect 470336 285008 470352 285072
rect 470416 285008 470432 285072
rect 470496 285008 470512 285072
rect 470576 285008 470592 285072
rect 470656 285008 470672 285072
rect 470736 285008 470752 285072
rect 470816 285008 470854 285072
rect 470234 267485 470854 285008
rect 470234 267421 470272 267485
rect 470336 267421 470352 267485
rect 470416 267421 470432 267485
rect 470496 267421 470512 267485
rect 470576 267421 470592 267485
rect 470656 267421 470672 267485
rect 470736 267421 470752 267485
rect 470816 267421 470854 267485
rect 470234 267405 470854 267421
rect 470234 267341 470272 267405
rect 470336 267341 470352 267405
rect 470416 267341 470432 267405
rect 470496 267341 470512 267405
rect 470576 267341 470592 267405
rect 470656 267341 470672 267405
rect 470736 267341 470752 267405
rect 470816 267341 470854 267405
rect 470234 267325 470854 267341
rect 470234 267261 470272 267325
rect 470336 267261 470352 267325
rect 470416 267261 470432 267325
rect 470496 267261 470512 267325
rect 470576 267261 470592 267325
rect 470656 267261 470672 267325
rect 470736 267261 470752 267325
rect 470816 267261 470854 267325
rect 470234 267245 470854 267261
rect 470234 267181 470272 267245
rect 470336 267181 470352 267245
rect 470416 267181 470432 267245
rect 470496 267181 470512 267245
rect 470576 267181 470592 267245
rect 470656 267181 470672 267245
rect 470736 267181 470752 267245
rect 470816 267181 470854 267245
rect 470234 265312 470854 267181
rect 470234 265248 470272 265312
rect 470336 265248 470352 265312
rect 470416 265248 470432 265312
rect 470496 265248 470512 265312
rect 470576 265248 470592 265312
rect 470656 265248 470672 265312
rect 470736 265248 470752 265312
rect 470816 265248 470854 265312
rect 470234 265232 470854 265248
rect 470234 265168 470272 265232
rect 470336 265168 470352 265232
rect 470416 265168 470432 265232
rect 470496 265168 470512 265232
rect 470576 265168 470592 265232
rect 470656 265168 470672 265232
rect 470736 265168 470752 265232
rect 470816 265168 470854 265232
rect 470234 265152 470854 265168
rect 470234 265088 470272 265152
rect 470336 265088 470352 265152
rect 470416 265088 470432 265152
rect 470496 265088 470512 265152
rect 470576 265088 470592 265152
rect 470656 265088 470672 265152
rect 470736 265088 470752 265152
rect 470816 265088 470854 265152
rect 470234 265072 470854 265088
rect 470234 265008 470272 265072
rect 470336 265008 470352 265072
rect 470416 265008 470432 265072
rect 470496 265008 470512 265072
rect 470576 265008 470592 265072
rect 470656 265008 470672 265072
rect 470736 265008 470752 265072
rect 470816 265008 470854 265072
rect 470234 255894 470854 265008
rect 470234 255658 470266 255894
rect 470502 255658 470586 255894
rect 470822 255658 470854 255894
rect 470234 255574 470854 255658
rect 470234 255338 470266 255574
rect 470502 255338 470586 255574
rect 470822 255338 470854 255574
rect 470234 219894 470854 255338
rect 470234 219658 470266 219894
rect 470502 219658 470586 219894
rect 470822 219658 470854 219894
rect 470234 219574 470854 219658
rect 470234 219338 470266 219574
rect 470502 219338 470586 219574
rect 470822 219338 470854 219574
rect 470234 183894 470854 219338
rect 470234 183658 470266 183894
rect 470502 183658 470586 183894
rect 470822 183658 470854 183894
rect 470234 183574 470854 183658
rect 470234 183338 470266 183574
rect 470502 183338 470586 183574
rect 470822 183338 470854 183574
rect 470234 147894 470854 183338
rect 470234 147658 470266 147894
rect 470502 147658 470586 147894
rect 470822 147658 470854 147894
rect 470234 147574 470854 147658
rect 470234 147338 470266 147574
rect 470502 147338 470586 147574
rect 470822 147338 470854 147574
rect 470234 111894 470854 147338
rect 470234 111658 470266 111894
rect 470502 111658 470586 111894
rect 470822 111658 470854 111894
rect 470234 111574 470854 111658
rect 470234 111338 470266 111574
rect 470502 111338 470586 111574
rect 470822 111338 470854 111574
rect 470234 75894 470854 111338
rect 470234 75658 470266 75894
rect 470502 75658 470586 75894
rect 470822 75658 470854 75894
rect 470234 75574 470854 75658
rect 470234 75338 470266 75574
rect 470502 75338 470586 75574
rect 470822 75338 470854 75574
rect 470234 39894 470854 75338
rect 470234 39658 470266 39894
rect 470502 39658 470586 39894
rect 470822 39658 470854 39894
rect 470234 39574 470854 39658
rect 470234 39338 470266 39574
rect 470502 39338 470586 39574
rect 470822 39338 470854 39574
rect 470234 3894 470854 39338
rect 470234 3658 470266 3894
rect 470502 3658 470586 3894
rect 470822 3658 470854 3894
rect 470234 3574 470854 3658
rect 470234 3338 470266 3574
rect 470502 3338 470586 3574
rect 470822 3338 470854 3574
rect 470234 -1306 470854 3338
rect 470234 -1542 470266 -1306
rect 470502 -1542 470586 -1306
rect 470822 -1542 470854 -1306
rect 470234 -1626 470854 -1542
rect 470234 -1862 470266 -1626
rect 470502 -1862 470586 -1626
rect 470822 -1862 470854 -1626
rect 470234 -7654 470854 -1862
rect 471474 706758 472094 711590
rect 471474 706522 471506 706758
rect 471742 706522 471826 706758
rect 472062 706522 472094 706758
rect 471474 706438 472094 706522
rect 471474 706202 471506 706438
rect 471742 706202 471826 706438
rect 472062 706202 472094 706438
rect 471474 689134 472094 706202
rect 471474 688898 471506 689134
rect 471742 688898 471826 689134
rect 472062 688898 472094 689134
rect 471474 688814 472094 688898
rect 471474 688578 471506 688814
rect 471742 688578 471826 688814
rect 472062 688578 472094 688814
rect 471474 653134 472094 688578
rect 471474 652898 471506 653134
rect 471742 652898 471826 653134
rect 472062 652898 472094 653134
rect 471474 652814 472094 652898
rect 471474 652578 471506 652814
rect 471742 652578 471826 652814
rect 472062 652578 472094 652814
rect 471474 617134 472094 652578
rect 471474 616898 471506 617134
rect 471742 616898 471826 617134
rect 472062 616898 472094 617134
rect 471474 616814 472094 616898
rect 471474 616578 471506 616814
rect 471742 616578 471826 616814
rect 472062 616578 472094 616814
rect 471474 581134 472094 616578
rect 471474 580898 471506 581134
rect 471742 580898 471826 581134
rect 472062 580898 472094 581134
rect 471474 580814 472094 580898
rect 471474 580578 471506 580814
rect 471742 580578 471826 580814
rect 472062 580578 472094 580814
rect 471474 545134 472094 580578
rect 471474 544898 471506 545134
rect 471742 544898 471826 545134
rect 472062 544898 472094 545134
rect 471474 544814 472094 544898
rect 471474 544578 471506 544814
rect 471742 544578 471826 544814
rect 472062 544578 472094 544814
rect 471474 509134 472094 544578
rect 471474 508898 471506 509134
rect 471742 508898 471826 509134
rect 472062 508898 472094 509134
rect 471474 508814 472094 508898
rect 471474 508578 471506 508814
rect 471742 508578 471826 508814
rect 472062 508578 472094 508814
rect 471474 473134 472094 508578
rect 471474 472898 471506 473134
rect 471742 472898 471826 473134
rect 472062 472898 472094 473134
rect 471474 472814 472094 472898
rect 471474 472578 471506 472814
rect 471742 472578 471826 472814
rect 472062 472578 472094 472814
rect 471474 437134 472094 472578
rect 471474 436898 471506 437134
rect 471742 436898 471826 437134
rect 472062 436898 472094 437134
rect 471474 436814 472094 436898
rect 471474 436578 471506 436814
rect 471742 436578 471826 436814
rect 472062 436578 472094 436814
rect 471474 401134 472094 436578
rect 471474 400898 471506 401134
rect 471742 400898 471826 401134
rect 472062 400898 472094 401134
rect 471474 400814 472094 400898
rect 471474 400578 471506 400814
rect 471742 400578 471826 400814
rect 472062 400578 472094 400814
rect 471474 365134 472094 400578
rect 471474 364898 471506 365134
rect 471742 364898 471826 365134
rect 472062 364898 472094 365134
rect 471474 364814 472094 364898
rect 471474 364578 471506 364814
rect 471742 364578 471826 364814
rect 472062 364578 472094 364814
rect 471474 329134 472094 364578
rect 472714 707718 473334 711590
rect 472714 707482 472746 707718
rect 472982 707482 473066 707718
rect 473302 707482 473334 707718
rect 472714 707398 473334 707482
rect 472714 707162 472746 707398
rect 472982 707162 473066 707398
rect 473302 707162 473334 707398
rect 472714 690374 473334 707162
rect 472714 690138 472746 690374
rect 472982 690138 473066 690374
rect 473302 690138 473334 690374
rect 472714 690054 473334 690138
rect 472714 689818 472746 690054
rect 472982 689818 473066 690054
rect 473302 689818 473334 690054
rect 472714 654374 473334 689818
rect 472714 654138 472746 654374
rect 472982 654138 473066 654374
rect 473302 654138 473334 654374
rect 472714 654054 473334 654138
rect 472714 653818 472746 654054
rect 472982 653818 473066 654054
rect 473302 653818 473334 654054
rect 472714 618374 473334 653818
rect 472714 618138 472746 618374
rect 472982 618138 473066 618374
rect 473302 618138 473334 618374
rect 472714 618054 473334 618138
rect 472714 617818 472746 618054
rect 472982 617818 473066 618054
rect 473302 617818 473334 618054
rect 472714 582374 473334 617818
rect 472714 582138 472746 582374
rect 472982 582138 473066 582374
rect 473302 582138 473334 582374
rect 472714 582054 473334 582138
rect 472714 581818 472746 582054
rect 472982 581818 473066 582054
rect 473302 581818 473334 582054
rect 472714 546374 473334 581818
rect 472714 546138 472746 546374
rect 472982 546138 473066 546374
rect 473302 546138 473334 546374
rect 472714 546054 473334 546138
rect 472714 545818 472746 546054
rect 472982 545818 473066 546054
rect 473302 545818 473334 546054
rect 472714 510374 473334 545818
rect 472714 510138 472746 510374
rect 472982 510138 473066 510374
rect 473302 510138 473334 510374
rect 472714 510054 473334 510138
rect 472714 509818 472746 510054
rect 472982 509818 473066 510054
rect 473302 509818 473334 510054
rect 472714 474374 473334 509818
rect 472714 474138 472746 474374
rect 472982 474138 473066 474374
rect 473302 474138 473334 474374
rect 472714 474054 473334 474138
rect 472714 473818 472746 474054
rect 472982 473818 473066 474054
rect 473302 473818 473334 474054
rect 472714 438374 473334 473818
rect 473954 708678 474574 711590
rect 473954 708442 473986 708678
rect 474222 708442 474306 708678
rect 474542 708442 474574 708678
rect 473954 708358 474574 708442
rect 473954 708122 473986 708358
rect 474222 708122 474306 708358
rect 474542 708122 474574 708358
rect 473954 691614 474574 708122
rect 473954 691378 473986 691614
rect 474222 691378 474306 691614
rect 474542 691378 474574 691614
rect 473954 691294 474574 691378
rect 473954 691058 473986 691294
rect 474222 691058 474306 691294
rect 474542 691058 474574 691294
rect 473954 655614 474574 691058
rect 473954 655378 473986 655614
rect 474222 655378 474306 655614
rect 474542 655378 474574 655614
rect 473954 655294 474574 655378
rect 473954 655058 473986 655294
rect 474222 655058 474306 655294
rect 474542 655058 474574 655294
rect 473954 619614 474574 655058
rect 473954 619378 473986 619614
rect 474222 619378 474306 619614
rect 474542 619378 474574 619614
rect 473954 619294 474574 619378
rect 473954 619058 473986 619294
rect 474222 619058 474306 619294
rect 474542 619058 474574 619294
rect 473954 583614 474574 619058
rect 473954 583378 473986 583614
rect 474222 583378 474306 583614
rect 474542 583378 474574 583614
rect 473954 583294 474574 583378
rect 473954 583058 473986 583294
rect 474222 583058 474306 583294
rect 474542 583058 474574 583294
rect 473954 547614 474574 583058
rect 473954 547378 473986 547614
rect 474222 547378 474306 547614
rect 474542 547378 474574 547614
rect 473954 547294 474574 547378
rect 473954 547058 473986 547294
rect 474222 547058 474306 547294
rect 474542 547058 474574 547294
rect 473954 511614 474574 547058
rect 473954 511378 473986 511614
rect 474222 511378 474306 511614
rect 474542 511378 474574 511614
rect 473954 511294 474574 511378
rect 473954 511058 473986 511294
rect 474222 511058 474306 511294
rect 474542 511058 474574 511294
rect 473954 475614 474574 511058
rect 473954 475378 473986 475614
rect 474222 475378 474306 475614
rect 474542 475378 474574 475614
rect 473954 475294 474574 475378
rect 473954 475058 473986 475294
rect 474222 475058 474306 475294
rect 474542 475058 474574 475294
rect 473675 449716 473741 449717
rect 473675 449652 473676 449716
rect 473740 449652 473741 449716
rect 473675 449651 473741 449652
rect 472714 438138 472746 438374
rect 472982 438138 473066 438374
rect 473302 438138 473334 438374
rect 472714 438054 473334 438138
rect 472714 437818 472746 438054
rect 472982 437818 473066 438054
rect 473302 437818 473334 438054
rect 472714 402374 473334 437818
rect 473678 431901 473738 449651
rect 473954 439614 474574 475058
rect 473954 439378 473986 439614
rect 474222 439378 474306 439614
rect 474542 439378 474574 439614
rect 473954 439294 474574 439378
rect 473954 439058 473986 439294
rect 474222 439058 474306 439294
rect 474542 439058 474574 439294
rect 473675 431900 473741 431901
rect 473675 431836 473676 431900
rect 473740 431836 473741 431900
rect 473675 431835 473741 431836
rect 473678 410957 473738 431835
rect 473675 410956 473741 410957
rect 473675 410892 473676 410956
rect 473740 410892 473741 410956
rect 473675 410891 473741 410892
rect 472714 402138 472746 402374
rect 472982 402138 473066 402374
rect 473302 402138 473334 402374
rect 472714 402054 473334 402138
rect 472714 401818 472746 402054
rect 472982 401818 473066 402054
rect 473302 401818 473334 402054
rect 472714 366374 473334 401818
rect 473678 392053 473738 410891
rect 473954 403614 474574 439058
rect 473954 403378 473986 403614
rect 474222 403378 474306 403614
rect 474542 403378 474574 403614
rect 473954 403294 474574 403378
rect 473954 403058 473986 403294
rect 474222 403058 474306 403294
rect 474542 403058 474574 403294
rect 473675 392052 473741 392053
rect 473675 391988 473676 392052
rect 473740 391988 473741 392052
rect 473675 391987 473741 391988
rect 472714 366138 472746 366374
rect 472982 366138 473066 366374
rect 473302 366138 473334 366374
rect 472714 366054 473334 366138
rect 472714 365818 472746 366054
rect 472982 365818 473066 366054
rect 473302 365818 473334 366054
rect 472714 359060 473334 365818
rect 473954 367614 474574 403058
rect 475194 709638 475814 711590
rect 475194 709402 475226 709638
rect 475462 709402 475546 709638
rect 475782 709402 475814 709638
rect 475194 709318 475814 709402
rect 475194 709082 475226 709318
rect 475462 709082 475546 709318
rect 475782 709082 475814 709318
rect 475194 692854 475814 709082
rect 475194 692618 475226 692854
rect 475462 692618 475546 692854
rect 475782 692618 475814 692854
rect 475194 692534 475814 692618
rect 475194 692298 475226 692534
rect 475462 692298 475546 692534
rect 475782 692298 475814 692534
rect 475194 656854 475814 692298
rect 475194 656618 475226 656854
rect 475462 656618 475546 656854
rect 475782 656618 475814 656854
rect 475194 656534 475814 656618
rect 475194 656298 475226 656534
rect 475462 656298 475546 656534
rect 475782 656298 475814 656534
rect 475194 620854 475814 656298
rect 475194 620618 475226 620854
rect 475462 620618 475546 620854
rect 475782 620618 475814 620854
rect 475194 620534 475814 620618
rect 475194 620298 475226 620534
rect 475462 620298 475546 620534
rect 475782 620298 475814 620534
rect 475194 584854 475814 620298
rect 475194 584618 475226 584854
rect 475462 584618 475546 584854
rect 475782 584618 475814 584854
rect 475194 584534 475814 584618
rect 475194 584298 475226 584534
rect 475462 584298 475546 584534
rect 475782 584298 475814 584534
rect 475194 548854 475814 584298
rect 475194 548618 475226 548854
rect 475462 548618 475546 548854
rect 475782 548618 475814 548854
rect 475194 548534 475814 548618
rect 475194 548298 475226 548534
rect 475462 548298 475546 548534
rect 475782 548298 475814 548534
rect 475194 512854 475814 548298
rect 475194 512618 475226 512854
rect 475462 512618 475546 512854
rect 475782 512618 475814 512854
rect 475194 512534 475814 512618
rect 475194 512298 475226 512534
rect 475462 512298 475546 512534
rect 475782 512298 475814 512534
rect 475194 476854 475814 512298
rect 475194 476618 475226 476854
rect 475462 476618 475546 476854
rect 475782 476618 475814 476854
rect 475194 476534 475814 476618
rect 475194 476298 475226 476534
rect 475462 476298 475546 476534
rect 475782 476298 475814 476534
rect 475194 440854 475814 476298
rect 475194 440618 475226 440854
rect 475462 440618 475546 440854
rect 475782 440618 475814 440854
rect 475194 440534 475814 440618
rect 475194 440298 475226 440534
rect 475462 440298 475546 440534
rect 475782 440298 475814 440534
rect 475194 404854 475814 440298
rect 475194 404618 475226 404854
rect 475462 404618 475546 404854
rect 475782 404618 475814 404854
rect 475194 404534 475814 404618
rect 475194 404298 475226 404534
rect 475462 404298 475546 404534
rect 475782 404298 475814 404534
rect 474963 392052 475029 392053
rect 474963 391988 474964 392052
rect 475028 391988 475029 392052
rect 474963 391987 475029 391988
rect 474966 389333 475026 391987
rect 474963 389332 475029 389333
rect 474963 389268 474964 389332
rect 475028 389268 475029 389332
rect 474963 389267 475029 389268
rect 473954 367378 473986 367614
rect 474222 367378 474306 367614
rect 474542 367378 474574 367614
rect 473954 367294 474574 367378
rect 473954 367058 473986 367294
rect 474222 367058 474306 367294
rect 474542 367058 474574 367294
rect 473954 359060 474574 367058
rect 474966 357509 475026 389267
rect 475194 368854 475814 404298
rect 475194 368618 475226 368854
rect 475462 368618 475546 368854
rect 475782 368618 475814 368854
rect 475194 368534 475814 368618
rect 475194 368298 475226 368534
rect 475462 368298 475546 368534
rect 475782 368298 475814 368534
rect 475194 359060 475814 368298
rect 476434 710598 477054 711590
rect 476434 710362 476466 710598
rect 476702 710362 476786 710598
rect 477022 710362 477054 710598
rect 476434 710278 477054 710362
rect 476434 710042 476466 710278
rect 476702 710042 476786 710278
rect 477022 710042 477054 710278
rect 476434 694094 477054 710042
rect 476434 693858 476466 694094
rect 476702 693858 476786 694094
rect 477022 693858 477054 694094
rect 476434 693774 477054 693858
rect 476434 693538 476466 693774
rect 476702 693538 476786 693774
rect 477022 693538 477054 693774
rect 476434 658094 477054 693538
rect 476434 657858 476466 658094
rect 476702 657858 476786 658094
rect 477022 657858 477054 658094
rect 476434 657774 477054 657858
rect 476434 657538 476466 657774
rect 476702 657538 476786 657774
rect 477022 657538 477054 657774
rect 476434 622094 477054 657538
rect 476434 621858 476466 622094
rect 476702 621858 476786 622094
rect 477022 621858 477054 622094
rect 476434 621774 477054 621858
rect 476434 621538 476466 621774
rect 476702 621538 476786 621774
rect 477022 621538 477054 621774
rect 476434 586094 477054 621538
rect 476434 585858 476466 586094
rect 476702 585858 476786 586094
rect 477022 585858 477054 586094
rect 476434 585774 477054 585858
rect 476434 585538 476466 585774
rect 476702 585538 476786 585774
rect 477022 585538 477054 585774
rect 476434 550094 477054 585538
rect 476434 549858 476466 550094
rect 476702 549858 476786 550094
rect 477022 549858 477054 550094
rect 476434 549774 477054 549858
rect 476434 549538 476466 549774
rect 476702 549538 476786 549774
rect 477022 549538 477054 549774
rect 476434 514094 477054 549538
rect 476434 513858 476466 514094
rect 476702 513858 476786 514094
rect 477022 513858 477054 514094
rect 476434 513774 477054 513858
rect 476434 513538 476466 513774
rect 476702 513538 476786 513774
rect 477022 513538 477054 513774
rect 476434 478094 477054 513538
rect 476434 477858 476466 478094
rect 476702 477858 476786 478094
rect 477022 477858 477054 478094
rect 476434 477774 477054 477858
rect 476434 477538 476466 477774
rect 476702 477538 476786 477774
rect 477022 477538 477054 477774
rect 476434 442094 477054 477538
rect 476434 441858 476466 442094
rect 476702 441858 476786 442094
rect 477022 441858 477054 442094
rect 476434 441774 477054 441858
rect 476434 441538 476466 441774
rect 476702 441538 476786 441774
rect 477022 441538 477054 441774
rect 476434 406094 477054 441538
rect 476434 405858 476466 406094
rect 476702 405858 476786 406094
rect 477022 405858 477054 406094
rect 476434 405774 477054 405858
rect 476434 405538 476466 405774
rect 476702 405538 476786 405774
rect 477022 405538 477054 405774
rect 476434 370094 477054 405538
rect 476434 369858 476466 370094
rect 476702 369858 476786 370094
rect 477022 369858 477054 370094
rect 476434 369774 477054 369858
rect 476434 369538 476466 369774
rect 476702 369538 476786 369774
rect 477022 369538 477054 369774
rect 476434 359060 477054 369538
rect 477674 711558 478294 711590
rect 477674 711322 477706 711558
rect 477942 711322 478026 711558
rect 478262 711322 478294 711558
rect 477674 711238 478294 711322
rect 477674 711002 477706 711238
rect 477942 711002 478026 711238
rect 478262 711002 478294 711238
rect 477674 695334 478294 711002
rect 477674 695098 477706 695334
rect 477942 695098 478026 695334
rect 478262 695098 478294 695334
rect 477674 695014 478294 695098
rect 477674 694778 477706 695014
rect 477942 694778 478026 695014
rect 478262 694778 478294 695014
rect 477674 659334 478294 694778
rect 477674 659098 477706 659334
rect 477942 659098 478026 659334
rect 478262 659098 478294 659334
rect 477674 659014 478294 659098
rect 477674 658778 477706 659014
rect 477942 658778 478026 659014
rect 478262 658778 478294 659014
rect 477674 623334 478294 658778
rect 477674 623098 477706 623334
rect 477942 623098 478026 623334
rect 478262 623098 478294 623334
rect 477674 623014 478294 623098
rect 477674 622778 477706 623014
rect 477942 622778 478026 623014
rect 478262 622778 478294 623014
rect 477674 587334 478294 622778
rect 477674 587098 477706 587334
rect 477942 587098 478026 587334
rect 478262 587098 478294 587334
rect 477674 587014 478294 587098
rect 477674 586778 477706 587014
rect 477942 586778 478026 587014
rect 478262 586778 478294 587014
rect 477674 551334 478294 586778
rect 477674 551098 477706 551334
rect 477942 551098 478026 551334
rect 478262 551098 478294 551334
rect 477674 551014 478294 551098
rect 477674 550778 477706 551014
rect 477942 550778 478026 551014
rect 478262 550778 478294 551014
rect 477674 515334 478294 550778
rect 477674 515098 477706 515334
rect 477942 515098 478026 515334
rect 478262 515098 478294 515334
rect 477674 515014 478294 515098
rect 477674 514778 477706 515014
rect 477942 514778 478026 515014
rect 478262 514778 478294 515014
rect 477674 479334 478294 514778
rect 477674 479098 477706 479334
rect 477942 479098 478026 479334
rect 478262 479098 478294 479334
rect 477674 479014 478294 479098
rect 477674 478778 477706 479014
rect 477942 478778 478026 479014
rect 478262 478778 478294 479014
rect 477674 443334 478294 478778
rect 504994 704838 505614 711590
rect 504994 704602 505026 704838
rect 505262 704602 505346 704838
rect 505582 704602 505614 704838
rect 504994 704518 505614 704602
rect 504994 704282 505026 704518
rect 505262 704282 505346 704518
rect 505582 704282 505614 704518
rect 504994 686654 505614 704282
rect 504994 686418 505026 686654
rect 505262 686418 505346 686654
rect 505582 686418 505614 686654
rect 504994 686334 505614 686418
rect 504994 686098 505026 686334
rect 505262 686098 505346 686334
rect 505582 686098 505614 686334
rect 504994 650654 505614 686098
rect 504994 650418 505026 650654
rect 505262 650418 505346 650654
rect 505582 650418 505614 650654
rect 504994 650334 505614 650418
rect 504994 650098 505026 650334
rect 505262 650098 505346 650334
rect 505582 650098 505614 650334
rect 504994 614654 505614 650098
rect 504994 614418 505026 614654
rect 505262 614418 505346 614654
rect 505582 614418 505614 614654
rect 504994 614334 505614 614418
rect 504994 614098 505026 614334
rect 505262 614098 505346 614334
rect 505582 614098 505614 614334
rect 504994 578654 505614 614098
rect 504994 578418 505026 578654
rect 505262 578418 505346 578654
rect 505582 578418 505614 578654
rect 504994 578334 505614 578418
rect 504994 578098 505026 578334
rect 505262 578098 505346 578334
rect 505582 578098 505614 578334
rect 504994 542654 505614 578098
rect 504994 542418 505026 542654
rect 505262 542418 505346 542654
rect 505582 542418 505614 542654
rect 504994 542334 505614 542418
rect 504994 542098 505026 542334
rect 505262 542098 505346 542334
rect 505582 542098 505614 542334
rect 504994 506654 505614 542098
rect 504994 506418 505026 506654
rect 505262 506418 505346 506654
rect 505582 506418 505614 506654
rect 504994 506334 505614 506418
rect 504994 506098 505026 506334
rect 505262 506098 505346 506334
rect 505582 506098 505614 506334
rect 504994 470654 505614 506098
rect 504994 470418 505026 470654
rect 505262 470418 505346 470654
rect 505582 470418 505614 470654
rect 504994 470334 505614 470418
rect 504994 470098 505026 470334
rect 505262 470098 505346 470334
rect 505582 470098 505614 470334
rect 478459 450260 478525 450261
rect 478459 450196 478460 450260
rect 478524 450196 478525 450260
rect 478459 450195 478525 450196
rect 481219 450260 481285 450261
rect 481219 450196 481220 450260
rect 481284 450196 481285 450260
rect 481219 450195 481285 450196
rect 484163 450260 484229 450261
rect 484163 450196 484164 450260
rect 484228 450196 484229 450260
rect 484163 450195 484229 450196
rect 487843 450260 487909 450261
rect 487843 450196 487844 450260
rect 487908 450196 487909 450260
rect 487843 450195 487909 450196
rect 477674 443098 477706 443334
rect 477942 443098 478026 443334
rect 478262 443098 478294 443334
rect 477674 443014 478294 443098
rect 477674 442778 477706 443014
rect 477942 442778 478026 443014
rect 478262 442778 478294 443014
rect 477674 407334 478294 442778
rect 478462 431629 478522 450195
rect 481222 432173 481282 450195
rect 483611 432308 483677 432309
rect 483611 432244 483612 432308
rect 483676 432244 483677 432308
rect 483611 432243 483677 432244
rect 481219 432172 481285 432173
rect 481219 432108 481220 432172
rect 481284 432108 481285 432172
rect 481219 432107 481285 432108
rect 481222 431970 481282 432107
rect 481038 431910 481282 431970
rect 483614 431970 483674 432243
rect 484166 431970 484226 450195
rect 487846 441630 487906 450195
rect 483614 431910 484226 431970
rect 487662 441570 487906 441630
rect 478459 431628 478525 431629
rect 478459 431564 478460 431628
rect 478524 431564 478525 431628
rect 478459 431563 478525 431564
rect 478462 410141 478522 431563
rect 480115 427956 480181 427957
rect 480115 427892 480116 427956
rect 480180 427892 480181 427956
rect 480115 427891 480181 427892
rect 478459 410140 478525 410141
rect 478459 410076 478460 410140
rect 478524 410076 478525 410140
rect 478459 410075 478525 410076
rect 477674 407098 477706 407334
rect 477942 407098 478026 407334
rect 478262 407098 478294 407334
rect 477674 407014 478294 407098
rect 477674 406778 477706 407014
rect 477942 406778 478026 407014
rect 478262 406778 478294 407014
rect 477674 371334 478294 406778
rect 478462 402990 478522 410075
rect 480118 407557 480178 427891
rect 481038 422310 481098 431910
rect 483614 422310 483674 431910
rect 487662 431901 487722 441570
rect 504994 434654 505614 470098
rect 504994 434418 505026 434654
rect 505262 434418 505346 434654
rect 505582 434418 505614 434654
rect 504994 434334 505614 434418
rect 504994 434098 505026 434334
rect 505262 434098 505346 434334
rect 505582 434098 505614 434334
rect 487659 431900 487725 431901
rect 487659 431836 487660 431900
rect 487724 431836 487725 431900
rect 487659 431835 487725 431836
rect 486555 427956 486621 427957
rect 486555 427892 486556 427956
rect 486620 427892 486621 427956
rect 486555 427891 486621 427892
rect 481038 422250 481466 422310
rect 483614 422250 484226 422310
rect 481406 410141 481466 422250
rect 484166 410413 484226 422250
rect 484163 410412 484229 410413
rect 484163 410348 484164 410412
rect 484228 410348 484229 410412
rect 484163 410347 484229 410348
rect 481403 410140 481469 410141
rect 481403 410076 481404 410140
rect 481468 410076 481469 410140
rect 481403 410075 481469 410076
rect 480115 407556 480181 407557
rect 480115 407492 480116 407556
rect 480180 407492 480181 407556
rect 480115 407491 480181 407492
rect 478462 402930 478706 402990
rect 478646 389333 478706 402930
rect 481406 393330 481466 410075
rect 482875 407148 482941 407149
rect 482875 407084 482876 407148
rect 482940 407084 482941 407148
rect 482875 407083 482941 407084
rect 481406 393270 481834 393330
rect 481774 389469 481834 393270
rect 481771 389468 481837 389469
rect 481771 389404 481772 389468
rect 481836 389404 481837 389468
rect 481771 389403 481837 389404
rect 478643 389332 478709 389333
rect 478643 389268 478644 389332
rect 478708 389268 478709 389332
rect 478643 389267 478709 389268
rect 477674 371098 477706 371334
rect 477942 371098 478026 371334
rect 478262 371098 478294 371334
rect 477674 371014 478294 371098
rect 477674 370778 477706 371014
rect 477942 370778 478026 371014
rect 478262 370778 478294 371014
rect 477674 359060 478294 370778
rect 478646 358053 478706 389267
rect 481774 358053 481834 389403
rect 482878 370157 482938 407083
rect 484166 393330 484226 410347
rect 485635 407148 485701 407149
rect 485635 407084 485636 407148
rect 485700 407084 485701 407148
rect 485635 407083 485701 407084
rect 484166 393270 484962 393330
rect 484902 390298 484962 393270
rect 484899 390297 484965 390298
rect 484899 390233 484900 390297
rect 484964 390233 484965 390297
rect 484899 390232 484965 390233
rect 482875 370156 482941 370157
rect 482875 370092 482876 370156
rect 482940 370092 482941 370156
rect 482875 370091 482941 370092
rect 484902 358053 484962 390232
rect 478643 358052 478709 358053
rect 478643 357988 478644 358052
rect 478708 357988 478709 358052
rect 478643 357987 478709 357988
rect 481771 358052 481837 358053
rect 481771 357988 481772 358052
rect 481836 357988 481837 358052
rect 481771 357987 481837 357988
rect 484899 358052 484965 358053
rect 484899 357988 484900 358052
rect 484964 357988 484965 358052
rect 484899 357987 484965 357988
rect 474963 357508 475029 357509
rect 474963 357444 474964 357508
rect 475028 357444 475029 357508
rect 474963 357443 475029 357444
rect 474966 357370 475026 357443
rect 474966 357310 475394 357370
rect 475334 356690 475394 357310
rect 474966 356630 475394 356690
rect 471474 328898 471506 329134
rect 471742 328898 471826 329134
rect 472062 328898 472094 329134
rect 471474 328814 472094 328898
rect 471474 328578 471506 328814
rect 471742 328578 471826 328814
rect 472062 328578 472094 328814
rect 471474 293134 472094 328578
rect 471474 292898 471506 293134
rect 471742 292898 471826 293134
rect 472062 292898 472094 293134
rect 471474 292814 472094 292898
rect 471474 292578 471506 292814
rect 471742 292578 471826 292814
rect 472062 292578 472094 292814
rect 471474 257134 472094 292578
rect 472714 330374 473334 354615
rect 473675 343772 473741 343773
rect 473675 343708 473676 343772
rect 473740 343708 473741 343772
rect 473675 343707 473741 343708
rect 473678 340509 473738 343707
rect 473675 340508 473741 340509
rect 473675 340444 473676 340508
rect 473740 340444 473741 340508
rect 473675 340443 473741 340444
rect 472714 330138 472746 330374
rect 472982 330138 473066 330374
rect 473302 330138 473334 330374
rect 472714 330054 473334 330138
rect 472714 329818 472746 330054
rect 472982 329818 473066 330054
rect 473302 329818 473334 330054
rect 472714 294374 473334 329818
rect 473678 321333 473738 340443
rect 473954 331614 474574 354615
rect 474966 343773 475026 356630
rect 474963 343772 475029 343773
rect 474963 343708 474964 343772
rect 475028 343708 475029 343772
rect 474963 343707 475029 343708
rect 473954 331378 473986 331614
rect 474222 331378 474306 331614
rect 474542 331378 474574 331614
rect 473954 331294 474574 331378
rect 473954 331058 473986 331294
rect 474222 331058 474306 331294
rect 474542 331058 474574 331294
rect 473675 321332 473741 321333
rect 473675 321268 473676 321332
rect 473740 321268 473741 321332
rect 473675 321267 473741 321268
rect 473678 305965 473738 321267
rect 473675 305964 473741 305965
rect 473675 305900 473676 305964
rect 473740 305900 473741 305964
rect 473675 305899 473741 305900
rect 472714 294138 472746 294374
rect 472982 294138 473066 294374
rect 473302 294138 473334 294374
rect 472714 294054 473334 294138
rect 472714 293818 472746 294054
rect 472982 293818 473066 294054
rect 473302 293818 473334 294054
rect 472714 268060 473334 293818
rect 473678 289781 473738 305899
rect 473954 295614 474574 331058
rect 473954 295378 473986 295614
rect 474222 295378 474306 295614
rect 474542 295378 474574 295614
rect 473954 295294 474574 295378
rect 473954 295058 473986 295294
rect 474222 295058 474306 295294
rect 474542 295058 474574 295294
rect 473675 289780 473741 289781
rect 473675 289716 473676 289780
rect 473740 289716 473741 289780
rect 473675 289715 473741 289716
rect 473954 268060 474574 295058
rect 475194 332854 475814 354615
rect 475194 332618 475226 332854
rect 475462 332618 475546 332854
rect 475782 332618 475814 332854
rect 475194 332534 475814 332618
rect 475194 332298 475226 332534
rect 475462 332298 475546 332534
rect 475782 332298 475814 332534
rect 475194 296854 475814 332298
rect 475194 296618 475226 296854
rect 475462 296618 475546 296854
rect 475782 296618 475814 296854
rect 475194 296534 475814 296618
rect 475194 296298 475226 296534
rect 475462 296298 475546 296534
rect 475782 296298 475814 296534
rect 475194 268060 475814 296298
rect 476434 334094 477054 354615
rect 476434 333858 476466 334094
rect 476702 333858 476786 334094
rect 477022 333858 477054 334094
rect 476434 333774 477054 333858
rect 476434 333538 476466 333774
rect 476702 333538 476786 333774
rect 477022 333538 477054 333774
rect 476434 298094 477054 333538
rect 476434 297858 476466 298094
rect 476702 297858 476786 298094
rect 477022 297858 477054 298094
rect 476434 297774 477054 297858
rect 476434 297538 476466 297774
rect 476702 297538 476786 297774
rect 477022 297538 477054 297774
rect 476067 289780 476133 289781
rect 476067 289716 476068 289780
rect 476132 289716 476133 289780
rect 476067 289715 476133 289716
rect 476070 286653 476130 289715
rect 476067 286652 476133 286653
rect 476067 286588 476068 286652
rect 476132 286588 476133 286652
rect 476067 286587 476133 286588
rect 476070 267750 476130 286587
rect 476434 268060 477054 297538
rect 477674 335334 478294 354615
rect 478646 345030 478706 357987
rect 481774 354690 481834 357987
rect 484902 354690 484962 357987
rect 481590 354630 481834 354690
rect 484534 354630 484962 354690
rect 481590 345030 481650 354630
rect 484534 345030 484594 354630
rect 478462 344970 478706 345030
rect 481406 344970 481650 345030
rect 484166 344970 484594 345030
rect 478462 341053 478522 344970
rect 481406 341053 481466 344970
rect 484166 341053 484226 344970
rect 478459 341052 478525 341053
rect 478459 340988 478460 341052
rect 478524 340988 478525 341052
rect 478459 340987 478525 340988
rect 481403 341052 481469 341053
rect 481403 340988 481404 341052
rect 481468 340988 481469 341052
rect 481403 340987 481469 340988
rect 484163 341052 484229 341053
rect 484163 340988 484164 341052
rect 484228 340988 484229 341052
rect 484163 340987 484229 340988
rect 477674 335098 477706 335334
rect 477942 335098 478026 335334
rect 478262 335098 478294 335334
rect 477674 335014 478294 335098
rect 477674 334778 477706 335014
rect 477942 334778 478026 335014
rect 478262 334778 478294 335014
rect 477674 299334 478294 334778
rect 478462 325710 478522 340987
rect 481406 325710 481466 340987
rect 478462 325650 478706 325710
rect 481406 325650 481650 325710
rect 478646 320925 478706 325650
rect 481590 320925 481650 325650
rect 484166 321333 484226 340987
rect 485638 334117 485698 407083
rect 486558 335477 486618 427891
rect 487662 422310 487722 431835
rect 487662 422250 487906 422310
rect 487846 410141 487906 422250
rect 487843 410140 487909 410141
rect 487843 410076 487844 410140
rect 487908 410076 487909 410140
rect 487843 410075 487909 410076
rect 488395 410140 488461 410141
rect 488395 410076 488396 410140
rect 488460 410076 488461 410140
rect 488395 410075 488461 410076
rect 488398 390149 488458 410075
rect 504994 398654 505614 434098
rect 504994 398418 505026 398654
rect 505262 398418 505346 398654
rect 505582 398418 505614 398654
rect 504994 398334 505614 398418
rect 504994 398098 505026 398334
rect 505262 398098 505346 398334
rect 505582 398098 505614 398334
rect 488395 390148 488461 390149
rect 488395 390084 488396 390148
rect 488460 390084 488461 390148
rect 488395 390083 488461 390084
rect 486739 386476 486805 386477
rect 486739 386412 486740 386476
rect 486804 386412 486805 386476
rect 486739 386411 486805 386412
rect 486555 335476 486621 335477
rect 486555 335412 486556 335476
rect 486620 335412 486621 335476
rect 486555 335411 486621 335412
rect 485635 334116 485701 334117
rect 485635 334052 485636 334116
rect 485700 334052 485701 334116
rect 485635 334051 485701 334052
rect 486742 332757 486802 386411
rect 488398 358053 488458 390083
rect 504994 362654 505614 398098
rect 504994 362418 505026 362654
rect 505262 362418 505346 362654
rect 505582 362418 505614 362654
rect 504994 362334 505614 362418
rect 504994 362098 505026 362334
rect 505262 362098 505346 362334
rect 505582 362098 505614 362334
rect 488395 358052 488461 358053
rect 488395 357988 488396 358052
rect 488460 357988 488461 358052
rect 488395 357987 488461 357988
rect 488398 354690 488458 357987
rect 487662 354630 488458 354690
rect 487662 345030 487722 354630
rect 487662 344970 488090 345030
rect 488030 341053 488090 344970
rect 488027 341052 488093 341053
rect 488027 340988 488028 341052
rect 488092 340988 488093 341052
rect 488027 340987 488093 340988
rect 486739 332756 486805 332757
rect 486739 332692 486740 332756
rect 486804 332692 486805 332756
rect 486739 332691 486805 332692
rect 484163 321332 484229 321333
rect 484163 321268 484164 321332
rect 484228 321268 484229 321332
rect 484163 321267 484229 321268
rect 478643 320924 478709 320925
rect 478643 320860 478644 320924
rect 478708 320860 478709 320924
rect 478643 320859 478709 320860
rect 481587 320924 481653 320925
rect 481587 320860 481588 320924
rect 481652 320860 481653 320924
rect 481587 320859 481653 320860
rect 478646 306390 478706 320859
rect 481590 306390 481650 320859
rect 478646 306330 478890 306390
rect 478830 305693 478890 306330
rect 481590 306330 482202 306390
rect 481590 306101 481650 306330
rect 481587 306100 481653 306101
rect 481587 306036 481588 306100
rect 481652 306036 481653 306100
rect 481587 306035 481653 306036
rect 478827 305692 478893 305693
rect 478827 305628 478828 305692
rect 478892 305628 478893 305692
rect 478827 305627 478893 305628
rect 477674 299098 477706 299334
rect 477942 299098 478026 299334
rect 478262 299098 478294 299334
rect 477674 299014 478294 299098
rect 477674 298778 477706 299014
rect 477942 298778 478026 299014
rect 478262 298778 478294 299014
rect 477674 268060 478294 298778
rect 478830 287070 478890 305627
rect 482142 287070 482202 306330
rect 484166 305557 484226 321267
rect 488030 321061 488090 340987
rect 504994 326654 505614 362098
rect 504994 326418 505026 326654
rect 505262 326418 505346 326654
rect 505582 326418 505614 326654
rect 504994 326334 505614 326418
rect 504994 326098 505026 326334
rect 505262 326098 505346 326334
rect 505582 326098 505614 326334
rect 488027 321060 488093 321061
rect 488027 320996 488028 321060
rect 488092 320996 488093 321060
rect 488027 320995 488093 320996
rect 488030 316050 488090 320995
rect 487662 315990 488090 316050
rect 487662 306390 487722 315990
rect 487662 306373 488458 306390
rect 487659 306372 488458 306373
rect 487659 306308 487660 306372
rect 487724 306330 488458 306372
rect 487724 306308 487725 306330
rect 487659 306307 487725 306308
rect 484163 305556 484229 305557
rect 484163 305492 484164 305556
rect 484228 305492 484229 305556
rect 484163 305491 484229 305492
rect 484166 289781 484226 305491
rect 484163 289780 484229 289781
rect 484163 289716 484164 289780
rect 484228 289716 484229 289780
rect 484163 289715 484229 289716
rect 485819 289780 485885 289781
rect 485819 289716 485820 289780
rect 485884 289716 485885 289780
rect 485819 289715 485885 289716
rect 478830 287010 479074 287070
rect 482142 287010 482386 287070
rect 478830 286925 478890 287010
rect 478827 286924 478893 286925
rect 478827 286860 478828 286924
rect 478892 286860 478893 286924
rect 478827 286859 478893 286860
rect 476070 267690 476498 267750
rect 476438 265029 476498 267690
rect 479014 265981 479074 287010
rect 482326 285837 482386 287010
rect 485822 285837 485882 289715
rect 488398 288690 488458 306330
rect 504994 290654 505614 326098
rect 504994 290418 505026 290654
rect 505262 290418 505346 290654
rect 505582 290418 505614 290654
rect 504994 290334 505614 290418
rect 504994 290098 505026 290334
rect 505262 290098 505346 290334
rect 505582 290098 505614 290334
rect 488398 288630 488642 288690
rect 488582 286789 488642 288630
rect 488579 286788 488645 286789
rect 488579 286724 488580 286788
rect 488644 286724 488645 286788
rect 488579 286723 488645 286724
rect 482323 285836 482389 285837
rect 482323 285772 482324 285836
rect 482388 285772 482389 285836
rect 482323 285771 482389 285772
rect 482875 285836 482941 285837
rect 482875 285772 482876 285836
rect 482940 285772 482941 285836
rect 482875 285771 482941 285772
rect 485819 285836 485885 285837
rect 485819 285772 485820 285836
rect 485884 285772 485885 285836
rect 485819 285771 485885 285772
rect 479011 265980 479077 265981
rect 479011 265916 479012 265980
rect 479076 265916 479077 265980
rect 479011 265915 479077 265916
rect 482878 265029 482938 285771
rect 485822 265029 485882 285771
rect 488582 267750 488642 286723
rect 488582 267690 489194 267750
rect 489134 265573 489194 267690
rect 489131 265572 489197 265573
rect 489131 265508 489132 265572
rect 489196 265508 489197 265572
rect 489131 265507 489197 265508
rect 476435 265028 476501 265029
rect 476435 264964 476436 265028
rect 476500 264964 476501 265028
rect 476435 264963 476501 264964
rect 477355 265028 477421 265029
rect 477355 264964 477356 265028
rect 477420 264964 477421 265028
rect 477355 264963 477421 264964
rect 480115 265028 480181 265029
rect 480115 264964 480116 265028
rect 480180 264964 480181 265028
rect 480115 264963 480181 264964
rect 482875 265028 482941 265029
rect 482875 264964 482876 265028
rect 482940 264964 482941 265028
rect 482875 264963 482941 264964
rect 485819 265028 485885 265029
rect 485819 264964 485820 265028
rect 485884 264964 485885 265028
rect 485819 264963 485885 264964
rect 486371 265028 486437 265029
rect 486371 264964 486372 265028
rect 486436 264964 486437 265028
rect 486371 264963 486437 264964
rect 471474 256898 471506 257134
rect 471742 256898 471826 257134
rect 472062 256898 472094 257134
rect 471474 256814 472094 256898
rect 471474 256578 471506 256814
rect 471742 256578 471826 256814
rect 472062 256578 472094 256814
rect 471474 221134 472094 256578
rect 471474 220898 471506 221134
rect 471742 220898 471826 221134
rect 472062 220898 472094 221134
rect 471474 220814 472094 220898
rect 471474 220578 471506 220814
rect 471742 220578 471826 220814
rect 472062 220578 472094 220814
rect 471474 185134 472094 220578
rect 471474 184898 471506 185134
rect 471742 184898 471826 185134
rect 472062 184898 472094 185134
rect 471474 184814 472094 184898
rect 471474 184578 471506 184814
rect 471742 184578 471826 184814
rect 472062 184578 472094 184814
rect 471474 149134 472094 184578
rect 471474 148898 471506 149134
rect 471742 148898 471826 149134
rect 472062 148898 472094 149134
rect 471474 148814 472094 148898
rect 471474 148578 471506 148814
rect 471742 148578 471826 148814
rect 472062 148578 472094 148814
rect 471474 113134 472094 148578
rect 471474 112898 471506 113134
rect 471742 112898 471826 113134
rect 472062 112898 472094 113134
rect 471474 112814 472094 112898
rect 471474 112578 471506 112814
rect 471742 112578 471826 112814
rect 472062 112578 472094 112814
rect 471474 77134 472094 112578
rect 471474 76898 471506 77134
rect 471742 76898 471826 77134
rect 472062 76898 472094 77134
rect 471474 76814 472094 76898
rect 471474 76578 471506 76814
rect 471742 76578 471826 76814
rect 472062 76578 472094 76814
rect 471474 41134 472094 76578
rect 471474 40898 471506 41134
rect 471742 40898 471826 41134
rect 472062 40898 472094 41134
rect 471474 40814 472094 40898
rect 471474 40578 471506 40814
rect 471742 40578 471826 40814
rect 472062 40578 472094 40814
rect 471474 5134 472094 40578
rect 471474 4898 471506 5134
rect 471742 4898 471826 5134
rect 472062 4898 472094 5134
rect 471474 4814 472094 4898
rect 471474 4578 471506 4814
rect 471742 4578 471826 4814
rect 472062 4578 472094 4814
rect 471474 -2266 472094 4578
rect 471474 -2502 471506 -2266
rect 471742 -2502 471826 -2266
rect 472062 -2502 472094 -2266
rect 471474 -2586 472094 -2502
rect 471474 -2822 471506 -2586
rect 471742 -2822 471826 -2586
rect 472062 -2822 472094 -2586
rect 471474 -7654 472094 -2822
rect 472714 258374 473334 263615
rect 472714 258138 472746 258374
rect 472982 258138 473066 258374
rect 473302 258138 473334 258374
rect 472714 258054 473334 258138
rect 472714 257818 472746 258054
rect 472982 257818 473066 258054
rect 473302 257818 473334 258054
rect 472714 222374 473334 257818
rect 472714 222138 472746 222374
rect 472982 222138 473066 222374
rect 473302 222138 473334 222374
rect 472714 222054 473334 222138
rect 472714 221818 472746 222054
rect 472982 221818 473066 222054
rect 473302 221818 473334 222054
rect 472714 186374 473334 221818
rect 472714 186138 472746 186374
rect 472982 186138 473066 186374
rect 473302 186138 473334 186374
rect 472714 186054 473334 186138
rect 472714 185818 472746 186054
rect 472982 185818 473066 186054
rect 473302 185818 473334 186054
rect 472714 150374 473334 185818
rect 472714 150138 472746 150374
rect 472982 150138 473066 150374
rect 473302 150138 473334 150374
rect 472714 150054 473334 150138
rect 472714 149818 472746 150054
rect 472982 149818 473066 150054
rect 473302 149818 473334 150054
rect 472714 114374 473334 149818
rect 472714 114138 472746 114374
rect 472982 114138 473066 114374
rect 473302 114138 473334 114374
rect 472714 114054 473334 114138
rect 472714 113818 472746 114054
rect 472982 113818 473066 114054
rect 473302 113818 473334 114054
rect 472714 78374 473334 113818
rect 472714 78138 472746 78374
rect 472982 78138 473066 78374
rect 473302 78138 473334 78374
rect 472714 78054 473334 78138
rect 472714 77818 472746 78054
rect 472982 77818 473066 78054
rect 473302 77818 473334 78054
rect 472714 42374 473334 77818
rect 472714 42138 472746 42374
rect 472982 42138 473066 42374
rect 473302 42138 473334 42374
rect 472714 42054 473334 42138
rect 472714 41818 472746 42054
rect 472982 41818 473066 42054
rect 473302 41818 473334 42054
rect 472714 6374 473334 41818
rect 472714 6138 472746 6374
rect 472982 6138 473066 6374
rect 473302 6138 473334 6374
rect 472714 6054 473334 6138
rect 472714 5818 472746 6054
rect 472982 5818 473066 6054
rect 473302 5818 473334 6054
rect 472714 -3226 473334 5818
rect 472714 -3462 472746 -3226
rect 472982 -3462 473066 -3226
rect 473302 -3462 473334 -3226
rect 472714 -3546 473334 -3462
rect 472714 -3782 472746 -3546
rect 472982 -3782 473066 -3546
rect 473302 -3782 473334 -3546
rect 472714 -7654 473334 -3782
rect 473954 259614 474574 263615
rect 473954 259378 473986 259614
rect 474222 259378 474306 259614
rect 474542 259378 474574 259614
rect 473954 259294 474574 259378
rect 473954 259058 473986 259294
rect 474222 259058 474306 259294
rect 474542 259058 474574 259294
rect 473954 223614 474574 259058
rect 473954 223378 473986 223614
rect 474222 223378 474306 223614
rect 474542 223378 474574 223614
rect 473954 223294 474574 223378
rect 473954 223058 473986 223294
rect 474222 223058 474306 223294
rect 474542 223058 474574 223294
rect 473954 187614 474574 223058
rect 473954 187378 473986 187614
rect 474222 187378 474306 187614
rect 474542 187378 474574 187614
rect 473954 187294 474574 187378
rect 473954 187058 473986 187294
rect 474222 187058 474306 187294
rect 474542 187058 474574 187294
rect 473954 151614 474574 187058
rect 473954 151378 473986 151614
rect 474222 151378 474306 151614
rect 474542 151378 474574 151614
rect 473954 151294 474574 151378
rect 473954 151058 473986 151294
rect 474222 151058 474306 151294
rect 474542 151058 474574 151294
rect 473954 115614 474574 151058
rect 473954 115378 473986 115614
rect 474222 115378 474306 115614
rect 474542 115378 474574 115614
rect 473954 115294 474574 115378
rect 473954 115058 473986 115294
rect 474222 115058 474306 115294
rect 474542 115058 474574 115294
rect 473954 79614 474574 115058
rect 473954 79378 473986 79614
rect 474222 79378 474306 79614
rect 474542 79378 474574 79614
rect 473954 79294 474574 79378
rect 473954 79058 473986 79294
rect 474222 79058 474306 79294
rect 474542 79058 474574 79294
rect 473954 43614 474574 79058
rect 473954 43378 473986 43614
rect 474222 43378 474306 43614
rect 474542 43378 474574 43614
rect 473954 43294 474574 43378
rect 473954 43058 473986 43294
rect 474222 43058 474306 43294
rect 474542 43058 474574 43294
rect 473954 7614 474574 43058
rect 473954 7378 473986 7614
rect 474222 7378 474306 7614
rect 474542 7378 474574 7614
rect 473954 7294 474574 7378
rect 473954 7058 473986 7294
rect 474222 7058 474306 7294
rect 474542 7058 474574 7294
rect 473954 -4186 474574 7058
rect 473954 -4422 473986 -4186
rect 474222 -4422 474306 -4186
rect 474542 -4422 474574 -4186
rect 473954 -4506 474574 -4422
rect 473954 -4742 473986 -4506
rect 474222 -4742 474306 -4506
rect 474542 -4742 474574 -4506
rect 473954 -7654 474574 -4742
rect 475194 260854 475814 263615
rect 475194 260618 475226 260854
rect 475462 260618 475546 260854
rect 475782 260618 475814 260854
rect 475194 260534 475814 260618
rect 475194 260298 475226 260534
rect 475462 260298 475546 260534
rect 475782 260298 475814 260534
rect 475194 224854 475814 260298
rect 475194 224618 475226 224854
rect 475462 224618 475546 224854
rect 475782 224618 475814 224854
rect 475194 224534 475814 224618
rect 475194 224298 475226 224534
rect 475462 224298 475546 224534
rect 475782 224298 475814 224534
rect 475194 188854 475814 224298
rect 475194 188618 475226 188854
rect 475462 188618 475546 188854
rect 475782 188618 475814 188854
rect 475194 188534 475814 188618
rect 475194 188298 475226 188534
rect 475462 188298 475546 188534
rect 475782 188298 475814 188534
rect 475194 152854 475814 188298
rect 475194 152618 475226 152854
rect 475462 152618 475546 152854
rect 475782 152618 475814 152854
rect 475194 152534 475814 152618
rect 475194 152298 475226 152534
rect 475462 152298 475546 152534
rect 475782 152298 475814 152534
rect 475194 116854 475814 152298
rect 475194 116618 475226 116854
rect 475462 116618 475546 116854
rect 475782 116618 475814 116854
rect 475194 116534 475814 116618
rect 475194 116298 475226 116534
rect 475462 116298 475546 116534
rect 475782 116298 475814 116534
rect 475194 80854 475814 116298
rect 475194 80618 475226 80854
rect 475462 80618 475546 80854
rect 475782 80618 475814 80854
rect 475194 80534 475814 80618
rect 475194 80298 475226 80534
rect 475462 80298 475546 80534
rect 475782 80298 475814 80534
rect 475194 44854 475814 80298
rect 475194 44618 475226 44854
rect 475462 44618 475546 44854
rect 475782 44618 475814 44854
rect 475194 44534 475814 44618
rect 475194 44298 475226 44534
rect 475462 44298 475546 44534
rect 475782 44298 475814 44534
rect 475194 8854 475814 44298
rect 475194 8618 475226 8854
rect 475462 8618 475546 8854
rect 475782 8618 475814 8854
rect 475194 8534 475814 8618
rect 475194 8298 475226 8534
rect 475462 8298 475546 8534
rect 475782 8298 475814 8534
rect 475194 -5146 475814 8298
rect 475194 -5382 475226 -5146
rect 475462 -5382 475546 -5146
rect 475782 -5382 475814 -5146
rect 475194 -5466 475814 -5382
rect 475194 -5702 475226 -5466
rect 475462 -5702 475546 -5466
rect 475782 -5702 475814 -5466
rect 475194 -7654 475814 -5702
rect 476434 262094 477054 263615
rect 476434 261858 476466 262094
rect 476702 261858 476786 262094
rect 477022 261858 477054 262094
rect 476434 261774 477054 261858
rect 476434 261538 476466 261774
rect 476702 261538 476786 261774
rect 477022 261538 477054 261774
rect 476434 226094 477054 261538
rect 476434 225858 476466 226094
rect 476702 225858 476786 226094
rect 477022 225858 477054 226094
rect 476434 225774 477054 225858
rect 476434 225538 476466 225774
rect 476702 225538 476786 225774
rect 477022 225538 477054 225774
rect 476434 190094 477054 225538
rect 476434 189858 476466 190094
rect 476702 189858 476786 190094
rect 477022 189858 477054 190094
rect 476434 189774 477054 189858
rect 476434 189538 476466 189774
rect 476702 189538 476786 189774
rect 477022 189538 477054 189774
rect 476434 154094 477054 189538
rect 476434 153858 476466 154094
rect 476702 153858 476786 154094
rect 477022 153858 477054 154094
rect 476434 153774 477054 153858
rect 476434 153538 476466 153774
rect 476702 153538 476786 153774
rect 477022 153538 477054 153774
rect 476434 118094 477054 153538
rect 476434 117858 476466 118094
rect 476702 117858 476786 118094
rect 477022 117858 477054 118094
rect 476434 117774 477054 117858
rect 476434 117538 476466 117774
rect 476702 117538 476786 117774
rect 477022 117538 477054 117774
rect 476434 82094 477054 117538
rect 476434 81858 476466 82094
rect 476702 81858 476786 82094
rect 477022 81858 477054 82094
rect 476434 81774 477054 81858
rect 476434 81538 476466 81774
rect 476702 81538 476786 81774
rect 477022 81538 477054 81774
rect 476434 46094 477054 81538
rect 476434 45858 476466 46094
rect 476702 45858 476786 46094
rect 477022 45858 477054 46094
rect 476434 45774 477054 45858
rect 476434 45538 476466 45774
rect 476702 45538 476786 45774
rect 477022 45538 477054 45774
rect 476434 10094 477054 45538
rect 476434 9858 476466 10094
rect 476702 9858 476786 10094
rect 477022 9858 477054 10094
rect 476434 9774 477054 9858
rect 476434 9538 476466 9774
rect 476702 9538 476786 9774
rect 477022 9538 477054 9774
rect 476434 -6106 477054 9538
rect 477358 6629 477418 264963
rect 477674 263334 478294 263615
rect 477674 263098 477706 263334
rect 477942 263098 478026 263334
rect 478262 263098 478294 263334
rect 477674 263014 478294 263098
rect 477674 262778 477706 263014
rect 477942 262778 478026 263014
rect 478262 262778 478294 263014
rect 477674 227334 478294 262778
rect 477674 227098 477706 227334
rect 477942 227098 478026 227334
rect 478262 227098 478294 227334
rect 477674 227014 478294 227098
rect 477674 226778 477706 227014
rect 477942 226778 478026 227014
rect 478262 226778 478294 227014
rect 477674 191334 478294 226778
rect 477674 191098 477706 191334
rect 477942 191098 478026 191334
rect 478262 191098 478294 191334
rect 477674 191014 478294 191098
rect 477674 190778 477706 191014
rect 477942 190778 478026 191014
rect 478262 190778 478294 191014
rect 477674 155334 478294 190778
rect 477674 155098 477706 155334
rect 477942 155098 478026 155334
rect 478262 155098 478294 155334
rect 477674 155014 478294 155098
rect 477674 154778 477706 155014
rect 477942 154778 478026 155014
rect 478262 154778 478294 155014
rect 477674 119334 478294 154778
rect 477674 119098 477706 119334
rect 477942 119098 478026 119334
rect 478262 119098 478294 119334
rect 477674 119014 478294 119098
rect 477674 118778 477706 119014
rect 477942 118778 478026 119014
rect 478262 118778 478294 119014
rect 477674 83334 478294 118778
rect 477674 83098 477706 83334
rect 477942 83098 478026 83334
rect 478262 83098 478294 83334
rect 477674 83014 478294 83098
rect 477674 82778 477706 83014
rect 477942 82778 478026 83014
rect 478262 82778 478294 83014
rect 477674 47334 478294 82778
rect 477674 47098 477706 47334
rect 477942 47098 478026 47334
rect 478262 47098 478294 47334
rect 477674 47014 478294 47098
rect 477674 46778 477706 47014
rect 477942 46778 478026 47014
rect 478262 46778 478294 47014
rect 477674 11334 478294 46778
rect 480118 46341 480178 264963
rect 482878 86189 482938 264963
rect 486374 126037 486434 264963
rect 489134 165885 489194 265507
rect 504994 254654 505614 290098
rect 504994 254418 505026 254654
rect 505262 254418 505346 254654
rect 505582 254418 505614 254654
rect 504994 254334 505614 254418
rect 504994 254098 505026 254334
rect 505262 254098 505346 254334
rect 505582 254098 505614 254334
rect 504994 218654 505614 254098
rect 504994 218418 505026 218654
rect 505262 218418 505346 218654
rect 505582 218418 505614 218654
rect 504994 218334 505614 218418
rect 504994 218098 505026 218334
rect 505262 218098 505346 218334
rect 505582 218098 505614 218334
rect 504994 182654 505614 218098
rect 504994 182418 505026 182654
rect 505262 182418 505346 182654
rect 505582 182418 505614 182654
rect 504994 182334 505614 182418
rect 504994 182098 505026 182334
rect 505262 182098 505346 182334
rect 505582 182098 505614 182334
rect 489131 165884 489197 165885
rect 489131 165820 489132 165884
rect 489196 165820 489197 165884
rect 489131 165819 489197 165820
rect 504994 146654 505614 182098
rect 504994 146418 505026 146654
rect 505262 146418 505346 146654
rect 505582 146418 505614 146654
rect 504994 146334 505614 146418
rect 504994 146098 505026 146334
rect 505262 146098 505346 146334
rect 505582 146098 505614 146334
rect 486371 126036 486437 126037
rect 486371 125972 486372 126036
rect 486436 125972 486437 126036
rect 486371 125971 486437 125972
rect 504994 110654 505614 146098
rect 504994 110418 505026 110654
rect 505262 110418 505346 110654
rect 505582 110418 505614 110654
rect 504994 110334 505614 110418
rect 504994 110098 505026 110334
rect 505262 110098 505346 110334
rect 505582 110098 505614 110334
rect 482875 86188 482941 86189
rect 482875 86124 482876 86188
rect 482940 86124 482941 86188
rect 482875 86123 482941 86124
rect 504994 74654 505614 110098
rect 504994 74418 505026 74654
rect 505262 74418 505346 74654
rect 505582 74418 505614 74654
rect 504994 74334 505614 74418
rect 504994 74098 505026 74334
rect 505262 74098 505346 74334
rect 505582 74098 505614 74334
rect 480115 46340 480181 46341
rect 480115 46276 480116 46340
rect 480180 46276 480181 46340
rect 480115 46275 480181 46276
rect 477674 11098 477706 11334
rect 477942 11098 478026 11334
rect 478262 11098 478294 11334
rect 477674 11014 478294 11098
rect 477674 10778 477706 11014
rect 477942 10778 478026 11014
rect 478262 10778 478294 11014
rect 477355 6628 477421 6629
rect 477355 6564 477356 6628
rect 477420 6564 477421 6628
rect 477355 6563 477421 6564
rect 476434 -6342 476466 -6106
rect 476702 -6342 476786 -6106
rect 477022 -6342 477054 -6106
rect 476434 -6426 477054 -6342
rect 476434 -6662 476466 -6426
rect 476702 -6662 476786 -6426
rect 477022 -6662 477054 -6426
rect 476434 -7654 477054 -6662
rect 477674 -7066 478294 10778
rect 477674 -7302 477706 -7066
rect 477942 -7302 478026 -7066
rect 478262 -7302 478294 -7066
rect 477674 -7386 478294 -7302
rect 477674 -7622 477706 -7386
rect 477942 -7622 478026 -7386
rect 478262 -7622 478294 -7386
rect 477674 -7654 478294 -7622
rect 504994 38654 505614 74098
rect 504994 38418 505026 38654
rect 505262 38418 505346 38654
rect 505582 38418 505614 38654
rect 504994 38334 505614 38418
rect 504994 38098 505026 38334
rect 505262 38098 505346 38334
rect 505582 38098 505614 38334
rect 504994 2654 505614 38098
rect 504994 2418 505026 2654
rect 505262 2418 505346 2654
rect 505582 2418 505614 2654
rect 504994 2334 505614 2418
rect 504994 2098 505026 2334
rect 505262 2098 505346 2334
rect 505582 2098 505614 2334
rect 504994 -346 505614 2098
rect 504994 -582 505026 -346
rect 505262 -582 505346 -346
rect 505582 -582 505614 -346
rect 504994 -666 505614 -582
rect 504994 -902 505026 -666
rect 505262 -902 505346 -666
rect 505582 -902 505614 -666
rect 504994 -7654 505614 -902
rect 506234 705798 506854 711590
rect 506234 705562 506266 705798
rect 506502 705562 506586 705798
rect 506822 705562 506854 705798
rect 506234 705478 506854 705562
rect 506234 705242 506266 705478
rect 506502 705242 506586 705478
rect 506822 705242 506854 705478
rect 506234 687894 506854 705242
rect 506234 687658 506266 687894
rect 506502 687658 506586 687894
rect 506822 687658 506854 687894
rect 506234 687574 506854 687658
rect 506234 687338 506266 687574
rect 506502 687338 506586 687574
rect 506822 687338 506854 687574
rect 506234 651894 506854 687338
rect 506234 651658 506266 651894
rect 506502 651658 506586 651894
rect 506822 651658 506854 651894
rect 506234 651574 506854 651658
rect 506234 651338 506266 651574
rect 506502 651338 506586 651574
rect 506822 651338 506854 651574
rect 506234 615894 506854 651338
rect 506234 615658 506266 615894
rect 506502 615658 506586 615894
rect 506822 615658 506854 615894
rect 506234 615574 506854 615658
rect 506234 615338 506266 615574
rect 506502 615338 506586 615574
rect 506822 615338 506854 615574
rect 506234 579894 506854 615338
rect 506234 579658 506266 579894
rect 506502 579658 506586 579894
rect 506822 579658 506854 579894
rect 506234 579574 506854 579658
rect 506234 579338 506266 579574
rect 506502 579338 506586 579574
rect 506822 579338 506854 579574
rect 506234 543894 506854 579338
rect 506234 543658 506266 543894
rect 506502 543658 506586 543894
rect 506822 543658 506854 543894
rect 506234 543574 506854 543658
rect 506234 543338 506266 543574
rect 506502 543338 506586 543574
rect 506822 543338 506854 543574
rect 506234 507894 506854 543338
rect 506234 507658 506266 507894
rect 506502 507658 506586 507894
rect 506822 507658 506854 507894
rect 506234 507574 506854 507658
rect 506234 507338 506266 507574
rect 506502 507338 506586 507574
rect 506822 507338 506854 507574
rect 506234 471894 506854 507338
rect 506234 471658 506266 471894
rect 506502 471658 506586 471894
rect 506822 471658 506854 471894
rect 506234 471574 506854 471658
rect 506234 471338 506266 471574
rect 506502 471338 506586 471574
rect 506822 471338 506854 471574
rect 506234 435894 506854 471338
rect 506234 435658 506266 435894
rect 506502 435658 506586 435894
rect 506822 435658 506854 435894
rect 506234 435574 506854 435658
rect 506234 435338 506266 435574
rect 506502 435338 506586 435574
rect 506822 435338 506854 435574
rect 506234 399894 506854 435338
rect 506234 399658 506266 399894
rect 506502 399658 506586 399894
rect 506822 399658 506854 399894
rect 506234 399574 506854 399658
rect 506234 399338 506266 399574
rect 506502 399338 506586 399574
rect 506822 399338 506854 399574
rect 506234 363894 506854 399338
rect 506234 363658 506266 363894
rect 506502 363658 506586 363894
rect 506822 363658 506854 363894
rect 506234 363574 506854 363658
rect 506234 363338 506266 363574
rect 506502 363338 506586 363574
rect 506822 363338 506854 363574
rect 506234 327894 506854 363338
rect 506234 327658 506266 327894
rect 506502 327658 506586 327894
rect 506822 327658 506854 327894
rect 506234 327574 506854 327658
rect 506234 327338 506266 327574
rect 506502 327338 506586 327574
rect 506822 327338 506854 327574
rect 506234 291894 506854 327338
rect 506234 291658 506266 291894
rect 506502 291658 506586 291894
rect 506822 291658 506854 291894
rect 506234 291574 506854 291658
rect 506234 291338 506266 291574
rect 506502 291338 506586 291574
rect 506822 291338 506854 291574
rect 506234 255894 506854 291338
rect 506234 255658 506266 255894
rect 506502 255658 506586 255894
rect 506822 255658 506854 255894
rect 506234 255574 506854 255658
rect 506234 255338 506266 255574
rect 506502 255338 506586 255574
rect 506822 255338 506854 255574
rect 506234 219894 506854 255338
rect 506234 219658 506266 219894
rect 506502 219658 506586 219894
rect 506822 219658 506854 219894
rect 506234 219574 506854 219658
rect 506234 219338 506266 219574
rect 506502 219338 506586 219574
rect 506822 219338 506854 219574
rect 506234 183894 506854 219338
rect 506234 183658 506266 183894
rect 506502 183658 506586 183894
rect 506822 183658 506854 183894
rect 506234 183574 506854 183658
rect 506234 183338 506266 183574
rect 506502 183338 506586 183574
rect 506822 183338 506854 183574
rect 506234 147894 506854 183338
rect 506234 147658 506266 147894
rect 506502 147658 506586 147894
rect 506822 147658 506854 147894
rect 506234 147574 506854 147658
rect 506234 147338 506266 147574
rect 506502 147338 506586 147574
rect 506822 147338 506854 147574
rect 506234 111894 506854 147338
rect 506234 111658 506266 111894
rect 506502 111658 506586 111894
rect 506822 111658 506854 111894
rect 506234 111574 506854 111658
rect 506234 111338 506266 111574
rect 506502 111338 506586 111574
rect 506822 111338 506854 111574
rect 506234 75894 506854 111338
rect 506234 75658 506266 75894
rect 506502 75658 506586 75894
rect 506822 75658 506854 75894
rect 506234 75574 506854 75658
rect 506234 75338 506266 75574
rect 506502 75338 506586 75574
rect 506822 75338 506854 75574
rect 506234 39894 506854 75338
rect 506234 39658 506266 39894
rect 506502 39658 506586 39894
rect 506822 39658 506854 39894
rect 506234 39574 506854 39658
rect 506234 39338 506266 39574
rect 506502 39338 506586 39574
rect 506822 39338 506854 39574
rect 506234 3894 506854 39338
rect 506234 3658 506266 3894
rect 506502 3658 506586 3894
rect 506822 3658 506854 3894
rect 506234 3574 506854 3658
rect 506234 3338 506266 3574
rect 506502 3338 506586 3574
rect 506822 3338 506854 3574
rect 506234 -1306 506854 3338
rect 506234 -1542 506266 -1306
rect 506502 -1542 506586 -1306
rect 506822 -1542 506854 -1306
rect 506234 -1626 506854 -1542
rect 506234 -1862 506266 -1626
rect 506502 -1862 506586 -1626
rect 506822 -1862 506854 -1626
rect 506234 -7654 506854 -1862
rect 507474 706758 508094 711590
rect 507474 706522 507506 706758
rect 507742 706522 507826 706758
rect 508062 706522 508094 706758
rect 507474 706438 508094 706522
rect 507474 706202 507506 706438
rect 507742 706202 507826 706438
rect 508062 706202 508094 706438
rect 507474 689134 508094 706202
rect 507474 688898 507506 689134
rect 507742 688898 507826 689134
rect 508062 688898 508094 689134
rect 507474 688814 508094 688898
rect 507474 688578 507506 688814
rect 507742 688578 507826 688814
rect 508062 688578 508094 688814
rect 507474 653134 508094 688578
rect 507474 652898 507506 653134
rect 507742 652898 507826 653134
rect 508062 652898 508094 653134
rect 507474 652814 508094 652898
rect 507474 652578 507506 652814
rect 507742 652578 507826 652814
rect 508062 652578 508094 652814
rect 507474 617134 508094 652578
rect 507474 616898 507506 617134
rect 507742 616898 507826 617134
rect 508062 616898 508094 617134
rect 507474 616814 508094 616898
rect 507474 616578 507506 616814
rect 507742 616578 507826 616814
rect 508062 616578 508094 616814
rect 507474 581134 508094 616578
rect 507474 580898 507506 581134
rect 507742 580898 507826 581134
rect 508062 580898 508094 581134
rect 507474 580814 508094 580898
rect 507474 580578 507506 580814
rect 507742 580578 507826 580814
rect 508062 580578 508094 580814
rect 507474 545134 508094 580578
rect 507474 544898 507506 545134
rect 507742 544898 507826 545134
rect 508062 544898 508094 545134
rect 507474 544814 508094 544898
rect 507474 544578 507506 544814
rect 507742 544578 507826 544814
rect 508062 544578 508094 544814
rect 507474 509134 508094 544578
rect 507474 508898 507506 509134
rect 507742 508898 507826 509134
rect 508062 508898 508094 509134
rect 507474 508814 508094 508898
rect 507474 508578 507506 508814
rect 507742 508578 507826 508814
rect 508062 508578 508094 508814
rect 507474 473134 508094 508578
rect 507474 472898 507506 473134
rect 507742 472898 507826 473134
rect 508062 472898 508094 473134
rect 507474 472814 508094 472898
rect 507474 472578 507506 472814
rect 507742 472578 507826 472814
rect 508062 472578 508094 472814
rect 507474 437134 508094 472578
rect 507474 436898 507506 437134
rect 507742 436898 507826 437134
rect 508062 436898 508094 437134
rect 507474 436814 508094 436898
rect 507474 436578 507506 436814
rect 507742 436578 507826 436814
rect 508062 436578 508094 436814
rect 507474 401134 508094 436578
rect 507474 400898 507506 401134
rect 507742 400898 507826 401134
rect 508062 400898 508094 401134
rect 507474 400814 508094 400898
rect 507474 400578 507506 400814
rect 507742 400578 507826 400814
rect 508062 400578 508094 400814
rect 507474 365134 508094 400578
rect 507474 364898 507506 365134
rect 507742 364898 507826 365134
rect 508062 364898 508094 365134
rect 507474 364814 508094 364898
rect 507474 364578 507506 364814
rect 507742 364578 507826 364814
rect 508062 364578 508094 364814
rect 507474 329134 508094 364578
rect 507474 328898 507506 329134
rect 507742 328898 507826 329134
rect 508062 328898 508094 329134
rect 507474 328814 508094 328898
rect 507474 328578 507506 328814
rect 507742 328578 507826 328814
rect 508062 328578 508094 328814
rect 507474 293134 508094 328578
rect 507474 292898 507506 293134
rect 507742 292898 507826 293134
rect 508062 292898 508094 293134
rect 507474 292814 508094 292898
rect 507474 292578 507506 292814
rect 507742 292578 507826 292814
rect 508062 292578 508094 292814
rect 507474 257134 508094 292578
rect 507474 256898 507506 257134
rect 507742 256898 507826 257134
rect 508062 256898 508094 257134
rect 507474 256814 508094 256898
rect 507474 256578 507506 256814
rect 507742 256578 507826 256814
rect 508062 256578 508094 256814
rect 507474 221134 508094 256578
rect 507474 220898 507506 221134
rect 507742 220898 507826 221134
rect 508062 220898 508094 221134
rect 507474 220814 508094 220898
rect 507474 220578 507506 220814
rect 507742 220578 507826 220814
rect 508062 220578 508094 220814
rect 507474 185134 508094 220578
rect 507474 184898 507506 185134
rect 507742 184898 507826 185134
rect 508062 184898 508094 185134
rect 507474 184814 508094 184898
rect 507474 184578 507506 184814
rect 507742 184578 507826 184814
rect 508062 184578 508094 184814
rect 507474 149134 508094 184578
rect 507474 148898 507506 149134
rect 507742 148898 507826 149134
rect 508062 148898 508094 149134
rect 507474 148814 508094 148898
rect 507474 148578 507506 148814
rect 507742 148578 507826 148814
rect 508062 148578 508094 148814
rect 507474 113134 508094 148578
rect 507474 112898 507506 113134
rect 507742 112898 507826 113134
rect 508062 112898 508094 113134
rect 507474 112814 508094 112898
rect 507474 112578 507506 112814
rect 507742 112578 507826 112814
rect 508062 112578 508094 112814
rect 507474 77134 508094 112578
rect 507474 76898 507506 77134
rect 507742 76898 507826 77134
rect 508062 76898 508094 77134
rect 507474 76814 508094 76898
rect 507474 76578 507506 76814
rect 507742 76578 507826 76814
rect 508062 76578 508094 76814
rect 507474 41134 508094 76578
rect 507474 40898 507506 41134
rect 507742 40898 507826 41134
rect 508062 40898 508094 41134
rect 507474 40814 508094 40898
rect 507474 40578 507506 40814
rect 507742 40578 507826 40814
rect 508062 40578 508094 40814
rect 507474 5134 508094 40578
rect 507474 4898 507506 5134
rect 507742 4898 507826 5134
rect 508062 4898 508094 5134
rect 507474 4814 508094 4898
rect 507474 4578 507506 4814
rect 507742 4578 507826 4814
rect 508062 4578 508094 4814
rect 507474 -2266 508094 4578
rect 507474 -2502 507506 -2266
rect 507742 -2502 507826 -2266
rect 508062 -2502 508094 -2266
rect 507474 -2586 508094 -2502
rect 507474 -2822 507506 -2586
rect 507742 -2822 507826 -2586
rect 508062 -2822 508094 -2586
rect 507474 -7654 508094 -2822
rect 508714 707718 509334 711590
rect 508714 707482 508746 707718
rect 508982 707482 509066 707718
rect 509302 707482 509334 707718
rect 508714 707398 509334 707482
rect 508714 707162 508746 707398
rect 508982 707162 509066 707398
rect 509302 707162 509334 707398
rect 508714 690374 509334 707162
rect 508714 690138 508746 690374
rect 508982 690138 509066 690374
rect 509302 690138 509334 690374
rect 508714 690054 509334 690138
rect 508714 689818 508746 690054
rect 508982 689818 509066 690054
rect 509302 689818 509334 690054
rect 508714 654374 509334 689818
rect 508714 654138 508746 654374
rect 508982 654138 509066 654374
rect 509302 654138 509334 654374
rect 508714 654054 509334 654138
rect 508714 653818 508746 654054
rect 508982 653818 509066 654054
rect 509302 653818 509334 654054
rect 508714 618374 509334 653818
rect 508714 618138 508746 618374
rect 508982 618138 509066 618374
rect 509302 618138 509334 618374
rect 508714 618054 509334 618138
rect 508714 617818 508746 618054
rect 508982 617818 509066 618054
rect 509302 617818 509334 618054
rect 508714 582374 509334 617818
rect 508714 582138 508746 582374
rect 508982 582138 509066 582374
rect 509302 582138 509334 582374
rect 508714 582054 509334 582138
rect 508714 581818 508746 582054
rect 508982 581818 509066 582054
rect 509302 581818 509334 582054
rect 508714 546374 509334 581818
rect 508714 546138 508746 546374
rect 508982 546138 509066 546374
rect 509302 546138 509334 546374
rect 508714 546054 509334 546138
rect 508714 545818 508746 546054
rect 508982 545818 509066 546054
rect 509302 545818 509334 546054
rect 508714 510374 509334 545818
rect 508714 510138 508746 510374
rect 508982 510138 509066 510374
rect 509302 510138 509334 510374
rect 508714 510054 509334 510138
rect 508714 509818 508746 510054
rect 508982 509818 509066 510054
rect 509302 509818 509334 510054
rect 508714 474374 509334 509818
rect 508714 474138 508746 474374
rect 508982 474138 509066 474374
rect 509302 474138 509334 474374
rect 508714 474054 509334 474138
rect 508714 473818 508746 474054
rect 508982 473818 509066 474054
rect 509302 473818 509334 474054
rect 508714 438374 509334 473818
rect 508714 438138 508746 438374
rect 508982 438138 509066 438374
rect 509302 438138 509334 438374
rect 508714 438054 509334 438138
rect 508714 437818 508746 438054
rect 508982 437818 509066 438054
rect 509302 437818 509334 438054
rect 508714 402374 509334 437818
rect 508714 402138 508746 402374
rect 508982 402138 509066 402374
rect 509302 402138 509334 402374
rect 508714 402054 509334 402138
rect 508714 401818 508746 402054
rect 508982 401818 509066 402054
rect 509302 401818 509334 402054
rect 508714 366374 509334 401818
rect 508714 366138 508746 366374
rect 508982 366138 509066 366374
rect 509302 366138 509334 366374
rect 508714 366054 509334 366138
rect 508714 365818 508746 366054
rect 508982 365818 509066 366054
rect 509302 365818 509334 366054
rect 508714 330374 509334 365818
rect 508714 330138 508746 330374
rect 508982 330138 509066 330374
rect 509302 330138 509334 330374
rect 508714 330054 509334 330138
rect 508714 329818 508746 330054
rect 508982 329818 509066 330054
rect 509302 329818 509334 330054
rect 508714 294374 509334 329818
rect 508714 294138 508746 294374
rect 508982 294138 509066 294374
rect 509302 294138 509334 294374
rect 508714 294054 509334 294138
rect 508714 293818 508746 294054
rect 508982 293818 509066 294054
rect 509302 293818 509334 294054
rect 508714 258374 509334 293818
rect 508714 258138 508746 258374
rect 508982 258138 509066 258374
rect 509302 258138 509334 258374
rect 508714 258054 509334 258138
rect 508714 257818 508746 258054
rect 508982 257818 509066 258054
rect 509302 257818 509334 258054
rect 508714 222374 509334 257818
rect 508714 222138 508746 222374
rect 508982 222138 509066 222374
rect 509302 222138 509334 222374
rect 508714 222054 509334 222138
rect 508714 221818 508746 222054
rect 508982 221818 509066 222054
rect 509302 221818 509334 222054
rect 508714 186374 509334 221818
rect 508714 186138 508746 186374
rect 508982 186138 509066 186374
rect 509302 186138 509334 186374
rect 508714 186054 509334 186138
rect 508714 185818 508746 186054
rect 508982 185818 509066 186054
rect 509302 185818 509334 186054
rect 508714 150374 509334 185818
rect 508714 150138 508746 150374
rect 508982 150138 509066 150374
rect 509302 150138 509334 150374
rect 508714 150054 509334 150138
rect 508714 149818 508746 150054
rect 508982 149818 509066 150054
rect 509302 149818 509334 150054
rect 508714 114374 509334 149818
rect 508714 114138 508746 114374
rect 508982 114138 509066 114374
rect 509302 114138 509334 114374
rect 508714 114054 509334 114138
rect 508714 113818 508746 114054
rect 508982 113818 509066 114054
rect 509302 113818 509334 114054
rect 508714 78374 509334 113818
rect 508714 78138 508746 78374
rect 508982 78138 509066 78374
rect 509302 78138 509334 78374
rect 508714 78054 509334 78138
rect 508714 77818 508746 78054
rect 508982 77818 509066 78054
rect 509302 77818 509334 78054
rect 508714 42374 509334 77818
rect 508714 42138 508746 42374
rect 508982 42138 509066 42374
rect 509302 42138 509334 42374
rect 508714 42054 509334 42138
rect 508714 41818 508746 42054
rect 508982 41818 509066 42054
rect 509302 41818 509334 42054
rect 508714 6374 509334 41818
rect 508714 6138 508746 6374
rect 508982 6138 509066 6374
rect 509302 6138 509334 6374
rect 508714 6054 509334 6138
rect 508714 5818 508746 6054
rect 508982 5818 509066 6054
rect 509302 5818 509334 6054
rect 508714 -3226 509334 5818
rect 508714 -3462 508746 -3226
rect 508982 -3462 509066 -3226
rect 509302 -3462 509334 -3226
rect 508714 -3546 509334 -3462
rect 508714 -3782 508746 -3546
rect 508982 -3782 509066 -3546
rect 509302 -3782 509334 -3546
rect 508714 -7654 509334 -3782
rect 509954 708678 510574 711590
rect 509954 708442 509986 708678
rect 510222 708442 510306 708678
rect 510542 708442 510574 708678
rect 509954 708358 510574 708442
rect 509954 708122 509986 708358
rect 510222 708122 510306 708358
rect 510542 708122 510574 708358
rect 509954 691614 510574 708122
rect 509954 691378 509986 691614
rect 510222 691378 510306 691614
rect 510542 691378 510574 691614
rect 509954 691294 510574 691378
rect 509954 691058 509986 691294
rect 510222 691058 510306 691294
rect 510542 691058 510574 691294
rect 509954 655614 510574 691058
rect 509954 655378 509986 655614
rect 510222 655378 510306 655614
rect 510542 655378 510574 655614
rect 509954 655294 510574 655378
rect 509954 655058 509986 655294
rect 510222 655058 510306 655294
rect 510542 655058 510574 655294
rect 509954 619614 510574 655058
rect 509954 619378 509986 619614
rect 510222 619378 510306 619614
rect 510542 619378 510574 619614
rect 509954 619294 510574 619378
rect 509954 619058 509986 619294
rect 510222 619058 510306 619294
rect 510542 619058 510574 619294
rect 509954 583614 510574 619058
rect 509954 583378 509986 583614
rect 510222 583378 510306 583614
rect 510542 583378 510574 583614
rect 509954 583294 510574 583378
rect 509954 583058 509986 583294
rect 510222 583058 510306 583294
rect 510542 583058 510574 583294
rect 509954 547614 510574 583058
rect 509954 547378 509986 547614
rect 510222 547378 510306 547614
rect 510542 547378 510574 547614
rect 509954 547294 510574 547378
rect 509954 547058 509986 547294
rect 510222 547058 510306 547294
rect 510542 547058 510574 547294
rect 509954 511614 510574 547058
rect 509954 511378 509986 511614
rect 510222 511378 510306 511614
rect 510542 511378 510574 511614
rect 509954 511294 510574 511378
rect 509954 511058 509986 511294
rect 510222 511058 510306 511294
rect 510542 511058 510574 511294
rect 509954 475614 510574 511058
rect 509954 475378 509986 475614
rect 510222 475378 510306 475614
rect 510542 475378 510574 475614
rect 509954 475294 510574 475378
rect 509954 475058 509986 475294
rect 510222 475058 510306 475294
rect 510542 475058 510574 475294
rect 509954 439614 510574 475058
rect 509954 439378 509986 439614
rect 510222 439378 510306 439614
rect 510542 439378 510574 439614
rect 509954 439294 510574 439378
rect 509954 439058 509986 439294
rect 510222 439058 510306 439294
rect 510542 439058 510574 439294
rect 509954 403614 510574 439058
rect 509954 403378 509986 403614
rect 510222 403378 510306 403614
rect 510542 403378 510574 403614
rect 509954 403294 510574 403378
rect 509954 403058 509986 403294
rect 510222 403058 510306 403294
rect 510542 403058 510574 403294
rect 509954 367614 510574 403058
rect 509954 367378 509986 367614
rect 510222 367378 510306 367614
rect 510542 367378 510574 367614
rect 509954 367294 510574 367378
rect 509954 367058 509986 367294
rect 510222 367058 510306 367294
rect 510542 367058 510574 367294
rect 509954 331614 510574 367058
rect 509954 331378 509986 331614
rect 510222 331378 510306 331614
rect 510542 331378 510574 331614
rect 509954 331294 510574 331378
rect 509954 331058 509986 331294
rect 510222 331058 510306 331294
rect 510542 331058 510574 331294
rect 509954 295614 510574 331058
rect 509954 295378 509986 295614
rect 510222 295378 510306 295614
rect 510542 295378 510574 295614
rect 509954 295294 510574 295378
rect 509954 295058 509986 295294
rect 510222 295058 510306 295294
rect 510542 295058 510574 295294
rect 509954 259614 510574 295058
rect 509954 259378 509986 259614
rect 510222 259378 510306 259614
rect 510542 259378 510574 259614
rect 509954 259294 510574 259378
rect 509954 259058 509986 259294
rect 510222 259058 510306 259294
rect 510542 259058 510574 259294
rect 509954 223614 510574 259058
rect 509954 223378 509986 223614
rect 510222 223378 510306 223614
rect 510542 223378 510574 223614
rect 509954 223294 510574 223378
rect 509954 223058 509986 223294
rect 510222 223058 510306 223294
rect 510542 223058 510574 223294
rect 509954 187614 510574 223058
rect 509954 187378 509986 187614
rect 510222 187378 510306 187614
rect 510542 187378 510574 187614
rect 509954 187294 510574 187378
rect 509954 187058 509986 187294
rect 510222 187058 510306 187294
rect 510542 187058 510574 187294
rect 509954 151614 510574 187058
rect 509954 151378 509986 151614
rect 510222 151378 510306 151614
rect 510542 151378 510574 151614
rect 509954 151294 510574 151378
rect 509954 151058 509986 151294
rect 510222 151058 510306 151294
rect 510542 151058 510574 151294
rect 509954 115614 510574 151058
rect 509954 115378 509986 115614
rect 510222 115378 510306 115614
rect 510542 115378 510574 115614
rect 509954 115294 510574 115378
rect 509954 115058 509986 115294
rect 510222 115058 510306 115294
rect 510542 115058 510574 115294
rect 509954 79614 510574 115058
rect 509954 79378 509986 79614
rect 510222 79378 510306 79614
rect 510542 79378 510574 79614
rect 509954 79294 510574 79378
rect 509954 79058 509986 79294
rect 510222 79058 510306 79294
rect 510542 79058 510574 79294
rect 509954 43614 510574 79058
rect 509954 43378 509986 43614
rect 510222 43378 510306 43614
rect 510542 43378 510574 43614
rect 509954 43294 510574 43378
rect 509954 43058 509986 43294
rect 510222 43058 510306 43294
rect 510542 43058 510574 43294
rect 509954 7614 510574 43058
rect 509954 7378 509986 7614
rect 510222 7378 510306 7614
rect 510542 7378 510574 7614
rect 509954 7294 510574 7378
rect 509954 7058 509986 7294
rect 510222 7058 510306 7294
rect 510542 7058 510574 7294
rect 509954 -4186 510574 7058
rect 509954 -4422 509986 -4186
rect 510222 -4422 510306 -4186
rect 510542 -4422 510574 -4186
rect 509954 -4506 510574 -4422
rect 509954 -4742 509986 -4506
rect 510222 -4742 510306 -4506
rect 510542 -4742 510574 -4506
rect 509954 -7654 510574 -4742
rect 511194 709638 511814 711590
rect 511194 709402 511226 709638
rect 511462 709402 511546 709638
rect 511782 709402 511814 709638
rect 511194 709318 511814 709402
rect 511194 709082 511226 709318
rect 511462 709082 511546 709318
rect 511782 709082 511814 709318
rect 511194 692854 511814 709082
rect 511194 692618 511226 692854
rect 511462 692618 511546 692854
rect 511782 692618 511814 692854
rect 511194 692534 511814 692618
rect 511194 692298 511226 692534
rect 511462 692298 511546 692534
rect 511782 692298 511814 692534
rect 511194 656854 511814 692298
rect 511194 656618 511226 656854
rect 511462 656618 511546 656854
rect 511782 656618 511814 656854
rect 511194 656534 511814 656618
rect 511194 656298 511226 656534
rect 511462 656298 511546 656534
rect 511782 656298 511814 656534
rect 511194 620854 511814 656298
rect 511194 620618 511226 620854
rect 511462 620618 511546 620854
rect 511782 620618 511814 620854
rect 511194 620534 511814 620618
rect 511194 620298 511226 620534
rect 511462 620298 511546 620534
rect 511782 620298 511814 620534
rect 511194 584854 511814 620298
rect 511194 584618 511226 584854
rect 511462 584618 511546 584854
rect 511782 584618 511814 584854
rect 511194 584534 511814 584618
rect 511194 584298 511226 584534
rect 511462 584298 511546 584534
rect 511782 584298 511814 584534
rect 511194 548854 511814 584298
rect 511194 548618 511226 548854
rect 511462 548618 511546 548854
rect 511782 548618 511814 548854
rect 511194 548534 511814 548618
rect 511194 548298 511226 548534
rect 511462 548298 511546 548534
rect 511782 548298 511814 548534
rect 511194 512854 511814 548298
rect 511194 512618 511226 512854
rect 511462 512618 511546 512854
rect 511782 512618 511814 512854
rect 511194 512534 511814 512618
rect 511194 512298 511226 512534
rect 511462 512298 511546 512534
rect 511782 512298 511814 512534
rect 511194 476854 511814 512298
rect 511194 476618 511226 476854
rect 511462 476618 511546 476854
rect 511782 476618 511814 476854
rect 511194 476534 511814 476618
rect 511194 476298 511226 476534
rect 511462 476298 511546 476534
rect 511782 476298 511814 476534
rect 511194 440854 511814 476298
rect 511194 440618 511226 440854
rect 511462 440618 511546 440854
rect 511782 440618 511814 440854
rect 511194 440534 511814 440618
rect 511194 440298 511226 440534
rect 511462 440298 511546 440534
rect 511782 440298 511814 440534
rect 511194 404854 511814 440298
rect 511194 404618 511226 404854
rect 511462 404618 511546 404854
rect 511782 404618 511814 404854
rect 511194 404534 511814 404618
rect 511194 404298 511226 404534
rect 511462 404298 511546 404534
rect 511782 404298 511814 404534
rect 511194 368854 511814 404298
rect 511194 368618 511226 368854
rect 511462 368618 511546 368854
rect 511782 368618 511814 368854
rect 511194 368534 511814 368618
rect 511194 368298 511226 368534
rect 511462 368298 511546 368534
rect 511782 368298 511814 368534
rect 511194 332854 511814 368298
rect 511194 332618 511226 332854
rect 511462 332618 511546 332854
rect 511782 332618 511814 332854
rect 511194 332534 511814 332618
rect 511194 332298 511226 332534
rect 511462 332298 511546 332534
rect 511782 332298 511814 332534
rect 511194 296854 511814 332298
rect 511194 296618 511226 296854
rect 511462 296618 511546 296854
rect 511782 296618 511814 296854
rect 511194 296534 511814 296618
rect 511194 296298 511226 296534
rect 511462 296298 511546 296534
rect 511782 296298 511814 296534
rect 511194 260854 511814 296298
rect 511194 260618 511226 260854
rect 511462 260618 511546 260854
rect 511782 260618 511814 260854
rect 511194 260534 511814 260618
rect 511194 260298 511226 260534
rect 511462 260298 511546 260534
rect 511782 260298 511814 260534
rect 511194 224854 511814 260298
rect 511194 224618 511226 224854
rect 511462 224618 511546 224854
rect 511782 224618 511814 224854
rect 511194 224534 511814 224618
rect 511194 224298 511226 224534
rect 511462 224298 511546 224534
rect 511782 224298 511814 224534
rect 511194 188854 511814 224298
rect 511194 188618 511226 188854
rect 511462 188618 511546 188854
rect 511782 188618 511814 188854
rect 511194 188534 511814 188618
rect 511194 188298 511226 188534
rect 511462 188298 511546 188534
rect 511782 188298 511814 188534
rect 511194 152854 511814 188298
rect 511194 152618 511226 152854
rect 511462 152618 511546 152854
rect 511782 152618 511814 152854
rect 511194 152534 511814 152618
rect 511194 152298 511226 152534
rect 511462 152298 511546 152534
rect 511782 152298 511814 152534
rect 511194 116854 511814 152298
rect 511194 116618 511226 116854
rect 511462 116618 511546 116854
rect 511782 116618 511814 116854
rect 511194 116534 511814 116618
rect 511194 116298 511226 116534
rect 511462 116298 511546 116534
rect 511782 116298 511814 116534
rect 511194 80854 511814 116298
rect 511194 80618 511226 80854
rect 511462 80618 511546 80854
rect 511782 80618 511814 80854
rect 511194 80534 511814 80618
rect 511194 80298 511226 80534
rect 511462 80298 511546 80534
rect 511782 80298 511814 80534
rect 511194 44854 511814 80298
rect 511194 44618 511226 44854
rect 511462 44618 511546 44854
rect 511782 44618 511814 44854
rect 511194 44534 511814 44618
rect 511194 44298 511226 44534
rect 511462 44298 511546 44534
rect 511782 44298 511814 44534
rect 511194 8854 511814 44298
rect 511194 8618 511226 8854
rect 511462 8618 511546 8854
rect 511782 8618 511814 8854
rect 511194 8534 511814 8618
rect 511194 8298 511226 8534
rect 511462 8298 511546 8534
rect 511782 8298 511814 8534
rect 511194 -5146 511814 8298
rect 511194 -5382 511226 -5146
rect 511462 -5382 511546 -5146
rect 511782 -5382 511814 -5146
rect 511194 -5466 511814 -5382
rect 511194 -5702 511226 -5466
rect 511462 -5702 511546 -5466
rect 511782 -5702 511814 -5466
rect 511194 -7654 511814 -5702
rect 512434 710598 513054 711590
rect 512434 710362 512466 710598
rect 512702 710362 512786 710598
rect 513022 710362 513054 710598
rect 512434 710278 513054 710362
rect 512434 710042 512466 710278
rect 512702 710042 512786 710278
rect 513022 710042 513054 710278
rect 512434 694094 513054 710042
rect 512434 693858 512466 694094
rect 512702 693858 512786 694094
rect 513022 693858 513054 694094
rect 512434 693774 513054 693858
rect 512434 693538 512466 693774
rect 512702 693538 512786 693774
rect 513022 693538 513054 693774
rect 512434 658094 513054 693538
rect 512434 657858 512466 658094
rect 512702 657858 512786 658094
rect 513022 657858 513054 658094
rect 512434 657774 513054 657858
rect 512434 657538 512466 657774
rect 512702 657538 512786 657774
rect 513022 657538 513054 657774
rect 512434 622094 513054 657538
rect 512434 621858 512466 622094
rect 512702 621858 512786 622094
rect 513022 621858 513054 622094
rect 512434 621774 513054 621858
rect 512434 621538 512466 621774
rect 512702 621538 512786 621774
rect 513022 621538 513054 621774
rect 512434 586094 513054 621538
rect 512434 585858 512466 586094
rect 512702 585858 512786 586094
rect 513022 585858 513054 586094
rect 512434 585774 513054 585858
rect 512434 585538 512466 585774
rect 512702 585538 512786 585774
rect 513022 585538 513054 585774
rect 512434 550094 513054 585538
rect 512434 549858 512466 550094
rect 512702 549858 512786 550094
rect 513022 549858 513054 550094
rect 512434 549774 513054 549858
rect 512434 549538 512466 549774
rect 512702 549538 512786 549774
rect 513022 549538 513054 549774
rect 512434 514094 513054 549538
rect 512434 513858 512466 514094
rect 512702 513858 512786 514094
rect 513022 513858 513054 514094
rect 512434 513774 513054 513858
rect 512434 513538 512466 513774
rect 512702 513538 512786 513774
rect 513022 513538 513054 513774
rect 512434 478094 513054 513538
rect 512434 477858 512466 478094
rect 512702 477858 512786 478094
rect 513022 477858 513054 478094
rect 512434 477774 513054 477858
rect 512434 477538 512466 477774
rect 512702 477538 512786 477774
rect 513022 477538 513054 477774
rect 512434 442094 513054 477538
rect 512434 441858 512466 442094
rect 512702 441858 512786 442094
rect 513022 441858 513054 442094
rect 512434 441774 513054 441858
rect 512434 441538 512466 441774
rect 512702 441538 512786 441774
rect 513022 441538 513054 441774
rect 512434 406094 513054 441538
rect 512434 405858 512466 406094
rect 512702 405858 512786 406094
rect 513022 405858 513054 406094
rect 512434 405774 513054 405858
rect 512434 405538 512466 405774
rect 512702 405538 512786 405774
rect 513022 405538 513054 405774
rect 512434 370094 513054 405538
rect 512434 369858 512466 370094
rect 512702 369858 512786 370094
rect 513022 369858 513054 370094
rect 512434 369774 513054 369858
rect 512434 369538 512466 369774
rect 512702 369538 512786 369774
rect 513022 369538 513054 369774
rect 512434 334094 513054 369538
rect 512434 333858 512466 334094
rect 512702 333858 512786 334094
rect 513022 333858 513054 334094
rect 512434 333774 513054 333858
rect 512434 333538 512466 333774
rect 512702 333538 512786 333774
rect 513022 333538 513054 333774
rect 512434 298094 513054 333538
rect 512434 297858 512466 298094
rect 512702 297858 512786 298094
rect 513022 297858 513054 298094
rect 512434 297774 513054 297858
rect 512434 297538 512466 297774
rect 512702 297538 512786 297774
rect 513022 297538 513054 297774
rect 512434 262094 513054 297538
rect 512434 261858 512466 262094
rect 512702 261858 512786 262094
rect 513022 261858 513054 262094
rect 512434 261774 513054 261858
rect 512434 261538 512466 261774
rect 512702 261538 512786 261774
rect 513022 261538 513054 261774
rect 512434 226094 513054 261538
rect 512434 225858 512466 226094
rect 512702 225858 512786 226094
rect 513022 225858 513054 226094
rect 512434 225774 513054 225858
rect 512434 225538 512466 225774
rect 512702 225538 512786 225774
rect 513022 225538 513054 225774
rect 512434 190094 513054 225538
rect 512434 189858 512466 190094
rect 512702 189858 512786 190094
rect 513022 189858 513054 190094
rect 512434 189774 513054 189858
rect 512434 189538 512466 189774
rect 512702 189538 512786 189774
rect 513022 189538 513054 189774
rect 512434 154094 513054 189538
rect 512434 153858 512466 154094
rect 512702 153858 512786 154094
rect 513022 153858 513054 154094
rect 512434 153774 513054 153858
rect 512434 153538 512466 153774
rect 512702 153538 512786 153774
rect 513022 153538 513054 153774
rect 512434 118094 513054 153538
rect 512434 117858 512466 118094
rect 512702 117858 512786 118094
rect 513022 117858 513054 118094
rect 512434 117774 513054 117858
rect 512434 117538 512466 117774
rect 512702 117538 512786 117774
rect 513022 117538 513054 117774
rect 512434 82094 513054 117538
rect 512434 81858 512466 82094
rect 512702 81858 512786 82094
rect 513022 81858 513054 82094
rect 512434 81774 513054 81858
rect 512434 81538 512466 81774
rect 512702 81538 512786 81774
rect 513022 81538 513054 81774
rect 512434 46094 513054 81538
rect 512434 45858 512466 46094
rect 512702 45858 512786 46094
rect 513022 45858 513054 46094
rect 512434 45774 513054 45858
rect 512434 45538 512466 45774
rect 512702 45538 512786 45774
rect 513022 45538 513054 45774
rect 512434 10094 513054 45538
rect 512434 9858 512466 10094
rect 512702 9858 512786 10094
rect 513022 9858 513054 10094
rect 512434 9774 513054 9858
rect 512434 9538 512466 9774
rect 512702 9538 512786 9774
rect 513022 9538 513054 9774
rect 512434 -6106 513054 9538
rect 512434 -6342 512466 -6106
rect 512702 -6342 512786 -6106
rect 513022 -6342 513054 -6106
rect 512434 -6426 513054 -6342
rect 512434 -6662 512466 -6426
rect 512702 -6662 512786 -6426
rect 513022 -6662 513054 -6426
rect 512434 -7654 513054 -6662
rect 513674 711558 514294 711590
rect 513674 711322 513706 711558
rect 513942 711322 514026 711558
rect 514262 711322 514294 711558
rect 513674 711238 514294 711322
rect 513674 711002 513706 711238
rect 513942 711002 514026 711238
rect 514262 711002 514294 711238
rect 513674 695334 514294 711002
rect 513674 695098 513706 695334
rect 513942 695098 514026 695334
rect 514262 695098 514294 695334
rect 513674 695014 514294 695098
rect 513674 694778 513706 695014
rect 513942 694778 514026 695014
rect 514262 694778 514294 695014
rect 513674 659334 514294 694778
rect 513674 659098 513706 659334
rect 513942 659098 514026 659334
rect 514262 659098 514294 659334
rect 513674 659014 514294 659098
rect 513674 658778 513706 659014
rect 513942 658778 514026 659014
rect 514262 658778 514294 659014
rect 513674 623334 514294 658778
rect 513674 623098 513706 623334
rect 513942 623098 514026 623334
rect 514262 623098 514294 623334
rect 513674 623014 514294 623098
rect 513674 622778 513706 623014
rect 513942 622778 514026 623014
rect 514262 622778 514294 623014
rect 513674 587334 514294 622778
rect 513674 587098 513706 587334
rect 513942 587098 514026 587334
rect 514262 587098 514294 587334
rect 513674 587014 514294 587098
rect 513674 586778 513706 587014
rect 513942 586778 514026 587014
rect 514262 586778 514294 587014
rect 513674 551334 514294 586778
rect 513674 551098 513706 551334
rect 513942 551098 514026 551334
rect 514262 551098 514294 551334
rect 513674 551014 514294 551098
rect 513674 550778 513706 551014
rect 513942 550778 514026 551014
rect 514262 550778 514294 551014
rect 513674 515334 514294 550778
rect 513674 515098 513706 515334
rect 513942 515098 514026 515334
rect 514262 515098 514294 515334
rect 513674 515014 514294 515098
rect 513674 514778 513706 515014
rect 513942 514778 514026 515014
rect 514262 514778 514294 515014
rect 513674 479334 514294 514778
rect 513674 479098 513706 479334
rect 513942 479098 514026 479334
rect 514262 479098 514294 479334
rect 513674 479014 514294 479098
rect 513674 478778 513706 479014
rect 513942 478778 514026 479014
rect 514262 478778 514294 479014
rect 513674 443334 514294 478778
rect 540994 704838 541614 711590
rect 540994 704602 541026 704838
rect 541262 704602 541346 704838
rect 541582 704602 541614 704838
rect 540994 704518 541614 704602
rect 540994 704282 541026 704518
rect 541262 704282 541346 704518
rect 541582 704282 541614 704518
rect 540994 686654 541614 704282
rect 540994 686418 541026 686654
rect 541262 686418 541346 686654
rect 541582 686418 541614 686654
rect 540994 686334 541614 686418
rect 540994 686098 541026 686334
rect 541262 686098 541346 686334
rect 541582 686098 541614 686334
rect 540994 650654 541614 686098
rect 540994 650418 541026 650654
rect 541262 650418 541346 650654
rect 541582 650418 541614 650654
rect 540994 650334 541614 650418
rect 540994 650098 541026 650334
rect 541262 650098 541346 650334
rect 541582 650098 541614 650334
rect 540994 614654 541614 650098
rect 540994 614418 541026 614654
rect 541262 614418 541346 614654
rect 541582 614418 541614 614654
rect 540994 614334 541614 614418
rect 540994 614098 541026 614334
rect 541262 614098 541346 614334
rect 541582 614098 541614 614334
rect 540994 578654 541614 614098
rect 540994 578418 541026 578654
rect 541262 578418 541346 578654
rect 541582 578418 541614 578654
rect 540994 578334 541614 578418
rect 540994 578098 541026 578334
rect 541262 578098 541346 578334
rect 541582 578098 541614 578334
rect 540994 542654 541614 578098
rect 540994 542418 541026 542654
rect 541262 542418 541346 542654
rect 541582 542418 541614 542654
rect 540994 542334 541614 542418
rect 540994 542098 541026 542334
rect 541262 542098 541346 542334
rect 541582 542098 541614 542334
rect 540994 506654 541614 542098
rect 540994 506418 541026 506654
rect 541262 506418 541346 506654
rect 541582 506418 541614 506654
rect 540994 506334 541614 506418
rect 540994 506098 541026 506334
rect 541262 506098 541346 506334
rect 541582 506098 541614 506334
rect 540994 470654 541614 506098
rect 540994 470418 541026 470654
rect 541262 470418 541346 470654
rect 541582 470418 541614 470654
rect 540994 470334 541614 470418
rect 540994 470098 541026 470334
rect 541262 470098 541346 470334
rect 541582 470098 541614 470334
rect 540994 445572 541614 470098
rect 542234 705798 542854 711590
rect 542234 705562 542266 705798
rect 542502 705562 542586 705798
rect 542822 705562 542854 705798
rect 542234 705478 542854 705562
rect 542234 705242 542266 705478
rect 542502 705242 542586 705478
rect 542822 705242 542854 705478
rect 542234 687894 542854 705242
rect 542234 687658 542266 687894
rect 542502 687658 542586 687894
rect 542822 687658 542854 687894
rect 542234 687574 542854 687658
rect 542234 687338 542266 687574
rect 542502 687338 542586 687574
rect 542822 687338 542854 687574
rect 542234 651894 542854 687338
rect 542234 651658 542266 651894
rect 542502 651658 542586 651894
rect 542822 651658 542854 651894
rect 542234 651574 542854 651658
rect 542234 651338 542266 651574
rect 542502 651338 542586 651574
rect 542822 651338 542854 651574
rect 542234 615894 542854 651338
rect 542234 615658 542266 615894
rect 542502 615658 542586 615894
rect 542822 615658 542854 615894
rect 542234 615574 542854 615658
rect 542234 615338 542266 615574
rect 542502 615338 542586 615574
rect 542822 615338 542854 615574
rect 542234 579894 542854 615338
rect 542234 579658 542266 579894
rect 542502 579658 542586 579894
rect 542822 579658 542854 579894
rect 542234 579574 542854 579658
rect 542234 579338 542266 579574
rect 542502 579338 542586 579574
rect 542822 579338 542854 579574
rect 542234 543894 542854 579338
rect 542234 543658 542266 543894
rect 542502 543658 542586 543894
rect 542822 543658 542854 543894
rect 542234 543574 542854 543658
rect 542234 543338 542266 543574
rect 542502 543338 542586 543574
rect 542822 543338 542854 543574
rect 542234 507894 542854 543338
rect 542234 507658 542266 507894
rect 542502 507658 542586 507894
rect 542822 507658 542854 507894
rect 542234 507574 542854 507658
rect 542234 507338 542266 507574
rect 542502 507338 542586 507574
rect 542822 507338 542854 507574
rect 542234 471894 542854 507338
rect 542234 471658 542266 471894
rect 542502 471658 542586 471894
rect 542822 471658 542854 471894
rect 542234 471574 542854 471658
rect 542234 471338 542266 471574
rect 542502 471338 542586 471574
rect 542822 471338 542854 471574
rect 542234 445572 542854 471338
rect 543474 706758 544094 711590
rect 543474 706522 543506 706758
rect 543742 706522 543826 706758
rect 544062 706522 544094 706758
rect 543474 706438 544094 706522
rect 543474 706202 543506 706438
rect 543742 706202 543826 706438
rect 544062 706202 544094 706438
rect 543474 689134 544094 706202
rect 543474 688898 543506 689134
rect 543742 688898 543826 689134
rect 544062 688898 544094 689134
rect 543474 688814 544094 688898
rect 543474 688578 543506 688814
rect 543742 688578 543826 688814
rect 544062 688578 544094 688814
rect 543474 653134 544094 688578
rect 543474 652898 543506 653134
rect 543742 652898 543826 653134
rect 544062 652898 544094 653134
rect 543474 652814 544094 652898
rect 543474 652578 543506 652814
rect 543742 652578 543826 652814
rect 544062 652578 544094 652814
rect 543474 617134 544094 652578
rect 543474 616898 543506 617134
rect 543742 616898 543826 617134
rect 544062 616898 544094 617134
rect 543474 616814 544094 616898
rect 543474 616578 543506 616814
rect 543742 616578 543826 616814
rect 544062 616578 544094 616814
rect 543474 581134 544094 616578
rect 543474 580898 543506 581134
rect 543742 580898 543826 581134
rect 544062 580898 544094 581134
rect 543474 580814 544094 580898
rect 543474 580578 543506 580814
rect 543742 580578 543826 580814
rect 544062 580578 544094 580814
rect 543474 545134 544094 580578
rect 543474 544898 543506 545134
rect 543742 544898 543826 545134
rect 544062 544898 544094 545134
rect 543474 544814 544094 544898
rect 543474 544578 543506 544814
rect 543742 544578 543826 544814
rect 544062 544578 544094 544814
rect 543474 509134 544094 544578
rect 543474 508898 543506 509134
rect 543742 508898 543826 509134
rect 544062 508898 544094 509134
rect 543474 508814 544094 508898
rect 543474 508578 543506 508814
rect 543742 508578 543826 508814
rect 544062 508578 544094 508814
rect 543474 473134 544094 508578
rect 543474 472898 543506 473134
rect 543742 472898 543826 473134
rect 544062 472898 544094 473134
rect 543474 472814 544094 472898
rect 543474 472578 543506 472814
rect 543742 472578 543826 472814
rect 544062 472578 544094 472814
rect 543474 445572 544094 472578
rect 544714 707718 545334 711590
rect 544714 707482 544746 707718
rect 544982 707482 545066 707718
rect 545302 707482 545334 707718
rect 544714 707398 545334 707482
rect 544714 707162 544746 707398
rect 544982 707162 545066 707398
rect 545302 707162 545334 707398
rect 544714 690374 545334 707162
rect 544714 690138 544746 690374
rect 544982 690138 545066 690374
rect 545302 690138 545334 690374
rect 544714 690054 545334 690138
rect 544714 689818 544746 690054
rect 544982 689818 545066 690054
rect 545302 689818 545334 690054
rect 544714 654374 545334 689818
rect 544714 654138 544746 654374
rect 544982 654138 545066 654374
rect 545302 654138 545334 654374
rect 544714 654054 545334 654138
rect 544714 653818 544746 654054
rect 544982 653818 545066 654054
rect 545302 653818 545334 654054
rect 544714 618374 545334 653818
rect 544714 618138 544746 618374
rect 544982 618138 545066 618374
rect 545302 618138 545334 618374
rect 544714 618054 545334 618138
rect 544714 617818 544746 618054
rect 544982 617818 545066 618054
rect 545302 617818 545334 618054
rect 544714 582374 545334 617818
rect 544714 582138 544746 582374
rect 544982 582138 545066 582374
rect 545302 582138 545334 582374
rect 544714 582054 545334 582138
rect 544714 581818 544746 582054
rect 544982 581818 545066 582054
rect 545302 581818 545334 582054
rect 544714 546374 545334 581818
rect 544714 546138 544746 546374
rect 544982 546138 545066 546374
rect 545302 546138 545334 546374
rect 544714 546054 545334 546138
rect 544714 545818 544746 546054
rect 544982 545818 545066 546054
rect 545302 545818 545334 546054
rect 544714 510374 545334 545818
rect 544714 510138 544746 510374
rect 544982 510138 545066 510374
rect 545302 510138 545334 510374
rect 544714 510054 545334 510138
rect 544714 509818 544746 510054
rect 544982 509818 545066 510054
rect 545302 509818 545334 510054
rect 544714 474374 545334 509818
rect 544714 474138 544746 474374
rect 544982 474138 545066 474374
rect 545302 474138 545334 474374
rect 544714 474054 545334 474138
rect 544714 473818 544746 474054
rect 544982 473818 545066 474054
rect 545302 473818 545334 474054
rect 544714 445572 545334 473818
rect 545954 708678 546574 711590
rect 545954 708442 545986 708678
rect 546222 708442 546306 708678
rect 546542 708442 546574 708678
rect 545954 708358 546574 708442
rect 545954 708122 545986 708358
rect 546222 708122 546306 708358
rect 546542 708122 546574 708358
rect 545954 691614 546574 708122
rect 545954 691378 545986 691614
rect 546222 691378 546306 691614
rect 546542 691378 546574 691614
rect 545954 691294 546574 691378
rect 545954 691058 545986 691294
rect 546222 691058 546306 691294
rect 546542 691058 546574 691294
rect 545954 655614 546574 691058
rect 545954 655378 545986 655614
rect 546222 655378 546306 655614
rect 546542 655378 546574 655614
rect 545954 655294 546574 655378
rect 545954 655058 545986 655294
rect 546222 655058 546306 655294
rect 546542 655058 546574 655294
rect 545954 619614 546574 655058
rect 545954 619378 545986 619614
rect 546222 619378 546306 619614
rect 546542 619378 546574 619614
rect 545954 619294 546574 619378
rect 545954 619058 545986 619294
rect 546222 619058 546306 619294
rect 546542 619058 546574 619294
rect 545954 583614 546574 619058
rect 545954 583378 545986 583614
rect 546222 583378 546306 583614
rect 546542 583378 546574 583614
rect 545954 583294 546574 583378
rect 545954 583058 545986 583294
rect 546222 583058 546306 583294
rect 546542 583058 546574 583294
rect 545954 547614 546574 583058
rect 545954 547378 545986 547614
rect 546222 547378 546306 547614
rect 546542 547378 546574 547614
rect 545954 547294 546574 547378
rect 545954 547058 545986 547294
rect 546222 547058 546306 547294
rect 546542 547058 546574 547294
rect 545954 511614 546574 547058
rect 545954 511378 545986 511614
rect 546222 511378 546306 511614
rect 546542 511378 546574 511614
rect 545954 511294 546574 511378
rect 545954 511058 545986 511294
rect 546222 511058 546306 511294
rect 546542 511058 546574 511294
rect 545954 475614 546574 511058
rect 545954 475378 545986 475614
rect 546222 475378 546306 475614
rect 546542 475378 546574 475614
rect 545954 475294 546574 475378
rect 545954 475058 545986 475294
rect 546222 475058 546306 475294
rect 546542 475058 546574 475294
rect 545954 445572 546574 475058
rect 547194 709638 547814 711590
rect 547194 709402 547226 709638
rect 547462 709402 547546 709638
rect 547782 709402 547814 709638
rect 547194 709318 547814 709402
rect 547194 709082 547226 709318
rect 547462 709082 547546 709318
rect 547782 709082 547814 709318
rect 547194 692854 547814 709082
rect 547194 692618 547226 692854
rect 547462 692618 547546 692854
rect 547782 692618 547814 692854
rect 547194 692534 547814 692618
rect 547194 692298 547226 692534
rect 547462 692298 547546 692534
rect 547782 692298 547814 692534
rect 547194 656854 547814 692298
rect 547194 656618 547226 656854
rect 547462 656618 547546 656854
rect 547782 656618 547814 656854
rect 547194 656534 547814 656618
rect 547194 656298 547226 656534
rect 547462 656298 547546 656534
rect 547782 656298 547814 656534
rect 547194 620854 547814 656298
rect 547194 620618 547226 620854
rect 547462 620618 547546 620854
rect 547782 620618 547814 620854
rect 547194 620534 547814 620618
rect 547194 620298 547226 620534
rect 547462 620298 547546 620534
rect 547782 620298 547814 620534
rect 547194 584854 547814 620298
rect 547194 584618 547226 584854
rect 547462 584618 547546 584854
rect 547782 584618 547814 584854
rect 547194 584534 547814 584618
rect 547194 584298 547226 584534
rect 547462 584298 547546 584534
rect 547782 584298 547814 584534
rect 547194 548854 547814 584298
rect 547194 548618 547226 548854
rect 547462 548618 547546 548854
rect 547782 548618 547814 548854
rect 547194 548534 547814 548618
rect 547194 548298 547226 548534
rect 547462 548298 547546 548534
rect 547782 548298 547814 548534
rect 547194 512854 547814 548298
rect 547194 512618 547226 512854
rect 547462 512618 547546 512854
rect 547782 512618 547814 512854
rect 547194 512534 547814 512618
rect 547194 512298 547226 512534
rect 547462 512298 547546 512534
rect 547782 512298 547814 512534
rect 547194 476854 547814 512298
rect 547194 476618 547226 476854
rect 547462 476618 547546 476854
rect 547782 476618 547814 476854
rect 547194 476534 547814 476618
rect 547194 476298 547226 476534
rect 547462 476298 547546 476534
rect 547782 476298 547814 476534
rect 541571 445092 541637 445093
rect 541571 445028 541572 445092
rect 541636 445028 541637 445092
rect 541571 445027 541637 445028
rect 544331 445092 544397 445093
rect 544331 445028 544332 445092
rect 544396 445028 544397 445092
rect 544331 445027 544397 445028
rect 513674 443098 513706 443334
rect 513942 443098 514026 443334
rect 514262 443098 514294 443334
rect 513674 443014 514294 443098
rect 513674 442778 513706 443014
rect 513942 442778 514026 443014
rect 514262 442778 514294 443014
rect 513674 407334 514294 442778
rect 540876 435894 541196 435926
rect 540876 435658 540918 435894
rect 541154 435658 541196 435894
rect 540876 435574 541196 435658
rect 540876 435338 540918 435574
rect 541154 435338 541196 435574
rect 540876 435306 541196 435338
rect 539910 434654 540230 434686
rect 539910 434418 539952 434654
rect 540188 434418 540230 434654
rect 539910 434334 540230 434418
rect 539910 434098 539952 434334
rect 540188 434098 540230 434334
rect 539910 434066 540230 434098
rect 541574 409325 541634 445027
rect 542808 435894 543128 435926
rect 542808 435658 542850 435894
rect 543086 435658 543128 435894
rect 542808 435574 543128 435658
rect 542808 435338 542850 435574
rect 543086 435338 543128 435574
rect 542808 435306 543128 435338
rect 541842 434654 542162 434686
rect 541842 434418 541884 434654
rect 542120 434418 542162 434654
rect 541842 434334 542162 434418
rect 541842 434098 541884 434334
rect 542120 434098 542162 434334
rect 541842 434066 542162 434098
rect 543774 434654 544094 434686
rect 543774 434418 543816 434654
rect 544052 434418 544094 434654
rect 543774 434334 544094 434418
rect 543774 434098 543816 434334
rect 544052 434098 544094 434334
rect 543774 434066 544094 434098
rect 544334 409325 544394 445027
rect 547194 440854 547814 476298
rect 547194 440618 547226 440854
rect 547462 440618 547546 440854
rect 547782 440618 547814 440854
rect 547194 440534 547814 440618
rect 547194 440298 547226 440534
rect 547462 440298 547546 440534
rect 547782 440298 547814 440534
rect 544740 435894 545060 435926
rect 544740 435658 544782 435894
rect 545018 435658 545060 435894
rect 544740 435574 545060 435658
rect 544740 435338 544782 435574
rect 545018 435338 545060 435574
rect 544740 435306 545060 435338
rect 546672 435894 546992 435926
rect 546672 435658 546714 435894
rect 546950 435658 546992 435894
rect 546672 435574 546992 435658
rect 546672 435338 546714 435574
rect 546950 435338 546992 435574
rect 546672 435306 546992 435338
rect 545706 434654 546026 434686
rect 545706 434418 545748 434654
rect 545984 434418 546026 434654
rect 545706 434334 546026 434418
rect 545706 434098 545748 434334
rect 545984 434098 546026 434334
rect 545706 434066 546026 434098
rect 541571 409324 541637 409325
rect 541571 409260 541572 409324
rect 541636 409260 541637 409324
rect 541571 409259 541637 409260
rect 544331 409324 544397 409325
rect 544331 409260 544332 409324
rect 544396 409260 544397 409324
rect 544331 409259 544397 409260
rect 513674 407098 513706 407334
rect 513942 407098 514026 407334
rect 514262 407098 514294 407334
rect 513674 407014 514294 407098
rect 513674 406778 513706 407014
rect 513942 406778 514026 407014
rect 514262 406778 514294 407014
rect 513674 371334 514294 406778
rect 540876 399894 541196 399926
rect 540876 399658 540918 399894
rect 541154 399658 541196 399894
rect 540876 399574 541196 399658
rect 540876 399338 540918 399574
rect 541154 399338 541196 399574
rect 540876 399306 541196 399338
rect 539910 398654 540230 398686
rect 539910 398418 539952 398654
rect 540188 398418 540230 398654
rect 539910 398334 540230 398418
rect 539910 398098 539952 398334
rect 540188 398098 540230 398334
rect 539910 398066 540230 398098
rect 541574 373149 541634 409259
rect 542808 399894 543128 399926
rect 542808 399658 542850 399894
rect 543086 399658 543128 399894
rect 542808 399574 543128 399658
rect 542808 399338 542850 399574
rect 543086 399338 543128 399574
rect 542808 399306 543128 399338
rect 541842 398654 542162 398686
rect 541842 398418 541884 398654
rect 542120 398418 542162 398654
rect 541842 398334 542162 398418
rect 541842 398098 541884 398334
rect 542120 398098 542162 398334
rect 541842 398066 542162 398098
rect 543774 398654 544094 398686
rect 543774 398418 543816 398654
rect 544052 398418 544094 398654
rect 543774 398334 544094 398418
rect 543774 398098 543816 398334
rect 544052 398098 544094 398334
rect 543774 398066 544094 398098
rect 544334 383670 544394 409259
rect 547194 404854 547814 440298
rect 547194 404618 547226 404854
rect 547462 404618 547546 404854
rect 547782 404618 547814 404854
rect 547194 404534 547814 404618
rect 547194 404298 547226 404534
rect 547462 404298 547546 404534
rect 547782 404298 547814 404534
rect 544740 399894 545060 399926
rect 544740 399658 544782 399894
rect 545018 399658 545060 399894
rect 544740 399574 545060 399658
rect 544740 399338 544782 399574
rect 545018 399338 545060 399574
rect 544740 399306 545060 399338
rect 546672 399894 546992 399926
rect 546672 399658 546714 399894
rect 546950 399658 546992 399894
rect 546672 399574 546992 399658
rect 546672 399338 546714 399574
rect 546950 399338 546992 399574
rect 546672 399306 546992 399338
rect 545706 398654 546026 398686
rect 545706 398418 545748 398654
rect 545984 398418 546026 398654
rect 545706 398334 546026 398418
rect 545706 398098 545748 398334
rect 545984 398098 546026 398334
rect 545706 398066 546026 398098
rect 544334 383610 544578 383670
rect 544518 373421 544578 383610
rect 544515 373420 544581 373421
rect 544515 373356 544516 373420
rect 544580 373356 544581 373420
rect 544515 373355 544581 373356
rect 541571 373148 541637 373149
rect 541571 373084 541572 373148
rect 541636 373084 541637 373148
rect 541571 373083 541637 373084
rect 513674 371098 513706 371334
rect 513942 371098 514026 371334
rect 514262 371098 514294 371334
rect 513674 371014 514294 371098
rect 513674 370778 513706 371014
rect 513942 370778 514026 371014
rect 514262 370778 514294 371014
rect 513674 335334 514294 370778
rect 540876 363894 541196 363926
rect 540876 363658 540918 363894
rect 541154 363658 541196 363894
rect 540876 363574 541196 363658
rect 540876 363338 540918 363574
rect 541154 363338 541196 363574
rect 540876 363306 541196 363338
rect 539910 362654 540230 362686
rect 539910 362418 539952 362654
rect 540188 362418 540230 362654
rect 539910 362334 540230 362418
rect 539910 362098 539952 362334
rect 540188 362098 540230 362334
rect 539910 362066 540230 362098
rect 541574 339557 541634 373083
rect 542808 363894 543128 363926
rect 542808 363658 542850 363894
rect 543086 363658 543128 363894
rect 542808 363574 543128 363658
rect 542808 363338 542850 363574
rect 543086 363338 543128 363574
rect 542808 363306 543128 363338
rect 541842 362654 542162 362686
rect 541842 362418 541884 362654
rect 542120 362418 542162 362654
rect 541842 362334 542162 362418
rect 541842 362098 541884 362334
rect 542120 362098 542162 362334
rect 541842 362066 542162 362098
rect 543774 362654 544094 362686
rect 543774 362418 543816 362654
rect 544052 362418 544094 362654
rect 543774 362334 544094 362418
rect 543774 362098 543816 362334
rect 544052 362098 544094 362334
rect 543774 362066 544094 362098
rect 544518 354690 544578 373355
rect 547194 368854 547814 404298
rect 547194 368618 547226 368854
rect 547462 368618 547546 368854
rect 547782 368618 547814 368854
rect 547194 368534 547814 368618
rect 547194 368298 547226 368534
rect 547462 368298 547546 368534
rect 547782 368298 547814 368534
rect 544740 363894 545060 363926
rect 544740 363658 544782 363894
rect 545018 363658 545060 363894
rect 544740 363574 545060 363658
rect 544740 363338 544782 363574
rect 545018 363338 545060 363574
rect 544740 363306 545060 363338
rect 546672 363894 546992 363926
rect 546672 363658 546714 363894
rect 546950 363658 546992 363894
rect 546672 363574 546992 363658
rect 546672 363338 546714 363574
rect 546950 363338 546992 363574
rect 546672 363306 546992 363338
rect 545706 362654 546026 362686
rect 545706 362418 545748 362654
rect 545984 362418 546026 362654
rect 545706 362334 546026 362418
rect 545706 362098 545748 362334
rect 545984 362098 546026 362334
rect 545706 362066 546026 362098
rect 544334 354630 544578 354690
rect 544334 351933 544394 354630
rect 544331 351932 544397 351933
rect 544331 351868 544332 351932
rect 544396 351868 544397 351932
rect 544331 351867 544397 351868
rect 544334 339557 544394 351867
rect 541571 339556 541637 339557
rect 541571 339492 541572 339556
rect 541636 339492 541637 339556
rect 541571 339491 541637 339492
rect 544331 339556 544397 339557
rect 544331 339492 544332 339556
rect 544396 339492 544397 339556
rect 544331 339491 544397 339492
rect 513674 335098 513706 335334
rect 513942 335098 514026 335334
rect 514262 335098 514294 335334
rect 513674 335014 514294 335098
rect 513674 334778 513706 335014
rect 513942 334778 514026 335014
rect 514262 334778 514294 335014
rect 513674 299334 514294 334778
rect 540876 327894 541196 327926
rect 540876 327658 540918 327894
rect 541154 327658 541196 327894
rect 540876 327574 541196 327658
rect 540876 327338 540918 327574
rect 541154 327338 541196 327574
rect 540876 327306 541196 327338
rect 539910 326654 540230 326686
rect 539910 326418 539952 326654
rect 540188 326418 540230 326654
rect 539910 326334 540230 326418
rect 539910 326098 539952 326334
rect 540188 326098 540230 326334
rect 539910 326066 540230 326098
rect 541574 303653 541634 339491
rect 542808 327894 543128 327926
rect 542808 327658 542850 327894
rect 543086 327658 543128 327894
rect 542808 327574 543128 327658
rect 542808 327338 542850 327574
rect 543086 327338 543128 327574
rect 542808 327306 543128 327338
rect 541842 326654 542162 326686
rect 541842 326418 541884 326654
rect 542120 326418 542162 326654
rect 541842 326334 542162 326418
rect 541842 326098 541884 326334
rect 542120 326098 542162 326334
rect 541842 326066 542162 326098
rect 543774 326654 544094 326686
rect 543774 326418 543816 326654
rect 544052 326418 544094 326654
rect 543774 326334 544094 326418
rect 543774 326098 543816 326334
rect 544052 326098 544094 326334
rect 543774 326066 544094 326098
rect 544334 303789 544394 339491
rect 547194 332854 547814 368298
rect 547194 332618 547226 332854
rect 547462 332618 547546 332854
rect 547782 332618 547814 332854
rect 547194 332534 547814 332618
rect 547194 332298 547226 332534
rect 547462 332298 547546 332534
rect 547782 332298 547814 332534
rect 544740 327894 545060 327926
rect 544740 327658 544782 327894
rect 545018 327658 545060 327894
rect 544740 327574 545060 327658
rect 544740 327338 544782 327574
rect 545018 327338 545060 327574
rect 544740 327306 545060 327338
rect 546672 327894 546992 327926
rect 546672 327658 546714 327894
rect 546950 327658 546992 327894
rect 546672 327574 546992 327658
rect 546672 327338 546714 327574
rect 546950 327338 546992 327574
rect 546672 327306 546992 327338
rect 545706 326654 546026 326686
rect 545706 326418 545748 326654
rect 545984 326418 546026 326654
rect 545706 326334 546026 326418
rect 545706 326098 545748 326334
rect 545984 326098 546026 326334
rect 545706 326066 546026 326098
rect 544331 303788 544397 303789
rect 544331 303724 544332 303788
rect 544396 303724 544397 303788
rect 544331 303723 544397 303724
rect 541571 303652 541637 303653
rect 541571 303588 541572 303652
rect 541636 303588 541637 303652
rect 541571 303587 541637 303588
rect 513674 299098 513706 299334
rect 513942 299098 514026 299334
rect 514262 299098 514294 299334
rect 513674 299014 514294 299098
rect 513674 298778 513706 299014
rect 513942 298778 514026 299014
rect 514262 298778 514294 299014
rect 513674 263334 514294 298778
rect 547194 296854 547814 332298
rect 547194 296618 547226 296854
rect 547462 296618 547546 296854
rect 547782 296618 547814 296854
rect 547194 296534 547814 296618
rect 547194 296298 547226 296534
rect 547462 296298 547546 296534
rect 547782 296298 547814 296534
rect 540876 291894 541196 291926
rect 540876 291658 540918 291894
rect 541154 291658 541196 291894
rect 540876 291574 541196 291658
rect 540876 291338 540918 291574
rect 541154 291338 541196 291574
rect 540876 291306 541196 291338
rect 542808 291894 543128 291926
rect 542808 291658 542850 291894
rect 543086 291658 543128 291894
rect 542808 291574 543128 291658
rect 542808 291338 542850 291574
rect 543086 291338 543128 291574
rect 542808 291306 543128 291338
rect 544740 291894 545060 291926
rect 544740 291658 544782 291894
rect 545018 291658 545060 291894
rect 544740 291574 545060 291658
rect 544740 291338 544782 291574
rect 545018 291338 545060 291574
rect 544740 291306 545060 291338
rect 546672 291894 546992 291926
rect 546672 291658 546714 291894
rect 546950 291658 546992 291894
rect 546672 291574 546992 291658
rect 546672 291338 546714 291574
rect 546950 291338 546992 291574
rect 546672 291306 546992 291338
rect 539910 290654 540230 290686
rect 539910 290418 539952 290654
rect 540188 290418 540230 290654
rect 539910 290334 540230 290418
rect 539910 290098 539952 290334
rect 540188 290098 540230 290334
rect 539910 290066 540230 290098
rect 541842 290654 542162 290686
rect 541842 290418 541884 290654
rect 542120 290418 542162 290654
rect 541842 290334 542162 290418
rect 541842 290098 541884 290334
rect 542120 290098 542162 290334
rect 541842 290066 542162 290098
rect 543774 290654 544094 290686
rect 543774 290418 543816 290654
rect 544052 290418 544094 290654
rect 543774 290334 544094 290418
rect 543774 290098 543816 290334
rect 544052 290098 544094 290334
rect 543774 290066 544094 290098
rect 545706 290654 546026 290686
rect 545706 290418 545748 290654
rect 545984 290418 546026 290654
rect 545706 290334 546026 290418
rect 545706 290098 545748 290334
rect 545984 290098 546026 290334
rect 545706 290066 546026 290098
rect 513674 263098 513706 263334
rect 513942 263098 514026 263334
rect 514262 263098 514294 263334
rect 513674 263014 514294 263098
rect 513674 262778 513706 263014
rect 513942 262778 514026 263014
rect 514262 262778 514294 263014
rect 513674 227334 514294 262778
rect 513674 227098 513706 227334
rect 513942 227098 514026 227334
rect 514262 227098 514294 227334
rect 513674 227014 514294 227098
rect 513674 226778 513706 227014
rect 513942 226778 514026 227014
rect 514262 226778 514294 227014
rect 513674 191334 514294 226778
rect 513674 191098 513706 191334
rect 513942 191098 514026 191334
rect 514262 191098 514294 191334
rect 513674 191014 514294 191098
rect 513674 190778 513706 191014
rect 513942 190778 514026 191014
rect 514262 190778 514294 191014
rect 513674 155334 514294 190778
rect 513674 155098 513706 155334
rect 513942 155098 514026 155334
rect 514262 155098 514294 155334
rect 513674 155014 514294 155098
rect 513674 154778 513706 155014
rect 513942 154778 514026 155014
rect 514262 154778 514294 155014
rect 513674 119334 514294 154778
rect 513674 119098 513706 119334
rect 513942 119098 514026 119334
rect 514262 119098 514294 119334
rect 513674 119014 514294 119098
rect 513674 118778 513706 119014
rect 513942 118778 514026 119014
rect 514262 118778 514294 119014
rect 513674 83334 514294 118778
rect 513674 83098 513706 83334
rect 513942 83098 514026 83334
rect 514262 83098 514294 83334
rect 513674 83014 514294 83098
rect 513674 82778 513706 83014
rect 513942 82778 514026 83014
rect 514262 82778 514294 83014
rect 513674 47334 514294 82778
rect 513674 47098 513706 47334
rect 513942 47098 514026 47334
rect 514262 47098 514294 47334
rect 513674 47014 514294 47098
rect 513674 46778 513706 47014
rect 513942 46778 514026 47014
rect 514262 46778 514294 47014
rect 513674 11334 514294 46778
rect 513674 11098 513706 11334
rect 513942 11098 514026 11334
rect 514262 11098 514294 11334
rect 513674 11014 514294 11098
rect 513674 10778 513706 11014
rect 513942 10778 514026 11014
rect 514262 10778 514294 11014
rect 513674 -7066 514294 10778
rect 513674 -7302 513706 -7066
rect 513942 -7302 514026 -7066
rect 514262 -7302 514294 -7066
rect 513674 -7386 514294 -7302
rect 513674 -7622 513706 -7386
rect 513942 -7622 514026 -7386
rect 514262 -7622 514294 -7386
rect 513674 -7654 514294 -7622
rect 540994 254654 541614 279788
rect 540994 254418 541026 254654
rect 541262 254418 541346 254654
rect 541582 254418 541614 254654
rect 540994 254334 541614 254418
rect 540994 254098 541026 254334
rect 541262 254098 541346 254334
rect 541582 254098 541614 254334
rect 540994 218654 541614 254098
rect 540994 218418 541026 218654
rect 541262 218418 541346 218654
rect 541582 218418 541614 218654
rect 540994 218334 541614 218418
rect 540994 218098 541026 218334
rect 541262 218098 541346 218334
rect 541582 218098 541614 218334
rect 540994 182654 541614 218098
rect 540994 182418 541026 182654
rect 541262 182418 541346 182654
rect 541582 182418 541614 182654
rect 540994 182334 541614 182418
rect 540994 182098 541026 182334
rect 541262 182098 541346 182334
rect 541582 182098 541614 182334
rect 540994 146654 541614 182098
rect 540994 146418 541026 146654
rect 541262 146418 541346 146654
rect 541582 146418 541614 146654
rect 540994 146334 541614 146418
rect 540994 146098 541026 146334
rect 541262 146098 541346 146334
rect 541582 146098 541614 146334
rect 540994 110654 541614 146098
rect 540994 110418 541026 110654
rect 541262 110418 541346 110654
rect 541582 110418 541614 110654
rect 540994 110334 541614 110418
rect 540994 110098 541026 110334
rect 541262 110098 541346 110334
rect 541582 110098 541614 110334
rect 540994 74654 541614 110098
rect 540994 74418 541026 74654
rect 541262 74418 541346 74654
rect 541582 74418 541614 74654
rect 540994 74334 541614 74418
rect 540994 74098 541026 74334
rect 541262 74098 541346 74334
rect 541582 74098 541614 74334
rect 540994 38654 541614 74098
rect 540994 38418 541026 38654
rect 541262 38418 541346 38654
rect 541582 38418 541614 38654
rect 540994 38334 541614 38418
rect 540994 38098 541026 38334
rect 541262 38098 541346 38334
rect 541582 38098 541614 38334
rect 540994 2654 541614 38098
rect 540994 2418 541026 2654
rect 541262 2418 541346 2654
rect 541582 2418 541614 2654
rect 540994 2334 541614 2418
rect 540994 2098 541026 2334
rect 541262 2098 541346 2334
rect 541582 2098 541614 2334
rect 540994 -346 541614 2098
rect 540994 -582 541026 -346
rect 541262 -582 541346 -346
rect 541582 -582 541614 -346
rect 540994 -666 541614 -582
rect 540994 -902 541026 -666
rect 541262 -902 541346 -666
rect 541582 -902 541614 -666
rect 540994 -7654 541614 -902
rect 542234 255894 542854 279788
rect 542234 255658 542266 255894
rect 542502 255658 542586 255894
rect 542822 255658 542854 255894
rect 542234 255574 542854 255658
rect 542234 255338 542266 255574
rect 542502 255338 542586 255574
rect 542822 255338 542854 255574
rect 542234 219894 542854 255338
rect 542234 219658 542266 219894
rect 542502 219658 542586 219894
rect 542822 219658 542854 219894
rect 542234 219574 542854 219658
rect 542234 219338 542266 219574
rect 542502 219338 542586 219574
rect 542822 219338 542854 219574
rect 542234 183894 542854 219338
rect 542234 183658 542266 183894
rect 542502 183658 542586 183894
rect 542822 183658 542854 183894
rect 542234 183574 542854 183658
rect 542234 183338 542266 183574
rect 542502 183338 542586 183574
rect 542822 183338 542854 183574
rect 542234 147894 542854 183338
rect 542234 147658 542266 147894
rect 542502 147658 542586 147894
rect 542822 147658 542854 147894
rect 542234 147574 542854 147658
rect 542234 147338 542266 147574
rect 542502 147338 542586 147574
rect 542822 147338 542854 147574
rect 542234 111894 542854 147338
rect 542234 111658 542266 111894
rect 542502 111658 542586 111894
rect 542822 111658 542854 111894
rect 542234 111574 542854 111658
rect 542234 111338 542266 111574
rect 542502 111338 542586 111574
rect 542822 111338 542854 111574
rect 542234 75894 542854 111338
rect 542234 75658 542266 75894
rect 542502 75658 542586 75894
rect 542822 75658 542854 75894
rect 542234 75574 542854 75658
rect 542234 75338 542266 75574
rect 542502 75338 542586 75574
rect 542822 75338 542854 75574
rect 542234 39894 542854 75338
rect 542234 39658 542266 39894
rect 542502 39658 542586 39894
rect 542822 39658 542854 39894
rect 542234 39574 542854 39658
rect 542234 39338 542266 39574
rect 542502 39338 542586 39574
rect 542822 39338 542854 39574
rect 542234 3894 542854 39338
rect 542234 3658 542266 3894
rect 542502 3658 542586 3894
rect 542822 3658 542854 3894
rect 542234 3574 542854 3658
rect 542234 3338 542266 3574
rect 542502 3338 542586 3574
rect 542822 3338 542854 3574
rect 542234 -1306 542854 3338
rect 542234 -1542 542266 -1306
rect 542502 -1542 542586 -1306
rect 542822 -1542 542854 -1306
rect 542234 -1626 542854 -1542
rect 542234 -1862 542266 -1626
rect 542502 -1862 542586 -1626
rect 542822 -1862 542854 -1626
rect 542234 -7654 542854 -1862
rect 543474 257134 544094 279788
rect 543474 256898 543506 257134
rect 543742 256898 543826 257134
rect 544062 256898 544094 257134
rect 543474 256814 544094 256898
rect 543474 256578 543506 256814
rect 543742 256578 543826 256814
rect 544062 256578 544094 256814
rect 543474 221134 544094 256578
rect 543474 220898 543506 221134
rect 543742 220898 543826 221134
rect 544062 220898 544094 221134
rect 543474 220814 544094 220898
rect 543474 220578 543506 220814
rect 543742 220578 543826 220814
rect 544062 220578 544094 220814
rect 543474 185134 544094 220578
rect 543474 184898 543506 185134
rect 543742 184898 543826 185134
rect 544062 184898 544094 185134
rect 543474 184814 544094 184898
rect 543474 184578 543506 184814
rect 543742 184578 543826 184814
rect 544062 184578 544094 184814
rect 543474 149134 544094 184578
rect 543474 148898 543506 149134
rect 543742 148898 543826 149134
rect 544062 148898 544094 149134
rect 543474 148814 544094 148898
rect 543474 148578 543506 148814
rect 543742 148578 543826 148814
rect 544062 148578 544094 148814
rect 543474 113134 544094 148578
rect 543474 112898 543506 113134
rect 543742 112898 543826 113134
rect 544062 112898 544094 113134
rect 543474 112814 544094 112898
rect 543474 112578 543506 112814
rect 543742 112578 543826 112814
rect 544062 112578 544094 112814
rect 543474 77134 544094 112578
rect 543474 76898 543506 77134
rect 543742 76898 543826 77134
rect 544062 76898 544094 77134
rect 543474 76814 544094 76898
rect 543474 76578 543506 76814
rect 543742 76578 543826 76814
rect 544062 76578 544094 76814
rect 543474 41134 544094 76578
rect 543474 40898 543506 41134
rect 543742 40898 543826 41134
rect 544062 40898 544094 41134
rect 543474 40814 544094 40898
rect 543474 40578 543506 40814
rect 543742 40578 543826 40814
rect 544062 40578 544094 40814
rect 543474 5134 544094 40578
rect 543474 4898 543506 5134
rect 543742 4898 543826 5134
rect 544062 4898 544094 5134
rect 543474 4814 544094 4898
rect 543474 4578 543506 4814
rect 543742 4578 543826 4814
rect 544062 4578 544094 4814
rect 543474 -2266 544094 4578
rect 543474 -2502 543506 -2266
rect 543742 -2502 543826 -2266
rect 544062 -2502 544094 -2266
rect 543474 -2586 544094 -2502
rect 543474 -2822 543506 -2586
rect 543742 -2822 543826 -2586
rect 544062 -2822 544094 -2586
rect 543474 -7654 544094 -2822
rect 544714 258374 545334 279788
rect 544714 258138 544746 258374
rect 544982 258138 545066 258374
rect 545302 258138 545334 258374
rect 544714 258054 545334 258138
rect 544714 257818 544746 258054
rect 544982 257818 545066 258054
rect 545302 257818 545334 258054
rect 544714 222374 545334 257818
rect 544714 222138 544746 222374
rect 544982 222138 545066 222374
rect 545302 222138 545334 222374
rect 544714 222054 545334 222138
rect 544714 221818 544746 222054
rect 544982 221818 545066 222054
rect 545302 221818 545334 222054
rect 544714 186374 545334 221818
rect 544714 186138 544746 186374
rect 544982 186138 545066 186374
rect 545302 186138 545334 186374
rect 544714 186054 545334 186138
rect 544714 185818 544746 186054
rect 544982 185818 545066 186054
rect 545302 185818 545334 186054
rect 544714 150374 545334 185818
rect 544714 150138 544746 150374
rect 544982 150138 545066 150374
rect 545302 150138 545334 150374
rect 544714 150054 545334 150138
rect 544714 149818 544746 150054
rect 544982 149818 545066 150054
rect 545302 149818 545334 150054
rect 544714 114374 545334 149818
rect 544714 114138 544746 114374
rect 544982 114138 545066 114374
rect 545302 114138 545334 114374
rect 544714 114054 545334 114138
rect 544714 113818 544746 114054
rect 544982 113818 545066 114054
rect 545302 113818 545334 114054
rect 544714 78374 545334 113818
rect 544714 78138 544746 78374
rect 544982 78138 545066 78374
rect 545302 78138 545334 78374
rect 544714 78054 545334 78138
rect 544714 77818 544746 78054
rect 544982 77818 545066 78054
rect 545302 77818 545334 78054
rect 544714 42374 545334 77818
rect 544714 42138 544746 42374
rect 544982 42138 545066 42374
rect 545302 42138 545334 42374
rect 544714 42054 545334 42138
rect 544714 41818 544746 42054
rect 544982 41818 545066 42054
rect 545302 41818 545334 42054
rect 544714 6374 545334 41818
rect 544714 6138 544746 6374
rect 544982 6138 545066 6374
rect 545302 6138 545334 6374
rect 544714 6054 545334 6138
rect 544714 5818 544746 6054
rect 544982 5818 545066 6054
rect 545302 5818 545334 6054
rect 544714 -3226 545334 5818
rect 544714 -3462 544746 -3226
rect 544982 -3462 545066 -3226
rect 545302 -3462 545334 -3226
rect 544714 -3546 545334 -3462
rect 544714 -3782 544746 -3546
rect 544982 -3782 545066 -3546
rect 545302 -3782 545334 -3546
rect 544714 -7654 545334 -3782
rect 545954 259614 546574 279788
rect 545954 259378 545986 259614
rect 546222 259378 546306 259614
rect 546542 259378 546574 259614
rect 545954 259294 546574 259378
rect 545954 259058 545986 259294
rect 546222 259058 546306 259294
rect 546542 259058 546574 259294
rect 545954 223614 546574 259058
rect 545954 223378 545986 223614
rect 546222 223378 546306 223614
rect 546542 223378 546574 223614
rect 545954 223294 546574 223378
rect 545954 223058 545986 223294
rect 546222 223058 546306 223294
rect 546542 223058 546574 223294
rect 545954 187614 546574 223058
rect 545954 187378 545986 187614
rect 546222 187378 546306 187614
rect 546542 187378 546574 187614
rect 545954 187294 546574 187378
rect 545954 187058 545986 187294
rect 546222 187058 546306 187294
rect 546542 187058 546574 187294
rect 545954 151614 546574 187058
rect 545954 151378 545986 151614
rect 546222 151378 546306 151614
rect 546542 151378 546574 151614
rect 545954 151294 546574 151378
rect 545954 151058 545986 151294
rect 546222 151058 546306 151294
rect 546542 151058 546574 151294
rect 545954 115614 546574 151058
rect 545954 115378 545986 115614
rect 546222 115378 546306 115614
rect 546542 115378 546574 115614
rect 545954 115294 546574 115378
rect 545954 115058 545986 115294
rect 546222 115058 546306 115294
rect 546542 115058 546574 115294
rect 545954 79614 546574 115058
rect 545954 79378 545986 79614
rect 546222 79378 546306 79614
rect 546542 79378 546574 79614
rect 545954 79294 546574 79378
rect 545954 79058 545986 79294
rect 546222 79058 546306 79294
rect 546542 79058 546574 79294
rect 545954 43614 546574 79058
rect 545954 43378 545986 43614
rect 546222 43378 546306 43614
rect 546542 43378 546574 43614
rect 545954 43294 546574 43378
rect 545954 43058 545986 43294
rect 546222 43058 546306 43294
rect 546542 43058 546574 43294
rect 545954 7614 546574 43058
rect 545954 7378 545986 7614
rect 546222 7378 546306 7614
rect 546542 7378 546574 7614
rect 545954 7294 546574 7378
rect 545954 7058 545986 7294
rect 546222 7058 546306 7294
rect 546542 7058 546574 7294
rect 545954 -4186 546574 7058
rect 545954 -4422 545986 -4186
rect 546222 -4422 546306 -4186
rect 546542 -4422 546574 -4186
rect 545954 -4506 546574 -4422
rect 545954 -4742 545986 -4506
rect 546222 -4742 546306 -4506
rect 546542 -4742 546574 -4506
rect 545954 -7654 546574 -4742
rect 547194 260854 547814 296298
rect 547194 260618 547226 260854
rect 547462 260618 547546 260854
rect 547782 260618 547814 260854
rect 547194 260534 547814 260618
rect 547194 260298 547226 260534
rect 547462 260298 547546 260534
rect 547782 260298 547814 260534
rect 547194 224854 547814 260298
rect 547194 224618 547226 224854
rect 547462 224618 547546 224854
rect 547782 224618 547814 224854
rect 547194 224534 547814 224618
rect 547194 224298 547226 224534
rect 547462 224298 547546 224534
rect 547782 224298 547814 224534
rect 547194 188854 547814 224298
rect 547194 188618 547226 188854
rect 547462 188618 547546 188854
rect 547782 188618 547814 188854
rect 547194 188534 547814 188618
rect 547194 188298 547226 188534
rect 547462 188298 547546 188534
rect 547782 188298 547814 188534
rect 547194 152854 547814 188298
rect 547194 152618 547226 152854
rect 547462 152618 547546 152854
rect 547782 152618 547814 152854
rect 547194 152534 547814 152618
rect 547194 152298 547226 152534
rect 547462 152298 547546 152534
rect 547782 152298 547814 152534
rect 547194 116854 547814 152298
rect 547194 116618 547226 116854
rect 547462 116618 547546 116854
rect 547782 116618 547814 116854
rect 547194 116534 547814 116618
rect 547194 116298 547226 116534
rect 547462 116298 547546 116534
rect 547782 116298 547814 116534
rect 547194 80854 547814 116298
rect 547194 80618 547226 80854
rect 547462 80618 547546 80854
rect 547782 80618 547814 80854
rect 547194 80534 547814 80618
rect 547194 80298 547226 80534
rect 547462 80298 547546 80534
rect 547782 80298 547814 80534
rect 547194 44854 547814 80298
rect 547194 44618 547226 44854
rect 547462 44618 547546 44854
rect 547782 44618 547814 44854
rect 547194 44534 547814 44618
rect 547194 44298 547226 44534
rect 547462 44298 547546 44534
rect 547782 44298 547814 44534
rect 547194 8854 547814 44298
rect 547194 8618 547226 8854
rect 547462 8618 547546 8854
rect 547782 8618 547814 8854
rect 547194 8534 547814 8618
rect 547194 8298 547226 8534
rect 547462 8298 547546 8534
rect 547782 8298 547814 8534
rect 547194 -5146 547814 8298
rect 547194 -5382 547226 -5146
rect 547462 -5382 547546 -5146
rect 547782 -5382 547814 -5146
rect 547194 -5466 547814 -5382
rect 547194 -5702 547226 -5466
rect 547462 -5702 547546 -5466
rect 547782 -5702 547814 -5466
rect 547194 -7654 547814 -5702
rect 548434 710598 549054 711590
rect 548434 710362 548466 710598
rect 548702 710362 548786 710598
rect 549022 710362 549054 710598
rect 548434 710278 549054 710362
rect 548434 710042 548466 710278
rect 548702 710042 548786 710278
rect 549022 710042 549054 710278
rect 548434 694094 549054 710042
rect 548434 693858 548466 694094
rect 548702 693858 548786 694094
rect 549022 693858 549054 694094
rect 548434 693774 549054 693858
rect 548434 693538 548466 693774
rect 548702 693538 548786 693774
rect 549022 693538 549054 693774
rect 548434 658094 549054 693538
rect 548434 657858 548466 658094
rect 548702 657858 548786 658094
rect 549022 657858 549054 658094
rect 548434 657774 549054 657858
rect 548434 657538 548466 657774
rect 548702 657538 548786 657774
rect 549022 657538 549054 657774
rect 548434 622094 549054 657538
rect 548434 621858 548466 622094
rect 548702 621858 548786 622094
rect 549022 621858 549054 622094
rect 548434 621774 549054 621858
rect 548434 621538 548466 621774
rect 548702 621538 548786 621774
rect 549022 621538 549054 621774
rect 548434 586094 549054 621538
rect 548434 585858 548466 586094
rect 548702 585858 548786 586094
rect 549022 585858 549054 586094
rect 548434 585774 549054 585858
rect 548434 585538 548466 585774
rect 548702 585538 548786 585774
rect 549022 585538 549054 585774
rect 548434 550094 549054 585538
rect 548434 549858 548466 550094
rect 548702 549858 548786 550094
rect 549022 549858 549054 550094
rect 548434 549774 549054 549858
rect 548434 549538 548466 549774
rect 548702 549538 548786 549774
rect 549022 549538 549054 549774
rect 548434 514094 549054 549538
rect 548434 513858 548466 514094
rect 548702 513858 548786 514094
rect 549022 513858 549054 514094
rect 548434 513774 549054 513858
rect 548434 513538 548466 513774
rect 548702 513538 548786 513774
rect 549022 513538 549054 513774
rect 548434 478094 549054 513538
rect 548434 477858 548466 478094
rect 548702 477858 548786 478094
rect 549022 477858 549054 478094
rect 548434 477774 549054 477858
rect 548434 477538 548466 477774
rect 548702 477538 548786 477774
rect 549022 477538 549054 477774
rect 548434 442094 549054 477538
rect 548434 441858 548466 442094
rect 548702 441858 548786 442094
rect 549022 441858 549054 442094
rect 548434 441774 549054 441858
rect 548434 441538 548466 441774
rect 548702 441538 548786 441774
rect 549022 441538 549054 441774
rect 548434 406094 549054 441538
rect 549674 711558 550294 711590
rect 549674 711322 549706 711558
rect 549942 711322 550026 711558
rect 550262 711322 550294 711558
rect 549674 711238 550294 711322
rect 549674 711002 549706 711238
rect 549942 711002 550026 711238
rect 550262 711002 550294 711238
rect 549674 695334 550294 711002
rect 549674 695098 549706 695334
rect 549942 695098 550026 695334
rect 550262 695098 550294 695334
rect 549674 695014 550294 695098
rect 549674 694778 549706 695014
rect 549942 694778 550026 695014
rect 550262 694778 550294 695014
rect 549674 659334 550294 694778
rect 549674 659098 549706 659334
rect 549942 659098 550026 659334
rect 550262 659098 550294 659334
rect 549674 659014 550294 659098
rect 549674 658778 549706 659014
rect 549942 658778 550026 659014
rect 550262 658778 550294 659014
rect 549674 623334 550294 658778
rect 549674 623098 549706 623334
rect 549942 623098 550026 623334
rect 550262 623098 550294 623334
rect 549674 623014 550294 623098
rect 549674 622778 549706 623014
rect 549942 622778 550026 623014
rect 550262 622778 550294 623014
rect 549674 587334 550294 622778
rect 549674 587098 549706 587334
rect 549942 587098 550026 587334
rect 550262 587098 550294 587334
rect 549674 587014 550294 587098
rect 549674 586778 549706 587014
rect 549942 586778 550026 587014
rect 550262 586778 550294 587014
rect 549674 551334 550294 586778
rect 549674 551098 549706 551334
rect 549942 551098 550026 551334
rect 550262 551098 550294 551334
rect 549674 551014 550294 551098
rect 549674 550778 549706 551014
rect 549942 550778 550026 551014
rect 550262 550778 550294 551014
rect 549674 515334 550294 550778
rect 549674 515098 549706 515334
rect 549942 515098 550026 515334
rect 550262 515098 550294 515334
rect 549674 515014 550294 515098
rect 549674 514778 549706 515014
rect 549942 514778 550026 515014
rect 550262 514778 550294 515014
rect 549674 479334 550294 514778
rect 549674 479098 549706 479334
rect 549942 479098 550026 479334
rect 550262 479098 550294 479334
rect 549674 479014 550294 479098
rect 549674 478778 549706 479014
rect 549942 478778 550026 479014
rect 550262 478778 550294 479014
rect 549674 443334 550294 478778
rect 549674 443098 549706 443334
rect 549942 443098 550026 443334
rect 550262 443098 550294 443334
rect 549674 443014 550294 443098
rect 549674 442778 549706 443014
rect 549942 442778 550026 443014
rect 550262 442778 550294 443014
rect 549299 434756 549365 434757
rect 549299 434692 549300 434756
rect 549364 434692 549365 434756
rect 549299 434691 549365 434692
rect 548434 405858 548466 406094
rect 548702 405858 548786 406094
rect 549022 405858 549054 406094
rect 548434 405774 549054 405858
rect 548434 405538 548466 405774
rect 548702 405538 548786 405774
rect 549022 405538 549054 405774
rect 548434 370094 549054 405538
rect 549302 398309 549362 434691
rect 549674 407334 550294 442778
rect 549674 407098 549706 407334
rect 549942 407098 550026 407334
rect 550262 407098 550294 407334
rect 549674 407014 550294 407098
rect 549674 406778 549706 407014
rect 549942 406778 550026 407014
rect 550262 406778 550294 407014
rect 549299 398308 549365 398309
rect 549299 398244 549300 398308
rect 549364 398244 549365 398308
rect 549299 398243 549365 398244
rect 548434 369858 548466 370094
rect 548702 369858 548786 370094
rect 549022 369858 549054 370094
rect 548434 369774 549054 369858
rect 548434 369538 548466 369774
rect 548702 369538 548786 369774
rect 549022 369538 549054 369774
rect 548434 334094 549054 369538
rect 549302 362813 549362 398243
rect 549674 371334 550294 406778
rect 549674 371098 549706 371334
rect 549942 371098 550026 371334
rect 550262 371098 550294 371334
rect 549674 371014 550294 371098
rect 549674 370778 549706 371014
rect 549942 370778 550026 371014
rect 550262 370778 550294 371014
rect 549299 362812 549365 362813
rect 549299 362748 549300 362812
rect 549364 362748 549365 362812
rect 549299 362747 549365 362748
rect 548434 333858 548466 334094
rect 548702 333858 548786 334094
rect 549022 333858 549054 334094
rect 548434 333774 549054 333858
rect 548434 333538 548466 333774
rect 548702 333538 548786 333774
rect 549022 333538 549054 333774
rect 548434 298094 549054 333538
rect 549302 326773 549362 362747
rect 549674 335334 550294 370778
rect 549674 335098 549706 335334
rect 549942 335098 550026 335334
rect 550262 335098 550294 335334
rect 549674 335014 550294 335098
rect 549674 334778 549706 335014
rect 549942 334778 550026 335014
rect 550262 334778 550294 335014
rect 549299 326772 549365 326773
rect 549299 326708 549300 326772
rect 549364 326708 549365 326772
rect 549299 326707 549365 326708
rect 548434 297858 548466 298094
rect 548702 297858 548786 298094
rect 549022 297858 549054 298094
rect 548434 297774 549054 297858
rect 548434 297538 548466 297774
rect 548702 297538 548786 297774
rect 549022 297538 549054 297774
rect 548434 262094 549054 297538
rect 549302 290733 549362 326707
rect 549674 299334 550294 334778
rect 549674 299098 549706 299334
rect 549942 299098 550026 299334
rect 550262 299098 550294 299334
rect 549674 299014 550294 299098
rect 549674 298778 549706 299014
rect 549942 298778 550026 299014
rect 550262 298778 550294 299014
rect 549299 290732 549365 290733
rect 549299 290668 549300 290732
rect 549364 290668 549365 290732
rect 549299 290667 549365 290668
rect 548434 261858 548466 262094
rect 548702 261858 548786 262094
rect 549022 261858 549054 262094
rect 548434 261774 549054 261858
rect 548434 261538 548466 261774
rect 548702 261538 548786 261774
rect 549022 261538 549054 261774
rect 548434 226094 549054 261538
rect 548434 225858 548466 226094
rect 548702 225858 548786 226094
rect 549022 225858 549054 226094
rect 548434 225774 549054 225858
rect 548434 225538 548466 225774
rect 548702 225538 548786 225774
rect 549022 225538 549054 225774
rect 548434 190094 549054 225538
rect 548434 189858 548466 190094
rect 548702 189858 548786 190094
rect 549022 189858 549054 190094
rect 548434 189774 549054 189858
rect 548434 189538 548466 189774
rect 548702 189538 548786 189774
rect 549022 189538 549054 189774
rect 548434 154094 549054 189538
rect 548434 153858 548466 154094
rect 548702 153858 548786 154094
rect 549022 153858 549054 154094
rect 548434 153774 549054 153858
rect 548434 153538 548466 153774
rect 548702 153538 548786 153774
rect 549022 153538 549054 153774
rect 548434 118094 549054 153538
rect 548434 117858 548466 118094
rect 548702 117858 548786 118094
rect 549022 117858 549054 118094
rect 548434 117774 549054 117858
rect 548434 117538 548466 117774
rect 548702 117538 548786 117774
rect 549022 117538 549054 117774
rect 548434 82094 549054 117538
rect 548434 81858 548466 82094
rect 548702 81858 548786 82094
rect 549022 81858 549054 82094
rect 548434 81774 549054 81858
rect 548434 81538 548466 81774
rect 548702 81538 548786 81774
rect 549022 81538 549054 81774
rect 548434 46094 549054 81538
rect 548434 45858 548466 46094
rect 548702 45858 548786 46094
rect 549022 45858 549054 46094
rect 548434 45774 549054 45858
rect 548434 45538 548466 45774
rect 548702 45538 548786 45774
rect 549022 45538 549054 45774
rect 548434 10094 549054 45538
rect 549302 19821 549362 290667
rect 549674 263334 550294 298778
rect 549674 263098 549706 263334
rect 549942 263098 550026 263334
rect 550262 263098 550294 263334
rect 549674 263014 550294 263098
rect 549674 262778 549706 263014
rect 549942 262778 550026 263014
rect 550262 262778 550294 263014
rect 549674 227334 550294 262778
rect 549674 227098 549706 227334
rect 549942 227098 550026 227334
rect 550262 227098 550294 227334
rect 549674 227014 550294 227098
rect 549674 226778 549706 227014
rect 549942 226778 550026 227014
rect 550262 226778 550294 227014
rect 549674 191334 550294 226778
rect 549674 191098 549706 191334
rect 549942 191098 550026 191334
rect 550262 191098 550294 191334
rect 549674 191014 550294 191098
rect 549674 190778 549706 191014
rect 549942 190778 550026 191014
rect 550262 190778 550294 191014
rect 549674 155334 550294 190778
rect 549674 155098 549706 155334
rect 549942 155098 550026 155334
rect 550262 155098 550294 155334
rect 549674 155014 550294 155098
rect 549674 154778 549706 155014
rect 549942 154778 550026 155014
rect 550262 154778 550294 155014
rect 549674 119334 550294 154778
rect 549674 119098 549706 119334
rect 549942 119098 550026 119334
rect 550262 119098 550294 119334
rect 549674 119014 550294 119098
rect 549674 118778 549706 119014
rect 549942 118778 550026 119014
rect 550262 118778 550294 119014
rect 549674 83334 550294 118778
rect 549674 83098 549706 83334
rect 549942 83098 550026 83334
rect 550262 83098 550294 83334
rect 549674 83014 550294 83098
rect 549674 82778 549706 83014
rect 549942 82778 550026 83014
rect 550262 82778 550294 83014
rect 549674 47334 550294 82778
rect 549674 47098 549706 47334
rect 549942 47098 550026 47334
rect 550262 47098 550294 47334
rect 549674 47014 550294 47098
rect 549674 46778 549706 47014
rect 549942 46778 550026 47014
rect 550262 46778 550294 47014
rect 549299 19820 549365 19821
rect 549299 19756 549300 19820
rect 549364 19756 549365 19820
rect 549299 19755 549365 19756
rect 548434 9858 548466 10094
rect 548702 9858 548786 10094
rect 549022 9858 549054 10094
rect 548434 9774 549054 9858
rect 548434 9538 548466 9774
rect 548702 9538 548786 9774
rect 549022 9538 549054 9774
rect 548434 -6106 549054 9538
rect 548434 -6342 548466 -6106
rect 548702 -6342 548786 -6106
rect 549022 -6342 549054 -6106
rect 548434 -6426 549054 -6342
rect 548434 -6662 548466 -6426
rect 548702 -6662 548786 -6426
rect 549022 -6662 549054 -6426
rect 548434 -7654 549054 -6662
rect 549674 11334 550294 46778
rect 549674 11098 549706 11334
rect 549942 11098 550026 11334
rect 550262 11098 550294 11334
rect 549674 11014 550294 11098
rect 549674 10778 549706 11014
rect 549942 10778 550026 11014
rect 550262 10778 550294 11014
rect 549674 -7066 550294 10778
rect 549674 -7302 549706 -7066
rect 549942 -7302 550026 -7066
rect 550262 -7302 550294 -7066
rect 549674 -7386 550294 -7302
rect 549674 -7622 549706 -7386
rect 549942 -7622 550026 -7386
rect 550262 -7622 550294 -7386
rect 549674 -7654 550294 -7622
rect 576994 704838 577614 711590
rect 576994 704602 577026 704838
rect 577262 704602 577346 704838
rect 577582 704602 577614 704838
rect 576994 704518 577614 704602
rect 576994 704282 577026 704518
rect 577262 704282 577346 704518
rect 577582 704282 577614 704518
rect 576994 686654 577614 704282
rect 576994 686418 577026 686654
rect 577262 686418 577346 686654
rect 577582 686418 577614 686654
rect 576994 686334 577614 686418
rect 576994 686098 577026 686334
rect 577262 686098 577346 686334
rect 577582 686098 577614 686334
rect 576994 650654 577614 686098
rect 576994 650418 577026 650654
rect 577262 650418 577346 650654
rect 577582 650418 577614 650654
rect 576994 650334 577614 650418
rect 576994 650098 577026 650334
rect 577262 650098 577346 650334
rect 577582 650098 577614 650334
rect 576994 614654 577614 650098
rect 576994 614418 577026 614654
rect 577262 614418 577346 614654
rect 577582 614418 577614 614654
rect 576994 614334 577614 614418
rect 576994 614098 577026 614334
rect 577262 614098 577346 614334
rect 577582 614098 577614 614334
rect 576994 578654 577614 614098
rect 576994 578418 577026 578654
rect 577262 578418 577346 578654
rect 577582 578418 577614 578654
rect 576994 578334 577614 578418
rect 576994 578098 577026 578334
rect 577262 578098 577346 578334
rect 577582 578098 577614 578334
rect 576994 542654 577614 578098
rect 576994 542418 577026 542654
rect 577262 542418 577346 542654
rect 577582 542418 577614 542654
rect 576994 542334 577614 542418
rect 576994 542098 577026 542334
rect 577262 542098 577346 542334
rect 577582 542098 577614 542334
rect 576994 506654 577614 542098
rect 576994 506418 577026 506654
rect 577262 506418 577346 506654
rect 577582 506418 577614 506654
rect 576994 506334 577614 506418
rect 576994 506098 577026 506334
rect 577262 506098 577346 506334
rect 577582 506098 577614 506334
rect 576994 470654 577614 506098
rect 576994 470418 577026 470654
rect 577262 470418 577346 470654
rect 577582 470418 577614 470654
rect 576994 470334 577614 470418
rect 576994 470098 577026 470334
rect 577262 470098 577346 470334
rect 577582 470098 577614 470334
rect 576994 434654 577614 470098
rect 576994 434418 577026 434654
rect 577262 434418 577346 434654
rect 577582 434418 577614 434654
rect 576994 434334 577614 434418
rect 576994 434098 577026 434334
rect 577262 434098 577346 434334
rect 577582 434098 577614 434334
rect 576994 398654 577614 434098
rect 576994 398418 577026 398654
rect 577262 398418 577346 398654
rect 577582 398418 577614 398654
rect 576994 398334 577614 398418
rect 576994 398098 577026 398334
rect 577262 398098 577346 398334
rect 577582 398098 577614 398334
rect 576994 362654 577614 398098
rect 576994 362418 577026 362654
rect 577262 362418 577346 362654
rect 577582 362418 577614 362654
rect 576994 362334 577614 362418
rect 576994 362098 577026 362334
rect 577262 362098 577346 362334
rect 577582 362098 577614 362334
rect 576994 326654 577614 362098
rect 576994 326418 577026 326654
rect 577262 326418 577346 326654
rect 577582 326418 577614 326654
rect 576994 326334 577614 326418
rect 576994 326098 577026 326334
rect 577262 326098 577346 326334
rect 577582 326098 577614 326334
rect 576994 290654 577614 326098
rect 576994 290418 577026 290654
rect 577262 290418 577346 290654
rect 577582 290418 577614 290654
rect 576994 290334 577614 290418
rect 576994 290098 577026 290334
rect 577262 290098 577346 290334
rect 577582 290098 577614 290334
rect 576994 254654 577614 290098
rect 576994 254418 577026 254654
rect 577262 254418 577346 254654
rect 577582 254418 577614 254654
rect 576994 254334 577614 254418
rect 576994 254098 577026 254334
rect 577262 254098 577346 254334
rect 577582 254098 577614 254334
rect 576994 218654 577614 254098
rect 576994 218418 577026 218654
rect 577262 218418 577346 218654
rect 577582 218418 577614 218654
rect 576994 218334 577614 218418
rect 576994 218098 577026 218334
rect 577262 218098 577346 218334
rect 577582 218098 577614 218334
rect 576994 182654 577614 218098
rect 576994 182418 577026 182654
rect 577262 182418 577346 182654
rect 577582 182418 577614 182654
rect 576994 182334 577614 182418
rect 576994 182098 577026 182334
rect 577262 182098 577346 182334
rect 577582 182098 577614 182334
rect 576994 146654 577614 182098
rect 576994 146418 577026 146654
rect 577262 146418 577346 146654
rect 577582 146418 577614 146654
rect 576994 146334 577614 146418
rect 576994 146098 577026 146334
rect 577262 146098 577346 146334
rect 577582 146098 577614 146334
rect 576994 110654 577614 146098
rect 576994 110418 577026 110654
rect 577262 110418 577346 110654
rect 577582 110418 577614 110654
rect 576994 110334 577614 110418
rect 576994 110098 577026 110334
rect 577262 110098 577346 110334
rect 577582 110098 577614 110334
rect 576994 74654 577614 110098
rect 576994 74418 577026 74654
rect 577262 74418 577346 74654
rect 577582 74418 577614 74654
rect 576994 74334 577614 74418
rect 576994 74098 577026 74334
rect 577262 74098 577346 74334
rect 577582 74098 577614 74334
rect 576994 38654 577614 74098
rect 576994 38418 577026 38654
rect 577262 38418 577346 38654
rect 577582 38418 577614 38654
rect 576994 38334 577614 38418
rect 576994 38098 577026 38334
rect 577262 38098 577346 38334
rect 577582 38098 577614 38334
rect 576994 2654 577614 38098
rect 576994 2418 577026 2654
rect 577262 2418 577346 2654
rect 577582 2418 577614 2654
rect 576994 2334 577614 2418
rect 576994 2098 577026 2334
rect 577262 2098 577346 2334
rect 577582 2098 577614 2334
rect 576994 -346 577614 2098
rect 576994 -582 577026 -346
rect 577262 -582 577346 -346
rect 577582 -582 577614 -346
rect 576994 -666 577614 -582
rect 576994 -902 577026 -666
rect 577262 -902 577346 -666
rect 577582 -902 577614 -666
rect 576994 -7654 577614 -902
rect 578234 705798 578854 711590
rect 578234 705562 578266 705798
rect 578502 705562 578586 705798
rect 578822 705562 578854 705798
rect 578234 705478 578854 705562
rect 578234 705242 578266 705478
rect 578502 705242 578586 705478
rect 578822 705242 578854 705478
rect 578234 687894 578854 705242
rect 578234 687658 578266 687894
rect 578502 687658 578586 687894
rect 578822 687658 578854 687894
rect 578234 687574 578854 687658
rect 578234 687338 578266 687574
rect 578502 687338 578586 687574
rect 578822 687338 578854 687574
rect 578234 651894 578854 687338
rect 578234 651658 578266 651894
rect 578502 651658 578586 651894
rect 578822 651658 578854 651894
rect 578234 651574 578854 651658
rect 578234 651338 578266 651574
rect 578502 651338 578586 651574
rect 578822 651338 578854 651574
rect 578234 615894 578854 651338
rect 578234 615658 578266 615894
rect 578502 615658 578586 615894
rect 578822 615658 578854 615894
rect 578234 615574 578854 615658
rect 578234 615338 578266 615574
rect 578502 615338 578586 615574
rect 578822 615338 578854 615574
rect 578234 579894 578854 615338
rect 578234 579658 578266 579894
rect 578502 579658 578586 579894
rect 578822 579658 578854 579894
rect 578234 579574 578854 579658
rect 578234 579338 578266 579574
rect 578502 579338 578586 579574
rect 578822 579338 578854 579574
rect 578234 543894 578854 579338
rect 578234 543658 578266 543894
rect 578502 543658 578586 543894
rect 578822 543658 578854 543894
rect 578234 543574 578854 543658
rect 578234 543338 578266 543574
rect 578502 543338 578586 543574
rect 578822 543338 578854 543574
rect 578234 507894 578854 543338
rect 578234 507658 578266 507894
rect 578502 507658 578586 507894
rect 578822 507658 578854 507894
rect 578234 507574 578854 507658
rect 578234 507338 578266 507574
rect 578502 507338 578586 507574
rect 578822 507338 578854 507574
rect 578234 471894 578854 507338
rect 578234 471658 578266 471894
rect 578502 471658 578586 471894
rect 578822 471658 578854 471894
rect 578234 471574 578854 471658
rect 578234 471338 578266 471574
rect 578502 471338 578586 471574
rect 578822 471338 578854 471574
rect 578234 435894 578854 471338
rect 578234 435658 578266 435894
rect 578502 435658 578586 435894
rect 578822 435658 578854 435894
rect 578234 435574 578854 435658
rect 578234 435338 578266 435574
rect 578502 435338 578586 435574
rect 578822 435338 578854 435574
rect 578234 399894 578854 435338
rect 578234 399658 578266 399894
rect 578502 399658 578586 399894
rect 578822 399658 578854 399894
rect 578234 399574 578854 399658
rect 578234 399338 578266 399574
rect 578502 399338 578586 399574
rect 578822 399338 578854 399574
rect 578234 363894 578854 399338
rect 578234 363658 578266 363894
rect 578502 363658 578586 363894
rect 578822 363658 578854 363894
rect 578234 363574 578854 363658
rect 578234 363338 578266 363574
rect 578502 363338 578586 363574
rect 578822 363338 578854 363574
rect 578234 327894 578854 363338
rect 578234 327658 578266 327894
rect 578502 327658 578586 327894
rect 578822 327658 578854 327894
rect 578234 327574 578854 327658
rect 578234 327338 578266 327574
rect 578502 327338 578586 327574
rect 578822 327338 578854 327574
rect 578234 291894 578854 327338
rect 578234 291658 578266 291894
rect 578502 291658 578586 291894
rect 578822 291658 578854 291894
rect 578234 291574 578854 291658
rect 578234 291338 578266 291574
rect 578502 291338 578586 291574
rect 578822 291338 578854 291574
rect 578234 255894 578854 291338
rect 578234 255658 578266 255894
rect 578502 255658 578586 255894
rect 578822 255658 578854 255894
rect 578234 255574 578854 255658
rect 578234 255338 578266 255574
rect 578502 255338 578586 255574
rect 578822 255338 578854 255574
rect 578234 219894 578854 255338
rect 578234 219658 578266 219894
rect 578502 219658 578586 219894
rect 578822 219658 578854 219894
rect 578234 219574 578854 219658
rect 578234 219338 578266 219574
rect 578502 219338 578586 219574
rect 578822 219338 578854 219574
rect 578234 183894 578854 219338
rect 578234 183658 578266 183894
rect 578502 183658 578586 183894
rect 578822 183658 578854 183894
rect 578234 183574 578854 183658
rect 578234 183338 578266 183574
rect 578502 183338 578586 183574
rect 578822 183338 578854 183574
rect 578234 147894 578854 183338
rect 578234 147658 578266 147894
rect 578502 147658 578586 147894
rect 578822 147658 578854 147894
rect 578234 147574 578854 147658
rect 578234 147338 578266 147574
rect 578502 147338 578586 147574
rect 578822 147338 578854 147574
rect 578234 111894 578854 147338
rect 578234 111658 578266 111894
rect 578502 111658 578586 111894
rect 578822 111658 578854 111894
rect 578234 111574 578854 111658
rect 578234 111338 578266 111574
rect 578502 111338 578586 111574
rect 578822 111338 578854 111574
rect 578234 75894 578854 111338
rect 578234 75658 578266 75894
rect 578502 75658 578586 75894
rect 578822 75658 578854 75894
rect 578234 75574 578854 75658
rect 578234 75338 578266 75574
rect 578502 75338 578586 75574
rect 578822 75338 578854 75574
rect 578234 39894 578854 75338
rect 578234 39658 578266 39894
rect 578502 39658 578586 39894
rect 578822 39658 578854 39894
rect 578234 39574 578854 39658
rect 578234 39338 578266 39574
rect 578502 39338 578586 39574
rect 578822 39338 578854 39574
rect 578234 3894 578854 39338
rect 578234 3658 578266 3894
rect 578502 3658 578586 3894
rect 578822 3658 578854 3894
rect 578234 3574 578854 3658
rect 578234 3338 578266 3574
rect 578502 3338 578586 3574
rect 578822 3338 578854 3574
rect 578234 -1306 578854 3338
rect 578234 -1542 578266 -1306
rect 578502 -1542 578586 -1306
rect 578822 -1542 578854 -1306
rect 578234 -1626 578854 -1542
rect 578234 -1862 578266 -1626
rect 578502 -1862 578586 -1626
rect 578822 -1862 578854 -1626
rect 578234 -7654 578854 -1862
rect 579474 706758 580094 711590
rect 579474 706522 579506 706758
rect 579742 706522 579826 706758
rect 580062 706522 580094 706758
rect 579474 706438 580094 706522
rect 579474 706202 579506 706438
rect 579742 706202 579826 706438
rect 580062 706202 580094 706438
rect 579474 689134 580094 706202
rect 579474 688898 579506 689134
rect 579742 688898 579826 689134
rect 580062 688898 580094 689134
rect 579474 688814 580094 688898
rect 579474 688578 579506 688814
rect 579742 688578 579826 688814
rect 580062 688578 580094 688814
rect 579474 653134 580094 688578
rect 579474 652898 579506 653134
rect 579742 652898 579826 653134
rect 580062 652898 580094 653134
rect 579474 652814 580094 652898
rect 579474 652578 579506 652814
rect 579742 652578 579826 652814
rect 580062 652578 580094 652814
rect 579474 617134 580094 652578
rect 579474 616898 579506 617134
rect 579742 616898 579826 617134
rect 580062 616898 580094 617134
rect 579474 616814 580094 616898
rect 579474 616578 579506 616814
rect 579742 616578 579826 616814
rect 580062 616578 580094 616814
rect 579474 581134 580094 616578
rect 579474 580898 579506 581134
rect 579742 580898 579826 581134
rect 580062 580898 580094 581134
rect 579474 580814 580094 580898
rect 579474 580578 579506 580814
rect 579742 580578 579826 580814
rect 580062 580578 580094 580814
rect 579474 545134 580094 580578
rect 579474 544898 579506 545134
rect 579742 544898 579826 545134
rect 580062 544898 580094 545134
rect 579474 544814 580094 544898
rect 579474 544578 579506 544814
rect 579742 544578 579826 544814
rect 580062 544578 580094 544814
rect 579474 509134 580094 544578
rect 579474 508898 579506 509134
rect 579742 508898 579826 509134
rect 580062 508898 580094 509134
rect 579474 508814 580094 508898
rect 579474 508578 579506 508814
rect 579742 508578 579826 508814
rect 580062 508578 580094 508814
rect 579474 473134 580094 508578
rect 579474 472898 579506 473134
rect 579742 472898 579826 473134
rect 580062 472898 580094 473134
rect 579474 472814 580094 472898
rect 579474 472578 579506 472814
rect 579742 472578 579826 472814
rect 580062 472578 580094 472814
rect 579474 437134 580094 472578
rect 579474 436898 579506 437134
rect 579742 436898 579826 437134
rect 580062 436898 580094 437134
rect 579474 436814 580094 436898
rect 579474 436578 579506 436814
rect 579742 436578 579826 436814
rect 580062 436578 580094 436814
rect 579474 401134 580094 436578
rect 579474 400898 579506 401134
rect 579742 400898 579826 401134
rect 580062 400898 580094 401134
rect 579474 400814 580094 400898
rect 579474 400578 579506 400814
rect 579742 400578 579826 400814
rect 580062 400578 580094 400814
rect 579474 365134 580094 400578
rect 579474 364898 579506 365134
rect 579742 364898 579826 365134
rect 580062 364898 580094 365134
rect 579474 364814 580094 364898
rect 579474 364578 579506 364814
rect 579742 364578 579826 364814
rect 580062 364578 580094 364814
rect 579474 329134 580094 364578
rect 579474 328898 579506 329134
rect 579742 328898 579826 329134
rect 580062 328898 580094 329134
rect 579474 328814 580094 328898
rect 579474 328578 579506 328814
rect 579742 328578 579826 328814
rect 580062 328578 580094 328814
rect 579474 293134 580094 328578
rect 579474 292898 579506 293134
rect 579742 292898 579826 293134
rect 580062 292898 580094 293134
rect 579474 292814 580094 292898
rect 579474 292578 579506 292814
rect 579742 292578 579826 292814
rect 580062 292578 580094 292814
rect 579474 257134 580094 292578
rect 579474 256898 579506 257134
rect 579742 256898 579826 257134
rect 580062 256898 580094 257134
rect 579474 256814 580094 256898
rect 579474 256578 579506 256814
rect 579742 256578 579826 256814
rect 580062 256578 580094 256814
rect 579474 221134 580094 256578
rect 579474 220898 579506 221134
rect 579742 220898 579826 221134
rect 580062 220898 580094 221134
rect 579474 220814 580094 220898
rect 579474 220578 579506 220814
rect 579742 220578 579826 220814
rect 580062 220578 580094 220814
rect 579474 185134 580094 220578
rect 579474 184898 579506 185134
rect 579742 184898 579826 185134
rect 580062 184898 580094 185134
rect 579474 184814 580094 184898
rect 579474 184578 579506 184814
rect 579742 184578 579826 184814
rect 580062 184578 580094 184814
rect 579474 149134 580094 184578
rect 579474 148898 579506 149134
rect 579742 148898 579826 149134
rect 580062 148898 580094 149134
rect 579474 148814 580094 148898
rect 579474 148578 579506 148814
rect 579742 148578 579826 148814
rect 580062 148578 580094 148814
rect 579474 113134 580094 148578
rect 579474 112898 579506 113134
rect 579742 112898 579826 113134
rect 580062 112898 580094 113134
rect 579474 112814 580094 112898
rect 579474 112578 579506 112814
rect 579742 112578 579826 112814
rect 580062 112578 580094 112814
rect 579474 77134 580094 112578
rect 579474 76898 579506 77134
rect 579742 76898 579826 77134
rect 580062 76898 580094 77134
rect 579474 76814 580094 76898
rect 579474 76578 579506 76814
rect 579742 76578 579826 76814
rect 580062 76578 580094 76814
rect 579474 41134 580094 76578
rect 579474 40898 579506 41134
rect 579742 40898 579826 41134
rect 580062 40898 580094 41134
rect 579474 40814 580094 40898
rect 579474 40578 579506 40814
rect 579742 40578 579826 40814
rect 580062 40578 580094 40814
rect 579474 5134 580094 40578
rect 579474 4898 579506 5134
rect 579742 4898 579826 5134
rect 580062 4898 580094 5134
rect 579474 4814 580094 4898
rect 579474 4578 579506 4814
rect 579742 4578 579826 4814
rect 580062 4578 580094 4814
rect 579474 -2266 580094 4578
rect 579474 -2502 579506 -2266
rect 579742 -2502 579826 -2266
rect 580062 -2502 580094 -2266
rect 579474 -2586 580094 -2502
rect 579474 -2822 579506 -2586
rect 579742 -2822 579826 -2586
rect 580062 -2822 580094 -2586
rect 579474 -7654 580094 -2822
rect 580714 707718 581334 711590
rect 580714 707482 580746 707718
rect 580982 707482 581066 707718
rect 581302 707482 581334 707718
rect 580714 707398 581334 707482
rect 580714 707162 580746 707398
rect 580982 707162 581066 707398
rect 581302 707162 581334 707398
rect 580714 690374 581334 707162
rect 580714 690138 580746 690374
rect 580982 690138 581066 690374
rect 581302 690138 581334 690374
rect 580714 690054 581334 690138
rect 580714 689818 580746 690054
rect 580982 689818 581066 690054
rect 581302 689818 581334 690054
rect 580714 654374 581334 689818
rect 580714 654138 580746 654374
rect 580982 654138 581066 654374
rect 581302 654138 581334 654374
rect 580714 654054 581334 654138
rect 580714 653818 580746 654054
rect 580982 653818 581066 654054
rect 581302 653818 581334 654054
rect 580714 618374 581334 653818
rect 580714 618138 580746 618374
rect 580982 618138 581066 618374
rect 581302 618138 581334 618374
rect 580714 618054 581334 618138
rect 580714 617818 580746 618054
rect 580982 617818 581066 618054
rect 581302 617818 581334 618054
rect 580714 582374 581334 617818
rect 580714 582138 580746 582374
rect 580982 582138 581066 582374
rect 581302 582138 581334 582374
rect 580714 582054 581334 582138
rect 580714 581818 580746 582054
rect 580982 581818 581066 582054
rect 581302 581818 581334 582054
rect 580714 546374 581334 581818
rect 580714 546138 580746 546374
rect 580982 546138 581066 546374
rect 581302 546138 581334 546374
rect 580714 546054 581334 546138
rect 580714 545818 580746 546054
rect 580982 545818 581066 546054
rect 581302 545818 581334 546054
rect 580714 510374 581334 545818
rect 580714 510138 580746 510374
rect 580982 510138 581066 510374
rect 581302 510138 581334 510374
rect 580714 510054 581334 510138
rect 580714 509818 580746 510054
rect 580982 509818 581066 510054
rect 581302 509818 581334 510054
rect 580714 474374 581334 509818
rect 580714 474138 580746 474374
rect 580982 474138 581066 474374
rect 581302 474138 581334 474374
rect 580714 474054 581334 474138
rect 580714 473818 580746 474054
rect 580982 473818 581066 474054
rect 581302 473818 581334 474054
rect 580714 438374 581334 473818
rect 580714 438138 580746 438374
rect 580982 438138 581066 438374
rect 581302 438138 581334 438374
rect 580714 438054 581334 438138
rect 580714 437818 580746 438054
rect 580982 437818 581066 438054
rect 581302 437818 581334 438054
rect 580714 402374 581334 437818
rect 580714 402138 580746 402374
rect 580982 402138 581066 402374
rect 581302 402138 581334 402374
rect 580714 402054 581334 402138
rect 580714 401818 580746 402054
rect 580982 401818 581066 402054
rect 581302 401818 581334 402054
rect 580714 366374 581334 401818
rect 580714 366138 580746 366374
rect 580982 366138 581066 366374
rect 581302 366138 581334 366374
rect 580714 366054 581334 366138
rect 580714 365818 580746 366054
rect 580982 365818 581066 366054
rect 581302 365818 581334 366054
rect 580714 330374 581334 365818
rect 580714 330138 580746 330374
rect 580982 330138 581066 330374
rect 581302 330138 581334 330374
rect 580714 330054 581334 330138
rect 580714 329818 580746 330054
rect 580982 329818 581066 330054
rect 581302 329818 581334 330054
rect 580714 294374 581334 329818
rect 580714 294138 580746 294374
rect 580982 294138 581066 294374
rect 581302 294138 581334 294374
rect 580714 294054 581334 294138
rect 580714 293818 580746 294054
rect 580982 293818 581066 294054
rect 581302 293818 581334 294054
rect 580714 258374 581334 293818
rect 580714 258138 580746 258374
rect 580982 258138 581066 258374
rect 581302 258138 581334 258374
rect 580714 258054 581334 258138
rect 580714 257818 580746 258054
rect 580982 257818 581066 258054
rect 581302 257818 581334 258054
rect 580714 222374 581334 257818
rect 580714 222138 580746 222374
rect 580982 222138 581066 222374
rect 581302 222138 581334 222374
rect 580714 222054 581334 222138
rect 580714 221818 580746 222054
rect 580982 221818 581066 222054
rect 581302 221818 581334 222054
rect 580714 186374 581334 221818
rect 580714 186138 580746 186374
rect 580982 186138 581066 186374
rect 581302 186138 581334 186374
rect 580714 186054 581334 186138
rect 580714 185818 580746 186054
rect 580982 185818 581066 186054
rect 581302 185818 581334 186054
rect 580714 150374 581334 185818
rect 580714 150138 580746 150374
rect 580982 150138 581066 150374
rect 581302 150138 581334 150374
rect 580714 150054 581334 150138
rect 580714 149818 580746 150054
rect 580982 149818 581066 150054
rect 581302 149818 581334 150054
rect 580714 114374 581334 149818
rect 580714 114138 580746 114374
rect 580982 114138 581066 114374
rect 581302 114138 581334 114374
rect 580714 114054 581334 114138
rect 580714 113818 580746 114054
rect 580982 113818 581066 114054
rect 581302 113818 581334 114054
rect 580714 78374 581334 113818
rect 580714 78138 580746 78374
rect 580982 78138 581066 78374
rect 581302 78138 581334 78374
rect 580714 78054 581334 78138
rect 580714 77818 580746 78054
rect 580982 77818 581066 78054
rect 581302 77818 581334 78054
rect 580714 42374 581334 77818
rect 580714 42138 580746 42374
rect 580982 42138 581066 42374
rect 581302 42138 581334 42374
rect 580714 42054 581334 42138
rect 580714 41818 580746 42054
rect 580982 41818 581066 42054
rect 581302 41818 581334 42054
rect 580714 6374 581334 41818
rect 580714 6138 580746 6374
rect 580982 6138 581066 6374
rect 581302 6138 581334 6374
rect 580714 6054 581334 6138
rect 580714 5818 580746 6054
rect 580982 5818 581066 6054
rect 581302 5818 581334 6054
rect 580714 -3226 581334 5818
rect 580714 -3462 580746 -3226
rect 580982 -3462 581066 -3226
rect 581302 -3462 581334 -3226
rect 580714 -3546 581334 -3462
rect 580714 -3782 580746 -3546
rect 580982 -3782 581066 -3546
rect 581302 -3782 581334 -3546
rect 580714 -7654 581334 -3782
rect 581954 708678 582574 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 581954 708442 581986 708678
rect 582222 708442 582306 708678
rect 582542 708442 582574 708678
rect 581954 708358 582574 708442
rect 581954 708122 581986 708358
rect 582222 708122 582306 708358
rect 582542 708122 582574 708358
rect 581954 691614 582574 708122
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581954 691378 581986 691614
rect 582222 691378 582306 691614
rect 582542 691378 582574 691614
rect 581954 691294 582574 691378
rect 581954 691058 581986 691294
rect 582222 691058 582306 691294
rect 582542 691058 582574 691294
rect 581954 655614 582574 691058
rect 581954 655378 581986 655614
rect 582222 655378 582306 655614
rect 582542 655378 582574 655614
rect 581954 655294 582574 655378
rect 581954 655058 581986 655294
rect 582222 655058 582306 655294
rect 582542 655058 582574 655294
rect 581954 619614 582574 655058
rect 581954 619378 581986 619614
rect 582222 619378 582306 619614
rect 582542 619378 582574 619614
rect 581954 619294 582574 619378
rect 581954 619058 581986 619294
rect 582222 619058 582306 619294
rect 582542 619058 582574 619294
rect 581954 583614 582574 619058
rect 581954 583378 581986 583614
rect 582222 583378 582306 583614
rect 582542 583378 582574 583614
rect 581954 583294 582574 583378
rect 581954 583058 581986 583294
rect 582222 583058 582306 583294
rect 582542 583058 582574 583294
rect 581954 547614 582574 583058
rect 581954 547378 581986 547614
rect 582222 547378 582306 547614
rect 582542 547378 582574 547614
rect 581954 547294 582574 547378
rect 581954 547058 581986 547294
rect 582222 547058 582306 547294
rect 582542 547058 582574 547294
rect 581954 511614 582574 547058
rect 581954 511378 581986 511614
rect 582222 511378 582306 511614
rect 582542 511378 582574 511614
rect 581954 511294 582574 511378
rect 581954 511058 581986 511294
rect 582222 511058 582306 511294
rect 582542 511058 582574 511294
rect 581954 475614 582574 511058
rect 581954 475378 581986 475614
rect 582222 475378 582306 475614
rect 582542 475378 582574 475614
rect 581954 475294 582574 475378
rect 581954 475058 581986 475294
rect 582222 475058 582306 475294
rect 582542 475058 582574 475294
rect 581954 439614 582574 475058
rect 581954 439378 581986 439614
rect 582222 439378 582306 439614
rect 582542 439378 582574 439614
rect 581954 439294 582574 439378
rect 581954 439058 581986 439294
rect 582222 439058 582306 439294
rect 582542 439058 582574 439294
rect 581954 403614 582574 439058
rect 581954 403378 581986 403614
rect 582222 403378 582306 403614
rect 582542 403378 582574 403614
rect 581954 403294 582574 403378
rect 581954 403058 581986 403294
rect 582222 403058 582306 403294
rect 582542 403058 582574 403294
rect 581954 367614 582574 403058
rect 581954 367378 581986 367614
rect 582222 367378 582306 367614
rect 582542 367378 582574 367614
rect 581954 367294 582574 367378
rect 581954 367058 581986 367294
rect 582222 367058 582306 367294
rect 582542 367058 582574 367294
rect 581954 331614 582574 367058
rect 581954 331378 581986 331614
rect 582222 331378 582306 331614
rect 582542 331378 582574 331614
rect 581954 331294 582574 331378
rect 581954 331058 581986 331294
rect 582222 331058 582306 331294
rect 582542 331058 582574 331294
rect 581954 295614 582574 331058
rect 581954 295378 581986 295614
rect 582222 295378 582306 295614
rect 582542 295378 582574 295614
rect 581954 295294 582574 295378
rect 581954 295058 581986 295294
rect 582222 295058 582306 295294
rect 582542 295058 582574 295294
rect 581954 259614 582574 295058
rect 581954 259378 581986 259614
rect 582222 259378 582306 259614
rect 582542 259378 582574 259614
rect 581954 259294 582574 259378
rect 581954 259058 581986 259294
rect 582222 259058 582306 259294
rect 582542 259058 582574 259294
rect 581954 223614 582574 259058
rect 581954 223378 581986 223614
rect 582222 223378 582306 223614
rect 582542 223378 582574 223614
rect 581954 223294 582574 223378
rect 581954 223058 581986 223294
rect 582222 223058 582306 223294
rect 582542 223058 582574 223294
rect 581954 187614 582574 223058
rect 581954 187378 581986 187614
rect 582222 187378 582306 187614
rect 582542 187378 582574 187614
rect 581954 187294 582574 187378
rect 581954 187058 581986 187294
rect 582222 187058 582306 187294
rect 582542 187058 582574 187294
rect 581954 151614 582574 187058
rect 581954 151378 581986 151614
rect 582222 151378 582306 151614
rect 582542 151378 582574 151614
rect 581954 151294 582574 151378
rect 581954 151058 581986 151294
rect 582222 151058 582306 151294
rect 582542 151058 582574 151294
rect 581954 115614 582574 151058
rect 581954 115378 581986 115614
rect 582222 115378 582306 115614
rect 582542 115378 582574 115614
rect 581954 115294 582574 115378
rect 581954 115058 581986 115294
rect 582222 115058 582306 115294
rect 582542 115058 582574 115294
rect 581954 79614 582574 115058
rect 581954 79378 581986 79614
rect 582222 79378 582306 79614
rect 582542 79378 582574 79614
rect 581954 79294 582574 79378
rect 581954 79058 581986 79294
rect 582222 79058 582306 79294
rect 582542 79058 582574 79294
rect 581954 43614 582574 79058
rect 581954 43378 581986 43614
rect 582222 43378 582306 43614
rect 582542 43378 582574 43614
rect 581954 43294 582574 43378
rect 581954 43058 581986 43294
rect 582222 43058 582306 43294
rect 582542 43058 582574 43294
rect 581954 7614 582574 43058
rect 581954 7378 581986 7614
rect 582222 7378 582306 7614
rect 582542 7378 582574 7614
rect 581954 7294 582574 7378
rect 581954 7058 581986 7294
rect 582222 7058 582306 7294
rect 582542 7058 582574 7294
rect 581954 -4186 582574 7058
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 686654 585930 704282
rect 585310 686418 585342 686654
rect 585578 686418 585662 686654
rect 585898 686418 585930 686654
rect 585310 686334 585930 686418
rect 585310 686098 585342 686334
rect 585578 686098 585662 686334
rect 585898 686098 585930 686334
rect 585310 650654 585930 686098
rect 585310 650418 585342 650654
rect 585578 650418 585662 650654
rect 585898 650418 585930 650654
rect 585310 650334 585930 650418
rect 585310 650098 585342 650334
rect 585578 650098 585662 650334
rect 585898 650098 585930 650334
rect 585310 614654 585930 650098
rect 585310 614418 585342 614654
rect 585578 614418 585662 614654
rect 585898 614418 585930 614654
rect 585310 614334 585930 614418
rect 585310 614098 585342 614334
rect 585578 614098 585662 614334
rect 585898 614098 585930 614334
rect 585310 578654 585930 614098
rect 585310 578418 585342 578654
rect 585578 578418 585662 578654
rect 585898 578418 585930 578654
rect 585310 578334 585930 578418
rect 585310 578098 585342 578334
rect 585578 578098 585662 578334
rect 585898 578098 585930 578334
rect 585310 542654 585930 578098
rect 585310 542418 585342 542654
rect 585578 542418 585662 542654
rect 585898 542418 585930 542654
rect 585310 542334 585930 542418
rect 585310 542098 585342 542334
rect 585578 542098 585662 542334
rect 585898 542098 585930 542334
rect 585310 506654 585930 542098
rect 585310 506418 585342 506654
rect 585578 506418 585662 506654
rect 585898 506418 585930 506654
rect 585310 506334 585930 506418
rect 585310 506098 585342 506334
rect 585578 506098 585662 506334
rect 585898 506098 585930 506334
rect 585310 470654 585930 506098
rect 585310 470418 585342 470654
rect 585578 470418 585662 470654
rect 585898 470418 585930 470654
rect 585310 470334 585930 470418
rect 585310 470098 585342 470334
rect 585578 470098 585662 470334
rect 585898 470098 585930 470334
rect 585310 434654 585930 470098
rect 585310 434418 585342 434654
rect 585578 434418 585662 434654
rect 585898 434418 585930 434654
rect 585310 434334 585930 434418
rect 585310 434098 585342 434334
rect 585578 434098 585662 434334
rect 585898 434098 585930 434334
rect 585310 398654 585930 434098
rect 585310 398418 585342 398654
rect 585578 398418 585662 398654
rect 585898 398418 585930 398654
rect 585310 398334 585930 398418
rect 585310 398098 585342 398334
rect 585578 398098 585662 398334
rect 585898 398098 585930 398334
rect 585310 362654 585930 398098
rect 585310 362418 585342 362654
rect 585578 362418 585662 362654
rect 585898 362418 585930 362654
rect 585310 362334 585930 362418
rect 585310 362098 585342 362334
rect 585578 362098 585662 362334
rect 585898 362098 585930 362334
rect 585310 326654 585930 362098
rect 585310 326418 585342 326654
rect 585578 326418 585662 326654
rect 585898 326418 585930 326654
rect 585310 326334 585930 326418
rect 585310 326098 585342 326334
rect 585578 326098 585662 326334
rect 585898 326098 585930 326334
rect 585310 290654 585930 326098
rect 585310 290418 585342 290654
rect 585578 290418 585662 290654
rect 585898 290418 585930 290654
rect 585310 290334 585930 290418
rect 585310 290098 585342 290334
rect 585578 290098 585662 290334
rect 585898 290098 585930 290334
rect 585310 254654 585930 290098
rect 585310 254418 585342 254654
rect 585578 254418 585662 254654
rect 585898 254418 585930 254654
rect 585310 254334 585930 254418
rect 585310 254098 585342 254334
rect 585578 254098 585662 254334
rect 585898 254098 585930 254334
rect 585310 218654 585930 254098
rect 585310 218418 585342 218654
rect 585578 218418 585662 218654
rect 585898 218418 585930 218654
rect 585310 218334 585930 218418
rect 585310 218098 585342 218334
rect 585578 218098 585662 218334
rect 585898 218098 585930 218334
rect 585310 182654 585930 218098
rect 585310 182418 585342 182654
rect 585578 182418 585662 182654
rect 585898 182418 585930 182654
rect 585310 182334 585930 182418
rect 585310 182098 585342 182334
rect 585578 182098 585662 182334
rect 585898 182098 585930 182334
rect 585310 146654 585930 182098
rect 585310 146418 585342 146654
rect 585578 146418 585662 146654
rect 585898 146418 585930 146654
rect 585310 146334 585930 146418
rect 585310 146098 585342 146334
rect 585578 146098 585662 146334
rect 585898 146098 585930 146334
rect 585310 110654 585930 146098
rect 585310 110418 585342 110654
rect 585578 110418 585662 110654
rect 585898 110418 585930 110654
rect 585310 110334 585930 110418
rect 585310 110098 585342 110334
rect 585578 110098 585662 110334
rect 585898 110098 585930 110334
rect 585310 74654 585930 110098
rect 585310 74418 585342 74654
rect 585578 74418 585662 74654
rect 585898 74418 585930 74654
rect 585310 74334 585930 74418
rect 585310 74098 585342 74334
rect 585578 74098 585662 74334
rect 585898 74098 585930 74334
rect 585310 38654 585930 74098
rect 585310 38418 585342 38654
rect 585578 38418 585662 38654
rect 585898 38418 585930 38654
rect 585310 38334 585930 38418
rect 585310 38098 585342 38334
rect 585578 38098 585662 38334
rect 585898 38098 585930 38334
rect 585310 2654 585930 38098
rect 585310 2418 585342 2654
rect 585578 2418 585662 2654
rect 585898 2418 585930 2654
rect 585310 2334 585930 2418
rect 585310 2098 585342 2334
rect 585578 2098 585662 2334
rect 585898 2098 585930 2334
rect 585310 -346 585930 2098
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 687894 586890 705242
rect 586270 687658 586302 687894
rect 586538 687658 586622 687894
rect 586858 687658 586890 687894
rect 586270 687574 586890 687658
rect 586270 687338 586302 687574
rect 586538 687338 586622 687574
rect 586858 687338 586890 687574
rect 586270 651894 586890 687338
rect 586270 651658 586302 651894
rect 586538 651658 586622 651894
rect 586858 651658 586890 651894
rect 586270 651574 586890 651658
rect 586270 651338 586302 651574
rect 586538 651338 586622 651574
rect 586858 651338 586890 651574
rect 586270 615894 586890 651338
rect 586270 615658 586302 615894
rect 586538 615658 586622 615894
rect 586858 615658 586890 615894
rect 586270 615574 586890 615658
rect 586270 615338 586302 615574
rect 586538 615338 586622 615574
rect 586858 615338 586890 615574
rect 586270 579894 586890 615338
rect 586270 579658 586302 579894
rect 586538 579658 586622 579894
rect 586858 579658 586890 579894
rect 586270 579574 586890 579658
rect 586270 579338 586302 579574
rect 586538 579338 586622 579574
rect 586858 579338 586890 579574
rect 586270 543894 586890 579338
rect 586270 543658 586302 543894
rect 586538 543658 586622 543894
rect 586858 543658 586890 543894
rect 586270 543574 586890 543658
rect 586270 543338 586302 543574
rect 586538 543338 586622 543574
rect 586858 543338 586890 543574
rect 586270 507894 586890 543338
rect 586270 507658 586302 507894
rect 586538 507658 586622 507894
rect 586858 507658 586890 507894
rect 586270 507574 586890 507658
rect 586270 507338 586302 507574
rect 586538 507338 586622 507574
rect 586858 507338 586890 507574
rect 586270 471894 586890 507338
rect 586270 471658 586302 471894
rect 586538 471658 586622 471894
rect 586858 471658 586890 471894
rect 586270 471574 586890 471658
rect 586270 471338 586302 471574
rect 586538 471338 586622 471574
rect 586858 471338 586890 471574
rect 586270 435894 586890 471338
rect 586270 435658 586302 435894
rect 586538 435658 586622 435894
rect 586858 435658 586890 435894
rect 586270 435574 586890 435658
rect 586270 435338 586302 435574
rect 586538 435338 586622 435574
rect 586858 435338 586890 435574
rect 586270 399894 586890 435338
rect 586270 399658 586302 399894
rect 586538 399658 586622 399894
rect 586858 399658 586890 399894
rect 586270 399574 586890 399658
rect 586270 399338 586302 399574
rect 586538 399338 586622 399574
rect 586858 399338 586890 399574
rect 586270 363894 586890 399338
rect 586270 363658 586302 363894
rect 586538 363658 586622 363894
rect 586858 363658 586890 363894
rect 586270 363574 586890 363658
rect 586270 363338 586302 363574
rect 586538 363338 586622 363574
rect 586858 363338 586890 363574
rect 586270 327894 586890 363338
rect 586270 327658 586302 327894
rect 586538 327658 586622 327894
rect 586858 327658 586890 327894
rect 586270 327574 586890 327658
rect 586270 327338 586302 327574
rect 586538 327338 586622 327574
rect 586858 327338 586890 327574
rect 586270 291894 586890 327338
rect 586270 291658 586302 291894
rect 586538 291658 586622 291894
rect 586858 291658 586890 291894
rect 586270 291574 586890 291658
rect 586270 291338 586302 291574
rect 586538 291338 586622 291574
rect 586858 291338 586890 291574
rect 586270 255894 586890 291338
rect 586270 255658 586302 255894
rect 586538 255658 586622 255894
rect 586858 255658 586890 255894
rect 586270 255574 586890 255658
rect 586270 255338 586302 255574
rect 586538 255338 586622 255574
rect 586858 255338 586890 255574
rect 586270 219894 586890 255338
rect 586270 219658 586302 219894
rect 586538 219658 586622 219894
rect 586858 219658 586890 219894
rect 586270 219574 586890 219658
rect 586270 219338 586302 219574
rect 586538 219338 586622 219574
rect 586858 219338 586890 219574
rect 586270 183894 586890 219338
rect 586270 183658 586302 183894
rect 586538 183658 586622 183894
rect 586858 183658 586890 183894
rect 586270 183574 586890 183658
rect 586270 183338 586302 183574
rect 586538 183338 586622 183574
rect 586858 183338 586890 183574
rect 586270 147894 586890 183338
rect 586270 147658 586302 147894
rect 586538 147658 586622 147894
rect 586858 147658 586890 147894
rect 586270 147574 586890 147658
rect 586270 147338 586302 147574
rect 586538 147338 586622 147574
rect 586858 147338 586890 147574
rect 586270 111894 586890 147338
rect 586270 111658 586302 111894
rect 586538 111658 586622 111894
rect 586858 111658 586890 111894
rect 586270 111574 586890 111658
rect 586270 111338 586302 111574
rect 586538 111338 586622 111574
rect 586858 111338 586890 111574
rect 586270 75894 586890 111338
rect 586270 75658 586302 75894
rect 586538 75658 586622 75894
rect 586858 75658 586890 75894
rect 586270 75574 586890 75658
rect 586270 75338 586302 75574
rect 586538 75338 586622 75574
rect 586858 75338 586890 75574
rect 586270 39894 586890 75338
rect 586270 39658 586302 39894
rect 586538 39658 586622 39894
rect 586858 39658 586890 39894
rect 586270 39574 586890 39658
rect 586270 39338 586302 39574
rect 586538 39338 586622 39574
rect 586858 39338 586890 39574
rect 586270 3894 586890 39338
rect 586270 3658 586302 3894
rect 586538 3658 586622 3894
rect 586858 3658 586890 3894
rect 586270 3574 586890 3658
rect 586270 3338 586302 3574
rect 586538 3338 586622 3574
rect 586858 3338 586890 3574
rect 586270 -1306 586890 3338
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 689134 587850 706202
rect 587230 688898 587262 689134
rect 587498 688898 587582 689134
rect 587818 688898 587850 689134
rect 587230 688814 587850 688898
rect 587230 688578 587262 688814
rect 587498 688578 587582 688814
rect 587818 688578 587850 688814
rect 587230 653134 587850 688578
rect 587230 652898 587262 653134
rect 587498 652898 587582 653134
rect 587818 652898 587850 653134
rect 587230 652814 587850 652898
rect 587230 652578 587262 652814
rect 587498 652578 587582 652814
rect 587818 652578 587850 652814
rect 587230 617134 587850 652578
rect 587230 616898 587262 617134
rect 587498 616898 587582 617134
rect 587818 616898 587850 617134
rect 587230 616814 587850 616898
rect 587230 616578 587262 616814
rect 587498 616578 587582 616814
rect 587818 616578 587850 616814
rect 587230 581134 587850 616578
rect 587230 580898 587262 581134
rect 587498 580898 587582 581134
rect 587818 580898 587850 581134
rect 587230 580814 587850 580898
rect 587230 580578 587262 580814
rect 587498 580578 587582 580814
rect 587818 580578 587850 580814
rect 587230 545134 587850 580578
rect 587230 544898 587262 545134
rect 587498 544898 587582 545134
rect 587818 544898 587850 545134
rect 587230 544814 587850 544898
rect 587230 544578 587262 544814
rect 587498 544578 587582 544814
rect 587818 544578 587850 544814
rect 587230 509134 587850 544578
rect 587230 508898 587262 509134
rect 587498 508898 587582 509134
rect 587818 508898 587850 509134
rect 587230 508814 587850 508898
rect 587230 508578 587262 508814
rect 587498 508578 587582 508814
rect 587818 508578 587850 508814
rect 587230 473134 587850 508578
rect 587230 472898 587262 473134
rect 587498 472898 587582 473134
rect 587818 472898 587850 473134
rect 587230 472814 587850 472898
rect 587230 472578 587262 472814
rect 587498 472578 587582 472814
rect 587818 472578 587850 472814
rect 587230 437134 587850 472578
rect 587230 436898 587262 437134
rect 587498 436898 587582 437134
rect 587818 436898 587850 437134
rect 587230 436814 587850 436898
rect 587230 436578 587262 436814
rect 587498 436578 587582 436814
rect 587818 436578 587850 436814
rect 587230 401134 587850 436578
rect 587230 400898 587262 401134
rect 587498 400898 587582 401134
rect 587818 400898 587850 401134
rect 587230 400814 587850 400898
rect 587230 400578 587262 400814
rect 587498 400578 587582 400814
rect 587818 400578 587850 400814
rect 587230 365134 587850 400578
rect 587230 364898 587262 365134
rect 587498 364898 587582 365134
rect 587818 364898 587850 365134
rect 587230 364814 587850 364898
rect 587230 364578 587262 364814
rect 587498 364578 587582 364814
rect 587818 364578 587850 364814
rect 587230 329134 587850 364578
rect 587230 328898 587262 329134
rect 587498 328898 587582 329134
rect 587818 328898 587850 329134
rect 587230 328814 587850 328898
rect 587230 328578 587262 328814
rect 587498 328578 587582 328814
rect 587818 328578 587850 328814
rect 587230 293134 587850 328578
rect 587230 292898 587262 293134
rect 587498 292898 587582 293134
rect 587818 292898 587850 293134
rect 587230 292814 587850 292898
rect 587230 292578 587262 292814
rect 587498 292578 587582 292814
rect 587818 292578 587850 292814
rect 587230 257134 587850 292578
rect 587230 256898 587262 257134
rect 587498 256898 587582 257134
rect 587818 256898 587850 257134
rect 587230 256814 587850 256898
rect 587230 256578 587262 256814
rect 587498 256578 587582 256814
rect 587818 256578 587850 256814
rect 587230 221134 587850 256578
rect 587230 220898 587262 221134
rect 587498 220898 587582 221134
rect 587818 220898 587850 221134
rect 587230 220814 587850 220898
rect 587230 220578 587262 220814
rect 587498 220578 587582 220814
rect 587818 220578 587850 220814
rect 587230 185134 587850 220578
rect 587230 184898 587262 185134
rect 587498 184898 587582 185134
rect 587818 184898 587850 185134
rect 587230 184814 587850 184898
rect 587230 184578 587262 184814
rect 587498 184578 587582 184814
rect 587818 184578 587850 184814
rect 587230 149134 587850 184578
rect 587230 148898 587262 149134
rect 587498 148898 587582 149134
rect 587818 148898 587850 149134
rect 587230 148814 587850 148898
rect 587230 148578 587262 148814
rect 587498 148578 587582 148814
rect 587818 148578 587850 148814
rect 587230 113134 587850 148578
rect 587230 112898 587262 113134
rect 587498 112898 587582 113134
rect 587818 112898 587850 113134
rect 587230 112814 587850 112898
rect 587230 112578 587262 112814
rect 587498 112578 587582 112814
rect 587818 112578 587850 112814
rect 587230 77134 587850 112578
rect 587230 76898 587262 77134
rect 587498 76898 587582 77134
rect 587818 76898 587850 77134
rect 587230 76814 587850 76898
rect 587230 76578 587262 76814
rect 587498 76578 587582 76814
rect 587818 76578 587850 76814
rect 587230 41134 587850 76578
rect 587230 40898 587262 41134
rect 587498 40898 587582 41134
rect 587818 40898 587850 41134
rect 587230 40814 587850 40898
rect 587230 40578 587262 40814
rect 587498 40578 587582 40814
rect 587818 40578 587850 40814
rect 587230 5134 587850 40578
rect 587230 4898 587262 5134
rect 587498 4898 587582 5134
rect 587818 4898 587850 5134
rect 587230 4814 587850 4898
rect 587230 4578 587262 4814
rect 587498 4578 587582 4814
rect 587818 4578 587850 4814
rect 587230 -2266 587850 4578
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 690374 588810 707162
rect 588190 690138 588222 690374
rect 588458 690138 588542 690374
rect 588778 690138 588810 690374
rect 588190 690054 588810 690138
rect 588190 689818 588222 690054
rect 588458 689818 588542 690054
rect 588778 689818 588810 690054
rect 588190 654374 588810 689818
rect 588190 654138 588222 654374
rect 588458 654138 588542 654374
rect 588778 654138 588810 654374
rect 588190 654054 588810 654138
rect 588190 653818 588222 654054
rect 588458 653818 588542 654054
rect 588778 653818 588810 654054
rect 588190 618374 588810 653818
rect 588190 618138 588222 618374
rect 588458 618138 588542 618374
rect 588778 618138 588810 618374
rect 588190 618054 588810 618138
rect 588190 617818 588222 618054
rect 588458 617818 588542 618054
rect 588778 617818 588810 618054
rect 588190 582374 588810 617818
rect 588190 582138 588222 582374
rect 588458 582138 588542 582374
rect 588778 582138 588810 582374
rect 588190 582054 588810 582138
rect 588190 581818 588222 582054
rect 588458 581818 588542 582054
rect 588778 581818 588810 582054
rect 588190 546374 588810 581818
rect 588190 546138 588222 546374
rect 588458 546138 588542 546374
rect 588778 546138 588810 546374
rect 588190 546054 588810 546138
rect 588190 545818 588222 546054
rect 588458 545818 588542 546054
rect 588778 545818 588810 546054
rect 588190 510374 588810 545818
rect 588190 510138 588222 510374
rect 588458 510138 588542 510374
rect 588778 510138 588810 510374
rect 588190 510054 588810 510138
rect 588190 509818 588222 510054
rect 588458 509818 588542 510054
rect 588778 509818 588810 510054
rect 588190 474374 588810 509818
rect 588190 474138 588222 474374
rect 588458 474138 588542 474374
rect 588778 474138 588810 474374
rect 588190 474054 588810 474138
rect 588190 473818 588222 474054
rect 588458 473818 588542 474054
rect 588778 473818 588810 474054
rect 588190 438374 588810 473818
rect 588190 438138 588222 438374
rect 588458 438138 588542 438374
rect 588778 438138 588810 438374
rect 588190 438054 588810 438138
rect 588190 437818 588222 438054
rect 588458 437818 588542 438054
rect 588778 437818 588810 438054
rect 588190 402374 588810 437818
rect 588190 402138 588222 402374
rect 588458 402138 588542 402374
rect 588778 402138 588810 402374
rect 588190 402054 588810 402138
rect 588190 401818 588222 402054
rect 588458 401818 588542 402054
rect 588778 401818 588810 402054
rect 588190 366374 588810 401818
rect 588190 366138 588222 366374
rect 588458 366138 588542 366374
rect 588778 366138 588810 366374
rect 588190 366054 588810 366138
rect 588190 365818 588222 366054
rect 588458 365818 588542 366054
rect 588778 365818 588810 366054
rect 588190 330374 588810 365818
rect 588190 330138 588222 330374
rect 588458 330138 588542 330374
rect 588778 330138 588810 330374
rect 588190 330054 588810 330138
rect 588190 329818 588222 330054
rect 588458 329818 588542 330054
rect 588778 329818 588810 330054
rect 588190 294374 588810 329818
rect 588190 294138 588222 294374
rect 588458 294138 588542 294374
rect 588778 294138 588810 294374
rect 588190 294054 588810 294138
rect 588190 293818 588222 294054
rect 588458 293818 588542 294054
rect 588778 293818 588810 294054
rect 588190 258374 588810 293818
rect 588190 258138 588222 258374
rect 588458 258138 588542 258374
rect 588778 258138 588810 258374
rect 588190 258054 588810 258138
rect 588190 257818 588222 258054
rect 588458 257818 588542 258054
rect 588778 257818 588810 258054
rect 588190 222374 588810 257818
rect 588190 222138 588222 222374
rect 588458 222138 588542 222374
rect 588778 222138 588810 222374
rect 588190 222054 588810 222138
rect 588190 221818 588222 222054
rect 588458 221818 588542 222054
rect 588778 221818 588810 222054
rect 588190 186374 588810 221818
rect 588190 186138 588222 186374
rect 588458 186138 588542 186374
rect 588778 186138 588810 186374
rect 588190 186054 588810 186138
rect 588190 185818 588222 186054
rect 588458 185818 588542 186054
rect 588778 185818 588810 186054
rect 588190 150374 588810 185818
rect 588190 150138 588222 150374
rect 588458 150138 588542 150374
rect 588778 150138 588810 150374
rect 588190 150054 588810 150138
rect 588190 149818 588222 150054
rect 588458 149818 588542 150054
rect 588778 149818 588810 150054
rect 588190 114374 588810 149818
rect 588190 114138 588222 114374
rect 588458 114138 588542 114374
rect 588778 114138 588810 114374
rect 588190 114054 588810 114138
rect 588190 113818 588222 114054
rect 588458 113818 588542 114054
rect 588778 113818 588810 114054
rect 588190 78374 588810 113818
rect 588190 78138 588222 78374
rect 588458 78138 588542 78374
rect 588778 78138 588810 78374
rect 588190 78054 588810 78138
rect 588190 77818 588222 78054
rect 588458 77818 588542 78054
rect 588778 77818 588810 78054
rect 588190 42374 588810 77818
rect 588190 42138 588222 42374
rect 588458 42138 588542 42374
rect 588778 42138 588810 42374
rect 588190 42054 588810 42138
rect 588190 41818 588222 42054
rect 588458 41818 588542 42054
rect 588778 41818 588810 42054
rect 588190 6374 588810 41818
rect 588190 6138 588222 6374
rect 588458 6138 588542 6374
rect 588778 6138 588810 6374
rect 588190 6054 588810 6138
rect 588190 5818 588222 6054
rect 588458 5818 588542 6054
rect 588778 5818 588810 6054
rect 588190 -3226 588810 5818
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 691614 589770 708122
rect 589150 691378 589182 691614
rect 589418 691378 589502 691614
rect 589738 691378 589770 691614
rect 589150 691294 589770 691378
rect 589150 691058 589182 691294
rect 589418 691058 589502 691294
rect 589738 691058 589770 691294
rect 589150 655614 589770 691058
rect 589150 655378 589182 655614
rect 589418 655378 589502 655614
rect 589738 655378 589770 655614
rect 589150 655294 589770 655378
rect 589150 655058 589182 655294
rect 589418 655058 589502 655294
rect 589738 655058 589770 655294
rect 589150 619614 589770 655058
rect 589150 619378 589182 619614
rect 589418 619378 589502 619614
rect 589738 619378 589770 619614
rect 589150 619294 589770 619378
rect 589150 619058 589182 619294
rect 589418 619058 589502 619294
rect 589738 619058 589770 619294
rect 589150 583614 589770 619058
rect 589150 583378 589182 583614
rect 589418 583378 589502 583614
rect 589738 583378 589770 583614
rect 589150 583294 589770 583378
rect 589150 583058 589182 583294
rect 589418 583058 589502 583294
rect 589738 583058 589770 583294
rect 589150 547614 589770 583058
rect 589150 547378 589182 547614
rect 589418 547378 589502 547614
rect 589738 547378 589770 547614
rect 589150 547294 589770 547378
rect 589150 547058 589182 547294
rect 589418 547058 589502 547294
rect 589738 547058 589770 547294
rect 589150 511614 589770 547058
rect 589150 511378 589182 511614
rect 589418 511378 589502 511614
rect 589738 511378 589770 511614
rect 589150 511294 589770 511378
rect 589150 511058 589182 511294
rect 589418 511058 589502 511294
rect 589738 511058 589770 511294
rect 589150 475614 589770 511058
rect 589150 475378 589182 475614
rect 589418 475378 589502 475614
rect 589738 475378 589770 475614
rect 589150 475294 589770 475378
rect 589150 475058 589182 475294
rect 589418 475058 589502 475294
rect 589738 475058 589770 475294
rect 589150 439614 589770 475058
rect 589150 439378 589182 439614
rect 589418 439378 589502 439614
rect 589738 439378 589770 439614
rect 589150 439294 589770 439378
rect 589150 439058 589182 439294
rect 589418 439058 589502 439294
rect 589738 439058 589770 439294
rect 589150 403614 589770 439058
rect 589150 403378 589182 403614
rect 589418 403378 589502 403614
rect 589738 403378 589770 403614
rect 589150 403294 589770 403378
rect 589150 403058 589182 403294
rect 589418 403058 589502 403294
rect 589738 403058 589770 403294
rect 589150 367614 589770 403058
rect 589150 367378 589182 367614
rect 589418 367378 589502 367614
rect 589738 367378 589770 367614
rect 589150 367294 589770 367378
rect 589150 367058 589182 367294
rect 589418 367058 589502 367294
rect 589738 367058 589770 367294
rect 589150 331614 589770 367058
rect 589150 331378 589182 331614
rect 589418 331378 589502 331614
rect 589738 331378 589770 331614
rect 589150 331294 589770 331378
rect 589150 331058 589182 331294
rect 589418 331058 589502 331294
rect 589738 331058 589770 331294
rect 589150 295614 589770 331058
rect 589150 295378 589182 295614
rect 589418 295378 589502 295614
rect 589738 295378 589770 295614
rect 589150 295294 589770 295378
rect 589150 295058 589182 295294
rect 589418 295058 589502 295294
rect 589738 295058 589770 295294
rect 589150 259614 589770 295058
rect 589150 259378 589182 259614
rect 589418 259378 589502 259614
rect 589738 259378 589770 259614
rect 589150 259294 589770 259378
rect 589150 259058 589182 259294
rect 589418 259058 589502 259294
rect 589738 259058 589770 259294
rect 589150 223614 589770 259058
rect 589150 223378 589182 223614
rect 589418 223378 589502 223614
rect 589738 223378 589770 223614
rect 589150 223294 589770 223378
rect 589150 223058 589182 223294
rect 589418 223058 589502 223294
rect 589738 223058 589770 223294
rect 589150 187614 589770 223058
rect 589150 187378 589182 187614
rect 589418 187378 589502 187614
rect 589738 187378 589770 187614
rect 589150 187294 589770 187378
rect 589150 187058 589182 187294
rect 589418 187058 589502 187294
rect 589738 187058 589770 187294
rect 589150 151614 589770 187058
rect 589150 151378 589182 151614
rect 589418 151378 589502 151614
rect 589738 151378 589770 151614
rect 589150 151294 589770 151378
rect 589150 151058 589182 151294
rect 589418 151058 589502 151294
rect 589738 151058 589770 151294
rect 589150 115614 589770 151058
rect 589150 115378 589182 115614
rect 589418 115378 589502 115614
rect 589738 115378 589770 115614
rect 589150 115294 589770 115378
rect 589150 115058 589182 115294
rect 589418 115058 589502 115294
rect 589738 115058 589770 115294
rect 589150 79614 589770 115058
rect 589150 79378 589182 79614
rect 589418 79378 589502 79614
rect 589738 79378 589770 79614
rect 589150 79294 589770 79378
rect 589150 79058 589182 79294
rect 589418 79058 589502 79294
rect 589738 79058 589770 79294
rect 589150 43614 589770 79058
rect 589150 43378 589182 43614
rect 589418 43378 589502 43614
rect 589738 43378 589770 43614
rect 589150 43294 589770 43378
rect 589150 43058 589182 43294
rect 589418 43058 589502 43294
rect 589738 43058 589770 43294
rect 589150 7614 589770 43058
rect 589150 7378 589182 7614
rect 589418 7378 589502 7614
rect 589738 7378 589770 7614
rect 589150 7294 589770 7378
rect 589150 7058 589182 7294
rect 589418 7058 589502 7294
rect 589738 7058 589770 7294
rect 581954 -4422 581986 -4186
rect 582222 -4422 582306 -4186
rect 582542 -4422 582574 -4186
rect 581954 -4506 582574 -4422
rect 581954 -4742 581986 -4506
rect 582222 -4742 582306 -4506
rect 582542 -4742 582574 -4506
rect 581954 -7654 582574 -4742
rect 589150 -4186 589770 7058
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 692854 590730 709082
rect 590110 692618 590142 692854
rect 590378 692618 590462 692854
rect 590698 692618 590730 692854
rect 590110 692534 590730 692618
rect 590110 692298 590142 692534
rect 590378 692298 590462 692534
rect 590698 692298 590730 692534
rect 590110 656854 590730 692298
rect 590110 656618 590142 656854
rect 590378 656618 590462 656854
rect 590698 656618 590730 656854
rect 590110 656534 590730 656618
rect 590110 656298 590142 656534
rect 590378 656298 590462 656534
rect 590698 656298 590730 656534
rect 590110 620854 590730 656298
rect 590110 620618 590142 620854
rect 590378 620618 590462 620854
rect 590698 620618 590730 620854
rect 590110 620534 590730 620618
rect 590110 620298 590142 620534
rect 590378 620298 590462 620534
rect 590698 620298 590730 620534
rect 590110 584854 590730 620298
rect 590110 584618 590142 584854
rect 590378 584618 590462 584854
rect 590698 584618 590730 584854
rect 590110 584534 590730 584618
rect 590110 584298 590142 584534
rect 590378 584298 590462 584534
rect 590698 584298 590730 584534
rect 590110 548854 590730 584298
rect 590110 548618 590142 548854
rect 590378 548618 590462 548854
rect 590698 548618 590730 548854
rect 590110 548534 590730 548618
rect 590110 548298 590142 548534
rect 590378 548298 590462 548534
rect 590698 548298 590730 548534
rect 590110 512854 590730 548298
rect 590110 512618 590142 512854
rect 590378 512618 590462 512854
rect 590698 512618 590730 512854
rect 590110 512534 590730 512618
rect 590110 512298 590142 512534
rect 590378 512298 590462 512534
rect 590698 512298 590730 512534
rect 590110 476854 590730 512298
rect 590110 476618 590142 476854
rect 590378 476618 590462 476854
rect 590698 476618 590730 476854
rect 590110 476534 590730 476618
rect 590110 476298 590142 476534
rect 590378 476298 590462 476534
rect 590698 476298 590730 476534
rect 590110 440854 590730 476298
rect 590110 440618 590142 440854
rect 590378 440618 590462 440854
rect 590698 440618 590730 440854
rect 590110 440534 590730 440618
rect 590110 440298 590142 440534
rect 590378 440298 590462 440534
rect 590698 440298 590730 440534
rect 590110 404854 590730 440298
rect 590110 404618 590142 404854
rect 590378 404618 590462 404854
rect 590698 404618 590730 404854
rect 590110 404534 590730 404618
rect 590110 404298 590142 404534
rect 590378 404298 590462 404534
rect 590698 404298 590730 404534
rect 590110 368854 590730 404298
rect 590110 368618 590142 368854
rect 590378 368618 590462 368854
rect 590698 368618 590730 368854
rect 590110 368534 590730 368618
rect 590110 368298 590142 368534
rect 590378 368298 590462 368534
rect 590698 368298 590730 368534
rect 590110 332854 590730 368298
rect 590110 332618 590142 332854
rect 590378 332618 590462 332854
rect 590698 332618 590730 332854
rect 590110 332534 590730 332618
rect 590110 332298 590142 332534
rect 590378 332298 590462 332534
rect 590698 332298 590730 332534
rect 590110 296854 590730 332298
rect 590110 296618 590142 296854
rect 590378 296618 590462 296854
rect 590698 296618 590730 296854
rect 590110 296534 590730 296618
rect 590110 296298 590142 296534
rect 590378 296298 590462 296534
rect 590698 296298 590730 296534
rect 590110 260854 590730 296298
rect 590110 260618 590142 260854
rect 590378 260618 590462 260854
rect 590698 260618 590730 260854
rect 590110 260534 590730 260618
rect 590110 260298 590142 260534
rect 590378 260298 590462 260534
rect 590698 260298 590730 260534
rect 590110 224854 590730 260298
rect 590110 224618 590142 224854
rect 590378 224618 590462 224854
rect 590698 224618 590730 224854
rect 590110 224534 590730 224618
rect 590110 224298 590142 224534
rect 590378 224298 590462 224534
rect 590698 224298 590730 224534
rect 590110 188854 590730 224298
rect 590110 188618 590142 188854
rect 590378 188618 590462 188854
rect 590698 188618 590730 188854
rect 590110 188534 590730 188618
rect 590110 188298 590142 188534
rect 590378 188298 590462 188534
rect 590698 188298 590730 188534
rect 590110 152854 590730 188298
rect 590110 152618 590142 152854
rect 590378 152618 590462 152854
rect 590698 152618 590730 152854
rect 590110 152534 590730 152618
rect 590110 152298 590142 152534
rect 590378 152298 590462 152534
rect 590698 152298 590730 152534
rect 590110 116854 590730 152298
rect 590110 116618 590142 116854
rect 590378 116618 590462 116854
rect 590698 116618 590730 116854
rect 590110 116534 590730 116618
rect 590110 116298 590142 116534
rect 590378 116298 590462 116534
rect 590698 116298 590730 116534
rect 590110 80854 590730 116298
rect 590110 80618 590142 80854
rect 590378 80618 590462 80854
rect 590698 80618 590730 80854
rect 590110 80534 590730 80618
rect 590110 80298 590142 80534
rect 590378 80298 590462 80534
rect 590698 80298 590730 80534
rect 590110 44854 590730 80298
rect 590110 44618 590142 44854
rect 590378 44618 590462 44854
rect 590698 44618 590730 44854
rect 590110 44534 590730 44618
rect 590110 44298 590142 44534
rect 590378 44298 590462 44534
rect 590698 44298 590730 44534
rect 590110 8854 590730 44298
rect 590110 8618 590142 8854
rect 590378 8618 590462 8854
rect 590698 8618 590730 8854
rect 590110 8534 590730 8618
rect 590110 8298 590142 8534
rect 590378 8298 590462 8534
rect 590698 8298 590730 8534
rect 590110 -5146 590730 8298
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 694094 591690 710042
rect 591070 693858 591102 694094
rect 591338 693858 591422 694094
rect 591658 693858 591690 694094
rect 591070 693774 591690 693858
rect 591070 693538 591102 693774
rect 591338 693538 591422 693774
rect 591658 693538 591690 693774
rect 591070 658094 591690 693538
rect 591070 657858 591102 658094
rect 591338 657858 591422 658094
rect 591658 657858 591690 658094
rect 591070 657774 591690 657858
rect 591070 657538 591102 657774
rect 591338 657538 591422 657774
rect 591658 657538 591690 657774
rect 591070 622094 591690 657538
rect 591070 621858 591102 622094
rect 591338 621858 591422 622094
rect 591658 621858 591690 622094
rect 591070 621774 591690 621858
rect 591070 621538 591102 621774
rect 591338 621538 591422 621774
rect 591658 621538 591690 621774
rect 591070 586094 591690 621538
rect 591070 585858 591102 586094
rect 591338 585858 591422 586094
rect 591658 585858 591690 586094
rect 591070 585774 591690 585858
rect 591070 585538 591102 585774
rect 591338 585538 591422 585774
rect 591658 585538 591690 585774
rect 591070 550094 591690 585538
rect 591070 549858 591102 550094
rect 591338 549858 591422 550094
rect 591658 549858 591690 550094
rect 591070 549774 591690 549858
rect 591070 549538 591102 549774
rect 591338 549538 591422 549774
rect 591658 549538 591690 549774
rect 591070 514094 591690 549538
rect 591070 513858 591102 514094
rect 591338 513858 591422 514094
rect 591658 513858 591690 514094
rect 591070 513774 591690 513858
rect 591070 513538 591102 513774
rect 591338 513538 591422 513774
rect 591658 513538 591690 513774
rect 591070 478094 591690 513538
rect 591070 477858 591102 478094
rect 591338 477858 591422 478094
rect 591658 477858 591690 478094
rect 591070 477774 591690 477858
rect 591070 477538 591102 477774
rect 591338 477538 591422 477774
rect 591658 477538 591690 477774
rect 591070 442094 591690 477538
rect 591070 441858 591102 442094
rect 591338 441858 591422 442094
rect 591658 441858 591690 442094
rect 591070 441774 591690 441858
rect 591070 441538 591102 441774
rect 591338 441538 591422 441774
rect 591658 441538 591690 441774
rect 591070 406094 591690 441538
rect 591070 405858 591102 406094
rect 591338 405858 591422 406094
rect 591658 405858 591690 406094
rect 591070 405774 591690 405858
rect 591070 405538 591102 405774
rect 591338 405538 591422 405774
rect 591658 405538 591690 405774
rect 591070 370094 591690 405538
rect 591070 369858 591102 370094
rect 591338 369858 591422 370094
rect 591658 369858 591690 370094
rect 591070 369774 591690 369858
rect 591070 369538 591102 369774
rect 591338 369538 591422 369774
rect 591658 369538 591690 369774
rect 591070 334094 591690 369538
rect 591070 333858 591102 334094
rect 591338 333858 591422 334094
rect 591658 333858 591690 334094
rect 591070 333774 591690 333858
rect 591070 333538 591102 333774
rect 591338 333538 591422 333774
rect 591658 333538 591690 333774
rect 591070 298094 591690 333538
rect 591070 297858 591102 298094
rect 591338 297858 591422 298094
rect 591658 297858 591690 298094
rect 591070 297774 591690 297858
rect 591070 297538 591102 297774
rect 591338 297538 591422 297774
rect 591658 297538 591690 297774
rect 591070 262094 591690 297538
rect 591070 261858 591102 262094
rect 591338 261858 591422 262094
rect 591658 261858 591690 262094
rect 591070 261774 591690 261858
rect 591070 261538 591102 261774
rect 591338 261538 591422 261774
rect 591658 261538 591690 261774
rect 591070 226094 591690 261538
rect 591070 225858 591102 226094
rect 591338 225858 591422 226094
rect 591658 225858 591690 226094
rect 591070 225774 591690 225858
rect 591070 225538 591102 225774
rect 591338 225538 591422 225774
rect 591658 225538 591690 225774
rect 591070 190094 591690 225538
rect 591070 189858 591102 190094
rect 591338 189858 591422 190094
rect 591658 189858 591690 190094
rect 591070 189774 591690 189858
rect 591070 189538 591102 189774
rect 591338 189538 591422 189774
rect 591658 189538 591690 189774
rect 591070 154094 591690 189538
rect 591070 153858 591102 154094
rect 591338 153858 591422 154094
rect 591658 153858 591690 154094
rect 591070 153774 591690 153858
rect 591070 153538 591102 153774
rect 591338 153538 591422 153774
rect 591658 153538 591690 153774
rect 591070 118094 591690 153538
rect 591070 117858 591102 118094
rect 591338 117858 591422 118094
rect 591658 117858 591690 118094
rect 591070 117774 591690 117858
rect 591070 117538 591102 117774
rect 591338 117538 591422 117774
rect 591658 117538 591690 117774
rect 591070 82094 591690 117538
rect 591070 81858 591102 82094
rect 591338 81858 591422 82094
rect 591658 81858 591690 82094
rect 591070 81774 591690 81858
rect 591070 81538 591102 81774
rect 591338 81538 591422 81774
rect 591658 81538 591690 81774
rect 591070 46094 591690 81538
rect 591070 45858 591102 46094
rect 591338 45858 591422 46094
rect 591658 45858 591690 46094
rect 591070 45774 591690 45858
rect 591070 45538 591102 45774
rect 591338 45538 591422 45774
rect 591658 45538 591690 45774
rect 591070 10094 591690 45538
rect 591070 9858 591102 10094
rect 591338 9858 591422 10094
rect 591658 9858 591690 10094
rect 591070 9774 591690 9858
rect 591070 9538 591102 9774
rect 591338 9538 591422 9774
rect 591658 9538 591690 9774
rect 591070 -6106 591690 9538
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 695334 592650 711002
rect 592030 695098 592062 695334
rect 592298 695098 592382 695334
rect 592618 695098 592650 695334
rect 592030 695014 592650 695098
rect 592030 694778 592062 695014
rect 592298 694778 592382 695014
rect 592618 694778 592650 695014
rect 592030 659334 592650 694778
rect 592030 659098 592062 659334
rect 592298 659098 592382 659334
rect 592618 659098 592650 659334
rect 592030 659014 592650 659098
rect 592030 658778 592062 659014
rect 592298 658778 592382 659014
rect 592618 658778 592650 659014
rect 592030 623334 592650 658778
rect 592030 623098 592062 623334
rect 592298 623098 592382 623334
rect 592618 623098 592650 623334
rect 592030 623014 592650 623098
rect 592030 622778 592062 623014
rect 592298 622778 592382 623014
rect 592618 622778 592650 623014
rect 592030 587334 592650 622778
rect 592030 587098 592062 587334
rect 592298 587098 592382 587334
rect 592618 587098 592650 587334
rect 592030 587014 592650 587098
rect 592030 586778 592062 587014
rect 592298 586778 592382 587014
rect 592618 586778 592650 587014
rect 592030 551334 592650 586778
rect 592030 551098 592062 551334
rect 592298 551098 592382 551334
rect 592618 551098 592650 551334
rect 592030 551014 592650 551098
rect 592030 550778 592062 551014
rect 592298 550778 592382 551014
rect 592618 550778 592650 551014
rect 592030 515334 592650 550778
rect 592030 515098 592062 515334
rect 592298 515098 592382 515334
rect 592618 515098 592650 515334
rect 592030 515014 592650 515098
rect 592030 514778 592062 515014
rect 592298 514778 592382 515014
rect 592618 514778 592650 515014
rect 592030 479334 592650 514778
rect 592030 479098 592062 479334
rect 592298 479098 592382 479334
rect 592618 479098 592650 479334
rect 592030 479014 592650 479098
rect 592030 478778 592062 479014
rect 592298 478778 592382 479014
rect 592618 478778 592650 479014
rect 592030 443334 592650 478778
rect 592030 443098 592062 443334
rect 592298 443098 592382 443334
rect 592618 443098 592650 443334
rect 592030 443014 592650 443098
rect 592030 442778 592062 443014
rect 592298 442778 592382 443014
rect 592618 442778 592650 443014
rect 592030 407334 592650 442778
rect 592030 407098 592062 407334
rect 592298 407098 592382 407334
rect 592618 407098 592650 407334
rect 592030 407014 592650 407098
rect 592030 406778 592062 407014
rect 592298 406778 592382 407014
rect 592618 406778 592650 407014
rect 592030 371334 592650 406778
rect 592030 371098 592062 371334
rect 592298 371098 592382 371334
rect 592618 371098 592650 371334
rect 592030 371014 592650 371098
rect 592030 370778 592062 371014
rect 592298 370778 592382 371014
rect 592618 370778 592650 371014
rect 592030 335334 592650 370778
rect 592030 335098 592062 335334
rect 592298 335098 592382 335334
rect 592618 335098 592650 335334
rect 592030 335014 592650 335098
rect 592030 334778 592062 335014
rect 592298 334778 592382 335014
rect 592618 334778 592650 335014
rect 592030 299334 592650 334778
rect 592030 299098 592062 299334
rect 592298 299098 592382 299334
rect 592618 299098 592650 299334
rect 592030 299014 592650 299098
rect 592030 298778 592062 299014
rect 592298 298778 592382 299014
rect 592618 298778 592650 299014
rect 592030 263334 592650 298778
rect 592030 263098 592062 263334
rect 592298 263098 592382 263334
rect 592618 263098 592650 263334
rect 592030 263014 592650 263098
rect 592030 262778 592062 263014
rect 592298 262778 592382 263014
rect 592618 262778 592650 263014
rect 592030 227334 592650 262778
rect 592030 227098 592062 227334
rect 592298 227098 592382 227334
rect 592618 227098 592650 227334
rect 592030 227014 592650 227098
rect 592030 226778 592062 227014
rect 592298 226778 592382 227014
rect 592618 226778 592650 227014
rect 592030 191334 592650 226778
rect 592030 191098 592062 191334
rect 592298 191098 592382 191334
rect 592618 191098 592650 191334
rect 592030 191014 592650 191098
rect 592030 190778 592062 191014
rect 592298 190778 592382 191014
rect 592618 190778 592650 191014
rect 592030 155334 592650 190778
rect 592030 155098 592062 155334
rect 592298 155098 592382 155334
rect 592618 155098 592650 155334
rect 592030 155014 592650 155098
rect 592030 154778 592062 155014
rect 592298 154778 592382 155014
rect 592618 154778 592650 155014
rect 592030 119334 592650 154778
rect 592030 119098 592062 119334
rect 592298 119098 592382 119334
rect 592618 119098 592650 119334
rect 592030 119014 592650 119098
rect 592030 118778 592062 119014
rect 592298 118778 592382 119014
rect 592618 118778 592650 119014
rect 592030 83334 592650 118778
rect 592030 83098 592062 83334
rect 592298 83098 592382 83334
rect 592618 83098 592650 83334
rect 592030 83014 592650 83098
rect 592030 82778 592062 83014
rect 592298 82778 592382 83014
rect 592618 82778 592650 83014
rect 592030 47334 592650 82778
rect 592030 47098 592062 47334
rect 592298 47098 592382 47334
rect 592618 47098 592650 47334
rect 592030 47014 592650 47098
rect 592030 46778 592062 47014
rect 592298 46778 592382 47014
rect 592618 46778 592650 47014
rect 592030 11334 592650 46778
rect 592030 11098 592062 11334
rect 592298 11098 592382 11334
rect 592618 11098 592650 11334
rect 592030 11014 592650 11098
rect 592030 10778 592062 11014
rect 592298 10778 592382 11014
rect 592618 10778 592650 11014
rect 592030 -7066 592650 10778
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 695098 -8458 695334
rect -8374 695098 -8138 695334
rect -8694 694778 -8458 695014
rect -8374 694778 -8138 695014
rect -8694 659098 -8458 659334
rect -8374 659098 -8138 659334
rect -8694 658778 -8458 659014
rect -8374 658778 -8138 659014
rect -8694 623098 -8458 623334
rect -8374 623098 -8138 623334
rect -8694 622778 -8458 623014
rect -8374 622778 -8138 623014
rect -8694 587098 -8458 587334
rect -8374 587098 -8138 587334
rect -8694 586778 -8458 587014
rect -8374 586778 -8138 587014
rect -8694 551098 -8458 551334
rect -8374 551098 -8138 551334
rect -8694 550778 -8458 551014
rect -8374 550778 -8138 551014
rect -8694 515098 -8458 515334
rect -8374 515098 -8138 515334
rect -8694 514778 -8458 515014
rect -8374 514778 -8138 515014
rect -8694 479098 -8458 479334
rect -8374 479098 -8138 479334
rect -8694 478778 -8458 479014
rect -8374 478778 -8138 479014
rect -8694 443098 -8458 443334
rect -8374 443098 -8138 443334
rect -8694 442778 -8458 443014
rect -8374 442778 -8138 443014
rect -8694 407098 -8458 407334
rect -8374 407098 -8138 407334
rect -8694 406778 -8458 407014
rect -8374 406778 -8138 407014
rect -8694 371098 -8458 371334
rect -8374 371098 -8138 371334
rect -8694 370778 -8458 371014
rect -8374 370778 -8138 371014
rect -8694 335098 -8458 335334
rect -8374 335098 -8138 335334
rect -8694 334778 -8458 335014
rect -8374 334778 -8138 335014
rect -8694 299098 -8458 299334
rect -8374 299098 -8138 299334
rect -8694 298778 -8458 299014
rect -8374 298778 -8138 299014
rect -8694 263098 -8458 263334
rect -8374 263098 -8138 263334
rect -8694 262778 -8458 263014
rect -8374 262778 -8138 263014
rect -8694 227098 -8458 227334
rect -8374 227098 -8138 227334
rect -8694 226778 -8458 227014
rect -8374 226778 -8138 227014
rect -8694 191098 -8458 191334
rect -8374 191098 -8138 191334
rect -8694 190778 -8458 191014
rect -8374 190778 -8138 191014
rect -8694 155098 -8458 155334
rect -8374 155098 -8138 155334
rect -8694 154778 -8458 155014
rect -8374 154778 -8138 155014
rect -8694 119098 -8458 119334
rect -8374 119098 -8138 119334
rect -8694 118778 -8458 119014
rect -8374 118778 -8138 119014
rect -8694 83098 -8458 83334
rect -8374 83098 -8138 83334
rect -8694 82778 -8458 83014
rect -8374 82778 -8138 83014
rect -8694 47098 -8458 47334
rect -8374 47098 -8138 47334
rect -8694 46778 -8458 47014
rect -8374 46778 -8138 47014
rect -8694 11098 -8458 11334
rect -8374 11098 -8138 11334
rect -8694 10778 -8458 11014
rect -8374 10778 -8138 11014
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 693858 -7498 694094
rect -7414 693858 -7178 694094
rect -7734 693538 -7498 693774
rect -7414 693538 -7178 693774
rect -7734 657858 -7498 658094
rect -7414 657858 -7178 658094
rect -7734 657538 -7498 657774
rect -7414 657538 -7178 657774
rect -7734 621858 -7498 622094
rect -7414 621858 -7178 622094
rect -7734 621538 -7498 621774
rect -7414 621538 -7178 621774
rect -7734 585858 -7498 586094
rect -7414 585858 -7178 586094
rect -7734 585538 -7498 585774
rect -7414 585538 -7178 585774
rect -7734 549858 -7498 550094
rect -7414 549858 -7178 550094
rect -7734 549538 -7498 549774
rect -7414 549538 -7178 549774
rect -7734 513858 -7498 514094
rect -7414 513858 -7178 514094
rect -7734 513538 -7498 513774
rect -7414 513538 -7178 513774
rect -7734 477858 -7498 478094
rect -7414 477858 -7178 478094
rect -7734 477538 -7498 477774
rect -7414 477538 -7178 477774
rect -7734 441858 -7498 442094
rect -7414 441858 -7178 442094
rect -7734 441538 -7498 441774
rect -7414 441538 -7178 441774
rect -7734 405858 -7498 406094
rect -7414 405858 -7178 406094
rect -7734 405538 -7498 405774
rect -7414 405538 -7178 405774
rect -7734 369858 -7498 370094
rect -7414 369858 -7178 370094
rect -7734 369538 -7498 369774
rect -7414 369538 -7178 369774
rect -7734 333858 -7498 334094
rect -7414 333858 -7178 334094
rect -7734 333538 -7498 333774
rect -7414 333538 -7178 333774
rect -7734 297858 -7498 298094
rect -7414 297858 -7178 298094
rect -7734 297538 -7498 297774
rect -7414 297538 -7178 297774
rect -7734 261858 -7498 262094
rect -7414 261858 -7178 262094
rect -7734 261538 -7498 261774
rect -7414 261538 -7178 261774
rect -7734 225858 -7498 226094
rect -7414 225858 -7178 226094
rect -7734 225538 -7498 225774
rect -7414 225538 -7178 225774
rect -7734 189858 -7498 190094
rect -7414 189858 -7178 190094
rect -7734 189538 -7498 189774
rect -7414 189538 -7178 189774
rect -7734 153858 -7498 154094
rect -7414 153858 -7178 154094
rect -7734 153538 -7498 153774
rect -7414 153538 -7178 153774
rect -7734 117858 -7498 118094
rect -7414 117858 -7178 118094
rect -7734 117538 -7498 117774
rect -7414 117538 -7178 117774
rect -7734 81858 -7498 82094
rect -7414 81858 -7178 82094
rect -7734 81538 -7498 81774
rect -7414 81538 -7178 81774
rect -7734 45858 -7498 46094
rect -7414 45858 -7178 46094
rect -7734 45538 -7498 45774
rect -7414 45538 -7178 45774
rect -7734 9858 -7498 10094
rect -7414 9858 -7178 10094
rect -7734 9538 -7498 9774
rect -7414 9538 -7178 9774
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 692618 -6538 692854
rect -6454 692618 -6218 692854
rect -6774 692298 -6538 692534
rect -6454 692298 -6218 692534
rect -6774 656618 -6538 656854
rect -6454 656618 -6218 656854
rect -6774 656298 -6538 656534
rect -6454 656298 -6218 656534
rect -6774 620618 -6538 620854
rect -6454 620618 -6218 620854
rect -6774 620298 -6538 620534
rect -6454 620298 -6218 620534
rect -6774 584618 -6538 584854
rect -6454 584618 -6218 584854
rect -6774 584298 -6538 584534
rect -6454 584298 -6218 584534
rect -6774 548618 -6538 548854
rect -6454 548618 -6218 548854
rect -6774 548298 -6538 548534
rect -6454 548298 -6218 548534
rect -6774 512618 -6538 512854
rect -6454 512618 -6218 512854
rect -6774 512298 -6538 512534
rect -6454 512298 -6218 512534
rect -6774 476618 -6538 476854
rect -6454 476618 -6218 476854
rect -6774 476298 -6538 476534
rect -6454 476298 -6218 476534
rect -6774 440618 -6538 440854
rect -6454 440618 -6218 440854
rect -6774 440298 -6538 440534
rect -6454 440298 -6218 440534
rect -6774 404618 -6538 404854
rect -6454 404618 -6218 404854
rect -6774 404298 -6538 404534
rect -6454 404298 -6218 404534
rect -6774 368618 -6538 368854
rect -6454 368618 -6218 368854
rect -6774 368298 -6538 368534
rect -6454 368298 -6218 368534
rect -6774 332618 -6538 332854
rect -6454 332618 -6218 332854
rect -6774 332298 -6538 332534
rect -6454 332298 -6218 332534
rect -6774 296618 -6538 296854
rect -6454 296618 -6218 296854
rect -6774 296298 -6538 296534
rect -6454 296298 -6218 296534
rect -6774 260618 -6538 260854
rect -6454 260618 -6218 260854
rect -6774 260298 -6538 260534
rect -6454 260298 -6218 260534
rect -6774 224618 -6538 224854
rect -6454 224618 -6218 224854
rect -6774 224298 -6538 224534
rect -6454 224298 -6218 224534
rect -6774 188618 -6538 188854
rect -6454 188618 -6218 188854
rect -6774 188298 -6538 188534
rect -6454 188298 -6218 188534
rect -6774 152618 -6538 152854
rect -6454 152618 -6218 152854
rect -6774 152298 -6538 152534
rect -6454 152298 -6218 152534
rect -6774 116618 -6538 116854
rect -6454 116618 -6218 116854
rect -6774 116298 -6538 116534
rect -6454 116298 -6218 116534
rect -6774 80618 -6538 80854
rect -6454 80618 -6218 80854
rect -6774 80298 -6538 80534
rect -6454 80298 -6218 80534
rect -6774 44618 -6538 44854
rect -6454 44618 -6218 44854
rect -6774 44298 -6538 44534
rect -6454 44298 -6218 44534
rect -6774 8618 -6538 8854
rect -6454 8618 -6218 8854
rect -6774 8298 -6538 8534
rect -6454 8298 -6218 8534
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 691378 -5578 691614
rect -5494 691378 -5258 691614
rect -5814 691058 -5578 691294
rect -5494 691058 -5258 691294
rect -5814 655378 -5578 655614
rect -5494 655378 -5258 655614
rect -5814 655058 -5578 655294
rect -5494 655058 -5258 655294
rect -5814 619378 -5578 619614
rect -5494 619378 -5258 619614
rect -5814 619058 -5578 619294
rect -5494 619058 -5258 619294
rect -5814 583378 -5578 583614
rect -5494 583378 -5258 583614
rect -5814 583058 -5578 583294
rect -5494 583058 -5258 583294
rect -5814 547378 -5578 547614
rect -5494 547378 -5258 547614
rect -5814 547058 -5578 547294
rect -5494 547058 -5258 547294
rect -5814 511378 -5578 511614
rect -5494 511378 -5258 511614
rect -5814 511058 -5578 511294
rect -5494 511058 -5258 511294
rect -5814 475378 -5578 475614
rect -5494 475378 -5258 475614
rect -5814 475058 -5578 475294
rect -5494 475058 -5258 475294
rect -5814 439378 -5578 439614
rect -5494 439378 -5258 439614
rect -5814 439058 -5578 439294
rect -5494 439058 -5258 439294
rect -5814 403378 -5578 403614
rect -5494 403378 -5258 403614
rect -5814 403058 -5578 403294
rect -5494 403058 -5258 403294
rect -5814 367378 -5578 367614
rect -5494 367378 -5258 367614
rect -5814 367058 -5578 367294
rect -5494 367058 -5258 367294
rect -5814 331378 -5578 331614
rect -5494 331378 -5258 331614
rect -5814 331058 -5578 331294
rect -5494 331058 -5258 331294
rect -5814 295378 -5578 295614
rect -5494 295378 -5258 295614
rect -5814 295058 -5578 295294
rect -5494 295058 -5258 295294
rect -5814 259378 -5578 259614
rect -5494 259378 -5258 259614
rect -5814 259058 -5578 259294
rect -5494 259058 -5258 259294
rect -5814 223378 -5578 223614
rect -5494 223378 -5258 223614
rect -5814 223058 -5578 223294
rect -5494 223058 -5258 223294
rect -5814 187378 -5578 187614
rect -5494 187378 -5258 187614
rect -5814 187058 -5578 187294
rect -5494 187058 -5258 187294
rect -5814 151378 -5578 151614
rect -5494 151378 -5258 151614
rect -5814 151058 -5578 151294
rect -5494 151058 -5258 151294
rect -5814 115378 -5578 115614
rect -5494 115378 -5258 115614
rect -5814 115058 -5578 115294
rect -5494 115058 -5258 115294
rect -5814 79378 -5578 79614
rect -5494 79378 -5258 79614
rect -5814 79058 -5578 79294
rect -5494 79058 -5258 79294
rect -5814 43378 -5578 43614
rect -5494 43378 -5258 43614
rect -5814 43058 -5578 43294
rect -5494 43058 -5258 43294
rect -5814 7378 -5578 7614
rect -5494 7378 -5258 7614
rect -5814 7058 -5578 7294
rect -5494 7058 -5258 7294
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 690138 -4618 690374
rect -4534 690138 -4298 690374
rect -4854 689818 -4618 690054
rect -4534 689818 -4298 690054
rect -4854 654138 -4618 654374
rect -4534 654138 -4298 654374
rect -4854 653818 -4618 654054
rect -4534 653818 -4298 654054
rect -4854 618138 -4618 618374
rect -4534 618138 -4298 618374
rect -4854 617818 -4618 618054
rect -4534 617818 -4298 618054
rect -4854 582138 -4618 582374
rect -4534 582138 -4298 582374
rect -4854 581818 -4618 582054
rect -4534 581818 -4298 582054
rect -4854 546138 -4618 546374
rect -4534 546138 -4298 546374
rect -4854 545818 -4618 546054
rect -4534 545818 -4298 546054
rect -4854 510138 -4618 510374
rect -4534 510138 -4298 510374
rect -4854 509818 -4618 510054
rect -4534 509818 -4298 510054
rect -4854 474138 -4618 474374
rect -4534 474138 -4298 474374
rect -4854 473818 -4618 474054
rect -4534 473818 -4298 474054
rect -4854 438138 -4618 438374
rect -4534 438138 -4298 438374
rect -4854 437818 -4618 438054
rect -4534 437818 -4298 438054
rect -4854 402138 -4618 402374
rect -4534 402138 -4298 402374
rect -4854 401818 -4618 402054
rect -4534 401818 -4298 402054
rect -4854 366138 -4618 366374
rect -4534 366138 -4298 366374
rect -4854 365818 -4618 366054
rect -4534 365818 -4298 366054
rect -4854 330138 -4618 330374
rect -4534 330138 -4298 330374
rect -4854 329818 -4618 330054
rect -4534 329818 -4298 330054
rect -4854 294138 -4618 294374
rect -4534 294138 -4298 294374
rect -4854 293818 -4618 294054
rect -4534 293818 -4298 294054
rect -4854 258138 -4618 258374
rect -4534 258138 -4298 258374
rect -4854 257818 -4618 258054
rect -4534 257818 -4298 258054
rect -4854 222138 -4618 222374
rect -4534 222138 -4298 222374
rect -4854 221818 -4618 222054
rect -4534 221818 -4298 222054
rect -4854 186138 -4618 186374
rect -4534 186138 -4298 186374
rect -4854 185818 -4618 186054
rect -4534 185818 -4298 186054
rect -4854 150138 -4618 150374
rect -4534 150138 -4298 150374
rect -4854 149818 -4618 150054
rect -4534 149818 -4298 150054
rect -4854 114138 -4618 114374
rect -4534 114138 -4298 114374
rect -4854 113818 -4618 114054
rect -4534 113818 -4298 114054
rect -4854 78138 -4618 78374
rect -4534 78138 -4298 78374
rect -4854 77818 -4618 78054
rect -4534 77818 -4298 78054
rect -4854 42138 -4618 42374
rect -4534 42138 -4298 42374
rect -4854 41818 -4618 42054
rect -4534 41818 -4298 42054
rect -4854 6138 -4618 6374
rect -4534 6138 -4298 6374
rect -4854 5818 -4618 6054
rect -4534 5818 -4298 6054
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 688898 -3658 689134
rect -3574 688898 -3338 689134
rect -3894 688578 -3658 688814
rect -3574 688578 -3338 688814
rect -3894 652898 -3658 653134
rect -3574 652898 -3338 653134
rect -3894 652578 -3658 652814
rect -3574 652578 -3338 652814
rect -3894 616898 -3658 617134
rect -3574 616898 -3338 617134
rect -3894 616578 -3658 616814
rect -3574 616578 -3338 616814
rect -3894 580898 -3658 581134
rect -3574 580898 -3338 581134
rect -3894 580578 -3658 580814
rect -3574 580578 -3338 580814
rect -3894 544898 -3658 545134
rect -3574 544898 -3338 545134
rect -3894 544578 -3658 544814
rect -3574 544578 -3338 544814
rect -3894 508898 -3658 509134
rect -3574 508898 -3338 509134
rect -3894 508578 -3658 508814
rect -3574 508578 -3338 508814
rect -3894 472898 -3658 473134
rect -3574 472898 -3338 473134
rect -3894 472578 -3658 472814
rect -3574 472578 -3338 472814
rect -3894 436898 -3658 437134
rect -3574 436898 -3338 437134
rect -3894 436578 -3658 436814
rect -3574 436578 -3338 436814
rect -3894 400898 -3658 401134
rect -3574 400898 -3338 401134
rect -3894 400578 -3658 400814
rect -3574 400578 -3338 400814
rect -3894 364898 -3658 365134
rect -3574 364898 -3338 365134
rect -3894 364578 -3658 364814
rect -3574 364578 -3338 364814
rect -3894 328898 -3658 329134
rect -3574 328898 -3338 329134
rect -3894 328578 -3658 328814
rect -3574 328578 -3338 328814
rect -3894 292898 -3658 293134
rect -3574 292898 -3338 293134
rect -3894 292578 -3658 292814
rect -3574 292578 -3338 292814
rect -3894 256898 -3658 257134
rect -3574 256898 -3338 257134
rect -3894 256578 -3658 256814
rect -3574 256578 -3338 256814
rect -3894 220898 -3658 221134
rect -3574 220898 -3338 221134
rect -3894 220578 -3658 220814
rect -3574 220578 -3338 220814
rect -3894 184898 -3658 185134
rect -3574 184898 -3338 185134
rect -3894 184578 -3658 184814
rect -3574 184578 -3338 184814
rect -3894 148898 -3658 149134
rect -3574 148898 -3338 149134
rect -3894 148578 -3658 148814
rect -3574 148578 -3338 148814
rect -3894 112898 -3658 113134
rect -3574 112898 -3338 113134
rect -3894 112578 -3658 112814
rect -3574 112578 -3338 112814
rect -3894 76898 -3658 77134
rect -3574 76898 -3338 77134
rect -3894 76578 -3658 76814
rect -3574 76578 -3338 76814
rect -3894 40898 -3658 41134
rect -3574 40898 -3338 41134
rect -3894 40578 -3658 40814
rect -3574 40578 -3338 40814
rect -3894 4898 -3658 5134
rect -3574 4898 -3338 5134
rect -3894 4578 -3658 4814
rect -3574 4578 -3338 4814
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 687658 -2698 687894
rect -2614 687658 -2378 687894
rect -2934 687338 -2698 687574
rect -2614 687338 -2378 687574
rect -2934 651658 -2698 651894
rect -2614 651658 -2378 651894
rect -2934 651338 -2698 651574
rect -2614 651338 -2378 651574
rect -2934 615658 -2698 615894
rect -2614 615658 -2378 615894
rect -2934 615338 -2698 615574
rect -2614 615338 -2378 615574
rect -2934 579658 -2698 579894
rect -2614 579658 -2378 579894
rect -2934 579338 -2698 579574
rect -2614 579338 -2378 579574
rect -2934 543658 -2698 543894
rect -2614 543658 -2378 543894
rect -2934 543338 -2698 543574
rect -2614 543338 -2378 543574
rect -2934 507658 -2698 507894
rect -2614 507658 -2378 507894
rect -2934 507338 -2698 507574
rect -2614 507338 -2378 507574
rect -2934 471658 -2698 471894
rect -2614 471658 -2378 471894
rect -2934 471338 -2698 471574
rect -2614 471338 -2378 471574
rect -2934 435658 -2698 435894
rect -2614 435658 -2378 435894
rect -2934 435338 -2698 435574
rect -2614 435338 -2378 435574
rect -2934 399658 -2698 399894
rect -2614 399658 -2378 399894
rect -2934 399338 -2698 399574
rect -2614 399338 -2378 399574
rect -2934 363658 -2698 363894
rect -2614 363658 -2378 363894
rect -2934 363338 -2698 363574
rect -2614 363338 -2378 363574
rect -2934 327658 -2698 327894
rect -2614 327658 -2378 327894
rect -2934 327338 -2698 327574
rect -2614 327338 -2378 327574
rect -2934 291658 -2698 291894
rect -2614 291658 -2378 291894
rect -2934 291338 -2698 291574
rect -2614 291338 -2378 291574
rect -2934 255658 -2698 255894
rect -2614 255658 -2378 255894
rect -2934 255338 -2698 255574
rect -2614 255338 -2378 255574
rect -2934 219658 -2698 219894
rect -2614 219658 -2378 219894
rect -2934 219338 -2698 219574
rect -2614 219338 -2378 219574
rect -2934 183658 -2698 183894
rect -2614 183658 -2378 183894
rect -2934 183338 -2698 183574
rect -2614 183338 -2378 183574
rect -2934 147658 -2698 147894
rect -2614 147658 -2378 147894
rect -2934 147338 -2698 147574
rect -2614 147338 -2378 147574
rect -2934 111658 -2698 111894
rect -2614 111658 -2378 111894
rect -2934 111338 -2698 111574
rect -2614 111338 -2378 111574
rect -2934 75658 -2698 75894
rect -2614 75658 -2378 75894
rect -2934 75338 -2698 75574
rect -2614 75338 -2378 75574
rect -2934 39658 -2698 39894
rect -2614 39658 -2378 39894
rect -2934 39338 -2698 39574
rect -2614 39338 -2378 39574
rect -2934 3658 -2698 3894
rect -2614 3658 -2378 3894
rect -2934 3338 -2698 3574
rect -2614 3338 -2378 3574
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 686418 -1738 686654
rect -1654 686418 -1418 686654
rect -1974 686098 -1738 686334
rect -1654 686098 -1418 686334
rect -1974 650418 -1738 650654
rect -1654 650418 -1418 650654
rect -1974 650098 -1738 650334
rect -1654 650098 -1418 650334
rect -1974 614418 -1738 614654
rect -1654 614418 -1418 614654
rect -1974 614098 -1738 614334
rect -1654 614098 -1418 614334
rect -1974 578418 -1738 578654
rect -1654 578418 -1418 578654
rect -1974 578098 -1738 578334
rect -1654 578098 -1418 578334
rect -1974 542418 -1738 542654
rect -1654 542418 -1418 542654
rect -1974 542098 -1738 542334
rect -1654 542098 -1418 542334
rect -1974 506418 -1738 506654
rect -1654 506418 -1418 506654
rect -1974 506098 -1738 506334
rect -1654 506098 -1418 506334
rect -1974 470418 -1738 470654
rect -1654 470418 -1418 470654
rect -1974 470098 -1738 470334
rect -1654 470098 -1418 470334
rect -1974 434418 -1738 434654
rect -1654 434418 -1418 434654
rect -1974 434098 -1738 434334
rect -1654 434098 -1418 434334
rect -1974 398418 -1738 398654
rect -1654 398418 -1418 398654
rect -1974 398098 -1738 398334
rect -1654 398098 -1418 398334
rect -1974 362418 -1738 362654
rect -1654 362418 -1418 362654
rect -1974 362098 -1738 362334
rect -1654 362098 -1418 362334
rect -1974 326418 -1738 326654
rect -1654 326418 -1418 326654
rect -1974 326098 -1738 326334
rect -1654 326098 -1418 326334
rect -1974 290418 -1738 290654
rect -1654 290418 -1418 290654
rect -1974 290098 -1738 290334
rect -1654 290098 -1418 290334
rect -1974 254418 -1738 254654
rect -1654 254418 -1418 254654
rect -1974 254098 -1738 254334
rect -1654 254098 -1418 254334
rect -1974 218418 -1738 218654
rect -1654 218418 -1418 218654
rect -1974 218098 -1738 218334
rect -1654 218098 -1418 218334
rect -1974 182418 -1738 182654
rect -1654 182418 -1418 182654
rect -1974 182098 -1738 182334
rect -1654 182098 -1418 182334
rect -1974 146418 -1738 146654
rect -1654 146418 -1418 146654
rect -1974 146098 -1738 146334
rect -1654 146098 -1418 146334
rect -1974 110418 -1738 110654
rect -1654 110418 -1418 110654
rect -1974 110098 -1738 110334
rect -1654 110098 -1418 110334
rect -1974 74418 -1738 74654
rect -1654 74418 -1418 74654
rect -1974 74098 -1738 74334
rect -1654 74098 -1418 74334
rect -1974 38418 -1738 38654
rect -1654 38418 -1418 38654
rect -1974 38098 -1738 38334
rect -1654 38098 -1418 38334
rect -1974 2418 -1738 2654
rect -1654 2418 -1418 2654
rect -1974 2098 -1738 2334
rect -1654 2098 -1418 2334
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1026 704602 1262 704838
rect 1346 704602 1582 704838
rect 1026 704282 1262 704518
rect 1346 704282 1582 704518
rect 1026 686418 1262 686654
rect 1346 686418 1582 686654
rect 1026 686098 1262 686334
rect 1346 686098 1582 686334
rect 1026 650418 1262 650654
rect 1346 650418 1582 650654
rect 1026 650098 1262 650334
rect 1346 650098 1582 650334
rect 1026 614418 1262 614654
rect 1346 614418 1582 614654
rect 1026 614098 1262 614334
rect 1346 614098 1582 614334
rect 1026 578418 1262 578654
rect 1346 578418 1582 578654
rect 1026 578098 1262 578334
rect 1346 578098 1582 578334
rect 1026 542418 1262 542654
rect 1346 542418 1582 542654
rect 1026 542098 1262 542334
rect 1346 542098 1582 542334
rect 1026 506418 1262 506654
rect 1346 506418 1582 506654
rect 1026 506098 1262 506334
rect 1346 506098 1582 506334
rect 1026 470418 1262 470654
rect 1346 470418 1582 470654
rect 1026 470098 1262 470334
rect 1346 470098 1582 470334
rect 1026 434418 1262 434654
rect 1346 434418 1582 434654
rect 1026 434098 1262 434334
rect 1346 434098 1582 434334
rect 1026 398418 1262 398654
rect 1346 398418 1582 398654
rect 1026 398098 1262 398334
rect 1346 398098 1582 398334
rect 1026 362418 1262 362654
rect 1346 362418 1582 362654
rect 1026 362098 1262 362334
rect 1346 362098 1582 362334
rect 1026 326418 1262 326654
rect 1346 326418 1582 326654
rect 1026 326098 1262 326334
rect 1346 326098 1582 326334
rect 1026 290418 1262 290654
rect 1346 290418 1582 290654
rect 1026 290098 1262 290334
rect 1346 290098 1582 290334
rect 1026 254418 1262 254654
rect 1346 254418 1582 254654
rect 1026 254098 1262 254334
rect 1346 254098 1582 254334
rect 1026 218418 1262 218654
rect 1346 218418 1582 218654
rect 1026 218098 1262 218334
rect 1346 218098 1582 218334
rect 1026 182418 1262 182654
rect 1346 182418 1582 182654
rect 1026 182098 1262 182334
rect 1346 182098 1582 182334
rect 1026 146418 1262 146654
rect 1346 146418 1582 146654
rect 1026 146098 1262 146334
rect 1346 146098 1582 146334
rect 1026 110418 1262 110654
rect 1346 110418 1582 110654
rect 1026 110098 1262 110334
rect 1346 110098 1582 110334
rect 1026 74418 1262 74654
rect 1346 74418 1582 74654
rect 1026 74098 1262 74334
rect 1346 74098 1582 74334
rect 1026 38418 1262 38654
rect 1346 38418 1582 38654
rect 1026 38098 1262 38334
rect 1346 38098 1582 38334
rect 1026 2418 1262 2654
rect 1346 2418 1582 2654
rect 1026 2098 1262 2334
rect 1346 2098 1582 2334
rect 1026 -582 1262 -346
rect 1346 -582 1582 -346
rect 1026 -902 1262 -666
rect 1346 -902 1582 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 2266 705562 2502 705798
rect 2586 705562 2822 705798
rect 2266 705242 2502 705478
rect 2586 705242 2822 705478
rect 2266 687658 2502 687894
rect 2586 687658 2822 687894
rect 2266 687338 2502 687574
rect 2586 687338 2822 687574
rect 2266 651658 2502 651894
rect 2586 651658 2822 651894
rect 2266 651338 2502 651574
rect 2586 651338 2822 651574
rect 2266 615658 2502 615894
rect 2586 615658 2822 615894
rect 2266 615338 2502 615574
rect 2586 615338 2822 615574
rect 2266 579658 2502 579894
rect 2586 579658 2822 579894
rect 2266 579338 2502 579574
rect 2586 579338 2822 579574
rect 2266 543658 2502 543894
rect 2586 543658 2822 543894
rect 2266 543338 2502 543574
rect 2586 543338 2822 543574
rect 2266 507658 2502 507894
rect 2586 507658 2822 507894
rect 2266 507338 2502 507574
rect 2586 507338 2822 507574
rect 2266 471658 2502 471894
rect 2586 471658 2822 471894
rect 2266 471338 2502 471574
rect 2586 471338 2822 471574
rect 2266 435658 2502 435894
rect 2586 435658 2822 435894
rect 2266 435338 2502 435574
rect 2586 435338 2822 435574
rect 2266 399658 2502 399894
rect 2586 399658 2822 399894
rect 2266 399338 2502 399574
rect 2586 399338 2822 399574
rect 2266 363658 2502 363894
rect 2586 363658 2822 363894
rect 2266 363338 2502 363574
rect 2586 363338 2822 363574
rect 2266 327658 2502 327894
rect 2586 327658 2822 327894
rect 2266 327338 2502 327574
rect 2586 327338 2822 327574
rect 2266 291658 2502 291894
rect 2586 291658 2822 291894
rect 2266 291338 2502 291574
rect 2586 291338 2822 291574
rect 2266 255658 2502 255894
rect 2586 255658 2822 255894
rect 2266 255338 2502 255574
rect 2586 255338 2822 255574
rect 2266 219658 2502 219894
rect 2586 219658 2822 219894
rect 2266 219338 2502 219574
rect 2586 219338 2822 219574
rect 2266 183658 2502 183894
rect 2586 183658 2822 183894
rect 2266 183338 2502 183574
rect 2586 183338 2822 183574
rect 2266 147658 2502 147894
rect 2586 147658 2822 147894
rect 2266 147338 2502 147574
rect 2586 147338 2822 147574
rect 2266 111658 2502 111894
rect 2586 111658 2822 111894
rect 2266 111338 2502 111574
rect 2586 111338 2822 111574
rect 2266 75658 2502 75894
rect 2586 75658 2822 75894
rect 2266 75338 2502 75574
rect 2586 75338 2822 75574
rect 2266 39658 2502 39894
rect 2586 39658 2822 39894
rect 2266 39338 2502 39574
rect 2586 39338 2822 39574
rect 2266 3658 2502 3894
rect 2586 3658 2822 3894
rect 2266 3338 2502 3574
rect 2586 3338 2822 3574
rect 2266 -1542 2502 -1306
rect 2586 -1542 2822 -1306
rect 2266 -1862 2502 -1626
rect 2586 -1862 2822 -1626
rect 3506 706522 3742 706758
rect 3826 706522 4062 706758
rect 3506 706202 3742 706438
rect 3826 706202 4062 706438
rect 3506 688898 3742 689134
rect 3826 688898 4062 689134
rect 3506 688578 3742 688814
rect 3826 688578 4062 688814
rect 3506 652898 3742 653134
rect 3826 652898 4062 653134
rect 3506 652578 3742 652814
rect 3826 652578 4062 652814
rect 3506 616898 3742 617134
rect 3826 616898 4062 617134
rect 3506 616578 3742 616814
rect 3826 616578 4062 616814
rect 3506 580898 3742 581134
rect 3826 580898 4062 581134
rect 3506 580578 3742 580814
rect 3826 580578 4062 580814
rect 3506 544898 3742 545134
rect 3826 544898 4062 545134
rect 3506 544578 3742 544814
rect 3826 544578 4062 544814
rect 3506 508898 3742 509134
rect 3826 508898 4062 509134
rect 3506 508578 3742 508814
rect 3826 508578 4062 508814
rect 3506 472898 3742 473134
rect 3826 472898 4062 473134
rect 3506 472578 3742 472814
rect 3826 472578 4062 472814
rect 3506 436898 3742 437134
rect 3826 436898 4062 437134
rect 3506 436578 3742 436814
rect 3826 436578 4062 436814
rect 3506 400898 3742 401134
rect 3826 400898 4062 401134
rect 3506 400578 3742 400814
rect 3826 400578 4062 400814
rect 3506 364898 3742 365134
rect 3826 364898 4062 365134
rect 3506 364578 3742 364814
rect 3826 364578 4062 364814
rect 3506 328898 3742 329134
rect 3826 328898 4062 329134
rect 3506 328578 3742 328814
rect 3826 328578 4062 328814
rect 3506 292898 3742 293134
rect 3826 292898 4062 293134
rect 3506 292578 3742 292814
rect 3826 292578 4062 292814
rect 3506 256898 3742 257134
rect 3826 256898 4062 257134
rect 3506 256578 3742 256814
rect 3826 256578 4062 256814
rect 3506 220898 3742 221134
rect 3826 220898 4062 221134
rect 3506 220578 3742 220814
rect 3826 220578 4062 220814
rect 3506 184898 3742 185134
rect 3826 184898 4062 185134
rect 3506 184578 3742 184814
rect 3826 184578 4062 184814
rect 3506 148898 3742 149134
rect 3826 148898 4062 149134
rect 3506 148578 3742 148814
rect 3826 148578 4062 148814
rect 3506 112898 3742 113134
rect 3826 112898 4062 113134
rect 3506 112578 3742 112814
rect 3826 112578 4062 112814
rect 3506 76898 3742 77134
rect 3826 76898 4062 77134
rect 3506 76578 3742 76814
rect 3826 76578 4062 76814
rect 3506 40898 3742 41134
rect 3826 40898 4062 41134
rect 3506 40578 3742 40814
rect 3826 40578 4062 40814
rect 3506 4898 3742 5134
rect 3826 4898 4062 5134
rect 3506 4578 3742 4814
rect 3826 4578 4062 4814
rect 3506 -2502 3742 -2266
rect 3826 -2502 4062 -2266
rect 3506 -2822 3742 -2586
rect 3826 -2822 4062 -2586
rect 4746 707482 4982 707718
rect 5066 707482 5302 707718
rect 4746 707162 4982 707398
rect 5066 707162 5302 707398
rect 4746 690138 4982 690374
rect 5066 690138 5302 690374
rect 4746 689818 4982 690054
rect 5066 689818 5302 690054
rect 4746 654138 4982 654374
rect 5066 654138 5302 654374
rect 4746 653818 4982 654054
rect 5066 653818 5302 654054
rect 4746 618138 4982 618374
rect 5066 618138 5302 618374
rect 4746 617818 4982 618054
rect 5066 617818 5302 618054
rect 4746 582138 4982 582374
rect 5066 582138 5302 582374
rect 4746 581818 4982 582054
rect 5066 581818 5302 582054
rect 4746 546138 4982 546374
rect 5066 546138 5302 546374
rect 4746 545818 4982 546054
rect 5066 545818 5302 546054
rect 4746 510138 4982 510374
rect 5066 510138 5302 510374
rect 4746 509818 4982 510054
rect 5066 509818 5302 510054
rect 4746 474138 4982 474374
rect 5066 474138 5302 474374
rect 4746 473818 4982 474054
rect 5066 473818 5302 474054
rect 4746 438138 4982 438374
rect 5066 438138 5302 438374
rect 4746 437818 4982 438054
rect 5066 437818 5302 438054
rect 4746 402138 4982 402374
rect 5066 402138 5302 402374
rect 4746 401818 4982 402054
rect 5066 401818 5302 402054
rect 4746 366138 4982 366374
rect 5066 366138 5302 366374
rect 4746 365818 4982 366054
rect 5066 365818 5302 366054
rect 4746 330138 4982 330374
rect 5066 330138 5302 330374
rect 4746 329818 4982 330054
rect 5066 329818 5302 330054
rect 4746 294138 4982 294374
rect 5066 294138 5302 294374
rect 4746 293818 4982 294054
rect 5066 293818 5302 294054
rect 4746 258138 4982 258374
rect 5066 258138 5302 258374
rect 4746 257818 4982 258054
rect 5066 257818 5302 258054
rect 4746 222138 4982 222374
rect 5066 222138 5302 222374
rect 4746 221818 4982 222054
rect 5066 221818 5302 222054
rect 4746 186138 4982 186374
rect 5066 186138 5302 186374
rect 4746 185818 4982 186054
rect 5066 185818 5302 186054
rect 4746 150138 4982 150374
rect 5066 150138 5302 150374
rect 4746 149818 4982 150054
rect 5066 149818 5302 150054
rect 4746 114138 4982 114374
rect 5066 114138 5302 114374
rect 4746 113818 4982 114054
rect 5066 113818 5302 114054
rect 4746 78138 4982 78374
rect 5066 78138 5302 78374
rect 4746 77818 4982 78054
rect 5066 77818 5302 78054
rect 4746 42138 4982 42374
rect 5066 42138 5302 42374
rect 4746 41818 4982 42054
rect 5066 41818 5302 42054
rect 4746 6138 4982 6374
rect 5066 6138 5302 6374
rect 4746 5818 4982 6054
rect 5066 5818 5302 6054
rect 4746 -3462 4982 -3226
rect 5066 -3462 5302 -3226
rect 4746 -3782 4982 -3546
rect 5066 -3782 5302 -3546
rect 5986 708442 6222 708678
rect 6306 708442 6542 708678
rect 5986 708122 6222 708358
rect 6306 708122 6542 708358
rect 5986 691378 6222 691614
rect 6306 691378 6542 691614
rect 5986 691058 6222 691294
rect 6306 691058 6542 691294
rect 5986 655378 6222 655614
rect 6306 655378 6542 655614
rect 5986 655058 6222 655294
rect 6306 655058 6542 655294
rect 5986 619378 6222 619614
rect 6306 619378 6542 619614
rect 5986 619058 6222 619294
rect 6306 619058 6542 619294
rect 5986 583378 6222 583614
rect 6306 583378 6542 583614
rect 5986 583058 6222 583294
rect 6306 583058 6542 583294
rect 5986 547378 6222 547614
rect 6306 547378 6542 547614
rect 5986 547058 6222 547294
rect 6306 547058 6542 547294
rect 5986 511378 6222 511614
rect 6306 511378 6542 511614
rect 5986 511058 6222 511294
rect 6306 511058 6542 511294
rect 5986 475378 6222 475614
rect 6306 475378 6542 475614
rect 5986 475058 6222 475294
rect 6306 475058 6542 475294
rect 5986 439378 6222 439614
rect 6306 439378 6542 439614
rect 5986 439058 6222 439294
rect 6306 439058 6542 439294
rect 5986 403378 6222 403614
rect 6306 403378 6542 403614
rect 5986 403058 6222 403294
rect 6306 403058 6542 403294
rect 5986 367378 6222 367614
rect 6306 367378 6542 367614
rect 5986 367058 6222 367294
rect 6306 367058 6542 367294
rect 5986 331378 6222 331614
rect 6306 331378 6542 331614
rect 5986 331058 6222 331294
rect 6306 331058 6542 331294
rect 5986 295378 6222 295614
rect 6306 295378 6542 295614
rect 5986 295058 6222 295294
rect 6306 295058 6542 295294
rect 5986 259378 6222 259614
rect 6306 259378 6542 259614
rect 5986 259058 6222 259294
rect 6306 259058 6542 259294
rect 5986 223378 6222 223614
rect 6306 223378 6542 223614
rect 5986 223058 6222 223294
rect 6306 223058 6542 223294
rect 5986 187378 6222 187614
rect 6306 187378 6542 187614
rect 5986 187058 6222 187294
rect 6306 187058 6542 187294
rect 5986 151378 6222 151614
rect 6306 151378 6542 151614
rect 5986 151058 6222 151294
rect 6306 151058 6542 151294
rect 5986 115378 6222 115614
rect 6306 115378 6542 115614
rect 5986 115058 6222 115294
rect 6306 115058 6542 115294
rect 5986 79378 6222 79614
rect 6306 79378 6542 79614
rect 5986 79058 6222 79294
rect 6306 79058 6542 79294
rect 5986 43378 6222 43614
rect 6306 43378 6542 43614
rect 5986 43058 6222 43294
rect 6306 43058 6542 43294
rect 5986 7378 6222 7614
rect 6306 7378 6542 7614
rect 5986 7058 6222 7294
rect 6306 7058 6542 7294
rect 5986 -4422 6222 -4186
rect 6306 -4422 6542 -4186
rect 5986 -4742 6222 -4506
rect 6306 -4742 6542 -4506
rect 7226 709402 7462 709638
rect 7546 709402 7782 709638
rect 7226 709082 7462 709318
rect 7546 709082 7782 709318
rect 7226 692618 7462 692854
rect 7546 692618 7782 692854
rect 7226 692298 7462 692534
rect 7546 692298 7782 692534
rect 7226 656618 7462 656854
rect 7546 656618 7782 656854
rect 7226 656298 7462 656534
rect 7546 656298 7782 656534
rect 7226 620618 7462 620854
rect 7546 620618 7782 620854
rect 7226 620298 7462 620534
rect 7546 620298 7782 620534
rect 7226 584618 7462 584854
rect 7546 584618 7782 584854
rect 7226 584298 7462 584534
rect 7546 584298 7782 584534
rect 7226 548618 7462 548854
rect 7546 548618 7782 548854
rect 7226 548298 7462 548534
rect 7546 548298 7782 548534
rect 7226 512618 7462 512854
rect 7546 512618 7782 512854
rect 7226 512298 7462 512534
rect 7546 512298 7782 512534
rect 7226 476618 7462 476854
rect 7546 476618 7782 476854
rect 7226 476298 7462 476534
rect 7546 476298 7782 476534
rect 7226 440618 7462 440854
rect 7546 440618 7782 440854
rect 7226 440298 7462 440534
rect 7546 440298 7782 440534
rect 7226 404618 7462 404854
rect 7546 404618 7782 404854
rect 7226 404298 7462 404534
rect 7546 404298 7782 404534
rect 7226 368618 7462 368854
rect 7546 368618 7782 368854
rect 7226 368298 7462 368534
rect 7546 368298 7782 368534
rect 7226 332618 7462 332854
rect 7546 332618 7782 332854
rect 7226 332298 7462 332534
rect 7546 332298 7782 332534
rect 7226 296618 7462 296854
rect 7546 296618 7782 296854
rect 7226 296298 7462 296534
rect 7546 296298 7782 296534
rect 7226 260618 7462 260854
rect 7546 260618 7782 260854
rect 7226 260298 7462 260534
rect 7546 260298 7782 260534
rect 7226 224618 7462 224854
rect 7546 224618 7782 224854
rect 7226 224298 7462 224534
rect 7546 224298 7782 224534
rect 7226 188618 7462 188854
rect 7546 188618 7782 188854
rect 7226 188298 7462 188534
rect 7546 188298 7782 188534
rect 7226 152618 7462 152854
rect 7546 152618 7782 152854
rect 7226 152298 7462 152534
rect 7546 152298 7782 152534
rect 7226 116618 7462 116854
rect 7546 116618 7782 116854
rect 7226 116298 7462 116534
rect 7546 116298 7782 116534
rect 7226 80618 7462 80854
rect 7546 80618 7782 80854
rect 7226 80298 7462 80534
rect 7546 80298 7782 80534
rect 7226 44618 7462 44854
rect 7546 44618 7782 44854
rect 7226 44298 7462 44534
rect 7546 44298 7782 44534
rect 7226 8618 7462 8854
rect 7546 8618 7782 8854
rect 7226 8298 7462 8534
rect 7546 8298 7782 8534
rect 7226 -5382 7462 -5146
rect 7546 -5382 7782 -5146
rect 7226 -5702 7462 -5466
rect 7546 -5702 7782 -5466
rect 8466 710362 8702 710598
rect 8786 710362 9022 710598
rect 8466 710042 8702 710278
rect 8786 710042 9022 710278
rect 8466 693858 8702 694094
rect 8786 693858 9022 694094
rect 8466 693538 8702 693774
rect 8786 693538 9022 693774
rect 8466 657858 8702 658094
rect 8786 657858 9022 658094
rect 8466 657538 8702 657774
rect 8786 657538 9022 657774
rect 8466 621858 8702 622094
rect 8786 621858 9022 622094
rect 8466 621538 8702 621774
rect 8786 621538 9022 621774
rect 8466 585858 8702 586094
rect 8786 585858 9022 586094
rect 8466 585538 8702 585774
rect 8786 585538 9022 585774
rect 8466 549858 8702 550094
rect 8786 549858 9022 550094
rect 8466 549538 8702 549774
rect 8786 549538 9022 549774
rect 8466 513858 8702 514094
rect 8786 513858 9022 514094
rect 8466 513538 8702 513774
rect 8786 513538 9022 513774
rect 8466 477858 8702 478094
rect 8786 477858 9022 478094
rect 8466 477538 8702 477774
rect 8786 477538 9022 477774
rect 8466 441858 8702 442094
rect 8786 441858 9022 442094
rect 8466 441538 8702 441774
rect 8786 441538 9022 441774
rect 8466 405858 8702 406094
rect 8786 405858 9022 406094
rect 8466 405538 8702 405774
rect 8786 405538 9022 405774
rect 8466 369858 8702 370094
rect 8786 369858 9022 370094
rect 8466 369538 8702 369774
rect 8786 369538 9022 369774
rect 8466 333858 8702 334094
rect 8786 333858 9022 334094
rect 8466 333538 8702 333774
rect 8786 333538 9022 333774
rect 8466 297858 8702 298094
rect 8786 297858 9022 298094
rect 8466 297538 8702 297774
rect 8786 297538 9022 297774
rect 8466 261858 8702 262094
rect 8786 261858 9022 262094
rect 8466 261538 8702 261774
rect 8786 261538 9022 261774
rect 8466 225858 8702 226094
rect 8786 225858 9022 226094
rect 8466 225538 8702 225774
rect 8786 225538 9022 225774
rect 8466 189858 8702 190094
rect 8786 189858 9022 190094
rect 8466 189538 8702 189774
rect 8786 189538 9022 189774
rect 8466 153858 8702 154094
rect 8786 153858 9022 154094
rect 8466 153538 8702 153774
rect 8786 153538 9022 153774
rect 8466 117858 8702 118094
rect 8786 117858 9022 118094
rect 8466 117538 8702 117774
rect 8786 117538 9022 117774
rect 8466 81858 8702 82094
rect 8786 81858 9022 82094
rect 8466 81538 8702 81774
rect 8786 81538 9022 81774
rect 8466 45858 8702 46094
rect 8786 45858 9022 46094
rect 8466 45538 8702 45774
rect 8786 45538 9022 45774
rect 8466 9858 8702 10094
rect 8786 9858 9022 10094
rect 8466 9538 8702 9774
rect 8786 9538 9022 9774
rect 8466 -6342 8702 -6106
rect 8786 -6342 9022 -6106
rect 8466 -6662 8702 -6426
rect 8786 -6662 9022 -6426
rect 9706 711322 9942 711558
rect 10026 711322 10262 711558
rect 9706 711002 9942 711238
rect 10026 711002 10262 711238
rect 9706 695098 9942 695334
rect 10026 695098 10262 695334
rect 9706 694778 9942 695014
rect 10026 694778 10262 695014
rect 9706 659098 9942 659334
rect 10026 659098 10262 659334
rect 9706 658778 9942 659014
rect 10026 658778 10262 659014
rect 9706 623098 9942 623334
rect 10026 623098 10262 623334
rect 9706 622778 9942 623014
rect 10026 622778 10262 623014
rect 9706 587098 9942 587334
rect 10026 587098 10262 587334
rect 9706 586778 9942 587014
rect 10026 586778 10262 587014
rect 9706 551098 9942 551334
rect 10026 551098 10262 551334
rect 9706 550778 9942 551014
rect 10026 550778 10262 551014
rect 9706 515098 9942 515334
rect 10026 515098 10262 515334
rect 9706 514778 9942 515014
rect 10026 514778 10262 515014
rect 9706 479098 9942 479334
rect 10026 479098 10262 479334
rect 9706 478778 9942 479014
rect 10026 478778 10262 479014
rect 9706 443098 9942 443334
rect 10026 443098 10262 443334
rect 9706 442778 9942 443014
rect 10026 442778 10262 443014
rect 9706 407098 9942 407334
rect 10026 407098 10262 407334
rect 9706 406778 9942 407014
rect 10026 406778 10262 407014
rect 9706 371098 9942 371334
rect 10026 371098 10262 371334
rect 9706 370778 9942 371014
rect 10026 370778 10262 371014
rect 9706 335098 9942 335334
rect 10026 335098 10262 335334
rect 9706 334778 9942 335014
rect 10026 334778 10262 335014
rect 9706 299098 9942 299334
rect 10026 299098 10262 299334
rect 9706 298778 9942 299014
rect 10026 298778 10262 299014
rect 9706 263098 9942 263334
rect 10026 263098 10262 263334
rect 9706 262778 9942 263014
rect 10026 262778 10262 263014
rect 9706 227098 9942 227334
rect 10026 227098 10262 227334
rect 9706 226778 9942 227014
rect 10026 226778 10262 227014
rect 9706 191098 9942 191334
rect 10026 191098 10262 191334
rect 9706 190778 9942 191014
rect 10026 190778 10262 191014
rect 9706 155098 9942 155334
rect 10026 155098 10262 155334
rect 9706 154778 9942 155014
rect 10026 154778 10262 155014
rect 9706 119098 9942 119334
rect 10026 119098 10262 119334
rect 9706 118778 9942 119014
rect 10026 118778 10262 119014
rect 9706 83098 9942 83334
rect 10026 83098 10262 83334
rect 9706 82778 9942 83014
rect 10026 82778 10262 83014
rect 9706 47098 9942 47334
rect 10026 47098 10262 47334
rect 9706 46778 9942 47014
rect 10026 46778 10262 47014
rect 9706 11098 9942 11334
rect 10026 11098 10262 11334
rect 9706 10778 9942 11014
rect 10026 10778 10262 11014
rect 9706 -7302 9942 -7066
rect 10026 -7302 10262 -7066
rect 9706 -7622 9942 -7386
rect 10026 -7622 10262 -7386
rect 37026 704602 37262 704838
rect 37346 704602 37582 704838
rect 37026 704282 37262 704518
rect 37346 704282 37582 704518
rect 37026 686418 37262 686654
rect 37346 686418 37582 686654
rect 37026 686098 37262 686334
rect 37346 686098 37582 686334
rect 37026 650418 37262 650654
rect 37346 650418 37582 650654
rect 37026 650098 37262 650334
rect 37346 650098 37582 650334
rect 37026 614418 37262 614654
rect 37346 614418 37582 614654
rect 37026 614098 37262 614334
rect 37346 614098 37582 614334
rect 37026 578418 37262 578654
rect 37346 578418 37582 578654
rect 37026 578098 37262 578334
rect 37346 578098 37582 578334
rect 37026 542418 37262 542654
rect 37346 542418 37582 542654
rect 37026 542098 37262 542334
rect 37346 542098 37582 542334
rect 37026 506418 37262 506654
rect 37346 506418 37582 506654
rect 37026 506098 37262 506334
rect 37346 506098 37582 506334
rect 37026 470418 37262 470654
rect 37346 470418 37582 470654
rect 37026 470098 37262 470334
rect 37346 470098 37582 470334
rect 37026 434418 37262 434654
rect 37346 434418 37582 434654
rect 37026 434098 37262 434334
rect 37346 434098 37582 434334
rect 37026 398418 37262 398654
rect 37346 398418 37582 398654
rect 37026 398098 37262 398334
rect 37346 398098 37582 398334
rect 37026 362418 37262 362654
rect 37346 362418 37582 362654
rect 37026 362098 37262 362334
rect 37346 362098 37582 362334
rect 37026 326418 37262 326654
rect 37346 326418 37582 326654
rect 37026 326098 37262 326334
rect 37346 326098 37582 326334
rect 37026 290418 37262 290654
rect 37346 290418 37582 290654
rect 37026 290098 37262 290334
rect 37346 290098 37582 290334
rect 37026 254418 37262 254654
rect 37346 254418 37582 254654
rect 37026 254098 37262 254334
rect 37346 254098 37582 254334
rect 37026 218418 37262 218654
rect 37346 218418 37582 218654
rect 37026 218098 37262 218334
rect 37346 218098 37582 218334
rect 37026 182418 37262 182654
rect 37346 182418 37582 182654
rect 37026 182098 37262 182334
rect 37346 182098 37582 182334
rect 37026 146418 37262 146654
rect 37346 146418 37582 146654
rect 37026 146098 37262 146334
rect 37346 146098 37582 146334
rect 37026 110418 37262 110654
rect 37346 110418 37582 110654
rect 37026 110098 37262 110334
rect 37346 110098 37582 110334
rect 37026 74418 37262 74654
rect 37346 74418 37582 74654
rect 37026 74098 37262 74334
rect 37346 74098 37582 74334
rect 37026 38418 37262 38654
rect 37346 38418 37582 38654
rect 37026 38098 37262 38334
rect 37346 38098 37582 38334
rect 37026 2418 37262 2654
rect 37346 2418 37582 2654
rect 37026 2098 37262 2334
rect 37346 2098 37582 2334
rect 37026 -582 37262 -346
rect 37346 -582 37582 -346
rect 37026 -902 37262 -666
rect 37346 -902 37582 -666
rect 38266 705562 38502 705798
rect 38586 705562 38822 705798
rect 38266 705242 38502 705478
rect 38586 705242 38822 705478
rect 38266 687658 38502 687894
rect 38586 687658 38822 687894
rect 38266 687338 38502 687574
rect 38586 687338 38822 687574
rect 38266 651658 38502 651894
rect 38586 651658 38822 651894
rect 38266 651338 38502 651574
rect 38586 651338 38822 651574
rect 38266 615658 38502 615894
rect 38586 615658 38822 615894
rect 38266 615338 38502 615574
rect 38586 615338 38822 615574
rect 38266 579658 38502 579894
rect 38586 579658 38822 579894
rect 38266 579338 38502 579574
rect 38586 579338 38822 579574
rect 38266 543658 38502 543894
rect 38586 543658 38822 543894
rect 38266 543338 38502 543574
rect 38586 543338 38822 543574
rect 38266 507658 38502 507894
rect 38586 507658 38822 507894
rect 38266 507338 38502 507574
rect 38586 507338 38822 507574
rect 38266 471658 38502 471894
rect 38586 471658 38822 471894
rect 38266 471338 38502 471574
rect 38586 471338 38822 471574
rect 38266 435658 38502 435894
rect 38586 435658 38822 435894
rect 38266 435338 38502 435574
rect 38586 435338 38822 435574
rect 38266 399658 38502 399894
rect 38586 399658 38822 399894
rect 38266 399338 38502 399574
rect 38586 399338 38822 399574
rect 38266 363658 38502 363894
rect 38586 363658 38822 363894
rect 38266 363338 38502 363574
rect 38586 363338 38822 363574
rect 38266 327658 38502 327894
rect 38586 327658 38822 327894
rect 38266 327338 38502 327574
rect 38586 327338 38822 327574
rect 38266 291658 38502 291894
rect 38586 291658 38822 291894
rect 38266 291338 38502 291574
rect 38586 291338 38822 291574
rect 38266 255658 38502 255894
rect 38586 255658 38822 255894
rect 38266 255338 38502 255574
rect 38586 255338 38822 255574
rect 38266 219658 38502 219894
rect 38586 219658 38822 219894
rect 38266 219338 38502 219574
rect 38586 219338 38822 219574
rect 38266 183658 38502 183894
rect 38586 183658 38822 183894
rect 38266 183338 38502 183574
rect 38586 183338 38822 183574
rect 38266 147658 38502 147894
rect 38586 147658 38822 147894
rect 38266 147338 38502 147574
rect 38586 147338 38822 147574
rect 38266 111658 38502 111894
rect 38586 111658 38822 111894
rect 38266 111338 38502 111574
rect 38586 111338 38822 111574
rect 38266 75658 38502 75894
rect 38586 75658 38822 75894
rect 38266 75338 38502 75574
rect 38586 75338 38822 75574
rect 38266 39658 38502 39894
rect 38586 39658 38822 39894
rect 38266 39338 38502 39574
rect 38586 39338 38822 39574
rect 38266 3658 38502 3894
rect 38586 3658 38822 3894
rect 38266 3338 38502 3574
rect 38586 3338 38822 3574
rect 38266 -1542 38502 -1306
rect 38586 -1542 38822 -1306
rect 38266 -1862 38502 -1626
rect 38586 -1862 38822 -1626
rect 39506 706522 39742 706758
rect 39826 706522 40062 706758
rect 39506 706202 39742 706438
rect 39826 706202 40062 706438
rect 39506 688898 39742 689134
rect 39826 688898 40062 689134
rect 39506 688578 39742 688814
rect 39826 688578 40062 688814
rect 39506 652898 39742 653134
rect 39826 652898 40062 653134
rect 39506 652578 39742 652814
rect 39826 652578 40062 652814
rect 39506 616898 39742 617134
rect 39826 616898 40062 617134
rect 39506 616578 39742 616814
rect 39826 616578 40062 616814
rect 39506 580898 39742 581134
rect 39826 580898 40062 581134
rect 39506 580578 39742 580814
rect 39826 580578 40062 580814
rect 39506 544898 39742 545134
rect 39826 544898 40062 545134
rect 39506 544578 39742 544814
rect 39826 544578 40062 544814
rect 39506 508898 39742 509134
rect 39826 508898 40062 509134
rect 39506 508578 39742 508814
rect 39826 508578 40062 508814
rect 39506 472898 39742 473134
rect 39826 472898 40062 473134
rect 39506 472578 39742 472814
rect 39826 472578 40062 472814
rect 39506 436898 39742 437134
rect 39826 436898 40062 437134
rect 39506 436578 39742 436814
rect 39826 436578 40062 436814
rect 39506 400898 39742 401134
rect 39826 400898 40062 401134
rect 39506 400578 39742 400814
rect 39826 400578 40062 400814
rect 39506 364898 39742 365134
rect 39826 364898 40062 365134
rect 39506 364578 39742 364814
rect 39826 364578 40062 364814
rect 39506 328898 39742 329134
rect 39826 328898 40062 329134
rect 39506 328578 39742 328814
rect 39826 328578 40062 328814
rect 39506 292898 39742 293134
rect 39826 292898 40062 293134
rect 39506 292578 39742 292814
rect 39826 292578 40062 292814
rect 39506 256898 39742 257134
rect 39826 256898 40062 257134
rect 39506 256578 39742 256814
rect 39826 256578 40062 256814
rect 39506 220898 39742 221134
rect 39826 220898 40062 221134
rect 39506 220578 39742 220814
rect 39826 220578 40062 220814
rect 39506 184898 39742 185134
rect 39826 184898 40062 185134
rect 39506 184578 39742 184814
rect 39826 184578 40062 184814
rect 39506 148898 39742 149134
rect 39826 148898 40062 149134
rect 39506 148578 39742 148814
rect 39826 148578 40062 148814
rect 39506 112898 39742 113134
rect 39826 112898 40062 113134
rect 39506 112578 39742 112814
rect 39826 112578 40062 112814
rect 39506 76898 39742 77134
rect 39826 76898 40062 77134
rect 39506 76578 39742 76814
rect 39826 76578 40062 76814
rect 39506 40898 39742 41134
rect 39826 40898 40062 41134
rect 39506 40578 39742 40814
rect 39826 40578 40062 40814
rect 39506 4898 39742 5134
rect 39826 4898 40062 5134
rect 39506 4578 39742 4814
rect 39826 4578 40062 4814
rect 39506 -2502 39742 -2266
rect 39826 -2502 40062 -2266
rect 39506 -2822 39742 -2586
rect 39826 -2822 40062 -2586
rect 40746 707482 40982 707718
rect 41066 707482 41302 707718
rect 40746 707162 40982 707398
rect 41066 707162 41302 707398
rect 40746 690138 40982 690374
rect 41066 690138 41302 690374
rect 40746 689818 40982 690054
rect 41066 689818 41302 690054
rect 40746 654138 40982 654374
rect 41066 654138 41302 654374
rect 40746 653818 40982 654054
rect 41066 653818 41302 654054
rect 40746 618138 40982 618374
rect 41066 618138 41302 618374
rect 40746 617818 40982 618054
rect 41066 617818 41302 618054
rect 40746 582138 40982 582374
rect 41066 582138 41302 582374
rect 40746 581818 40982 582054
rect 41066 581818 41302 582054
rect 40746 546138 40982 546374
rect 41066 546138 41302 546374
rect 40746 545818 40982 546054
rect 41066 545818 41302 546054
rect 40746 510138 40982 510374
rect 41066 510138 41302 510374
rect 40746 509818 40982 510054
rect 41066 509818 41302 510054
rect 40746 474138 40982 474374
rect 41066 474138 41302 474374
rect 40746 473818 40982 474054
rect 41066 473818 41302 474054
rect 40746 438138 40982 438374
rect 41066 438138 41302 438374
rect 40746 437818 40982 438054
rect 41066 437818 41302 438054
rect 40746 402138 40982 402374
rect 41066 402138 41302 402374
rect 40746 401818 40982 402054
rect 41066 401818 41302 402054
rect 40746 366138 40982 366374
rect 41066 366138 41302 366374
rect 40746 365818 40982 366054
rect 41066 365818 41302 366054
rect 40746 330138 40982 330374
rect 41066 330138 41302 330374
rect 40746 329818 40982 330054
rect 41066 329818 41302 330054
rect 40746 294138 40982 294374
rect 41066 294138 41302 294374
rect 40746 293818 40982 294054
rect 41066 293818 41302 294054
rect 40746 258138 40982 258374
rect 41066 258138 41302 258374
rect 40746 257818 40982 258054
rect 41066 257818 41302 258054
rect 40746 222138 40982 222374
rect 41066 222138 41302 222374
rect 40746 221818 40982 222054
rect 41066 221818 41302 222054
rect 40746 186138 40982 186374
rect 41066 186138 41302 186374
rect 40746 185818 40982 186054
rect 41066 185818 41302 186054
rect 40746 150138 40982 150374
rect 41066 150138 41302 150374
rect 40746 149818 40982 150054
rect 41066 149818 41302 150054
rect 40746 114138 40982 114374
rect 41066 114138 41302 114374
rect 40746 113818 40982 114054
rect 41066 113818 41302 114054
rect 40746 78138 40982 78374
rect 41066 78138 41302 78374
rect 40746 77818 40982 78054
rect 41066 77818 41302 78054
rect 40746 42138 40982 42374
rect 41066 42138 41302 42374
rect 40746 41818 40982 42054
rect 41066 41818 41302 42054
rect 40746 6138 40982 6374
rect 41066 6138 41302 6374
rect 40746 5818 40982 6054
rect 41066 5818 41302 6054
rect 40746 -3462 40982 -3226
rect 41066 -3462 41302 -3226
rect 40746 -3782 40982 -3546
rect 41066 -3782 41302 -3546
rect 41986 708442 42222 708678
rect 42306 708442 42542 708678
rect 41986 708122 42222 708358
rect 42306 708122 42542 708358
rect 41986 691378 42222 691614
rect 42306 691378 42542 691614
rect 41986 691058 42222 691294
rect 42306 691058 42542 691294
rect 41986 655378 42222 655614
rect 42306 655378 42542 655614
rect 41986 655058 42222 655294
rect 42306 655058 42542 655294
rect 41986 619378 42222 619614
rect 42306 619378 42542 619614
rect 41986 619058 42222 619294
rect 42306 619058 42542 619294
rect 41986 583378 42222 583614
rect 42306 583378 42542 583614
rect 41986 583058 42222 583294
rect 42306 583058 42542 583294
rect 41986 547378 42222 547614
rect 42306 547378 42542 547614
rect 41986 547058 42222 547294
rect 42306 547058 42542 547294
rect 41986 511378 42222 511614
rect 42306 511378 42542 511614
rect 41986 511058 42222 511294
rect 42306 511058 42542 511294
rect 41986 475378 42222 475614
rect 42306 475378 42542 475614
rect 41986 475058 42222 475294
rect 42306 475058 42542 475294
rect 41986 439378 42222 439614
rect 42306 439378 42542 439614
rect 41986 439058 42222 439294
rect 42306 439058 42542 439294
rect 41986 403378 42222 403614
rect 42306 403378 42542 403614
rect 41986 403058 42222 403294
rect 42306 403058 42542 403294
rect 41986 367378 42222 367614
rect 42306 367378 42542 367614
rect 41986 367058 42222 367294
rect 42306 367058 42542 367294
rect 41986 331378 42222 331614
rect 42306 331378 42542 331614
rect 41986 331058 42222 331294
rect 42306 331058 42542 331294
rect 41986 295378 42222 295614
rect 42306 295378 42542 295614
rect 41986 295058 42222 295294
rect 42306 295058 42542 295294
rect 41986 259378 42222 259614
rect 42306 259378 42542 259614
rect 41986 259058 42222 259294
rect 42306 259058 42542 259294
rect 41986 223378 42222 223614
rect 42306 223378 42542 223614
rect 41986 223058 42222 223294
rect 42306 223058 42542 223294
rect 41986 187378 42222 187614
rect 42306 187378 42542 187614
rect 41986 187058 42222 187294
rect 42306 187058 42542 187294
rect 41986 151378 42222 151614
rect 42306 151378 42542 151614
rect 41986 151058 42222 151294
rect 42306 151058 42542 151294
rect 41986 115378 42222 115614
rect 42306 115378 42542 115614
rect 41986 115058 42222 115294
rect 42306 115058 42542 115294
rect 41986 79378 42222 79614
rect 42306 79378 42542 79614
rect 41986 79058 42222 79294
rect 42306 79058 42542 79294
rect 41986 43378 42222 43614
rect 42306 43378 42542 43614
rect 41986 43058 42222 43294
rect 42306 43058 42542 43294
rect 41986 7378 42222 7614
rect 42306 7378 42542 7614
rect 41986 7058 42222 7294
rect 42306 7058 42542 7294
rect 41986 -4422 42222 -4186
rect 42306 -4422 42542 -4186
rect 41986 -4742 42222 -4506
rect 42306 -4742 42542 -4506
rect 43226 709402 43462 709638
rect 43546 709402 43782 709638
rect 43226 709082 43462 709318
rect 43546 709082 43782 709318
rect 43226 692618 43462 692854
rect 43546 692618 43782 692854
rect 43226 692298 43462 692534
rect 43546 692298 43782 692534
rect 43226 656618 43462 656854
rect 43546 656618 43782 656854
rect 43226 656298 43462 656534
rect 43546 656298 43782 656534
rect 43226 620618 43462 620854
rect 43546 620618 43782 620854
rect 43226 620298 43462 620534
rect 43546 620298 43782 620534
rect 43226 584618 43462 584854
rect 43546 584618 43782 584854
rect 43226 584298 43462 584534
rect 43546 584298 43782 584534
rect 43226 548618 43462 548854
rect 43546 548618 43782 548854
rect 43226 548298 43462 548534
rect 43546 548298 43782 548534
rect 43226 512618 43462 512854
rect 43546 512618 43782 512854
rect 43226 512298 43462 512534
rect 43546 512298 43782 512534
rect 43226 476618 43462 476854
rect 43546 476618 43782 476854
rect 43226 476298 43462 476534
rect 43546 476298 43782 476534
rect 43226 440618 43462 440854
rect 43546 440618 43782 440854
rect 43226 440298 43462 440534
rect 43546 440298 43782 440534
rect 43226 404618 43462 404854
rect 43546 404618 43782 404854
rect 43226 404298 43462 404534
rect 43546 404298 43782 404534
rect 43226 368618 43462 368854
rect 43546 368618 43782 368854
rect 43226 368298 43462 368534
rect 43546 368298 43782 368534
rect 43226 332618 43462 332854
rect 43546 332618 43782 332854
rect 43226 332298 43462 332534
rect 43546 332298 43782 332534
rect 43226 296618 43462 296854
rect 43546 296618 43782 296854
rect 43226 296298 43462 296534
rect 43546 296298 43782 296534
rect 43226 260618 43462 260854
rect 43546 260618 43782 260854
rect 43226 260298 43462 260534
rect 43546 260298 43782 260534
rect 43226 224618 43462 224854
rect 43546 224618 43782 224854
rect 43226 224298 43462 224534
rect 43546 224298 43782 224534
rect 43226 188618 43462 188854
rect 43546 188618 43782 188854
rect 43226 188298 43462 188534
rect 43546 188298 43782 188534
rect 43226 152618 43462 152854
rect 43546 152618 43782 152854
rect 43226 152298 43462 152534
rect 43546 152298 43782 152534
rect 43226 116618 43462 116854
rect 43546 116618 43782 116854
rect 43226 116298 43462 116534
rect 43546 116298 43782 116534
rect 43226 80618 43462 80854
rect 43546 80618 43782 80854
rect 43226 80298 43462 80534
rect 43546 80298 43782 80534
rect 43226 44618 43462 44854
rect 43546 44618 43782 44854
rect 43226 44298 43462 44534
rect 43546 44298 43782 44534
rect 43226 8618 43462 8854
rect 43546 8618 43782 8854
rect 43226 8298 43462 8534
rect 43546 8298 43782 8534
rect 43226 -5382 43462 -5146
rect 43546 -5382 43782 -5146
rect 43226 -5702 43462 -5466
rect 43546 -5702 43782 -5466
rect 44466 710362 44702 710598
rect 44786 710362 45022 710598
rect 44466 710042 44702 710278
rect 44786 710042 45022 710278
rect 44466 693858 44702 694094
rect 44786 693858 45022 694094
rect 44466 693538 44702 693774
rect 44786 693538 45022 693774
rect 44466 657858 44702 658094
rect 44786 657858 45022 658094
rect 44466 657538 44702 657774
rect 44786 657538 45022 657774
rect 44466 621858 44702 622094
rect 44786 621858 45022 622094
rect 44466 621538 44702 621774
rect 44786 621538 45022 621774
rect 44466 585858 44702 586094
rect 44786 585858 45022 586094
rect 44466 585538 44702 585774
rect 44786 585538 45022 585774
rect 44466 549858 44702 550094
rect 44786 549858 45022 550094
rect 44466 549538 44702 549774
rect 44786 549538 45022 549774
rect 44466 513858 44702 514094
rect 44786 513858 45022 514094
rect 44466 513538 44702 513774
rect 44786 513538 45022 513774
rect 44466 477858 44702 478094
rect 44786 477858 45022 478094
rect 44466 477538 44702 477774
rect 44786 477538 45022 477774
rect 44466 441858 44702 442094
rect 44786 441858 45022 442094
rect 44466 441538 44702 441774
rect 44786 441538 45022 441774
rect 44466 405858 44702 406094
rect 44786 405858 45022 406094
rect 44466 405538 44702 405774
rect 44786 405538 45022 405774
rect 44466 369858 44702 370094
rect 44786 369858 45022 370094
rect 44466 369538 44702 369774
rect 44786 369538 45022 369774
rect 44466 333858 44702 334094
rect 44786 333858 45022 334094
rect 44466 333538 44702 333774
rect 44786 333538 45022 333774
rect 44466 297858 44702 298094
rect 44786 297858 45022 298094
rect 44466 297538 44702 297774
rect 44786 297538 45022 297774
rect 44466 261858 44702 262094
rect 44786 261858 45022 262094
rect 44466 261538 44702 261774
rect 44786 261538 45022 261774
rect 44466 225858 44702 226094
rect 44786 225858 45022 226094
rect 44466 225538 44702 225774
rect 44786 225538 45022 225774
rect 44466 189858 44702 190094
rect 44786 189858 45022 190094
rect 44466 189538 44702 189774
rect 44786 189538 45022 189774
rect 44466 153858 44702 154094
rect 44786 153858 45022 154094
rect 44466 153538 44702 153774
rect 44786 153538 45022 153774
rect 44466 117858 44702 118094
rect 44786 117858 45022 118094
rect 44466 117538 44702 117774
rect 44786 117538 45022 117774
rect 44466 81858 44702 82094
rect 44786 81858 45022 82094
rect 44466 81538 44702 81774
rect 44786 81538 45022 81774
rect 44466 45858 44702 46094
rect 44786 45858 45022 46094
rect 44466 45538 44702 45774
rect 44786 45538 45022 45774
rect 44466 9858 44702 10094
rect 44786 9858 45022 10094
rect 44466 9538 44702 9774
rect 44786 9538 45022 9774
rect 44466 -6342 44702 -6106
rect 44786 -6342 45022 -6106
rect 44466 -6662 44702 -6426
rect 44786 -6662 45022 -6426
rect 45706 711322 45942 711558
rect 46026 711322 46262 711558
rect 45706 711002 45942 711238
rect 46026 711002 46262 711238
rect 45706 695098 45942 695334
rect 46026 695098 46262 695334
rect 45706 694778 45942 695014
rect 46026 694778 46262 695014
rect 45706 659098 45942 659334
rect 46026 659098 46262 659334
rect 45706 658778 45942 659014
rect 46026 658778 46262 659014
rect 45706 623098 45942 623334
rect 46026 623098 46262 623334
rect 45706 622778 45942 623014
rect 46026 622778 46262 623014
rect 45706 587098 45942 587334
rect 46026 587098 46262 587334
rect 45706 586778 45942 587014
rect 46026 586778 46262 587014
rect 45706 551098 45942 551334
rect 46026 551098 46262 551334
rect 45706 550778 45942 551014
rect 46026 550778 46262 551014
rect 45706 515098 45942 515334
rect 46026 515098 46262 515334
rect 45706 514778 45942 515014
rect 46026 514778 46262 515014
rect 45706 479098 45942 479334
rect 46026 479098 46262 479334
rect 45706 478778 45942 479014
rect 46026 478778 46262 479014
rect 45706 443098 45942 443334
rect 46026 443098 46262 443334
rect 45706 442778 45942 443014
rect 46026 442778 46262 443014
rect 45706 407098 45942 407334
rect 46026 407098 46262 407334
rect 45706 406778 45942 407014
rect 46026 406778 46262 407014
rect 45706 371098 45942 371334
rect 46026 371098 46262 371334
rect 45706 370778 45942 371014
rect 46026 370778 46262 371014
rect 45706 335098 45942 335334
rect 46026 335098 46262 335334
rect 45706 334778 45942 335014
rect 46026 334778 46262 335014
rect 45706 299098 45942 299334
rect 46026 299098 46262 299334
rect 45706 298778 45942 299014
rect 46026 298778 46262 299014
rect 45706 263098 45942 263334
rect 46026 263098 46262 263334
rect 45706 262778 45942 263014
rect 46026 262778 46262 263014
rect 45706 227098 45942 227334
rect 46026 227098 46262 227334
rect 45706 226778 45942 227014
rect 46026 226778 46262 227014
rect 45706 191098 45942 191334
rect 46026 191098 46262 191334
rect 45706 190778 45942 191014
rect 46026 190778 46262 191014
rect 45706 155098 45942 155334
rect 46026 155098 46262 155334
rect 45706 154778 45942 155014
rect 46026 154778 46262 155014
rect 45706 119098 45942 119334
rect 46026 119098 46262 119334
rect 45706 118778 45942 119014
rect 46026 118778 46262 119014
rect 45706 83098 45942 83334
rect 46026 83098 46262 83334
rect 45706 82778 45942 83014
rect 46026 82778 46262 83014
rect 45706 47098 45942 47334
rect 46026 47098 46262 47334
rect 45706 46778 45942 47014
rect 46026 46778 46262 47014
rect 45706 11098 45942 11334
rect 46026 11098 46262 11334
rect 45706 10778 45942 11014
rect 46026 10778 46262 11014
rect 45706 -7302 45942 -7066
rect 46026 -7302 46262 -7066
rect 45706 -7622 45942 -7386
rect 46026 -7622 46262 -7386
rect 73026 704602 73262 704838
rect 73346 704602 73582 704838
rect 73026 704282 73262 704518
rect 73346 704282 73582 704518
rect 73026 686418 73262 686654
rect 73346 686418 73582 686654
rect 73026 686098 73262 686334
rect 73346 686098 73582 686334
rect 73026 650418 73262 650654
rect 73346 650418 73582 650654
rect 73026 650098 73262 650334
rect 73346 650098 73582 650334
rect 73026 614418 73262 614654
rect 73346 614418 73582 614654
rect 73026 614098 73262 614334
rect 73346 614098 73582 614334
rect 73026 578418 73262 578654
rect 73346 578418 73582 578654
rect 73026 578098 73262 578334
rect 73346 578098 73582 578334
rect 73026 542418 73262 542654
rect 73346 542418 73582 542654
rect 73026 542098 73262 542334
rect 73346 542098 73582 542334
rect 73026 506418 73262 506654
rect 73346 506418 73582 506654
rect 73026 506098 73262 506334
rect 73346 506098 73582 506334
rect 73026 470418 73262 470654
rect 73346 470418 73582 470654
rect 73026 470098 73262 470334
rect 73346 470098 73582 470334
rect 73026 434418 73262 434654
rect 73346 434418 73582 434654
rect 73026 434098 73262 434334
rect 73346 434098 73582 434334
rect 73026 398418 73262 398654
rect 73346 398418 73582 398654
rect 73026 398098 73262 398334
rect 73346 398098 73582 398334
rect 73026 362418 73262 362654
rect 73346 362418 73582 362654
rect 73026 362098 73262 362334
rect 73346 362098 73582 362334
rect 73026 326418 73262 326654
rect 73346 326418 73582 326654
rect 73026 326098 73262 326334
rect 73346 326098 73582 326334
rect 73026 290418 73262 290654
rect 73346 290418 73582 290654
rect 73026 290098 73262 290334
rect 73346 290098 73582 290334
rect 73026 254418 73262 254654
rect 73346 254418 73582 254654
rect 73026 254098 73262 254334
rect 73346 254098 73582 254334
rect 73026 218418 73262 218654
rect 73346 218418 73582 218654
rect 73026 218098 73262 218334
rect 73346 218098 73582 218334
rect 73026 182418 73262 182654
rect 73346 182418 73582 182654
rect 73026 182098 73262 182334
rect 73346 182098 73582 182334
rect 73026 146418 73262 146654
rect 73346 146418 73582 146654
rect 73026 146098 73262 146334
rect 73346 146098 73582 146334
rect 73026 110418 73262 110654
rect 73346 110418 73582 110654
rect 73026 110098 73262 110334
rect 73346 110098 73582 110334
rect 73026 74418 73262 74654
rect 73346 74418 73582 74654
rect 73026 74098 73262 74334
rect 73346 74098 73582 74334
rect 73026 38418 73262 38654
rect 73346 38418 73582 38654
rect 73026 38098 73262 38334
rect 73346 38098 73582 38334
rect 73026 2418 73262 2654
rect 73346 2418 73582 2654
rect 73026 2098 73262 2334
rect 73346 2098 73582 2334
rect 73026 -582 73262 -346
rect 73346 -582 73582 -346
rect 73026 -902 73262 -666
rect 73346 -902 73582 -666
rect 74266 705562 74502 705798
rect 74586 705562 74822 705798
rect 74266 705242 74502 705478
rect 74586 705242 74822 705478
rect 74266 687658 74502 687894
rect 74586 687658 74822 687894
rect 74266 687338 74502 687574
rect 74586 687338 74822 687574
rect 74266 651658 74502 651894
rect 74586 651658 74822 651894
rect 74266 651338 74502 651574
rect 74586 651338 74822 651574
rect 74266 615658 74502 615894
rect 74586 615658 74822 615894
rect 74266 615338 74502 615574
rect 74586 615338 74822 615574
rect 74266 579658 74502 579894
rect 74586 579658 74822 579894
rect 74266 579338 74502 579574
rect 74586 579338 74822 579574
rect 74266 543658 74502 543894
rect 74586 543658 74822 543894
rect 74266 543338 74502 543574
rect 74586 543338 74822 543574
rect 74266 507658 74502 507894
rect 74586 507658 74822 507894
rect 74266 507338 74502 507574
rect 74586 507338 74822 507574
rect 74266 471658 74502 471894
rect 74586 471658 74822 471894
rect 74266 471338 74502 471574
rect 74586 471338 74822 471574
rect 74266 435658 74502 435894
rect 74586 435658 74822 435894
rect 74266 435338 74502 435574
rect 74586 435338 74822 435574
rect 74266 399658 74502 399894
rect 74586 399658 74822 399894
rect 74266 399338 74502 399574
rect 74586 399338 74822 399574
rect 74266 363658 74502 363894
rect 74586 363658 74822 363894
rect 74266 363338 74502 363574
rect 74586 363338 74822 363574
rect 74266 327658 74502 327894
rect 74586 327658 74822 327894
rect 74266 327338 74502 327574
rect 74586 327338 74822 327574
rect 74266 291658 74502 291894
rect 74586 291658 74822 291894
rect 74266 291338 74502 291574
rect 74586 291338 74822 291574
rect 74266 255658 74502 255894
rect 74586 255658 74822 255894
rect 74266 255338 74502 255574
rect 74586 255338 74822 255574
rect 74266 219658 74502 219894
rect 74586 219658 74822 219894
rect 74266 219338 74502 219574
rect 74586 219338 74822 219574
rect 74266 183658 74502 183894
rect 74586 183658 74822 183894
rect 74266 183338 74502 183574
rect 74586 183338 74822 183574
rect 74266 147658 74502 147894
rect 74586 147658 74822 147894
rect 74266 147338 74502 147574
rect 74586 147338 74822 147574
rect 74266 111658 74502 111894
rect 74586 111658 74822 111894
rect 74266 111338 74502 111574
rect 74586 111338 74822 111574
rect 74266 75658 74502 75894
rect 74586 75658 74822 75894
rect 74266 75338 74502 75574
rect 74586 75338 74822 75574
rect 74266 39658 74502 39894
rect 74586 39658 74822 39894
rect 74266 39338 74502 39574
rect 74586 39338 74822 39574
rect 74266 3658 74502 3894
rect 74586 3658 74822 3894
rect 74266 3338 74502 3574
rect 74586 3338 74822 3574
rect 74266 -1542 74502 -1306
rect 74586 -1542 74822 -1306
rect 74266 -1862 74502 -1626
rect 74586 -1862 74822 -1626
rect 75506 706522 75742 706758
rect 75826 706522 76062 706758
rect 75506 706202 75742 706438
rect 75826 706202 76062 706438
rect 75506 688898 75742 689134
rect 75826 688898 76062 689134
rect 75506 688578 75742 688814
rect 75826 688578 76062 688814
rect 75506 652898 75742 653134
rect 75826 652898 76062 653134
rect 75506 652578 75742 652814
rect 75826 652578 76062 652814
rect 75506 616898 75742 617134
rect 75826 616898 76062 617134
rect 75506 616578 75742 616814
rect 75826 616578 76062 616814
rect 75506 580898 75742 581134
rect 75826 580898 76062 581134
rect 75506 580578 75742 580814
rect 75826 580578 76062 580814
rect 75506 544898 75742 545134
rect 75826 544898 76062 545134
rect 75506 544578 75742 544814
rect 75826 544578 76062 544814
rect 75506 508898 75742 509134
rect 75826 508898 76062 509134
rect 75506 508578 75742 508814
rect 75826 508578 76062 508814
rect 75506 472898 75742 473134
rect 75826 472898 76062 473134
rect 75506 472578 75742 472814
rect 75826 472578 76062 472814
rect 75506 436898 75742 437134
rect 75826 436898 76062 437134
rect 75506 436578 75742 436814
rect 75826 436578 76062 436814
rect 75506 400898 75742 401134
rect 75826 400898 76062 401134
rect 75506 400578 75742 400814
rect 75826 400578 76062 400814
rect 75506 364898 75742 365134
rect 75826 364898 76062 365134
rect 75506 364578 75742 364814
rect 75826 364578 76062 364814
rect 75506 328898 75742 329134
rect 75826 328898 76062 329134
rect 75506 328578 75742 328814
rect 75826 328578 76062 328814
rect 75506 292898 75742 293134
rect 75826 292898 76062 293134
rect 75506 292578 75742 292814
rect 75826 292578 76062 292814
rect 75506 256898 75742 257134
rect 75826 256898 76062 257134
rect 75506 256578 75742 256814
rect 75826 256578 76062 256814
rect 75506 220898 75742 221134
rect 75826 220898 76062 221134
rect 75506 220578 75742 220814
rect 75826 220578 76062 220814
rect 75506 184898 75742 185134
rect 75826 184898 76062 185134
rect 75506 184578 75742 184814
rect 75826 184578 76062 184814
rect 75506 148898 75742 149134
rect 75826 148898 76062 149134
rect 75506 148578 75742 148814
rect 75826 148578 76062 148814
rect 75506 112898 75742 113134
rect 75826 112898 76062 113134
rect 75506 112578 75742 112814
rect 75826 112578 76062 112814
rect 75506 76898 75742 77134
rect 75826 76898 76062 77134
rect 75506 76578 75742 76814
rect 75826 76578 76062 76814
rect 75506 40898 75742 41134
rect 75826 40898 76062 41134
rect 75506 40578 75742 40814
rect 75826 40578 76062 40814
rect 75506 4898 75742 5134
rect 75826 4898 76062 5134
rect 75506 4578 75742 4814
rect 75826 4578 76062 4814
rect 75506 -2502 75742 -2266
rect 75826 -2502 76062 -2266
rect 75506 -2822 75742 -2586
rect 75826 -2822 76062 -2586
rect 76746 707482 76982 707718
rect 77066 707482 77302 707718
rect 76746 707162 76982 707398
rect 77066 707162 77302 707398
rect 76746 690138 76982 690374
rect 77066 690138 77302 690374
rect 76746 689818 76982 690054
rect 77066 689818 77302 690054
rect 76746 654138 76982 654374
rect 77066 654138 77302 654374
rect 76746 653818 76982 654054
rect 77066 653818 77302 654054
rect 76746 618138 76982 618374
rect 77066 618138 77302 618374
rect 76746 617818 76982 618054
rect 77066 617818 77302 618054
rect 76746 582138 76982 582374
rect 77066 582138 77302 582374
rect 76746 581818 76982 582054
rect 77066 581818 77302 582054
rect 76746 546138 76982 546374
rect 77066 546138 77302 546374
rect 76746 545818 76982 546054
rect 77066 545818 77302 546054
rect 76746 510138 76982 510374
rect 77066 510138 77302 510374
rect 76746 509818 76982 510054
rect 77066 509818 77302 510054
rect 76746 474138 76982 474374
rect 77066 474138 77302 474374
rect 76746 473818 76982 474054
rect 77066 473818 77302 474054
rect 76746 438138 76982 438374
rect 77066 438138 77302 438374
rect 76746 437818 76982 438054
rect 77066 437818 77302 438054
rect 76746 402138 76982 402374
rect 77066 402138 77302 402374
rect 76746 401818 76982 402054
rect 77066 401818 77302 402054
rect 76746 366138 76982 366374
rect 77066 366138 77302 366374
rect 76746 365818 76982 366054
rect 77066 365818 77302 366054
rect 76746 330138 76982 330374
rect 77066 330138 77302 330374
rect 76746 329818 76982 330054
rect 77066 329818 77302 330054
rect 76746 294138 76982 294374
rect 77066 294138 77302 294374
rect 76746 293818 76982 294054
rect 77066 293818 77302 294054
rect 76746 258138 76982 258374
rect 77066 258138 77302 258374
rect 76746 257818 76982 258054
rect 77066 257818 77302 258054
rect 76746 222138 76982 222374
rect 77066 222138 77302 222374
rect 76746 221818 76982 222054
rect 77066 221818 77302 222054
rect 76746 186138 76982 186374
rect 77066 186138 77302 186374
rect 76746 185818 76982 186054
rect 77066 185818 77302 186054
rect 76746 150138 76982 150374
rect 77066 150138 77302 150374
rect 76746 149818 76982 150054
rect 77066 149818 77302 150054
rect 76746 114138 76982 114374
rect 77066 114138 77302 114374
rect 76746 113818 76982 114054
rect 77066 113818 77302 114054
rect 76746 78138 76982 78374
rect 77066 78138 77302 78374
rect 76746 77818 76982 78054
rect 77066 77818 77302 78054
rect 76746 42138 76982 42374
rect 77066 42138 77302 42374
rect 76746 41818 76982 42054
rect 77066 41818 77302 42054
rect 76746 6138 76982 6374
rect 77066 6138 77302 6374
rect 76746 5818 76982 6054
rect 77066 5818 77302 6054
rect 76746 -3462 76982 -3226
rect 77066 -3462 77302 -3226
rect 76746 -3782 76982 -3546
rect 77066 -3782 77302 -3546
rect 77986 708442 78222 708678
rect 78306 708442 78542 708678
rect 77986 708122 78222 708358
rect 78306 708122 78542 708358
rect 77986 691378 78222 691614
rect 78306 691378 78542 691614
rect 77986 691058 78222 691294
rect 78306 691058 78542 691294
rect 77986 655378 78222 655614
rect 78306 655378 78542 655614
rect 77986 655058 78222 655294
rect 78306 655058 78542 655294
rect 77986 619378 78222 619614
rect 78306 619378 78542 619614
rect 77986 619058 78222 619294
rect 78306 619058 78542 619294
rect 77986 583378 78222 583614
rect 78306 583378 78542 583614
rect 77986 583058 78222 583294
rect 78306 583058 78542 583294
rect 77986 547378 78222 547614
rect 78306 547378 78542 547614
rect 77986 547058 78222 547294
rect 78306 547058 78542 547294
rect 77986 511378 78222 511614
rect 78306 511378 78542 511614
rect 77986 511058 78222 511294
rect 78306 511058 78542 511294
rect 77986 475378 78222 475614
rect 78306 475378 78542 475614
rect 77986 475058 78222 475294
rect 78306 475058 78542 475294
rect 77986 439378 78222 439614
rect 78306 439378 78542 439614
rect 77986 439058 78222 439294
rect 78306 439058 78542 439294
rect 77986 403378 78222 403614
rect 78306 403378 78542 403614
rect 77986 403058 78222 403294
rect 78306 403058 78542 403294
rect 77986 367378 78222 367614
rect 78306 367378 78542 367614
rect 77986 367058 78222 367294
rect 78306 367058 78542 367294
rect 77986 331378 78222 331614
rect 78306 331378 78542 331614
rect 77986 331058 78222 331294
rect 78306 331058 78542 331294
rect 77986 295378 78222 295614
rect 78306 295378 78542 295614
rect 77986 295058 78222 295294
rect 78306 295058 78542 295294
rect 77986 259378 78222 259614
rect 78306 259378 78542 259614
rect 77986 259058 78222 259294
rect 78306 259058 78542 259294
rect 77986 223378 78222 223614
rect 78306 223378 78542 223614
rect 77986 223058 78222 223294
rect 78306 223058 78542 223294
rect 77986 187378 78222 187614
rect 78306 187378 78542 187614
rect 77986 187058 78222 187294
rect 78306 187058 78542 187294
rect 77986 151378 78222 151614
rect 78306 151378 78542 151614
rect 77986 151058 78222 151294
rect 78306 151058 78542 151294
rect 77986 115378 78222 115614
rect 78306 115378 78542 115614
rect 77986 115058 78222 115294
rect 78306 115058 78542 115294
rect 77986 79378 78222 79614
rect 78306 79378 78542 79614
rect 77986 79058 78222 79294
rect 78306 79058 78542 79294
rect 77986 43378 78222 43614
rect 78306 43378 78542 43614
rect 77986 43058 78222 43294
rect 78306 43058 78542 43294
rect 77986 7378 78222 7614
rect 78306 7378 78542 7614
rect 77986 7058 78222 7294
rect 78306 7058 78542 7294
rect 77986 -4422 78222 -4186
rect 78306 -4422 78542 -4186
rect 77986 -4742 78222 -4506
rect 78306 -4742 78542 -4506
rect 79226 709402 79462 709638
rect 79546 709402 79782 709638
rect 79226 709082 79462 709318
rect 79546 709082 79782 709318
rect 79226 692618 79462 692854
rect 79546 692618 79782 692854
rect 79226 692298 79462 692534
rect 79546 692298 79782 692534
rect 79226 656618 79462 656854
rect 79546 656618 79782 656854
rect 79226 656298 79462 656534
rect 79546 656298 79782 656534
rect 79226 620618 79462 620854
rect 79546 620618 79782 620854
rect 79226 620298 79462 620534
rect 79546 620298 79782 620534
rect 79226 584618 79462 584854
rect 79546 584618 79782 584854
rect 79226 584298 79462 584534
rect 79546 584298 79782 584534
rect 79226 548618 79462 548854
rect 79546 548618 79782 548854
rect 79226 548298 79462 548534
rect 79546 548298 79782 548534
rect 79226 512618 79462 512854
rect 79546 512618 79782 512854
rect 79226 512298 79462 512534
rect 79546 512298 79782 512534
rect 79226 476618 79462 476854
rect 79546 476618 79782 476854
rect 79226 476298 79462 476534
rect 79546 476298 79782 476534
rect 79226 440618 79462 440854
rect 79546 440618 79782 440854
rect 79226 440298 79462 440534
rect 79546 440298 79782 440534
rect 79226 404618 79462 404854
rect 79546 404618 79782 404854
rect 79226 404298 79462 404534
rect 79546 404298 79782 404534
rect 79226 368618 79462 368854
rect 79546 368618 79782 368854
rect 79226 368298 79462 368534
rect 79546 368298 79782 368534
rect 79226 332618 79462 332854
rect 79546 332618 79782 332854
rect 79226 332298 79462 332534
rect 79546 332298 79782 332534
rect 79226 296618 79462 296854
rect 79546 296618 79782 296854
rect 79226 296298 79462 296534
rect 79546 296298 79782 296534
rect 79226 260618 79462 260854
rect 79546 260618 79782 260854
rect 79226 260298 79462 260534
rect 79546 260298 79782 260534
rect 79226 224618 79462 224854
rect 79546 224618 79782 224854
rect 79226 224298 79462 224534
rect 79546 224298 79782 224534
rect 79226 188618 79462 188854
rect 79546 188618 79782 188854
rect 79226 188298 79462 188534
rect 79546 188298 79782 188534
rect 79226 152618 79462 152854
rect 79546 152618 79782 152854
rect 79226 152298 79462 152534
rect 79546 152298 79782 152534
rect 79226 116618 79462 116854
rect 79546 116618 79782 116854
rect 79226 116298 79462 116534
rect 79546 116298 79782 116534
rect 79226 80618 79462 80854
rect 79546 80618 79782 80854
rect 79226 80298 79462 80534
rect 79546 80298 79782 80534
rect 79226 44618 79462 44854
rect 79546 44618 79782 44854
rect 79226 44298 79462 44534
rect 79546 44298 79782 44534
rect 79226 8618 79462 8854
rect 79546 8618 79782 8854
rect 79226 8298 79462 8534
rect 79546 8298 79782 8534
rect 79226 -5382 79462 -5146
rect 79546 -5382 79782 -5146
rect 79226 -5702 79462 -5466
rect 79546 -5702 79782 -5466
rect 80466 710362 80702 710598
rect 80786 710362 81022 710598
rect 80466 710042 80702 710278
rect 80786 710042 81022 710278
rect 80466 693858 80702 694094
rect 80786 693858 81022 694094
rect 80466 693538 80702 693774
rect 80786 693538 81022 693774
rect 80466 657858 80702 658094
rect 80786 657858 81022 658094
rect 80466 657538 80702 657774
rect 80786 657538 81022 657774
rect 80466 621858 80702 622094
rect 80786 621858 81022 622094
rect 80466 621538 80702 621774
rect 80786 621538 81022 621774
rect 80466 585858 80702 586094
rect 80786 585858 81022 586094
rect 80466 585538 80702 585774
rect 80786 585538 81022 585774
rect 80466 549858 80702 550094
rect 80786 549858 81022 550094
rect 80466 549538 80702 549774
rect 80786 549538 81022 549774
rect 80466 513858 80702 514094
rect 80786 513858 81022 514094
rect 80466 513538 80702 513774
rect 80786 513538 81022 513774
rect 80466 477858 80702 478094
rect 80786 477858 81022 478094
rect 80466 477538 80702 477774
rect 80786 477538 81022 477774
rect 80466 441858 80702 442094
rect 80786 441858 81022 442094
rect 80466 441538 80702 441774
rect 80786 441538 81022 441774
rect 80466 405858 80702 406094
rect 80786 405858 81022 406094
rect 80466 405538 80702 405774
rect 80786 405538 81022 405774
rect 80466 369858 80702 370094
rect 80786 369858 81022 370094
rect 80466 369538 80702 369774
rect 80786 369538 81022 369774
rect 80466 333858 80702 334094
rect 80786 333858 81022 334094
rect 80466 333538 80702 333774
rect 80786 333538 81022 333774
rect 80466 297858 80702 298094
rect 80786 297858 81022 298094
rect 80466 297538 80702 297774
rect 80786 297538 81022 297774
rect 80466 261858 80702 262094
rect 80786 261858 81022 262094
rect 80466 261538 80702 261774
rect 80786 261538 81022 261774
rect 80466 225858 80702 226094
rect 80786 225858 81022 226094
rect 80466 225538 80702 225774
rect 80786 225538 81022 225774
rect 80466 189858 80702 190094
rect 80786 189858 81022 190094
rect 80466 189538 80702 189774
rect 80786 189538 81022 189774
rect 80466 153858 80702 154094
rect 80786 153858 81022 154094
rect 80466 153538 80702 153774
rect 80786 153538 81022 153774
rect 80466 117858 80702 118094
rect 80786 117858 81022 118094
rect 80466 117538 80702 117774
rect 80786 117538 81022 117774
rect 80466 81858 80702 82094
rect 80786 81858 81022 82094
rect 80466 81538 80702 81774
rect 80786 81538 81022 81774
rect 80466 45858 80702 46094
rect 80786 45858 81022 46094
rect 80466 45538 80702 45774
rect 80786 45538 81022 45774
rect 80466 9858 80702 10094
rect 80786 9858 81022 10094
rect 80466 9538 80702 9774
rect 80786 9538 81022 9774
rect 80466 -6342 80702 -6106
rect 80786 -6342 81022 -6106
rect 80466 -6662 80702 -6426
rect 80786 -6662 81022 -6426
rect 81706 711322 81942 711558
rect 82026 711322 82262 711558
rect 81706 711002 81942 711238
rect 82026 711002 82262 711238
rect 81706 695098 81942 695334
rect 82026 695098 82262 695334
rect 81706 694778 81942 695014
rect 82026 694778 82262 695014
rect 81706 659098 81942 659334
rect 82026 659098 82262 659334
rect 81706 658778 81942 659014
rect 82026 658778 82262 659014
rect 81706 623098 81942 623334
rect 82026 623098 82262 623334
rect 81706 622778 81942 623014
rect 82026 622778 82262 623014
rect 81706 587098 81942 587334
rect 82026 587098 82262 587334
rect 81706 586778 81942 587014
rect 82026 586778 82262 587014
rect 81706 551098 81942 551334
rect 82026 551098 82262 551334
rect 81706 550778 81942 551014
rect 82026 550778 82262 551014
rect 81706 515098 81942 515334
rect 82026 515098 82262 515334
rect 81706 514778 81942 515014
rect 82026 514778 82262 515014
rect 81706 479098 81942 479334
rect 82026 479098 82262 479334
rect 81706 478778 81942 479014
rect 82026 478778 82262 479014
rect 81706 443098 81942 443334
rect 82026 443098 82262 443334
rect 81706 442778 81942 443014
rect 82026 442778 82262 443014
rect 81706 407098 81942 407334
rect 82026 407098 82262 407334
rect 81706 406778 81942 407014
rect 82026 406778 82262 407014
rect 81706 371098 81942 371334
rect 82026 371098 82262 371334
rect 81706 370778 81942 371014
rect 82026 370778 82262 371014
rect 81706 335098 81942 335334
rect 82026 335098 82262 335334
rect 81706 334778 81942 335014
rect 82026 334778 82262 335014
rect 81706 299098 81942 299334
rect 82026 299098 82262 299334
rect 81706 298778 81942 299014
rect 82026 298778 82262 299014
rect 81706 263098 81942 263334
rect 82026 263098 82262 263334
rect 81706 262778 81942 263014
rect 82026 262778 82262 263014
rect 81706 227098 81942 227334
rect 82026 227098 82262 227334
rect 81706 226778 81942 227014
rect 82026 226778 82262 227014
rect 81706 191098 81942 191334
rect 82026 191098 82262 191334
rect 81706 190778 81942 191014
rect 82026 190778 82262 191014
rect 81706 155098 81942 155334
rect 82026 155098 82262 155334
rect 81706 154778 81942 155014
rect 82026 154778 82262 155014
rect 81706 119098 81942 119334
rect 82026 119098 82262 119334
rect 81706 118778 81942 119014
rect 82026 118778 82262 119014
rect 81706 83098 81942 83334
rect 82026 83098 82262 83334
rect 81706 82778 81942 83014
rect 82026 82778 82262 83014
rect 81706 47098 81942 47334
rect 82026 47098 82262 47334
rect 81706 46778 81942 47014
rect 82026 46778 82262 47014
rect 81706 11098 81942 11334
rect 82026 11098 82262 11334
rect 81706 10778 81942 11014
rect 82026 10778 82262 11014
rect 81706 -7302 81942 -7066
rect 82026 -7302 82262 -7066
rect 81706 -7622 81942 -7386
rect 82026 -7622 82262 -7386
rect 109026 704602 109262 704838
rect 109346 704602 109582 704838
rect 109026 704282 109262 704518
rect 109346 704282 109582 704518
rect 109026 686418 109262 686654
rect 109346 686418 109582 686654
rect 109026 686098 109262 686334
rect 109346 686098 109582 686334
rect 109026 650418 109262 650654
rect 109346 650418 109582 650654
rect 109026 650098 109262 650334
rect 109346 650098 109582 650334
rect 109026 614418 109262 614654
rect 109346 614418 109582 614654
rect 109026 614098 109262 614334
rect 109346 614098 109582 614334
rect 109026 578418 109262 578654
rect 109346 578418 109582 578654
rect 109026 578098 109262 578334
rect 109346 578098 109582 578334
rect 109026 542418 109262 542654
rect 109346 542418 109582 542654
rect 109026 542098 109262 542334
rect 109346 542098 109582 542334
rect 109026 506418 109262 506654
rect 109346 506418 109582 506654
rect 109026 506098 109262 506334
rect 109346 506098 109582 506334
rect 109026 470418 109262 470654
rect 109346 470418 109582 470654
rect 109026 470098 109262 470334
rect 109346 470098 109582 470334
rect 109026 434418 109262 434654
rect 109346 434418 109582 434654
rect 109026 434098 109262 434334
rect 109346 434098 109582 434334
rect 109026 398418 109262 398654
rect 109346 398418 109582 398654
rect 109026 398098 109262 398334
rect 109346 398098 109582 398334
rect 109026 362418 109262 362654
rect 109346 362418 109582 362654
rect 109026 362098 109262 362334
rect 109346 362098 109582 362334
rect 109026 326418 109262 326654
rect 109346 326418 109582 326654
rect 109026 326098 109262 326334
rect 109346 326098 109582 326334
rect 109026 290418 109262 290654
rect 109346 290418 109582 290654
rect 109026 290098 109262 290334
rect 109346 290098 109582 290334
rect 109026 254418 109262 254654
rect 109346 254418 109582 254654
rect 109026 254098 109262 254334
rect 109346 254098 109582 254334
rect 109026 218418 109262 218654
rect 109346 218418 109582 218654
rect 109026 218098 109262 218334
rect 109346 218098 109582 218334
rect 109026 182418 109262 182654
rect 109346 182418 109582 182654
rect 109026 182098 109262 182334
rect 109346 182098 109582 182334
rect 109026 146418 109262 146654
rect 109346 146418 109582 146654
rect 109026 146098 109262 146334
rect 109346 146098 109582 146334
rect 109026 110418 109262 110654
rect 109346 110418 109582 110654
rect 109026 110098 109262 110334
rect 109346 110098 109582 110334
rect 109026 74418 109262 74654
rect 109346 74418 109582 74654
rect 109026 74098 109262 74334
rect 109346 74098 109582 74334
rect 109026 38418 109262 38654
rect 109346 38418 109582 38654
rect 109026 38098 109262 38334
rect 109346 38098 109582 38334
rect 109026 2418 109262 2654
rect 109346 2418 109582 2654
rect 109026 2098 109262 2334
rect 109346 2098 109582 2334
rect 109026 -582 109262 -346
rect 109346 -582 109582 -346
rect 109026 -902 109262 -666
rect 109346 -902 109582 -666
rect 110266 705562 110502 705798
rect 110586 705562 110822 705798
rect 110266 705242 110502 705478
rect 110586 705242 110822 705478
rect 110266 687658 110502 687894
rect 110586 687658 110822 687894
rect 110266 687338 110502 687574
rect 110586 687338 110822 687574
rect 110266 651658 110502 651894
rect 110586 651658 110822 651894
rect 110266 651338 110502 651574
rect 110586 651338 110822 651574
rect 110266 615658 110502 615894
rect 110586 615658 110822 615894
rect 110266 615338 110502 615574
rect 110586 615338 110822 615574
rect 110266 579658 110502 579894
rect 110586 579658 110822 579894
rect 110266 579338 110502 579574
rect 110586 579338 110822 579574
rect 110266 543658 110502 543894
rect 110586 543658 110822 543894
rect 110266 543338 110502 543574
rect 110586 543338 110822 543574
rect 110266 507658 110502 507894
rect 110586 507658 110822 507894
rect 110266 507338 110502 507574
rect 110586 507338 110822 507574
rect 110266 471658 110502 471894
rect 110586 471658 110822 471894
rect 110266 471338 110502 471574
rect 110586 471338 110822 471574
rect 110266 435658 110502 435894
rect 110586 435658 110822 435894
rect 110266 435338 110502 435574
rect 110586 435338 110822 435574
rect 110266 399658 110502 399894
rect 110586 399658 110822 399894
rect 110266 399338 110502 399574
rect 110586 399338 110822 399574
rect 110266 363658 110502 363894
rect 110586 363658 110822 363894
rect 110266 363338 110502 363574
rect 110586 363338 110822 363574
rect 110266 327658 110502 327894
rect 110586 327658 110822 327894
rect 110266 327338 110502 327574
rect 110586 327338 110822 327574
rect 110266 291658 110502 291894
rect 110586 291658 110822 291894
rect 110266 291338 110502 291574
rect 110586 291338 110822 291574
rect 110266 255658 110502 255894
rect 110586 255658 110822 255894
rect 110266 255338 110502 255574
rect 110586 255338 110822 255574
rect 110266 219658 110502 219894
rect 110586 219658 110822 219894
rect 110266 219338 110502 219574
rect 110586 219338 110822 219574
rect 110266 183658 110502 183894
rect 110586 183658 110822 183894
rect 110266 183338 110502 183574
rect 110586 183338 110822 183574
rect 110266 147658 110502 147894
rect 110586 147658 110822 147894
rect 110266 147338 110502 147574
rect 110586 147338 110822 147574
rect 110266 111658 110502 111894
rect 110586 111658 110822 111894
rect 110266 111338 110502 111574
rect 110586 111338 110822 111574
rect 110266 75658 110502 75894
rect 110586 75658 110822 75894
rect 110266 75338 110502 75574
rect 110586 75338 110822 75574
rect 110266 39658 110502 39894
rect 110586 39658 110822 39894
rect 110266 39338 110502 39574
rect 110586 39338 110822 39574
rect 110266 3658 110502 3894
rect 110586 3658 110822 3894
rect 110266 3338 110502 3574
rect 110586 3338 110822 3574
rect 110266 -1542 110502 -1306
rect 110586 -1542 110822 -1306
rect 110266 -1862 110502 -1626
rect 110586 -1862 110822 -1626
rect 111506 706522 111742 706758
rect 111826 706522 112062 706758
rect 111506 706202 111742 706438
rect 111826 706202 112062 706438
rect 111506 688898 111742 689134
rect 111826 688898 112062 689134
rect 111506 688578 111742 688814
rect 111826 688578 112062 688814
rect 111506 652898 111742 653134
rect 111826 652898 112062 653134
rect 111506 652578 111742 652814
rect 111826 652578 112062 652814
rect 111506 616898 111742 617134
rect 111826 616898 112062 617134
rect 111506 616578 111742 616814
rect 111826 616578 112062 616814
rect 111506 580898 111742 581134
rect 111826 580898 112062 581134
rect 111506 580578 111742 580814
rect 111826 580578 112062 580814
rect 111506 544898 111742 545134
rect 111826 544898 112062 545134
rect 111506 544578 111742 544814
rect 111826 544578 112062 544814
rect 111506 508898 111742 509134
rect 111826 508898 112062 509134
rect 111506 508578 111742 508814
rect 111826 508578 112062 508814
rect 111506 472898 111742 473134
rect 111826 472898 112062 473134
rect 111506 472578 111742 472814
rect 111826 472578 112062 472814
rect 111506 436898 111742 437134
rect 111826 436898 112062 437134
rect 111506 436578 111742 436814
rect 111826 436578 112062 436814
rect 111506 400898 111742 401134
rect 111826 400898 112062 401134
rect 111506 400578 111742 400814
rect 111826 400578 112062 400814
rect 111506 364898 111742 365134
rect 111826 364898 112062 365134
rect 111506 364578 111742 364814
rect 111826 364578 112062 364814
rect 111506 328898 111742 329134
rect 111826 328898 112062 329134
rect 111506 328578 111742 328814
rect 111826 328578 112062 328814
rect 111506 292898 111742 293134
rect 111826 292898 112062 293134
rect 111506 292578 111742 292814
rect 111826 292578 112062 292814
rect 111506 256898 111742 257134
rect 111826 256898 112062 257134
rect 111506 256578 111742 256814
rect 111826 256578 112062 256814
rect 111506 220898 111742 221134
rect 111826 220898 112062 221134
rect 111506 220578 111742 220814
rect 111826 220578 112062 220814
rect 111506 184898 111742 185134
rect 111826 184898 112062 185134
rect 111506 184578 111742 184814
rect 111826 184578 112062 184814
rect 111506 148898 111742 149134
rect 111826 148898 112062 149134
rect 111506 148578 111742 148814
rect 111826 148578 112062 148814
rect 111506 112898 111742 113134
rect 111826 112898 112062 113134
rect 111506 112578 111742 112814
rect 111826 112578 112062 112814
rect 111506 76898 111742 77134
rect 111826 76898 112062 77134
rect 111506 76578 111742 76814
rect 111826 76578 112062 76814
rect 111506 40898 111742 41134
rect 111826 40898 112062 41134
rect 111506 40578 111742 40814
rect 111826 40578 112062 40814
rect 111506 4898 111742 5134
rect 111826 4898 112062 5134
rect 111506 4578 111742 4814
rect 111826 4578 112062 4814
rect 111506 -2502 111742 -2266
rect 111826 -2502 112062 -2266
rect 111506 -2822 111742 -2586
rect 111826 -2822 112062 -2586
rect 112746 707482 112982 707718
rect 113066 707482 113302 707718
rect 112746 707162 112982 707398
rect 113066 707162 113302 707398
rect 112746 690138 112982 690374
rect 113066 690138 113302 690374
rect 112746 689818 112982 690054
rect 113066 689818 113302 690054
rect 112746 654138 112982 654374
rect 113066 654138 113302 654374
rect 112746 653818 112982 654054
rect 113066 653818 113302 654054
rect 112746 618138 112982 618374
rect 113066 618138 113302 618374
rect 112746 617818 112982 618054
rect 113066 617818 113302 618054
rect 112746 582138 112982 582374
rect 113066 582138 113302 582374
rect 112746 581818 112982 582054
rect 113066 581818 113302 582054
rect 112746 546138 112982 546374
rect 113066 546138 113302 546374
rect 112746 545818 112982 546054
rect 113066 545818 113302 546054
rect 112746 510138 112982 510374
rect 113066 510138 113302 510374
rect 112746 509818 112982 510054
rect 113066 509818 113302 510054
rect 112746 474138 112982 474374
rect 113066 474138 113302 474374
rect 112746 473818 112982 474054
rect 113066 473818 113302 474054
rect 112746 438138 112982 438374
rect 113066 438138 113302 438374
rect 112746 437818 112982 438054
rect 113066 437818 113302 438054
rect 112746 402138 112982 402374
rect 113066 402138 113302 402374
rect 112746 401818 112982 402054
rect 113066 401818 113302 402054
rect 112746 366138 112982 366374
rect 113066 366138 113302 366374
rect 112746 365818 112982 366054
rect 113066 365818 113302 366054
rect 112746 330138 112982 330374
rect 113066 330138 113302 330374
rect 112746 329818 112982 330054
rect 113066 329818 113302 330054
rect 112746 294138 112982 294374
rect 113066 294138 113302 294374
rect 112746 293818 112982 294054
rect 113066 293818 113302 294054
rect 112746 258138 112982 258374
rect 113066 258138 113302 258374
rect 112746 257818 112982 258054
rect 113066 257818 113302 258054
rect 112746 222138 112982 222374
rect 113066 222138 113302 222374
rect 112746 221818 112982 222054
rect 113066 221818 113302 222054
rect 112746 186138 112982 186374
rect 113066 186138 113302 186374
rect 112746 185818 112982 186054
rect 113066 185818 113302 186054
rect 112746 150138 112982 150374
rect 113066 150138 113302 150374
rect 112746 149818 112982 150054
rect 113066 149818 113302 150054
rect 112746 114138 112982 114374
rect 113066 114138 113302 114374
rect 112746 113818 112982 114054
rect 113066 113818 113302 114054
rect 112746 78138 112982 78374
rect 113066 78138 113302 78374
rect 112746 77818 112982 78054
rect 113066 77818 113302 78054
rect 112746 42138 112982 42374
rect 113066 42138 113302 42374
rect 112746 41818 112982 42054
rect 113066 41818 113302 42054
rect 112746 6138 112982 6374
rect 113066 6138 113302 6374
rect 112746 5818 112982 6054
rect 113066 5818 113302 6054
rect 112746 -3462 112982 -3226
rect 113066 -3462 113302 -3226
rect 112746 -3782 112982 -3546
rect 113066 -3782 113302 -3546
rect 113986 708442 114222 708678
rect 114306 708442 114542 708678
rect 113986 708122 114222 708358
rect 114306 708122 114542 708358
rect 113986 691378 114222 691614
rect 114306 691378 114542 691614
rect 113986 691058 114222 691294
rect 114306 691058 114542 691294
rect 113986 655378 114222 655614
rect 114306 655378 114542 655614
rect 113986 655058 114222 655294
rect 114306 655058 114542 655294
rect 113986 619378 114222 619614
rect 114306 619378 114542 619614
rect 113986 619058 114222 619294
rect 114306 619058 114542 619294
rect 113986 583378 114222 583614
rect 114306 583378 114542 583614
rect 113986 583058 114222 583294
rect 114306 583058 114542 583294
rect 113986 547378 114222 547614
rect 114306 547378 114542 547614
rect 113986 547058 114222 547294
rect 114306 547058 114542 547294
rect 113986 511378 114222 511614
rect 114306 511378 114542 511614
rect 113986 511058 114222 511294
rect 114306 511058 114542 511294
rect 113986 475378 114222 475614
rect 114306 475378 114542 475614
rect 113986 475058 114222 475294
rect 114306 475058 114542 475294
rect 113986 439378 114222 439614
rect 114306 439378 114542 439614
rect 113986 439058 114222 439294
rect 114306 439058 114542 439294
rect 113986 403378 114222 403614
rect 114306 403378 114542 403614
rect 113986 403058 114222 403294
rect 114306 403058 114542 403294
rect 113986 367378 114222 367614
rect 114306 367378 114542 367614
rect 113986 367058 114222 367294
rect 114306 367058 114542 367294
rect 113986 331378 114222 331614
rect 114306 331378 114542 331614
rect 113986 331058 114222 331294
rect 114306 331058 114542 331294
rect 113986 295378 114222 295614
rect 114306 295378 114542 295614
rect 113986 295058 114222 295294
rect 114306 295058 114542 295294
rect 113986 259378 114222 259614
rect 114306 259378 114542 259614
rect 113986 259058 114222 259294
rect 114306 259058 114542 259294
rect 113986 223378 114222 223614
rect 114306 223378 114542 223614
rect 113986 223058 114222 223294
rect 114306 223058 114542 223294
rect 113986 187378 114222 187614
rect 114306 187378 114542 187614
rect 113986 187058 114222 187294
rect 114306 187058 114542 187294
rect 113986 151378 114222 151614
rect 114306 151378 114542 151614
rect 113986 151058 114222 151294
rect 114306 151058 114542 151294
rect 113986 115378 114222 115614
rect 114306 115378 114542 115614
rect 113986 115058 114222 115294
rect 114306 115058 114542 115294
rect 113986 79378 114222 79614
rect 114306 79378 114542 79614
rect 113986 79058 114222 79294
rect 114306 79058 114542 79294
rect 113986 43378 114222 43614
rect 114306 43378 114542 43614
rect 113986 43058 114222 43294
rect 114306 43058 114542 43294
rect 113986 7378 114222 7614
rect 114306 7378 114542 7614
rect 113986 7058 114222 7294
rect 114306 7058 114542 7294
rect 113986 -4422 114222 -4186
rect 114306 -4422 114542 -4186
rect 113986 -4742 114222 -4506
rect 114306 -4742 114542 -4506
rect 115226 709402 115462 709638
rect 115546 709402 115782 709638
rect 115226 709082 115462 709318
rect 115546 709082 115782 709318
rect 115226 692618 115462 692854
rect 115546 692618 115782 692854
rect 115226 692298 115462 692534
rect 115546 692298 115782 692534
rect 115226 656618 115462 656854
rect 115546 656618 115782 656854
rect 115226 656298 115462 656534
rect 115546 656298 115782 656534
rect 115226 620618 115462 620854
rect 115546 620618 115782 620854
rect 115226 620298 115462 620534
rect 115546 620298 115782 620534
rect 115226 584618 115462 584854
rect 115546 584618 115782 584854
rect 115226 584298 115462 584534
rect 115546 584298 115782 584534
rect 115226 548618 115462 548854
rect 115546 548618 115782 548854
rect 115226 548298 115462 548534
rect 115546 548298 115782 548534
rect 115226 512618 115462 512854
rect 115546 512618 115782 512854
rect 115226 512298 115462 512534
rect 115546 512298 115782 512534
rect 115226 476618 115462 476854
rect 115546 476618 115782 476854
rect 115226 476298 115462 476534
rect 115546 476298 115782 476534
rect 115226 440618 115462 440854
rect 115546 440618 115782 440854
rect 115226 440298 115462 440534
rect 115546 440298 115782 440534
rect 115226 404618 115462 404854
rect 115546 404618 115782 404854
rect 115226 404298 115462 404534
rect 115546 404298 115782 404534
rect 115226 368618 115462 368854
rect 115546 368618 115782 368854
rect 115226 368298 115462 368534
rect 115546 368298 115782 368534
rect 115226 332618 115462 332854
rect 115546 332618 115782 332854
rect 115226 332298 115462 332534
rect 115546 332298 115782 332534
rect 115226 296618 115462 296854
rect 115546 296618 115782 296854
rect 115226 296298 115462 296534
rect 115546 296298 115782 296534
rect 115226 260618 115462 260854
rect 115546 260618 115782 260854
rect 115226 260298 115462 260534
rect 115546 260298 115782 260534
rect 115226 224618 115462 224854
rect 115546 224618 115782 224854
rect 115226 224298 115462 224534
rect 115546 224298 115782 224534
rect 115226 188618 115462 188854
rect 115546 188618 115782 188854
rect 115226 188298 115462 188534
rect 115546 188298 115782 188534
rect 115226 152618 115462 152854
rect 115546 152618 115782 152854
rect 115226 152298 115462 152534
rect 115546 152298 115782 152534
rect 115226 116618 115462 116854
rect 115546 116618 115782 116854
rect 115226 116298 115462 116534
rect 115546 116298 115782 116534
rect 115226 80618 115462 80854
rect 115546 80618 115782 80854
rect 115226 80298 115462 80534
rect 115546 80298 115782 80534
rect 115226 44618 115462 44854
rect 115546 44618 115782 44854
rect 115226 44298 115462 44534
rect 115546 44298 115782 44534
rect 115226 8618 115462 8854
rect 115546 8618 115782 8854
rect 115226 8298 115462 8534
rect 115546 8298 115782 8534
rect 115226 -5382 115462 -5146
rect 115546 -5382 115782 -5146
rect 115226 -5702 115462 -5466
rect 115546 -5702 115782 -5466
rect 116466 710362 116702 710598
rect 116786 710362 117022 710598
rect 116466 710042 116702 710278
rect 116786 710042 117022 710278
rect 116466 693858 116702 694094
rect 116786 693858 117022 694094
rect 116466 693538 116702 693774
rect 116786 693538 117022 693774
rect 116466 657858 116702 658094
rect 116786 657858 117022 658094
rect 116466 657538 116702 657774
rect 116786 657538 117022 657774
rect 116466 621858 116702 622094
rect 116786 621858 117022 622094
rect 116466 621538 116702 621774
rect 116786 621538 117022 621774
rect 116466 585858 116702 586094
rect 116786 585858 117022 586094
rect 116466 585538 116702 585774
rect 116786 585538 117022 585774
rect 116466 549858 116702 550094
rect 116786 549858 117022 550094
rect 116466 549538 116702 549774
rect 116786 549538 117022 549774
rect 116466 513858 116702 514094
rect 116786 513858 117022 514094
rect 116466 513538 116702 513774
rect 116786 513538 117022 513774
rect 116466 477858 116702 478094
rect 116786 477858 117022 478094
rect 116466 477538 116702 477774
rect 116786 477538 117022 477774
rect 116466 441858 116702 442094
rect 116786 441858 117022 442094
rect 116466 441538 116702 441774
rect 116786 441538 117022 441774
rect 116466 405858 116702 406094
rect 116786 405858 117022 406094
rect 116466 405538 116702 405774
rect 116786 405538 117022 405774
rect 116466 369858 116702 370094
rect 116786 369858 117022 370094
rect 116466 369538 116702 369774
rect 116786 369538 117022 369774
rect 116466 333858 116702 334094
rect 116786 333858 117022 334094
rect 116466 333538 116702 333774
rect 116786 333538 117022 333774
rect 116466 297858 116702 298094
rect 116786 297858 117022 298094
rect 116466 297538 116702 297774
rect 116786 297538 117022 297774
rect 116466 261858 116702 262094
rect 116786 261858 117022 262094
rect 116466 261538 116702 261774
rect 116786 261538 117022 261774
rect 116466 225858 116702 226094
rect 116786 225858 117022 226094
rect 116466 225538 116702 225774
rect 116786 225538 117022 225774
rect 116466 189858 116702 190094
rect 116786 189858 117022 190094
rect 116466 189538 116702 189774
rect 116786 189538 117022 189774
rect 116466 153858 116702 154094
rect 116786 153858 117022 154094
rect 116466 153538 116702 153774
rect 116786 153538 117022 153774
rect 116466 117858 116702 118094
rect 116786 117858 117022 118094
rect 116466 117538 116702 117774
rect 116786 117538 117022 117774
rect 116466 81858 116702 82094
rect 116786 81858 117022 82094
rect 116466 81538 116702 81774
rect 116786 81538 117022 81774
rect 116466 45858 116702 46094
rect 116786 45858 117022 46094
rect 116466 45538 116702 45774
rect 116786 45538 117022 45774
rect 116466 9858 116702 10094
rect 116786 9858 117022 10094
rect 116466 9538 116702 9774
rect 116786 9538 117022 9774
rect 116466 -6342 116702 -6106
rect 116786 -6342 117022 -6106
rect 116466 -6662 116702 -6426
rect 116786 -6662 117022 -6426
rect 117706 711322 117942 711558
rect 118026 711322 118262 711558
rect 117706 711002 117942 711238
rect 118026 711002 118262 711238
rect 117706 695098 117942 695334
rect 118026 695098 118262 695334
rect 117706 694778 117942 695014
rect 118026 694778 118262 695014
rect 117706 659098 117942 659334
rect 118026 659098 118262 659334
rect 117706 658778 117942 659014
rect 118026 658778 118262 659014
rect 117706 623098 117942 623334
rect 118026 623098 118262 623334
rect 117706 622778 117942 623014
rect 118026 622778 118262 623014
rect 117706 587098 117942 587334
rect 118026 587098 118262 587334
rect 117706 586778 117942 587014
rect 118026 586778 118262 587014
rect 117706 551098 117942 551334
rect 118026 551098 118262 551334
rect 117706 550778 117942 551014
rect 118026 550778 118262 551014
rect 117706 515098 117942 515334
rect 118026 515098 118262 515334
rect 117706 514778 117942 515014
rect 118026 514778 118262 515014
rect 117706 479098 117942 479334
rect 118026 479098 118262 479334
rect 117706 478778 117942 479014
rect 118026 478778 118262 479014
rect 117706 443098 117942 443334
rect 118026 443098 118262 443334
rect 117706 442778 117942 443014
rect 118026 442778 118262 443014
rect 117706 407098 117942 407334
rect 118026 407098 118262 407334
rect 117706 406778 117942 407014
rect 118026 406778 118262 407014
rect 117706 371098 117942 371334
rect 118026 371098 118262 371334
rect 117706 370778 117942 371014
rect 118026 370778 118262 371014
rect 117706 335098 117942 335334
rect 118026 335098 118262 335334
rect 117706 334778 117942 335014
rect 118026 334778 118262 335014
rect 117706 299098 117942 299334
rect 118026 299098 118262 299334
rect 117706 298778 117942 299014
rect 118026 298778 118262 299014
rect 117706 263098 117942 263334
rect 118026 263098 118262 263334
rect 117706 262778 117942 263014
rect 118026 262778 118262 263014
rect 117706 227098 117942 227334
rect 118026 227098 118262 227334
rect 117706 226778 117942 227014
rect 118026 226778 118262 227014
rect 117706 191098 117942 191334
rect 118026 191098 118262 191334
rect 117706 190778 117942 191014
rect 118026 190778 118262 191014
rect 117706 155098 117942 155334
rect 118026 155098 118262 155334
rect 117706 154778 117942 155014
rect 118026 154778 118262 155014
rect 117706 119098 117942 119334
rect 118026 119098 118262 119334
rect 117706 118778 117942 119014
rect 118026 118778 118262 119014
rect 117706 83098 117942 83334
rect 118026 83098 118262 83334
rect 117706 82778 117942 83014
rect 118026 82778 118262 83014
rect 117706 47098 117942 47334
rect 118026 47098 118262 47334
rect 117706 46778 117942 47014
rect 118026 46778 118262 47014
rect 117706 11098 117942 11334
rect 118026 11098 118262 11334
rect 117706 10778 117942 11014
rect 118026 10778 118262 11014
rect 117706 -7302 117942 -7066
rect 118026 -7302 118262 -7066
rect 117706 -7622 117942 -7386
rect 118026 -7622 118262 -7386
rect 145026 704602 145262 704838
rect 145346 704602 145582 704838
rect 145026 704282 145262 704518
rect 145346 704282 145582 704518
rect 145026 686418 145262 686654
rect 145346 686418 145582 686654
rect 145026 686098 145262 686334
rect 145346 686098 145582 686334
rect 145026 650418 145262 650654
rect 145346 650418 145582 650654
rect 145026 650098 145262 650334
rect 145346 650098 145582 650334
rect 145026 614418 145262 614654
rect 145346 614418 145582 614654
rect 145026 614098 145262 614334
rect 145346 614098 145582 614334
rect 145026 578418 145262 578654
rect 145346 578418 145582 578654
rect 145026 578098 145262 578334
rect 145346 578098 145582 578334
rect 145026 542418 145262 542654
rect 145346 542418 145582 542654
rect 145026 542098 145262 542334
rect 145346 542098 145582 542334
rect 145026 506418 145262 506654
rect 145346 506418 145582 506654
rect 145026 506098 145262 506334
rect 145346 506098 145582 506334
rect 145026 470418 145262 470654
rect 145346 470418 145582 470654
rect 145026 470098 145262 470334
rect 145346 470098 145582 470334
rect 145026 434418 145262 434654
rect 145346 434418 145582 434654
rect 145026 434098 145262 434334
rect 145346 434098 145582 434334
rect 145026 398418 145262 398654
rect 145346 398418 145582 398654
rect 145026 398098 145262 398334
rect 145346 398098 145582 398334
rect 145026 362418 145262 362654
rect 145346 362418 145582 362654
rect 145026 362098 145262 362334
rect 145346 362098 145582 362334
rect 145026 326418 145262 326654
rect 145346 326418 145582 326654
rect 145026 326098 145262 326334
rect 145346 326098 145582 326334
rect 145026 290418 145262 290654
rect 145346 290418 145582 290654
rect 145026 290098 145262 290334
rect 145346 290098 145582 290334
rect 145026 254418 145262 254654
rect 145346 254418 145582 254654
rect 145026 254098 145262 254334
rect 145346 254098 145582 254334
rect 145026 218418 145262 218654
rect 145346 218418 145582 218654
rect 145026 218098 145262 218334
rect 145346 218098 145582 218334
rect 145026 182418 145262 182654
rect 145346 182418 145582 182654
rect 145026 182098 145262 182334
rect 145346 182098 145582 182334
rect 145026 146418 145262 146654
rect 145346 146418 145582 146654
rect 145026 146098 145262 146334
rect 145346 146098 145582 146334
rect 145026 110418 145262 110654
rect 145346 110418 145582 110654
rect 145026 110098 145262 110334
rect 145346 110098 145582 110334
rect 145026 74418 145262 74654
rect 145346 74418 145582 74654
rect 145026 74098 145262 74334
rect 145346 74098 145582 74334
rect 145026 38418 145262 38654
rect 145346 38418 145582 38654
rect 145026 38098 145262 38334
rect 145346 38098 145582 38334
rect 145026 2418 145262 2654
rect 145346 2418 145582 2654
rect 145026 2098 145262 2334
rect 145346 2098 145582 2334
rect 145026 -582 145262 -346
rect 145346 -582 145582 -346
rect 145026 -902 145262 -666
rect 145346 -902 145582 -666
rect 146266 705562 146502 705798
rect 146586 705562 146822 705798
rect 146266 705242 146502 705478
rect 146586 705242 146822 705478
rect 146266 687658 146502 687894
rect 146586 687658 146822 687894
rect 146266 687338 146502 687574
rect 146586 687338 146822 687574
rect 146266 651658 146502 651894
rect 146586 651658 146822 651894
rect 146266 651338 146502 651574
rect 146586 651338 146822 651574
rect 146266 615658 146502 615894
rect 146586 615658 146822 615894
rect 146266 615338 146502 615574
rect 146586 615338 146822 615574
rect 146266 579658 146502 579894
rect 146586 579658 146822 579894
rect 146266 579338 146502 579574
rect 146586 579338 146822 579574
rect 146266 543658 146502 543894
rect 146586 543658 146822 543894
rect 146266 543338 146502 543574
rect 146586 543338 146822 543574
rect 146266 507658 146502 507894
rect 146586 507658 146822 507894
rect 146266 507338 146502 507574
rect 146586 507338 146822 507574
rect 146266 471658 146502 471894
rect 146586 471658 146822 471894
rect 146266 471338 146502 471574
rect 146586 471338 146822 471574
rect 146266 435658 146502 435894
rect 146586 435658 146822 435894
rect 146266 435338 146502 435574
rect 146586 435338 146822 435574
rect 146266 399658 146502 399894
rect 146586 399658 146822 399894
rect 146266 399338 146502 399574
rect 146586 399338 146822 399574
rect 146266 363658 146502 363894
rect 146586 363658 146822 363894
rect 146266 363338 146502 363574
rect 146586 363338 146822 363574
rect 146266 327658 146502 327894
rect 146586 327658 146822 327894
rect 146266 327338 146502 327574
rect 146586 327338 146822 327574
rect 146266 291658 146502 291894
rect 146586 291658 146822 291894
rect 146266 291338 146502 291574
rect 146586 291338 146822 291574
rect 146266 255658 146502 255894
rect 146586 255658 146822 255894
rect 146266 255338 146502 255574
rect 146586 255338 146822 255574
rect 146266 219658 146502 219894
rect 146586 219658 146822 219894
rect 146266 219338 146502 219574
rect 146586 219338 146822 219574
rect 146266 183658 146502 183894
rect 146586 183658 146822 183894
rect 146266 183338 146502 183574
rect 146586 183338 146822 183574
rect 146266 147658 146502 147894
rect 146586 147658 146822 147894
rect 146266 147338 146502 147574
rect 146586 147338 146822 147574
rect 146266 111658 146502 111894
rect 146586 111658 146822 111894
rect 146266 111338 146502 111574
rect 146586 111338 146822 111574
rect 146266 75658 146502 75894
rect 146586 75658 146822 75894
rect 146266 75338 146502 75574
rect 146586 75338 146822 75574
rect 146266 39658 146502 39894
rect 146586 39658 146822 39894
rect 146266 39338 146502 39574
rect 146586 39338 146822 39574
rect 146266 3658 146502 3894
rect 146586 3658 146822 3894
rect 146266 3338 146502 3574
rect 146586 3338 146822 3574
rect 146266 -1542 146502 -1306
rect 146586 -1542 146822 -1306
rect 146266 -1862 146502 -1626
rect 146586 -1862 146822 -1626
rect 147506 706522 147742 706758
rect 147826 706522 148062 706758
rect 147506 706202 147742 706438
rect 147826 706202 148062 706438
rect 147506 688898 147742 689134
rect 147826 688898 148062 689134
rect 147506 688578 147742 688814
rect 147826 688578 148062 688814
rect 147506 652898 147742 653134
rect 147826 652898 148062 653134
rect 147506 652578 147742 652814
rect 147826 652578 148062 652814
rect 147506 616898 147742 617134
rect 147826 616898 148062 617134
rect 147506 616578 147742 616814
rect 147826 616578 148062 616814
rect 147506 580898 147742 581134
rect 147826 580898 148062 581134
rect 147506 580578 147742 580814
rect 147826 580578 148062 580814
rect 147506 544898 147742 545134
rect 147826 544898 148062 545134
rect 147506 544578 147742 544814
rect 147826 544578 148062 544814
rect 147506 508898 147742 509134
rect 147826 508898 148062 509134
rect 147506 508578 147742 508814
rect 147826 508578 148062 508814
rect 147506 472898 147742 473134
rect 147826 472898 148062 473134
rect 147506 472578 147742 472814
rect 147826 472578 148062 472814
rect 147506 436898 147742 437134
rect 147826 436898 148062 437134
rect 147506 436578 147742 436814
rect 147826 436578 148062 436814
rect 147506 400898 147742 401134
rect 147826 400898 148062 401134
rect 147506 400578 147742 400814
rect 147826 400578 148062 400814
rect 147506 364898 147742 365134
rect 147826 364898 148062 365134
rect 147506 364578 147742 364814
rect 147826 364578 148062 364814
rect 147506 328898 147742 329134
rect 147826 328898 148062 329134
rect 147506 328578 147742 328814
rect 147826 328578 148062 328814
rect 147506 292898 147742 293134
rect 147826 292898 148062 293134
rect 147506 292578 147742 292814
rect 147826 292578 148062 292814
rect 147506 256898 147742 257134
rect 147826 256898 148062 257134
rect 147506 256578 147742 256814
rect 147826 256578 148062 256814
rect 147506 220898 147742 221134
rect 147826 220898 148062 221134
rect 147506 220578 147742 220814
rect 147826 220578 148062 220814
rect 147506 184898 147742 185134
rect 147826 184898 148062 185134
rect 147506 184578 147742 184814
rect 147826 184578 148062 184814
rect 147506 148898 147742 149134
rect 147826 148898 148062 149134
rect 147506 148578 147742 148814
rect 147826 148578 148062 148814
rect 147506 112898 147742 113134
rect 147826 112898 148062 113134
rect 147506 112578 147742 112814
rect 147826 112578 148062 112814
rect 147506 76898 147742 77134
rect 147826 76898 148062 77134
rect 147506 76578 147742 76814
rect 147826 76578 148062 76814
rect 147506 40898 147742 41134
rect 147826 40898 148062 41134
rect 147506 40578 147742 40814
rect 147826 40578 148062 40814
rect 147506 4898 147742 5134
rect 147826 4898 148062 5134
rect 147506 4578 147742 4814
rect 147826 4578 148062 4814
rect 147506 -2502 147742 -2266
rect 147826 -2502 148062 -2266
rect 147506 -2822 147742 -2586
rect 147826 -2822 148062 -2586
rect 148746 707482 148982 707718
rect 149066 707482 149302 707718
rect 148746 707162 148982 707398
rect 149066 707162 149302 707398
rect 148746 690138 148982 690374
rect 149066 690138 149302 690374
rect 148746 689818 148982 690054
rect 149066 689818 149302 690054
rect 148746 654138 148982 654374
rect 149066 654138 149302 654374
rect 148746 653818 148982 654054
rect 149066 653818 149302 654054
rect 148746 618138 148982 618374
rect 149066 618138 149302 618374
rect 148746 617818 148982 618054
rect 149066 617818 149302 618054
rect 148746 582138 148982 582374
rect 149066 582138 149302 582374
rect 148746 581818 148982 582054
rect 149066 581818 149302 582054
rect 148746 546138 148982 546374
rect 149066 546138 149302 546374
rect 148746 545818 148982 546054
rect 149066 545818 149302 546054
rect 148746 510138 148982 510374
rect 149066 510138 149302 510374
rect 148746 509818 148982 510054
rect 149066 509818 149302 510054
rect 148746 474138 148982 474374
rect 149066 474138 149302 474374
rect 148746 473818 148982 474054
rect 149066 473818 149302 474054
rect 148746 438138 148982 438374
rect 149066 438138 149302 438374
rect 148746 437818 148982 438054
rect 149066 437818 149302 438054
rect 148746 402138 148982 402374
rect 149066 402138 149302 402374
rect 148746 401818 148982 402054
rect 149066 401818 149302 402054
rect 148746 366138 148982 366374
rect 149066 366138 149302 366374
rect 148746 365818 148982 366054
rect 149066 365818 149302 366054
rect 148746 330138 148982 330374
rect 149066 330138 149302 330374
rect 148746 329818 148982 330054
rect 149066 329818 149302 330054
rect 148746 294138 148982 294374
rect 149066 294138 149302 294374
rect 148746 293818 148982 294054
rect 149066 293818 149302 294054
rect 148746 258138 148982 258374
rect 149066 258138 149302 258374
rect 148746 257818 148982 258054
rect 149066 257818 149302 258054
rect 148746 222138 148982 222374
rect 149066 222138 149302 222374
rect 148746 221818 148982 222054
rect 149066 221818 149302 222054
rect 148746 186138 148982 186374
rect 149066 186138 149302 186374
rect 148746 185818 148982 186054
rect 149066 185818 149302 186054
rect 148746 150138 148982 150374
rect 149066 150138 149302 150374
rect 148746 149818 148982 150054
rect 149066 149818 149302 150054
rect 148746 114138 148982 114374
rect 149066 114138 149302 114374
rect 148746 113818 148982 114054
rect 149066 113818 149302 114054
rect 148746 78138 148982 78374
rect 149066 78138 149302 78374
rect 148746 77818 148982 78054
rect 149066 77818 149302 78054
rect 148746 42138 148982 42374
rect 149066 42138 149302 42374
rect 148746 41818 148982 42054
rect 149066 41818 149302 42054
rect 148746 6138 148982 6374
rect 149066 6138 149302 6374
rect 148746 5818 148982 6054
rect 149066 5818 149302 6054
rect 148746 -3462 148982 -3226
rect 149066 -3462 149302 -3226
rect 148746 -3782 148982 -3546
rect 149066 -3782 149302 -3546
rect 149986 708442 150222 708678
rect 150306 708442 150542 708678
rect 149986 708122 150222 708358
rect 150306 708122 150542 708358
rect 149986 691378 150222 691614
rect 150306 691378 150542 691614
rect 149986 691058 150222 691294
rect 150306 691058 150542 691294
rect 149986 655378 150222 655614
rect 150306 655378 150542 655614
rect 149986 655058 150222 655294
rect 150306 655058 150542 655294
rect 149986 619378 150222 619614
rect 150306 619378 150542 619614
rect 149986 619058 150222 619294
rect 150306 619058 150542 619294
rect 149986 583378 150222 583614
rect 150306 583378 150542 583614
rect 149986 583058 150222 583294
rect 150306 583058 150542 583294
rect 149986 547378 150222 547614
rect 150306 547378 150542 547614
rect 149986 547058 150222 547294
rect 150306 547058 150542 547294
rect 149986 511378 150222 511614
rect 150306 511378 150542 511614
rect 149986 511058 150222 511294
rect 150306 511058 150542 511294
rect 149986 475378 150222 475614
rect 150306 475378 150542 475614
rect 149986 475058 150222 475294
rect 150306 475058 150542 475294
rect 149986 439378 150222 439614
rect 150306 439378 150542 439614
rect 149986 439058 150222 439294
rect 150306 439058 150542 439294
rect 149986 403378 150222 403614
rect 150306 403378 150542 403614
rect 149986 403058 150222 403294
rect 150306 403058 150542 403294
rect 149986 367378 150222 367614
rect 150306 367378 150542 367614
rect 149986 367058 150222 367294
rect 150306 367058 150542 367294
rect 149986 331378 150222 331614
rect 150306 331378 150542 331614
rect 149986 331058 150222 331294
rect 150306 331058 150542 331294
rect 149986 295378 150222 295614
rect 150306 295378 150542 295614
rect 149986 295058 150222 295294
rect 150306 295058 150542 295294
rect 149986 259378 150222 259614
rect 150306 259378 150542 259614
rect 149986 259058 150222 259294
rect 150306 259058 150542 259294
rect 149986 223378 150222 223614
rect 150306 223378 150542 223614
rect 149986 223058 150222 223294
rect 150306 223058 150542 223294
rect 149986 187378 150222 187614
rect 150306 187378 150542 187614
rect 149986 187058 150222 187294
rect 150306 187058 150542 187294
rect 149986 151378 150222 151614
rect 150306 151378 150542 151614
rect 149986 151058 150222 151294
rect 150306 151058 150542 151294
rect 149986 115378 150222 115614
rect 150306 115378 150542 115614
rect 149986 115058 150222 115294
rect 150306 115058 150542 115294
rect 149986 79378 150222 79614
rect 150306 79378 150542 79614
rect 149986 79058 150222 79294
rect 150306 79058 150542 79294
rect 149986 43378 150222 43614
rect 150306 43378 150542 43614
rect 149986 43058 150222 43294
rect 150306 43058 150542 43294
rect 149986 7378 150222 7614
rect 150306 7378 150542 7614
rect 149986 7058 150222 7294
rect 150306 7058 150542 7294
rect 149986 -4422 150222 -4186
rect 150306 -4422 150542 -4186
rect 149986 -4742 150222 -4506
rect 150306 -4742 150542 -4506
rect 151226 709402 151462 709638
rect 151546 709402 151782 709638
rect 151226 709082 151462 709318
rect 151546 709082 151782 709318
rect 151226 692618 151462 692854
rect 151546 692618 151782 692854
rect 151226 692298 151462 692534
rect 151546 692298 151782 692534
rect 151226 656618 151462 656854
rect 151546 656618 151782 656854
rect 151226 656298 151462 656534
rect 151546 656298 151782 656534
rect 151226 620618 151462 620854
rect 151546 620618 151782 620854
rect 151226 620298 151462 620534
rect 151546 620298 151782 620534
rect 151226 584618 151462 584854
rect 151546 584618 151782 584854
rect 151226 584298 151462 584534
rect 151546 584298 151782 584534
rect 151226 548618 151462 548854
rect 151546 548618 151782 548854
rect 151226 548298 151462 548534
rect 151546 548298 151782 548534
rect 151226 512618 151462 512854
rect 151546 512618 151782 512854
rect 151226 512298 151462 512534
rect 151546 512298 151782 512534
rect 151226 476618 151462 476854
rect 151546 476618 151782 476854
rect 151226 476298 151462 476534
rect 151546 476298 151782 476534
rect 151226 440618 151462 440854
rect 151546 440618 151782 440854
rect 151226 440298 151462 440534
rect 151546 440298 151782 440534
rect 151226 404618 151462 404854
rect 151546 404618 151782 404854
rect 151226 404298 151462 404534
rect 151546 404298 151782 404534
rect 151226 368618 151462 368854
rect 151546 368618 151782 368854
rect 151226 368298 151462 368534
rect 151546 368298 151782 368534
rect 151226 332618 151462 332854
rect 151546 332618 151782 332854
rect 151226 332298 151462 332534
rect 151546 332298 151782 332534
rect 151226 296618 151462 296854
rect 151546 296618 151782 296854
rect 151226 296298 151462 296534
rect 151546 296298 151782 296534
rect 151226 260618 151462 260854
rect 151546 260618 151782 260854
rect 151226 260298 151462 260534
rect 151546 260298 151782 260534
rect 151226 224618 151462 224854
rect 151546 224618 151782 224854
rect 151226 224298 151462 224534
rect 151546 224298 151782 224534
rect 151226 188618 151462 188854
rect 151546 188618 151782 188854
rect 151226 188298 151462 188534
rect 151546 188298 151782 188534
rect 151226 152618 151462 152854
rect 151546 152618 151782 152854
rect 151226 152298 151462 152534
rect 151546 152298 151782 152534
rect 151226 116618 151462 116854
rect 151546 116618 151782 116854
rect 151226 116298 151462 116534
rect 151546 116298 151782 116534
rect 151226 80618 151462 80854
rect 151546 80618 151782 80854
rect 151226 80298 151462 80534
rect 151546 80298 151782 80534
rect 151226 44618 151462 44854
rect 151546 44618 151782 44854
rect 151226 44298 151462 44534
rect 151546 44298 151782 44534
rect 151226 8618 151462 8854
rect 151546 8618 151782 8854
rect 151226 8298 151462 8534
rect 151546 8298 151782 8534
rect 151226 -5382 151462 -5146
rect 151546 -5382 151782 -5146
rect 151226 -5702 151462 -5466
rect 151546 -5702 151782 -5466
rect 152466 710362 152702 710598
rect 152786 710362 153022 710598
rect 152466 710042 152702 710278
rect 152786 710042 153022 710278
rect 152466 693858 152702 694094
rect 152786 693858 153022 694094
rect 152466 693538 152702 693774
rect 152786 693538 153022 693774
rect 152466 657858 152702 658094
rect 152786 657858 153022 658094
rect 152466 657538 152702 657774
rect 152786 657538 153022 657774
rect 152466 621858 152702 622094
rect 152786 621858 153022 622094
rect 152466 621538 152702 621774
rect 152786 621538 153022 621774
rect 152466 585858 152702 586094
rect 152786 585858 153022 586094
rect 152466 585538 152702 585774
rect 152786 585538 153022 585774
rect 152466 549858 152702 550094
rect 152786 549858 153022 550094
rect 152466 549538 152702 549774
rect 152786 549538 153022 549774
rect 152466 513858 152702 514094
rect 152786 513858 153022 514094
rect 152466 513538 152702 513774
rect 152786 513538 153022 513774
rect 152466 477858 152702 478094
rect 152786 477858 153022 478094
rect 152466 477538 152702 477774
rect 152786 477538 153022 477774
rect 152466 441858 152702 442094
rect 152786 441858 153022 442094
rect 152466 441538 152702 441774
rect 152786 441538 153022 441774
rect 152466 405858 152702 406094
rect 152786 405858 153022 406094
rect 152466 405538 152702 405774
rect 152786 405538 153022 405774
rect 152466 369858 152702 370094
rect 152786 369858 153022 370094
rect 152466 369538 152702 369774
rect 152786 369538 153022 369774
rect 152466 333858 152702 334094
rect 152786 333858 153022 334094
rect 152466 333538 152702 333774
rect 152786 333538 153022 333774
rect 152466 297858 152702 298094
rect 152786 297858 153022 298094
rect 152466 297538 152702 297774
rect 152786 297538 153022 297774
rect 152466 261858 152702 262094
rect 152786 261858 153022 262094
rect 152466 261538 152702 261774
rect 152786 261538 153022 261774
rect 152466 225858 152702 226094
rect 152786 225858 153022 226094
rect 152466 225538 152702 225774
rect 152786 225538 153022 225774
rect 152466 189858 152702 190094
rect 152786 189858 153022 190094
rect 152466 189538 152702 189774
rect 152786 189538 153022 189774
rect 152466 153858 152702 154094
rect 152786 153858 153022 154094
rect 152466 153538 152702 153774
rect 152786 153538 153022 153774
rect 152466 117858 152702 118094
rect 152786 117858 153022 118094
rect 152466 117538 152702 117774
rect 152786 117538 153022 117774
rect 152466 81858 152702 82094
rect 152786 81858 153022 82094
rect 152466 81538 152702 81774
rect 152786 81538 153022 81774
rect 152466 45858 152702 46094
rect 152786 45858 153022 46094
rect 152466 45538 152702 45774
rect 152786 45538 153022 45774
rect 152466 9858 152702 10094
rect 152786 9858 153022 10094
rect 152466 9538 152702 9774
rect 152786 9538 153022 9774
rect 152466 -6342 152702 -6106
rect 152786 -6342 153022 -6106
rect 152466 -6662 152702 -6426
rect 152786 -6662 153022 -6426
rect 153706 711322 153942 711558
rect 154026 711322 154262 711558
rect 153706 711002 153942 711238
rect 154026 711002 154262 711238
rect 153706 695098 153942 695334
rect 154026 695098 154262 695334
rect 153706 694778 153942 695014
rect 154026 694778 154262 695014
rect 153706 659098 153942 659334
rect 154026 659098 154262 659334
rect 153706 658778 153942 659014
rect 154026 658778 154262 659014
rect 153706 623098 153942 623334
rect 154026 623098 154262 623334
rect 153706 622778 153942 623014
rect 154026 622778 154262 623014
rect 153706 587098 153942 587334
rect 154026 587098 154262 587334
rect 153706 586778 153942 587014
rect 154026 586778 154262 587014
rect 153706 551098 153942 551334
rect 154026 551098 154262 551334
rect 153706 550778 153942 551014
rect 154026 550778 154262 551014
rect 153706 515098 153942 515334
rect 154026 515098 154262 515334
rect 153706 514778 153942 515014
rect 154026 514778 154262 515014
rect 153706 479098 153942 479334
rect 154026 479098 154262 479334
rect 153706 478778 153942 479014
rect 154026 478778 154262 479014
rect 153706 443098 153942 443334
rect 154026 443098 154262 443334
rect 153706 442778 153942 443014
rect 154026 442778 154262 443014
rect 153706 407098 153942 407334
rect 154026 407098 154262 407334
rect 153706 406778 153942 407014
rect 154026 406778 154262 407014
rect 153706 371098 153942 371334
rect 154026 371098 154262 371334
rect 153706 370778 153942 371014
rect 154026 370778 154262 371014
rect 153706 335098 153942 335334
rect 154026 335098 154262 335334
rect 153706 334778 153942 335014
rect 154026 334778 154262 335014
rect 153706 299098 153942 299334
rect 154026 299098 154262 299334
rect 153706 298778 153942 299014
rect 154026 298778 154262 299014
rect 153706 263098 153942 263334
rect 154026 263098 154262 263334
rect 153706 262778 153942 263014
rect 154026 262778 154262 263014
rect 153706 227098 153942 227334
rect 154026 227098 154262 227334
rect 153706 226778 153942 227014
rect 154026 226778 154262 227014
rect 153706 191098 153942 191334
rect 154026 191098 154262 191334
rect 153706 190778 153942 191014
rect 154026 190778 154262 191014
rect 153706 155098 153942 155334
rect 154026 155098 154262 155334
rect 153706 154778 153942 155014
rect 154026 154778 154262 155014
rect 153706 119098 153942 119334
rect 154026 119098 154262 119334
rect 153706 118778 153942 119014
rect 154026 118778 154262 119014
rect 153706 83098 153942 83334
rect 154026 83098 154262 83334
rect 153706 82778 153942 83014
rect 154026 82778 154262 83014
rect 153706 47098 153942 47334
rect 154026 47098 154262 47334
rect 153706 46778 153942 47014
rect 154026 46778 154262 47014
rect 153706 11098 153942 11334
rect 154026 11098 154262 11334
rect 153706 10778 153942 11014
rect 154026 10778 154262 11014
rect 153706 -7302 153942 -7066
rect 154026 -7302 154262 -7066
rect 153706 -7622 153942 -7386
rect 154026 -7622 154262 -7386
rect 181026 704602 181262 704838
rect 181346 704602 181582 704838
rect 181026 704282 181262 704518
rect 181346 704282 181582 704518
rect 181026 686418 181262 686654
rect 181346 686418 181582 686654
rect 181026 686098 181262 686334
rect 181346 686098 181582 686334
rect 181026 650418 181262 650654
rect 181346 650418 181582 650654
rect 181026 650098 181262 650334
rect 181346 650098 181582 650334
rect 181026 614418 181262 614654
rect 181346 614418 181582 614654
rect 181026 614098 181262 614334
rect 181346 614098 181582 614334
rect 181026 578418 181262 578654
rect 181346 578418 181582 578654
rect 181026 578098 181262 578334
rect 181346 578098 181582 578334
rect 181026 542418 181262 542654
rect 181346 542418 181582 542654
rect 181026 542098 181262 542334
rect 181346 542098 181582 542334
rect 181026 506418 181262 506654
rect 181346 506418 181582 506654
rect 181026 506098 181262 506334
rect 181346 506098 181582 506334
rect 181026 470418 181262 470654
rect 181346 470418 181582 470654
rect 181026 470098 181262 470334
rect 181346 470098 181582 470334
rect 181026 434418 181262 434654
rect 181346 434418 181582 434654
rect 181026 434098 181262 434334
rect 181346 434098 181582 434334
rect 181026 398418 181262 398654
rect 181346 398418 181582 398654
rect 181026 398098 181262 398334
rect 181346 398098 181582 398334
rect 181026 362418 181262 362654
rect 181346 362418 181582 362654
rect 181026 362098 181262 362334
rect 181346 362098 181582 362334
rect 181026 326418 181262 326654
rect 181346 326418 181582 326654
rect 181026 326098 181262 326334
rect 181346 326098 181582 326334
rect 181026 290418 181262 290654
rect 181346 290418 181582 290654
rect 181026 290098 181262 290334
rect 181346 290098 181582 290334
rect 181026 254418 181262 254654
rect 181346 254418 181582 254654
rect 181026 254098 181262 254334
rect 181346 254098 181582 254334
rect 181026 218418 181262 218654
rect 181346 218418 181582 218654
rect 181026 218098 181262 218334
rect 181346 218098 181582 218334
rect 181026 182418 181262 182654
rect 181346 182418 181582 182654
rect 181026 182098 181262 182334
rect 181346 182098 181582 182334
rect 181026 146418 181262 146654
rect 181346 146418 181582 146654
rect 181026 146098 181262 146334
rect 181346 146098 181582 146334
rect 181026 110418 181262 110654
rect 181346 110418 181582 110654
rect 181026 110098 181262 110334
rect 181346 110098 181582 110334
rect 181026 74418 181262 74654
rect 181346 74418 181582 74654
rect 181026 74098 181262 74334
rect 181346 74098 181582 74334
rect 181026 38418 181262 38654
rect 181346 38418 181582 38654
rect 181026 38098 181262 38334
rect 181346 38098 181582 38334
rect 181026 2418 181262 2654
rect 181346 2418 181582 2654
rect 181026 2098 181262 2334
rect 181346 2098 181582 2334
rect 181026 -582 181262 -346
rect 181346 -582 181582 -346
rect 181026 -902 181262 -666
rect 181346 -902 181582 -666
rect 182266 705562 182502 705798
rect 182586 705562 182822 705798
rect 182266 705242 182502 705478
rect 182586 705242 182822 705478
rect 182266 687658 182502 687894
rect 182586 687658 182822 687894
rect 182266 687338 182502 687574
rect 182586 687338 182822 687574
rect 182266 651658 182502 651894
rect 182586 651658 182822 651894
rect 182266 651338 182502 651574
rect 182586 651338 182822 651574
rect 182266 615658 182502 615894
rect 182586 615658 182822 615894
rect 182266 615338 182502 615574
rect 182586 615338 182822 615574
rect 182266 579658 182502 579894
rect 182586 579658 182822 579894
rect 182266 579338 182502 579574
rect 182586 579338 182822 579574
rect 182266 543658 182502 543894
rect 182586 543658 182822 543894
rect 182266 543338 182502 543574
rect 182586 543338 182822 543574
rect 182266 507658 182502 507894
rect 182586 507658 182822 507894
rect 182266 507338 182502 507574
rect 182586 507338 182822 507574
rect 182266 471658 182502 471894
rect 182586 471658 182822 471894
rect 182266 471338 182502 471574
rect 182586 471338 182822 471574
rect 182266 435658 182502 435894
rect 182586 435658 182822 435894
rect 182266 435338 182502 435574
rect 182586 435338 182822 435574
rect 182266 399658 182502 399894
rect 182586 399658 182822 399894
rect 182266 399338 182502 399574
rect 182586 399338 182822 399574
rect 182266 363658 182502 363894
rect 182586 363658 182822 363894
rect 182266 363338 182502 363574
rect 182586 363338 182822 363574
rect 182266 327658 182502 327894
rect 182586 327658 182822 327894
rect 182266 327338 182502 327574
rect 182586 327338 182822 327574
rect 182266 291658 182502 291894
rect 182586 291658 182822 291894
rect 182266 291338 182502 291574
rect 182586 291338 182822 291574
rect 182266 255658 182502 255894
rect 182586 255658 182822 255894
rect 182266 255338 182502 255574
rect 182586 255338 182822 255574
rect 182266 219658 182502 219894
rect 182586 219658 182822 219894
rect 182266 219338 182502 219574
rect 182586 219338 182822 219574
rect 182266 183658 182502 183894
rect 182586 183658 182822 183894
rect 182266 183338 182502 183574
rect 182586 183338 182822 183574
rect 182266 147658 182502 147894
rect 182586 147658 182822 147894
rect 182266 147338 182502 147574
rect 182586 147338 182822 147574
rect 182266 111658 182502 111894
rect 182586 111658 182822 111894
rect 182266 111338 182502 111574
rect 182586 111338 182822 111574
rect 182266 75658 182502 75894
rect 182586 75658 182822 75894
rect 182266 75338 182502 75574
rect 182586 75338 182822 75574
rect 182266 39658 182502 39894
rect 182586 39658 182822 39894
rect 182266 39338 182502 39574
rect 182586 39338 182822 39574
rect 182266 3658 182502 3894
rect 182586 3658 182822 3894
rect 182266 3338 182502 3574
rect 182586 3338 182822 3574
rect 182266 -1542 182502 -1306
rect 182586 -1542 182822 -1306
rect 182266 -1862 182502 -1626
rect 182586 -1862 182822 -1626
rect 183506 706522 183742 706758
rect 183826 706522 184062 706758
rect 183506 706202 183742 706438
rect 183826 706202 184062 706438
rect 183506 688898 183742 689134
rect 183826 688898 184062 689134
rect 183506 688578 183742 688814
rect 183826 688578 184062 688814
rect 183506 652898 183742 653134
rect 183826 652898 184062 653134
rect 183506 652578 183742 652814
rect 183826 652578 184062 652814
rect 183506 616898 183742 617134
rect 183826 616898 184062 617134
rect 183506 616578 183742 616814
rect 183826 616578 184062 616814
rect 183506 580898 183742 581134
rect 183826 580898 184062 581134
rect 183506 580578 183742 580814
rect 183826 580578 184062 580814
rect 183506 544898 183742 545134
rect 183826 544898 184062 545134
rect 183506 544578 183742 544814
rect 183826 544578 184062 544814
rect 183506 508898 183742 509134
rect 183826 508898 184062 509134
rect 183506 508578 183742 508814
rect 183826 508578 184062 508814
rect 183506 472898 183742 473134
rect 183826 472898 184062 473134
rect 183506 472578 183742 472814
rect 183826 472578 184062 472814
rect 183506 436898 183742 437134
rect 183826 436898 184062 437134
rect 183506 436578 183742 436814
rect 183826 436578 184062 436814
rect 183506 400898 183742 401134
rect 183826 400898 184062 401134
rect 183506 400578 183742 400814
rect 183826 400578 184062 400814
rect 183506 364898 183742 365134
rect 183826 364898 184062 365134
rect 183506 364578 183742 364814
rect 183826 364578 184062 364814
rect 183506 328898 183742 329134
rect 183826 328898 184062 329134
rect 183506 328578 183742 328814
rect 183826 328578 184062 328814
rect 183506 292898 183742 293134
rect 183826 292898 184062 293134
rect 183506 292578 183742 292814
rect 183826 292578 184062 292814
rect 183506 256898 183742 257134
rect 183826 256898 184062 257134
rect 183506 256578 183742 256814
rect 183826 256578 184062 256814
rect 183506 220898 183742 221134
rect 183826 220898 184062 221134
rect 183506 220578 183742 220814
rect 183826 220578 184062 220814
rect 183506 184898 183742 185134
rect 183826 184898 184062 185134
rect 183506 184578 183742 184814
rect 183826 184578 184062 184814
rect 183506 148898 183742 149134
rect 183826 148898 184062 149134
rect 183506 148578 183742 148814
rect 183826 148578 184062 148814
rect 183506 112898 183742 113134
rect 183826 112898 184062 113134
rect 183506 112578 183742 112814
rect 183826 112578 184062 112814
rect 183506 76898 183742 77134
rect 183826 76898 184062 77134
rect 183506 76578 183742 76814
rect 183826 76578 184062 76814
rect 183506 40898 183742 41134
rect 183826 40898 184062 41134
rect 183506 40578 183742 40814
rect 183826 40578 184062 40814
rect 183506 4898 183742 5134
rect 183826 4898 184062 5134
rect 183506 4578 183742 4814
rect 183826 4578 184062 4814
rect 183506 -2502 183742 -2266
rect 183826 -2502 184062 -2266
rect 183506 -2822 183742 -2586
rect 183826 -2822 184062 -2586
rect 184746 707482 184982 707718
rect 185066 707482 185302 707718
rect 184746 707162 184982 707398
rect 185066 707162 185302 707398
rect 184746 690138 184982 690374
rect 185066 690138 185302 690374
rect 184746 689818 184982 690054
rect 185066 689818 185302 690054
rect 184746 654138 184982 654374
rect 185066 654138 185302 654374
rect 184746 653818 184982 654054
rect 185066 653818 185302 654054
rect 184746 618138 184982 618374
rect 185066 618138 185302 618374
rect 184746 617818 184982 618054
rect 185066 617818 185302 618054
rect 184746 582138 184982 582374
rect 185066 582138 185302 582374
rect 184746 581818 184982 582054
rect 185066 581818 185302 582054
rect 184746 546138 184982 546374
rect 185066 546138 185302 546374
rect 184746 545818 184982 546054
rect 185066 545818 185302 546054
rect 184746 510138 184982 510374
rect 185066 510138 185302 510374
rect 184746 509818 184982 510054
rect 185066 509818 185302 510054
rect 184746 474138 184982 474374
rect 185066 474138 185302 474374
rect 184746 473818 184982 474054
rect 185066 473818 185302 474054
rect 184746 438138 184982 438374
rect 185066 438138 185302 438374
rect 184746 437818 184982 438054
rect 185066 437818 185302 438054
rect 184746 402138 184982 402374
rect 185066 402138 185302 402374
rect 184746 401818 184982 402054
rect 185066 401818 185302 402054
rect 184746 366138 184982 366374
rect 185066 366138 185302 366374
rect 184746 365818 184982 366054
rect 185066 365818 185302 366054
rect 184746 330138 184982 330374
rect 185066 330138 185302 330374
rect 184746 329818 184982 330054
rect 185066 329818 185302 330054
rect 184746 294138 184982 294374
rect 185066 294138 185302 294374
rect 184746 293818 184982 294054
rect 185066 293818 185302 294054
rect 184746 258138 184982 258374
rect 185066 258138 185302 258374
rect 184746 257818 184982 258054
rect 185066 257818 185302 258054
rect 184746 222138 184982 222374
rect 185066 222138 185302 222374
rect 184746 221818 184982 222054
rect 185066 221818 185302 222054
rect 184746 186138 184982 186374
rect 185066 186138 185302 186374
rect 184746 185818 184982 186054
rect 185066 185818 185302 186054
rect 184746 150138 184982 150374
rect 185066 150138 185302 150374
rect 184746 149818 184982 150054
rect 185066 149818 185302 150054
rect 184746 114138 184982 114374
rect 185066 114138 185302 114374
rect 184746 113818 184982 114054
rect 185066 113818 185302 114054
rect 184746 78138 184982 78374
rect 185066 78138 185302 78374
rect 184746 77818 184982 78054
rect 185066 77818 185302 78054
rect 184746 42138 184982 42374
rect 185066 42138 185302 42374
rect 184746 41818 184982 42054
rect 185066 41818 185302 42054
rect 184746 6138 184982 6374
rect 185066 6138 185302 6374
rect 184746 5818 184982 6054
rect 185066 5818 185302 6054
rect 184746 -3462 184982 -3226
rect 185066 -3462 185302 -3226
rect 184746 -3782 184982 -3546
rect 185066 -3782 185302 -3546
rect 185986 708442 186222 708678
rect 186306 708442 186542 708678
rect 185986 708122 186222 708358
rect 186306 708122 186542 708358
rect 185986 691378 186222 691614
rect 186306 691378 186542 691614
rect 185986 691058 186222 691294
rect 186306 691058 186542 691294
rect 185986 655378 186222 655614
rect 186306 655378 186542 655614
rect 185986 655058 186222 655294
rect 186306 655058 186542 655294
rect 185986 619378 186222 619614
rect 186306 619378 186542 619614
rect 185986 619058 186222 619294
rect 186306 619058 186542 619294
rect 185986 583378 186222 583614
rect 186306 583378 186542 583614
rect 185986 583058 186222 583294
rect 186306 583058 186542 583294
rect 185986 547378 186222 547614
rect 186306 547378 186542 547614
rect 185986 547058 186222 547294
rect 186306 547058 186542 547294
rect 185986 511378 186222 511614
rect 186306 511378 186542 511614
rect 185986 511058 186222 511294
rect 186306 511058 186542 511294
rect 185986 475378 186222 475614
rect 186306 475378 186542 475614
rect 185986 475058 186222 475294
rect 186306 475058 186542 475294
rect 185986 439378 186222 439614
rect 186306 439378 186542 439614
rect 185986 439058 186222 439294
rect 186306 439058 186542 439294
rect 185986 403378 186222 403614
rect 186306 403378 186542 403614
rect 185986 403058 186222 403294
rect 186306 403058 186542 403294
rect 185986 367378 186222 367614
rect 186306 367378 186542 367614
rect 185986 367058 186222 367294
rect 186306 367058 186542 367294
rect 185986 331378 186222 331614
rect 186306 331378 186542 331614
rect 185986 331058 186222 331294
rect 186306 331058 186542 331294
rect 185986 295378 186222 295614
rect 186306 295378 186542 295614
rect 185986 295058 186222 295294
rect 186306 295058 186542 295294
rect 185986 259378 186222 259614
rect 186306 259378 186542 259614
rect 185986 259058 186222 259294
rect 186306 259058 186542 259294
rect 185986 223378 186222 223614
rect 186306 223378 186542 223614
rect 185986 223058 186222 223294
rect 186306 223058 186542 223294
rect 185986 187378 186222 187614
rect 186306 187378 186542 187614
rect 185986 187058 186222 187294
rect 186306 187058 186542 187294
rect 185986 151378 186222 151614
rect 186306 151378 186542 151614
rect 185986 151058 186222 151294
rect 186306 151058 186542 151294
rect 185986 115378 186222 115614
rect 186306 115378 186542 115614
rect 185986 115058 186222 115294
rect 186306 115058 186542 115294
rect 185986 79378 186222 79614
rect 186306 79378 186542 79614
rect 185986 79058 186222 79294
rect 186306 79058 186542 79294
rect 185986 43378 186222 43614
rect 186306 43378 186542 43614
rect 185986 43058 186222 43294
rect 186306 43058 186542 43294
rect 185986 7378 186222 7614
rect 186306 7378 186542 7614
rect 185986 7058 186222 7294
rect 186306 7058 186542 7294
rect 185986 -4422 186222 -4186
rect 186306 -4422 186542 -4186
rect 185986 -4742 186222 -4506
rect 186306 -4742 186542 -4506
rect 187226 709402 187462 709638
rect 187546 709402 187782 709638
rect 187226 709082 187462 709318
rect 187546 709082 187782 709318
rect 187226 692618 187462 692854
rect 187546 692618 187782 692854
rect 187226 692298 187462 692534
rect 187546 692298 187782 692534
rect 187226 656618 187462 656854
rect 187546 656618 187782 656854
rect 187226 656298 187462 656534
rect 187546 656298 187782 656534
rect 187226 620618 187462 620854
rect 187546 620618 187782 620854
rect 187226 620298 187462 620534
rect 187546 620298 187782 620534
rect 187226 584618 187462 584854
rect 187546 584618 187782 584854
rect 187226 584298 187462 584534
rect 187546 584298 187782 584534
rect 187226 548618 187462 548854
rect 187546 548618 187782 548854
rect 187226 548298 187462 548534
rect 187546 548298 187782 548534
rect 187226 512618 187462 512854
rect 187546 512618 187782 512854
rect 187226 512298 187462 512534
rect 187546 512298 187782 512534
rect 187226 476618 187462 476854
rect 187546 476618 187782 476854
rect 187226 476298 187462 476534
rect 187546 476298 187782 476534
rect 187226 440618 187462 440854
rect 187546 440618 187782 440854
rect 187226 440298 187462 440534
rect 187546 440298 187782 440534
rect 187226 404618 187462 404854
rect 187546 404618 187782 404854
rect 187226 404298 187462 404534
rect 187546 404298 187782 404534
rect 187226 368618 187462 368854
rect 187546 368618 187782 368854
rect 187226 368298 187462 368534
rect 187546 368298 187782 368534
rect 187226 332618 187462 332854
rect 187546 332618 187782 332854
rect 187226 332298 187462 332534
rect 187546 332298 187782 332534
rect 187226 296618 187462 296854
rect 187546 296618 187782 296854
rect 187226 296298 187462 296534
rect 187546 296298 187782 296534
rect 187226 260618 187462 260854
rect 187546 260618 187782 260854
rect 187226 260298 187462 260534
rect 187546 260298 187782 260534
rect 187226 224618 187462 224854
rect 187546 224618 187782 224854
rect 187226 224298 187462 224534
rect 187546 224298 187782 224534
rect 187226 188618 187462 188854
rect 187546 188618 187782 188854
rect 187226 188298 187462 188534
rect 187546 188298 187782 188534
rect 187226 152618 187462 152854
rect 187546 152618 187782 152854
rect 187226 152298 187462 152534
rect 187546 152298 187782 152534
rect 187226 116618 187462 116854
rect 187546 116618 187782 116854
rect 187226 116298 187462 116534
rect 187546 116298 187782 116534
rect 187226 80618 187462 80854
rect 187546 80618 187782 80854
rect 187226 80298 187462 80534
rect 187546 80298 187782 80534
rect 187226 44618 187462 44854
rect 187546 44618 187782 44854
rect 187226 44298 187462 44534
rect 187546 44298 187782 44534
rect 187226 8618 187462 8854
rect 187546 8618 187782 8854
rect 187226 8298 187462 8534
rect 187546 8298 187782 8534
rect 187226 -5382 187462 -5146
rect 187546 -5382 187782 -5146
rect 187226 -5702 187462 -5466
rect 187546 -5702 187782 -5466
rect 188466 710362 188702 710598
rect 188786 710362 189022 710598
rect 188466 710042 188702 710278
rect 188786 710042 189022 710278
rect 188466 693858 188702 694094
rect 188786 693858 189022 694094
rect 188466 693538 188702 693774
rect 188786 693538 189022 693774
rect 188466 657858 188702 658094
rect 188786 657858 189022 658094
rect 188466 657538 188702 657774
rect 188786 657538 189022 657774
rect 188466 621858 188702 622094
rect 188786 621858 189022 622094
rect 188466 621538 188702 621774
rect 188786 621538 189022 621774
rect 188466 585858 188702 586094
rect 188786 585858 189022 586094
rect 188466 585538 188702 585774
rect 188786 585538 189022 585774
rect 188466 549858 188702 550094
rect 188786 549858 189022 550094
rect 188466 549538 188702 549774
rect 188786 549538 189022 549774
rect 188466 513858 188702 514094
rect 188786 513858 189022 514094
rect 188466 513538 188702 513774
rect 188786 513538 189022 513774
rect 188466 477858 188702 478094
rect 188786 477858 189022 478094
rect 188466 477538 188702 477774
rect 188786 477538 189022 477774
rect 188466 441858 188702 442094
rect 188786 441858 189022 442094
rect 188466 441538 188702 441774
rect 188786 441538 189022 441774
rect 188466 405858 188702 406094
rect 188786 405858 189022 406094
rect 188466 405538 188702 405774
rect 188786 405538 189022 405774
rect 188466 369858 188702 370094
rect 188786 369858 189022 370094
rect 188466 369538 188702 369774
rect 188786 369538 189022 369774
rect 188466 333858 188702 334094
rect 188786 333858 189022 334094
rect 188466 333538 188702 333774
rect 188786 333538 189022 333774
rect 188466 297858 188702 298094
rect 188786 297858 189022 298094
rect 188466 297538 188702 297774
rect 188786 297538 189022 297774
rect 188466 261858 188702 262094
rect 188786 261858 189022 262094
rect 188466 261538 188702 261774
rect 188786 261538 189022 261774
rect 188466 225858 188702 226094
rect 188786 225858 189022 226094
rect 188466 225538 188702 225774
rect 188786 225538 189022 225774
rect 188466 189858 188702 190094
rect 188786 189858 189022 190094
rect 188466 189538 188702 189774
rect 188786 189538 189022 189774
rect 188466 153858 188702 154094
rect 188786 153858 189022 154094
rect 188466 153538 188702 153774
rect 188786 153538 189022 153774
rect 188466 117858 188702 118094
rect 188786 117858 189022 118094
rect 188466 117538 188702 117774
rect 188786 117538 189022 117774
rect 188466 81858 188702 82094
rect 188786 81858 189022 82094
rect 188466 81538 188702 81774
rect 188786 81538 189022 81774
rect 188466 45858 188702 46094
rect 188786 45858 189022 46094
rect 188466 45538 188702 45774
rect 188786 45538 189022 45774
rect 188466 9858 188702 10094
rect 188786 9858 189022 10094
rect 188466 9538 188702 9774
rect 188786 9538 189022 9774
rect 188466 -6342 188702 -6106
rect 188786 -6342 189022 -6106
rect 188466 -6662 188702 -6426
rect 188786 -6662 189022 -6426
rect 189706 711322 189942 711558
rect 190026 711322 190262 711558
rect 189706 711002 189942 711238
rect 190026 711002 190262 711238
rect 189706 695098 189942 695334
rect 190026 695098 190262 695334
rect 189706 694778 189942 695014
rect 190026 694778 190262 695014
rect 189706 659098 189942 659334
rect 190026 659098 190262 659334
rect 189706 658778 189942 659014
rect 190026 658778 190262 659014
rect 189706 623098 189942 623334
rect 190026 623098 190262 623334
rect 189706 622778 189942 623014
rect 190026 622778 190262 623014
rect 189706 587098 189942 587334
rect 190026 587098 190262 587334
rect 189706 586778 189942 587014
rect 190026 586778 190262 587014
rect 189706 551098 189942 551334
rect 190026 551098 190262 551334
rect 189706 550778 189942 551014
rect 190026 550778 190262 551014
rect 189706 515098 189942 515334
rect 190026 515098 190262 515334
rect 189706 514778 189942 515014
rect 190026 514778 190262 515014
rect 189706 479098 189942 479334
rect 190026 479098 190262 479334
rect 189706 478778 189942 479014
rect 190026 478778 190262 479014
rect 189706 443098 189942 443334
rect 190026 443098 190262 443334
rect 189706 442778 189942 443014
rect 190026 442778 190262 443014
rect 189706 407098 189942 407334
rect 190026 407098 190262 407334
rect 189706 406778 189942 407014
rect 190026 406778 190262 407014
rect 189706 371098 189942 371334
rect 190026 371098 190262 371334
rect 189706 370778 189942 371014
rect 190026 370778 190262 371014
rect 189706 335098 189942 335334
rect 190026 335098 190262 335334
rect 189706 334778 189942 335014
rect 190026 334778 190262 335014
rect 189706 299098 189942 299334
rect 190026 299098 190262 299334
rect 189706 298778 189942 299014
rect 190026 298778 190262 299014
rect 189706 263098 189942 263334
rect 190026 263098 190262 263334
rect 189706 262778 189942 263014
rect 190026 262778 190262 263014
rect 189706 227098 189942 227334
rect 190026 227098 190262 227334
rect 189706 226778 189942 227014
rect 190026 226778 190262 227014
rect 189706 191098 189942 191334
rect 190026 191098 190262 191334
rect 189706 190778 189942 191014
rect 190026 190778 190262 191014
rect 189706 155098 189942 155334
rect 190026 155098 190262 155334
rect 189706 154778 189942 155014
rect 190026 154778 190262 155014
rect 189706 119098 189942 119334
rect 190026 119098 190262 119334
rect 189706 118778 189942 119014
rect 190026 118778 190262 119014
rect 189706 83098 189942 83334
rect 190026 83098 190262 83334
rect 189706 82778 189942 83014
rect 190026 82778 190262 83014
rect 189706 47098 189942 47334
rect 190026 47098 190262 47334
rect 189706 46778 189942 47014
rect 190026 46778 190262 47014
rect 189706 11098 189942 11334
rect 190026 11098 190262 11334
rect 189706 10778 189942 11014
rect 190026 10778 190262 11014
rect 189706 -7302 189942 -7066
rect 190026 -7302 190262 -7066
rect 189706 -7622 189942 -7386
rect 190026 -7622 190262 -7386
rect 217026 704602 217262 704838
rect 217346 704602 217582 704838
rect 217026 704282 217262 704518
rect 217346 704282 217582 704518
rect 217026 686418 217262 686654
rect 217346 686418 217582 686654
rect 217026 686098 217262 686334
rect 217346 686098 217582 686334
rect 217026 650418 217262 650654
rect 217346 650418 217582 650654
rect 217026 650098 217262 650334
rect 217346 650098 217582 650334
rect 217026 614418 217262 614654
rect 217346 614418 217582 614654
rect 217026 614098 217262 614334
rect 217346 614098 217582 614334
rect 217026 578418 217262 578654
rect 217346 578418 217582 578654
rect 217026 578098 217262 578334
rect 217346 578098 217582 578334
rect 217026 542418 217262 542654
rect 217346 542418 217582 542654
rect 217026 542098 217262 542334
rect 217346 542098 217582 542334
rect 217026 506418 217262 506654
rect 217346 506418 217582 506654
rect 217026 506098 217262 506334
rect 217346 506098 217582 506334
rect 217026 470418 217262 470654
rect 217346 470418 217582 470654
rect 217026 470098 217262 470334
rect 217346 470098 217582 470334
rect 217026 434418 217262 434654
rect 217346 434418 217582 434654
rect 217026 434098 217262 434334
rect 217346 434098 217582 434334
rect 217026 398418 217262 398654
rect 217346 398418 217582 398654
rect 217026 398098 217262 398334
rect 217346 398098 217582 398334
rect 217026 362418 217262 362654
rect 217346 362418 217582 362654
rect 217026 362098 217262 362334
rect 217346 362098 217582 362334
rect 217026 326418 217262 326654
rect 217346 326418 217582 326654
rect 217026 326098 217262 326334
rect 217346 326098 217582 326334
rect 217026 290418 217262 290654
rect 217346 290418 217582 290654
rect 217026 290098 217262 290334
rect 217346 290098 217582 290334
rect 217026 254418 217262 254654
rect 217346 254418 217582 254654
rect 217026 254098 217262 254334
rect 217346 254098 217582 254334
rect 217026 218418 217262 218654
rect 217346 218418 217582 218654
rect 217026 218098 217262 218334
rect 217346 218098 217582 218334
rect 217026 182418 217262 182654
rect 217346 182418 217582 182654
rect 217026 182098 217262 182334
rect 217346 182098 217582 182334
rect 217026 146418 217262 146654
rect 217346 146418 217582 146654
rect 217026 146098 217262 146334
rect 217346 146098 217582 146334
rect 217026 110418 217262 110654
rect 217346 110418 217582 110654
rect 217026 110098 217262 110334
rect 217346 110098 217582 110334
rect 217026 74418 217262 74654
rect 217346 74418 217582 74654
rect 217026 74098 217262 74334
rect 217346 74098 217582 74334
rect 217026 38418 217262 38654
rect 217346 38418 217582 38654
rect 217026 38098 217262 38334
rect 217346 38098 217582 38334
rect 217026 2418 217262 2654
rect 217346 2418 217582 2654
rect 217026 2098 217262 2334
rect 217346 2098 217582 2334
rect 217026 -582 217262 -346
rect 217346 -582 217582 -346
rect 217026 -902 217262 -666
rect 217346 -902 217582 -666
rect 218266 705562 218502 705798
rect 218586 705562 218822 705798
rect 218266 705242 218502 705478
rect 218586 705242 218822 705478
rect 218266 687658 218502 687894
rect 218586 687658 218822 687894
rect 218266 687338 218502 687574
rect 218586 687338 218822 687574
rect 218266 651658 218502 651894
rect 218586 651658 218822 651894
rect 218266 651338 218502 651574
rect 218586 651338 218822 651574
rect 218266 615658 218502 615894
rect 218586 615658 218822 615894
rect 218266 615338 218502 615574
rect 218586 615338 218822 615574
rect 218266 579658 218502 579894
rect 218586 579658 218822 579894
rect 218266 579338 218502 579574
rect 218586 579338 218822 579574
rect 218266 543658 218502 543894
rect 218586 543658 218822 543894
rect 218266 543338 218502 543574
rect 218586 543338 218822 543574
rect 218266 507658 218502 507894
rect 218586 507658 218822 507894
rect 218266 507338 218502 507574
rect 218586 507338 218822 507574
rect 218266 471658 218502 471894
rect 218586 471658 218822 471894
rect 218266 471338 218502 471574
rect 218586 471338 218822 471574
rect 218266 435658 218502 435894
rect 218586 435658 218822 435894
rect 218266 435338 218502 435574
rect 218586 435338 218822 435574
rect 218266 399658 218502 399894
rect 218586 399658 218822 399894
rect 218266 399338 218502 399574
rect 218586 399338 218822 399574
rect 218266 363658 218502 363894
rect 218586 363658 218822 363894
rect 218266 363338 218502 363574
rect 218586 363338 218822 363574
rect 218266 327658 218502 327894
rect 218586 327658 218822 327894
rect 218266 327338 218502 327574
rect 218586 327338 218822 327574
rect 218266 291658 218502 291894
rect 218586 291658 218822 291894
rect 218266 291338 218502 291574
rect 218586 291338 218822 291574
rect 218266 255658 218502 255894
rect 218586 255658 218822 255894
rect 218266 255338 218502 255574
rect 218586 255338 218822 255574
rect 218266 219658 218502 219894
rect 218586 219658 218822 219894
rect 218266 219338 218502 219574
rect 218586 219338 218822 219574
rect 218266 183658 218502 183894
rect 218586 183658 218822 183894
rect 218266 183338 218502 183574
rect 218586 183338 218822 183574
rect 218266 147658 218502 147894
rect 218586 147658 218822 147894
rect 218266 147338 218502 147574
rect 218586 147338 218822 147574
rect 218266 111658 218502 111894
rect 218586 111658 218822 111894
rect 218266 111338 218502 111574
rect 218586 111338 218822 111574
rect 218266 75658 218502 75894
rect 218586 75658 218822 75894
rect 218266 75338 218502 75574
rect 218586 75338 218822 75574
rect 218266 39658 218502 39894
rect 218586 39658 218822 39894
rect 218266 39338 218502 39574
rect 218586 39338 218822 39574
rect 218266 3658 218502 3894
rect 218586 3658 218822 3894
rect 218266 3338 218502 3574
rect 218586 3338 218822 3574
rect 218266 -1542 218502 -1306
rect 218586 -1542 218822 -1306
rect 218266 -1862 218502 -1626
rect 218586 -1862 218822 -1626
rect 219506 706522 219742 706758
rect 219826 706522 220062 706758
rect 219506 706202 219742 706438
rect 219826 706202 220062 706438
rect 219506 688898 219742 689134
rect 219826 688898 220062 689134
rect 219506 688578 219742 688814
rect 219826 688578 220062 688814
rect 219506 652898 219742 653134
rect 219826 652898 220062 653134
rect 219506 652578 219742 652814
rect 219826 652578 220062 652814
rect 219506 616898 219742 617134
rect 219826 616898 220062 617134
rect 219506 616578 219742 616814
rect 219826 616578 220062 616814
rect 219506 580898 219742 581134
rect 219826 580898 220062 581134
rect 219506 580578 219742 580814
rect 219826 580578 220062 580814
rect 219506 544898 219742 545134
rect 219826 544898 220062 545134
rect 219506 544578 219742 544814
rect 219826 544578 220062 544814
rect 219506 508898 219742 509134
rect 219826 508898 220062 509134
rect 219506 508578 219742 508814
rect 219826 508578 220062 508814
rect 219506 472898 219742 473134
rect 219826 472898 220062 473134
rect 219506 472578 219742 472814
rect 219826 472578 220062 472814
rect 219506 436898 219742 437134
rect 219826 436898 220062 437134
rect 219506 436578 219742 436814
rect 219826 436578 220062 436814
rect 219506 400898 219742 401134
rect 219826 400898 220062 401134
rect 219506 400578 219742 400814
rect 219826 400578 220062 400814
rect 219506 364898 219742 365134
rect 219826 364898 220062 365134
rect 219506 364578 219742 364814
rect 219826 364578 220062 364814
rect 219506 328898 219742 329134
rect 219826 328898 220062 329134
rect 219506 328578 219742 328814
rect 219826 328578 220062 328814
rect 219506 292898 219742 293134
rect 219826 292898 220062 293134
rect 219506 292578 219742 292814
rect 219826 292578 220062 292814
rect 219506 256898 219742 257134
rect 219826 256898 220062 257134
rect 219506 256578 219742 256814
rect 219826 256578 220062 256814
rect 219506 220898 219742 221134
rect 219826 220898 220062 221134
rect 219506 220578 219742 220814
rect 219826 220578 220062 220814
rect 219506 184898 219742 185134
rect 219826 184898 220062 185134
rect 219506 184578 219742 184814
rect 219826 184578 220062 184814
rect 219506 148898 219742 149134
rect 219826 148898 220062 149134
rect 219506 148578 219742 148814
rect 219826 148578 220062 148814
rect 219506 112898 219742 113134
rect 219826 112898 220062 113134
rect 219506 112578 219742 112814
rect 219826 112578 220062 112814
rect 219506 76898 219742 77134
rect 219826 76898 220062 77134
rect 219506 76578 219742 76814
rect 219826 76578 220062 76814
rect 219506 40898 219742 41134
rect 219826 40898 220062 41134
rect 219506 40578 219742 40814
rect 219826 40578 220062 40814
rect 219506 4898 219742 5134
rect 219826 4898 220062 5134
rect 219506 4578 219742 4814
rect 219826 4578 220062 4814
rect 219506 -2502 219742 -2266
rect 219826 -2502 220062 -2266
rect 219506 -2822 219742 -2586
rect 219826 -2822 220062 -2586
rect 220746 707482 220982 707718
rect 221066 707482 221302 707718
rect 220746 707162 220982 707398
rect 221066 707162 221302 707398
rect 220746 690138 220982 690374
rect 221066 690138 221302 690374
rect 220746 689818 220982 690054
rect 221066 689818 221302 690054
rect 220746 654138 220982 654374
rect 221066 654138 221302 654374
rect 220746 653818 220982 654054
rect 221066 653818 221302 654054
rect 220746 618138 220982 618374
rect 221066 618138 221302 618374
rect 220746 617818 220982 618054
rect 221066 617818 221302 618054
rect 220746 582138 220982 582374
rect 221066 582138 221302 582374
rect 220746 581818 220982 582054
rect 221066 581818 221302 582054
rect 220746 546138 220982 546374
rect 221066 546138 221302 546374
rect 220746 545818 220982 546054
rect 221066 545818 221302 546054
rect 220746 510138 220982 510374
rect 221066 510138 221302 510374
rect 220746 509818 220982 510054
rect 221066 509818 221302 510054
rect 220746 474138 220982 474374
rect 221066 474138 221302 474374
rect 220746 473818 220982 474054
rect 221066 473818 221302 474054
rect 220746 438138 220982 438374
rect 221066 438138 221302 438374
rect 220746 437818 220982 438054
rect 221066 437818 221302 438054
rect 220746 402138 220982 402374
rect 221066 402138 221302 402374
rect 220746 401818 220982 402054
rect 221066 401818 221302 402054
rect 220746 366138 220982 366374
rect 221066 366138 221302 366374
rect 220746 365818 220982 366054
rect 221066 365818 221302 366054
rect 220746 330138 220982 330374
rect 221066 330138 221302 330374
rect 220746 329818 220982 330054
rect 221066 329818 221302 330054
rect 220746 294138 220982 294374
rect 221066 294138 221302 294374
rect 220746 293818 220982 294054
rect 221066 293818 221302 294054
rect 220746 258138 220982 258374
rect 221066 258138 221302 258374
rect 220746 257818 220982 258054
rect 221066 257818 221302 258054
rect 220746 222138 220982 222374
rect 221066 222138 221302 222374
rect 220746 221818 220982 222054
rect 221066 221818 221302 222054
rect 220746 186138 220982 186374
rect 221066 186138 221302 186374
rect 220746 185818 220982 186054
rect 221066 185818 221302 186054
rect 220746 150138 220982 150374
rect 221066 150138 221302 150374
rect 220746 149818 220982 150054
rect 221066 149818 221302 150054
rect 220746 114138 220982 114374
rect 221066 114138 221302 114374
rect 220746 113818 220982 114054
rect 221066 113818 221302 114054
rect 220746 78138 220982 78374
rect 221066 78138 221302 78374
rect 220746 77818 220982 78054
rect 221066 77818 221302 78054
rect 220746 42138 220982 42374
rect 221066 42138 221302 42374
rect 220746 41818 220982 42054
rect 221066 41818 221302 42054
rect 220746 6138 220982 6374
rect 221066 6138 221302 6374
rect 220746 5818 220982 6054
rect 221066 5818 221302 6054
rect 220746 -3462 220982 -3226
rect 221066 -3462 221302 -3226
rect 220746 -3782 220982 -3546
rect 221066 -3782 221302 -3546
rect 221986 708442 222222 708678
rect 222306 708442 222542 708678
rect 221986 708122 222222 708358
rect 222306 708122 222542 708358
rect 221986 691378 222222 691614
rect 222306 691378 222542 691614
rect 221986 691058 222222 691294
rect 222306 691058 222542 691294
rect 221986 655378 222222 655614
rect 222306 655378 222542 655614
rect 221986 655058 222222 655294
rect 222306 655058 222542 655294
rect 221986 619378 222222 619614
rect 222306 619378 222542 619614
rect 221986 619058 222222 619294
rect 222306 619058 222542 619294
rect 221986 583378 222222 583614
rect 222306 583378 222542 583614
rect 221986 583058 222222 583294
rect 222306 583058 222542 583294
rect 221986 547378 222222 547614
rect 222306 547378 222542 547614
rect 221986 547058 222222 547294
rect 222306 547058 222542 547294
rect 221986 511378 222222 511614
rect 222306 511378 222542 511614
rect 221986 511058 222222 511294
rect 222306 511058 222542 511294
rect 221986 475378 222222 475614
rect 222306 475378 222542 475614
rect 221986 475058 222222 475294
rect 222306 475058 222542 475294
rect 221986 439378 222222 439614
rect 222306 439378 222542 439614
rect 221986 439058 222222 439294
rect 222306 439058 222542 439294
rect 221986 403378 222222 403614
rect 222306 403378 222542 403614
rect 221986 403058 222222 403294
rect 222306 403058 222542 403294
rect 221986 367378 222222 367614
rect 222306 367378 222542 367614
rect 221986 367058 222222 367294
rect 222306 367058 222542 367294
rect 221986 331378 222222 331614
rect 222306 331378 222542 331614
rect 221986 331058 222222 331294
rect 222306 331058 222542 331294
rect 221986 295378 222222 295614
rect 222306 295378 222542 295614
rect 221986 295058 222222 295294
rect 222306 295058 222542 295294
rect 221986 259378 222222 259614
rect 222306 259378 222542 259614
rect 221986 259058 222222 259294
rect 222306 259058 222542 259294
rect 221986 223378 222222 223614
rect 222306 223378 222542 223614
rect 221986 223058 222222 223294
rect 222306 223058 222542 223294
rect 221986 187378 222222 187614
rect 222306 187378 222542 187614
rect 221986 187058 222222 187294
rect 222306 187058 222542 187294
rect 221986 151378 222222 151614
rect 222306 151378 222542 151614
rect 221986 151058 222222 151294
rect 222306 151058 222542 151294
rect 221986 115378 222222 115614
rect 222306 115378 222542 115614
rect 221986 115058 222222 115294
rect 222306 115058 222542 115294
rect 221986 79378 222222 79614
rect 222306 79378 222542 79614
rect 221986 79058 222222 79294
rect 222306 79058 222542 79294
rect 221986 43378 222222 43614
rect 222306 43378 222542 43614
rect 221986 43058 222222 43294
rect 222306 43058 222542 43294
rect 221986 7378 222222 7614
rect 222306 7378 222542 7614
rect 221986 7058 222222 7294
rect 222306 7058 222542 7294
rect 221986 -4422 222222 -4186
rect 222306 -4422 222542 -4186
rect 221986 -4742 222222 -4506
rect 222306 -4742 222542 -4506
rect 223226 709402 223462 709638
rect 223546 709402 223782 709638
rect 223226 709082 223462 709318
rect 223546 709082 223782 709318
rect 223226 692618 223462 692854
rect 223546 692618 223782 692854
rect 223226 692298 223462 692534
rect 223546 692298 223782 692534
rect 223226 656618 223462 656854
rect 223546 656618 223782 656854
rect 223226 656298 223462 656534
rect 223546 656298 223782 656534
rect 223226 620618 223462 620854
rect 223546 620618 223782 620854
rect 223226 620298 223462 620534
rect 223546 620298 223782 620534
rect 223226 584618 223462 584854
rect 223546 584618 223782 584854
rect 223226 584298 223462 584534
rect 223546 584298 223782 584534
rect 223226 548618 223462 548854
rect 223546 548618 223782 548854
rect 223226 548298 223462 548534
rect 223546 548298 223782 548534
rect 223226 512618 223462 512854
rect 223546 512618 223782 512854
rect 223226 512298 223462 512534
rect 223546 512298 223782 512534
rect 223226 476618 223462 476854
rect 223546 476618 223782 476854
rect 223226 476298 223462 476534
rect 223546 476298 223782 476534
rect 223226 440618 223462 440854
rect 223546 440618 223782 440854
rect 223226 440298 223462 440534
rect 223546 440298 223782 440534
rect 223226 404618 223462 404854
rect 223546 404618 223782 404854
rect 223226 404298 223462 404534
rect 223546 404298 223782 404534
rect 223226 368618 223462 368854
rect 223546 368618 223782 368854
rect 223226 368298 223462 368534
rect 223546 368298 223782 368534
rect 223226 332618 223462 332854
rect 223546 332618 223782 332854
rect 223226 332298 223462 332534
rect 223546 332298 223782 332534
rect 223226 296618 223462 296854
rect 223546 296618 223782 296854
rect 223226 296298 223462 296534
rect 223546 296298 223782 296534
rect 223226 260618 223462 260854
rect 223546 260618 223782 260854
rect 223226 260298 223462 260534
rect 223546 260298 223782 260534
rect 223226 224618 223462 224854
rect 223546 224618 223782 224854
rect 223226 224298 223462 224534
rect 223546 224298 223782 224534
rect 223226 188618 223462 188854
rect 223546 188618 223782 188854
rect 223226 188298 223462 188534
rect 223546 188298 223782 188534
rect 223226 152618 223462 152854
rect 223546 152618 223782 152854
rect 223226 152298 223462 152534
rect 223546 152298 223782 152534
rect 223226 116618 223462 116854
rect 223546 116618 223782 116854
rect 223226 116298 223462 116534
rect 223546 116298 223782 116534
rect 223226 80618 223462 80854
rect 223546 80618 223782 80854
rect 223226 80298 223462 80534
rect 223546 80298 223782 80534
rect 223226 44618 223462 44854
rect 223546 44618 223782 44854
rect 223226 44298 223462 44534
rect 223546 44298 223782 44534
rect 223226 8618 223462 8854
rect 223546 8618 223782 8854
rect 223226 8298 223462 8534
rect 223546 8298 223782 8534
rect 223226 -5382 223462 -5146
rect 223546 -5382 223782 -5146
rect 223226 -5702 223462 -5466
rect 223546 -5702 223782 -5466
rect 224466 710362 224702 710598
rect 224786 710362 225022 710598
rect 224466 710042 224702 710278
rect 224786 710042 225022 710278
rect 224466 693858 224702 694094
rect 224786 693858 225022 694094
rect 224466 693538 224702 693774
rect 224786 693538 225022 693774
rect 224466 657858 224702 658094
rect 224786 657858 225022 658094
rect 224466 657538 224702 657774
rect 224786 657538 225022 657774
rect 224466 621858 224702 622094
rect 224786 621858 225022 622094
rect 224466 621538 224702 621774
rect 224786 621538 225022 621774
rect 224466 585858 224702 586094
rect 224786 585858 225022 586094
rect 224466 585538 224702 585774
rect 224786 585538 225022 585774
rect 224466 549858 224702 550094
rect 224786 549858 225022 550094
rect 224466 549538 224702 549774
rect 224786 549538 225022 549774
rect 224466 513858 224702 514094
rect 224786 513858 225022 514094
rect 224466 513538 224702 513774
rect 224786 513538 225022 513774
rect 224466 477858 224702 478094
rect 224786 477858 225022 478094
rect 224466 477538 224702 477774
rect 224786 477538 225022 477774
rect 224466 441858 224702 442094
rect 224786 441858 225022 442094
rect 224466 441538 224702 441774
rect 224786 441538 225022 441774
rect 224466 405858 224702 406094
rect 224786 405858 225022 406094
rect 224466 405538 224702 405774
rect 224786 405538 225022 405774
rect 224466 369858 224702 370094
rect 224786 369858 225022 370094
rect 224466 369538 224702 369774
rect 224786 369538 225022 369774
rect 224466 333858 224702 334094
rect 224786 333858 225022 334094
rect 224466 333538 224702 333774
rect 224786 333538 225022 333774
rect 224466 297858 224702 298094
rect 224786 297858 225022 298094
rect 224466 297538 224702 297774
rect 224786 297538 225022 297774
rect 224466 261858 224702 262094
rect 224786 261858 225022 262094
rect 224466 261538 224702 261774
rect 224786 261538 225022 261774
rect 224466 225858 224702 226094
rect 224786 225858 225022 226094
rect 224466 225538 224702 225774
rect 224786 225538 225022 225774
rect 224466 189858 224702 190094
rect 224786 189858 225022 190094
rect 224466 189538 224702 189774
rect 224786 189538 225022 189774
rect 224466 153858 224702 154094
rect 224786 153858 225022 154094
rect 224466 153538 224702 153774
rect 224786 153538 225022 153774
rect 224466 117858 224702 118094
rect 224786 117858 225022 118094
rect 224466 117538 224702 117774
rect 224786 117538 225022 117774
rect 224466 81858 224702 82094
rect 224786 81858 225022 82094
rect 224466 81538 224702 81774
rect 224786 81538 225022 81774
rect 224466 45858 224702 46094
rect 224786 45858 225022 46094
rect 224466 45538 224702 45774
rect 224786 45538 225022 45774
rect 224466 9858 224702 10094
rect 224786 9858 225022 10094
rect 224466 9538 224702 9774
rect 224786 9538 225022 9774
rect 224466 -6342 224702 -6106
rect 224786 -6342 225022 -6106
rect 224466 -6662 224702 -6426
rect 224786 -6662 225022 -6426
rect 225706 711322 225942 711558
rect 226026 711322 226262 711558
rect 225706 711002 225942 711238
rect 226026 711002 226262 711238
rect 225706 695098 225942 695334
rect 226026 695098 226262 695334
rect 225706 694778 225942 695014
rect 226026 694778 226262 695014
rect 225706 659098 225942 659334
rect 226026 659098 226262 659334
rect 225706 658778 225942 659014
rect 226026 658778 226262 659014
rect 225706 623098 225942 623334
rect 226026 623098 226262 623334
rect 225706 622778 225942 623014
rect 226026 622778 226262 623014
rect 225706 587098 225942 587334
rect 226026 587098 226262 587334
rect 225706 586778 225942 587014
rect 226026 586778 226262 587014
rect 225706 551098 225942 551334
rect 226026 551098 226262 551334
rect 225706 550778 225942 551014
rect 226026 550778 226262 551014
rect 225706 515098 225942 515334
rect 226026 515098 226262 515334
rect 225706 514778 225942 515014
rect 226026 514778 226262 515014
rect 225706 479098 225942 479334
rect 226026 479098 226262 479334
rect 225706 478778 225942 479014
rect 226026 478778 226262 479014
rect 225706 443098 225942 443334
rect 226026 443098 226262 443334
rect 225706 442778 225942 443014
rect 226026 442778 226262 443014
rect 225706 407098 225942 407334
rect 226026 407098 226262 407334
rect 225706 406778 225942 407014
rect 226026 406778 226262 407014
rect 225706 371098 225942 371334
rect 226026 371098 226262 371334
rect 225706 370778 225942 371014
rect 226026 370778 226262 371014
rect 225706 335098 225942 335334
rect 226026 335098 226262 335334
rect 225706 334778 225942 335014
rect 226026 334778 226262 335014
rect 225706 299098 225942 299334
rect 226026 299098 226262 299334
rect 225706 298778 225942 299014
rect 226026 298778 226262 299014
rect 225706 263098 225942 263334
rect 226026 263098 226262 263334
rect 225706 262778 225942 263014
rect 226026 262778 226262 263014
rect 225706 227098 225942 227334
rect 226026 227098 226262 227334
rect 225706 226778 225942 227014
rect 226026 226778 226262 227014
rect 225706 191098 225942 191334
rect 226026 191098 226262 191334
rect 225706 190778 225942 191014
rect 226026 190778 226262 191014
rect 225706 155098 225942 155334
rect 226026 155098 226262 155334
rect 225706 154778 225942 155014
rect 226026 154778 226262 155014
rect 225706 119098 225942 119334
rect 226026 119098 226262 119334
rect 225706 118778 225942 119014
rect 226026 118778 226262 119014
rect 225706 83098 225942 83334
rect 226026 83098 226262 83334
rect 225706 82778 225942 83014
rect 226026 82778 226262 83014
rect 225706 47098 225942 47334
rect 226026 47098 226262 47334
rect 225706 46778 225942 47014
rect 226026 46778 226262 47014
rect 225706 11098 225942 11334
rect 226026 11098 226262 11334
rect 225706 10778 225942 11014
rect 226026 10778 226262 11014
rect 225706 -7302 225942 -7066
rect 226026 -7302 226262 -7066
rect 225706 -7622 225942 -7386
rect 226026 -7622 226262 -7386
rect 253026 704602 253262 704838
rect 253346 704602 253582 704838
rect 253026 704282 253262 704518
rect 253346 704282 253582 704518
rect 253026 686418 253262 686654
rect 253346 686418 253582 686654
rect 253026 686098 253262 686334
rect 253346 686098 253582 686334
rect 253026 650418 253262 650654
rect 253346 650418 253582 650654
rect 253026 650098 253262 650334
rect 253346 650098 253582 650334
rect 253026 614418 253262 614654
rect 253346 614418 253582 614654
rect 253026 614098 253262 614334
rect 253346 614098 253582 614334
rect 253026 578418 253262 578654
rect 253346 578418 253582 578654
rect 253026 578098 253262 578334
rect 253346 578098 253582 578334
rect 253026 542418 253262 542654
rect 253346 542418 253582 542654
rect 253026 542098 253262 542334
rect 253346 542098 253582 542334
rect 253026 506418 253262 506654
rect 253346 506418 253582 506654
rect 253026 506098 253262 506334
rect 253346 506098 253582 506334
rect 253026 470418 253262 470654
rect 253346 470418 253582 470654
rect 253026 470098 253262 470334
rect 253346 470098 253582 470334
rect 253026 434418 253262 434654
rect 253346 434418 253582 434654
rect 253026 434098 253262 434334
rect 253346 434098 253582 434334
rect 253026 398418 253262 398654
rect 253346 398418 253582 398654
rect 253026 398098 253262 398334
rect 253346 398098 253582 398334
rect 253026 362418 253262 362654
rect 253346 362418 253582 362654
rect 253026 362098 253262 362334
rect 253346 362098 253582 362334
rect 253026 326418 253262 326654
rect 253346 326418 253582 326654
rect 253026 326098 253262 326334
rect 253346 326098 253582 326334
rect 253026 290418 253262 290654
rect 253346 290418 253582 290654
rect 253026 290098 253262 290334
rect 253346 290098 253582 290334
rect 253026 254418 253262 254654
rect 253346 254418 253582 254654
rect 253026 254098 253262 254334
rect 253346 254098 253582 254334
rect 253026 218418 253262 218654
rect 253346 218418 253582 218654
rect 253026 218098 253262 218334
rect 253346 218098 253582 218334
rect 253026 182418 253262 182654
rect 253346 182418 253582 182654
rect 253026 182098 253262 182334
rect 253346 182098 253582 182334
rect 253026 146418 253262 146654
rect 253346 146418 253582 146654
rect 253026 146098 253262 146334
rect 253346 146098 253582 146334
rect 253026 110418 253262 110654
rect 253346 110418 253582 110654
rect 253026 110098 253262 110334
rect 253346 110098 253582 110334
rect 253026 74418 253262 74654
rect 253346 74418 253582 74654
rect 253026 74098 253262 74334
rect 253346 74098 253582 74334
rect 253026 38418 253262 38654
rect 253346 38418 253582 38654
rect 253026 38098 253262 38334
rect 253346 38098 253582 38334
rect 253026 2418 253262 2654
rect 253346 2418 253582 2654
rect 253026 2098 253262 2334
rect 253346 2098 253582 2334
rect 253026 -582 253262 -346
rect 253346 -582 253582 -346
rect 253026 -902 253262 -666
rect 253346 -902 253582 -666
rect 254266 705562 254502 705798
rect 254586 705562 254822 705798
rect 254266 705242 254502 705478
rect 254586 705242 254822 705478
rect 254266 687658 254502 687894
rect 254586 687658 254822 687894
rect 254266 687338 254502 687574
rect 254586 687338 254822 687574
rect 254266 651658 254502 651894
rect 254586 651658 254822 651894
rect 254266 651338 254502 651574
rect 254586 651338 254822 651574
rect 254266 615658 254502 615894
rect 254586 615658 254822 615894
rect 254266 615338 254502 615574
rect 254586 615338 254822 615574
rect 254266 579658 254502 579894
rect 254586 579658 254822 579894
rect 254266 579338 254502 579574
rect 254586 579338 254822 579574
rect 254266 543658 254502 543894
rect 254586 543658 254822 543894
rect 254266 543338 254502 543574
rect 254586 543338 254822 543574
rect 254266 507658 254502 507894
rect 254586 507658 254822 507894
rect 254266 507338 254502 507574
rect 254586 507338 254822 507574
rect 254266 471658 254502 471894
rect 254586 471658 254822 471894
rect 254266 471338 254502 471574
rect 254586 471338 254822 471574
rect 254266 435658 254502 435894
rect 254586 435658 254822 435894
rect 254266 435338 254502 435574
rect 254586 435338 254822 435574
rect 254266 399658 254502 399894
rect 254586 399658 254822 399894
rect 254266 399338 254502 399574
rect 254586 399338 254822 399574
rect 254266 363658 254502 363894
rect 254586 363658 254822 363894
rect 254266 363338 254502 363574
rect 254586 363338 254822 363574
rect 254266 327658 254502 327894
rect 254586 327658 254822 327894
rect 254266 327338 254502 327574
rect 254586 327338 254822 327574
rect 254266 291658 254502 291894
rect 254586 291658 254822 291894
rect 254266 291338 254502 291574
rect 254586 291338 254822 291574
rect 254266 255658 254502 255894
rect 254586 255658 254822 255894
rect 254266 255338 254502 255574
rect 254586 255338 254822 255574
rect 254266 219658 254502 219894
rect 254586 219658 254822 219894
rect 254266 219338 254502 219574
rect 254586 219338 254822 219574
rect 254266 183658 254502 183894
rect 254586 183658 254822 183894
rect 254266 183338 254502 183574
rect 254586 183338 254822 183574
rect 254266 147658 254502 147894
rect 254586 147658 254822 147894
rect 254266 147338 254502 147574
rect 254586 147338 254822 147574
rect 254266 111658 254502 111894
rect 254586 111658 254822 111894
rect 254266 111338 254502 111574
rect 254586 111338 254822 111574
rect 254266 75658 254502 75894
rect 254586 75658 254822 75894
rect 254266 75338 254502 75574
rect 254586 75338 254822 75574
rect 254266 39658 254502 39894
rect 254586 39658 254822 39894
rect 254266 39338 254502 39574
rect 254586 39338 254822 39574
rect 254266 3658 254502 3894
rect 254586 3658 254822 3894
rect 254266 3338 254502 3574
rect 254586 3338 254822 3574
rect 254266 -1542 254502 -1306
rect 254586 -1542 254822 -1306
rect 254266 -1862 254502 -1626
rect 254586 -1862 254822 -1626
rect 255506 706522 255742 706758
rect 255826 706522 256062 706758
rect 255506 706202 255742 706438
rect 255826 706202 256062 706438
rect 255506 688898 255742 689134
rect 255826 688898 256062 689134
rect 255506 688578 255742 688814
rect 255826 688578 256062 688814
rect 255506 652898 255742 653134
rect 255826 652898 256062 653134
rect 255506 652578 255742 652814
rect 255826 652578 256062 652814
rect 255506 616898 255742 617134
rect 255826 616898 256062 617134
rect 255506 616578 255742 616814
rect 255826 616578 256062 616814
rect 255506 580898 255742 581134
rect 255826 580898 256062 581134
rect 255506 580578 255742 580814
rect 255826 580578 256062 580814
rect 255506 544898 255742 545134
rect 255826 544898 256062 545134
rect 255506 544578 255742 544814
rect 255826 544578 256062 544814
rect 255506 508898 255742 509134
rect 255826 508898 256062 509134
rect 255506 508578 255742 508814
rect 255826 508578 256062 508814
rect 255506 472898 255742 473134
rect 255826 472898 256062 473134
rect 255506 472578 255742 472814
rect 255826 472578 256062 472814
rect 255506 436898 255742 437134
rect 255826 436898 256062 437134
rect 255506 436578 255742 436814
rect 255826 436578 256062 436814
rect 255506 400898 255742 401134
rect 255826 400898 256062 401134
rect 255506 400578 255742 400814
rect 255826 400578 256062 400814
rect 255506 364898 255742 365134
rect 255826 364898 256062 365134
rect 255506 364578 255742 364814
rect 255826 364578 256062 364814
rect 255506 328898 255742 329134
rect 255826 328898 256062 329134
rect 255506 328578 255742 328814
rect 255826 328578 256062 328814
rect 255506 292898 255742 293134
rect 255826 292898 256062 293134
rect 255506 292578 255742 292814
rect 255826 292578 256062 292814
rect 255506 256898 255742 257134
rect 255826 256898 256062 257134
rect 255506 256578 255742 256814
rect 255826 256578 256062 256814
rect 255506 220898 255742 221134
rect 255826 220898 256062 221134
rect 255506 220578 255742 220814
rect 255826 220578 256062 220814
rect 255506 184898 255742 185134
rect 255826 184898 256062 185134
rect 255506 184578 255742 184814
rect 255826 184578 256062 184814
rect 255506 148898 255742 149134
rect 255826 148898 256062 149134
rect 255506 148578 255742 148814
rect 255826 148578 256062 148814
rect 255506 112898 255742 113134
rect 255826 112898 256062 113134
rect 255506 112578 255742 112814
rect 255826 112578 256062 112814
rect 255506 76898 255742 77134
rect 255826 76898 256062 77134
rect 255506 76578 255742 76814
rect 255826 76578 256062 76814
rect 255506 40898 255742 41134
rect 255826 40898 256062 41134
rect 255506 40578 255742 40814
rect 255826 40578 256062 40814
rect 255506 4898 255742 5134
rect 255826 4898 256062 5134
rect 255506 4578 255742 4814
rect 255826 4578 256062 4814
rect 255506 -2502 255742 -2266
rect 255826 -2502 256062 -2266
rect 255506 -2822 255742 -2586
rect 255826 -2822 256062 -2586
rect 256746 707482 256982 707718
rect 257066 707482 257302 707718
rect 256746 707162 256982 707398
rect 257066 707162 257302 707398
rect 256746 690138 256982 690374
rect 257066 690138 257302 690374
rect 256746 689818 256982 690054
rect 257066 689818 257302 690054
rect 256746 654138 256982 654374
rect 257066 654138 257302 654374
rect 256746 653818 256982 654054
rect 257066 653818 257302 654054
rect 256746 618138 256982 618374
rect 257066 618138 257302 618374
rect 256746 617818 256982 618054
rect 257066 617818 257302 618054
rect 256746 582138 256982 582374
rect 257066 582138 257302 582374
rect 256746 581818 256982 582054
rect 257066 581818 257302 582054
rect 256746 546138 256982 546374
rect 257066 546138 257302 546374
rect 256746 545818 256982 546054
rect 257066 545818 257302 546054
rect 256746 510138 256982 510374
rect 257066 510138 257302 510374
rect 256746 509818 256982 510054
rect 257066 509818 257302 510054
rect 256746 474138 256982 474374
rect 257066 474138 257302 474374
rect 256746 473818 256982 474054
rect 257066 473818 257302 474054
rect 256746 438138 256982 438374
rect 257066 438138 257302 438374
rect 256746 437818 256982 438054
rect 257066 437818 257302 438054
rect 256746 402138 256982 402374
rect 257066 402138 257302 402374
rect 256746 401818 256982 402054
rect 257066 401818 257302 402054
rect 256746 366138 256982 366374
rect 257066 366138 257302 366374
rect 256746 365818 256982 366054
rect 257066 365818 257302 366054
rect 256746 330138 256982 330374
rect 257066 330138 257302 330374
rect 256746 329818 256982 330054
rect 257066 329818 257302 330054
rect 256746 294138 256982 294374
rect 257066 294138 257302 294374
rect 256746 293818 256982 294054
rect 257066 293818 257302 294054
rect 256746 258138 256982 258374
rect 257066 258138 257302 258374
rect 256746 257818 256982 258054
rect 257066 257818 257302 258054
rect 256746 222138 256982 222374
rect 257066 222138 257302 222374
rect 256746 221818 256982 222054
rect 257066 221818 257302 222054
rect 256746 186138 256982 186374
rect 257066 186138 257302 186374
rect 256746 185818 256982 186054
rect 257066 185818 257302 186054
rect 256746 150138 256982 150374
rect 257066 150138 257302 150374
rect 256746 149818 256982 150054
rect 257066 149818 257302 150054
rect 256746 114138 256982 114374
rect 257066 114138 257302 114374
rect 256746 113818 256982 114054
rect 257066 113818 257302 114054
rect 256746 78138 256982 78374
rect 257066 78138 257302 78374
rect 256746 77818 256982 78054
rect 257066 77818 257302 78054
rect 256746 42138 256982 42374
rect 257066 42138 257302 42374
rect 256746 41818 256982 42054
rect 257066 41818 257302 42054
rect 256746 6138 256982 6374
rect 257066 6138 257302 6374
rect 256746 5818 256982 6054
rect 257066 5818 257302 6054
rect 256746 -3462 256982 -3226
rect 257066 -3462 257302 -3226
rect 256746 -3782 256982 -3546
rect 257066 -3782 257302 -3546
rect 257986 708442 258222 708678
rect 258306 708442 258542 708678
rect 257986 708122 258222 708358
rect 258306 708122 258542 708358
rect 257986 691378 258222 691614
rect 258306 691378 258542 691614
rect 257986 691058 258222 691294
rect 258306 691058 258542 691294
rect 257986 655378 258222 655614
rect 258306 655378 258542 655614
rect 257986 655058 258222 655294
rect 258306 655058 258542 655294
rect 257986 619378 258222 619614
rect 258306 619378 258542 619614
rect 257986 619058 258222 619294
rect 258306 619058 258542 619294
rect 257986 583378 258222 583614
rect 258306 583378 258542 583614
rect 257986 583058 258222 583294
rect 258306 583058 258542 583294
rect 257986 547378 258222 547614
rect 258306 547378 258542 547614
rect 257986 547058 258222 547294
rect 258306 547058 258542 547294
rect 257986 511378 258222 511614
rect 258306 511378 258542 511614
rect 257986 511058 258222 511294
rect 258306 511058 258542 511294
rect 257986 475378 258222 475614
rect 258306 475378 258542 475614
rect 257986 475058 258222 475294
rect 258306 475058 258542 475294
rect 257986 439378 258222 439614
rect 258306 439378 258542 439614
rect 257986 439058 258222 439294
rect 258306 439058 258542 439294
rect 257986 403378 258222 403614
rect 258306 403378 258542 403614
rect 257986 403058 258222 403294
rect 258306 403058 258542 403294
rect 257986 367378 258222 367614
rect 258306 367378 258542 367614
rect 257986 367058 258222 367294
rect 258306 367058 258542 367294
rect 257986 331378 258222 331614
rect 258306 331378 258542 331614
rect 257986 331058 258222 331294
rect 258306 331058 258542 331294
rect 257986 295378 258222 295614
rect 258306 295378 258542 295614
rect 257986 295058 258222 295294
rect 258306 295058 258542 295294
rect 257986 259378 258222 259614
rect 258306 259378 258542 259614
rect 257986 259058 258222 259294
rect 258306 259058 258542 259294
rect 257986 223378 258222 223614
rect 258306 223378 258542 223614
rect 257986 223058 258222 223294
rect 258306 223058 258542 223294
rect 257986 187378 258222 187614
rect 258306 187378 258542 187614
rect 257986 187058 258222 187294
rect 258306 187058 258542 187294
rect 257986 151378 258222 151614
rect 258306 151378 258542 151614
rect 257986 151058 258222 151294
rect 258306 151058 258542 151294
rect 257986 115378 258222 115614
rect 258306 115378 258542 115614
rect 257986 115058 258222 115294
rect 258306 115058 258542 115294
rect 257986 79378 258222 79614
rect 258306 79378 258542 79614
rect 257986 79058 258222 79294
rect 258306 79058 258542 79294
rect 257986 43378 258222 43614
rect 258306 43378 258542 43614
rect 257986 43058 258222 43294
rect 258306 43058 258542 43294
rect 257986 7378 258222 7614
rect 258306 7378 258542 7614
rect 257986 7058 258222 7294
rect 258306 7058 258542 7294
rect 257986 -4422 258222 -4186
rect 258306 -4422 258542 -4186
rect 257986 -4742 258222 -4506
rect 258306 -4742 258542 -4506
rect 259226 709402 259462 709638
rect 259546 709402 259782 709638
rect 259226 709082 259462 709318
rect 259546 709082 259782 709318
rect 259226 692618 259462 692854
rect 259546 692618 259782 692854
rect 259226 692298 259462 692534
rect 259546 692298 259782 692534
rect 259226 656618 259462 656854
rect 259546 656618 259782 656854
rect 259226 656298 259462 656534
rect 259546 656298 259782 656534
rect 259226 620618 259462 620854
rect 259546 620618 259782 620854
rect 259226 620298 259462 620534
rect 259546 620298 259782 620534
rect 259226 584618 259462 584854
rect 259546 584618 259782 584854
rect 259226 584298 259462 584534
rect 259546 584298 259782 584534
rect 259226 548618 259462 548854
rect 259546 548618 259782 548854
rect 259226 548298 259462 548534
rect 259546 548298 259782 548534
rect 259226 512618 259462 512854
rect 259546 512618 259782 512854
rect 259226 512298 259462 512534
rect 259546 512298 259782 512534
rect 259226 476618 259462 476854
rect 259546 476618 259782 476854
rect 259226 476298 259462 476534
rect 259546 476298 259782 476534
rect 259226 440618 259462 440854
rect 259546 440618 259782 440854
rect 259226 440298 259462 440534
rect 259546 440298 259782 440534
rect 259226 404618 259462 404854
rect 259546 404618 259782 404854
rect 259226 404298 259462 404534
rect 259546 404298 259782 404534
rect 259226 368618 259462 368854
rect 259546 368618 259782 368854
rect 259226 368298 259462 368534
rect 259546 368298 259782 368534
rect 259226 332618 259462 332854
rect 259546 332618 259782 332854
rect 259226 332298 259462 332534
rect 259546 332298 259782 332534
rect 259226 296618 259462 296854
rect 259546 296618 259782 296854
rect 259226 296298 259462 296534
rect 259546 296298 259782 296534
rect 259226 260618 259462 260854
rect 259546 260618 259782 260854
rect 259226 260298 259462 260534
rect 259546 260298 259782 260534
rect 259226 224618 259462 224854
rect 259546 224618 259782 224854
rect 259226 224298 259462 224534
rect 259546 224298 259782 224534
rect 259226 188618 259462 188854
rect 259546 188618 259782 188854
rect 259226 188298 259462 188534
rect 259546 188298 259782 188534
rect 259226 152618 259462 152854
rect 259546 152618 259782 152854
rect 259226 152298 259462 152534
rect 259546 152298 259782 152534
rect 259226 116618 259462 116854
rect 259546 116618 259782 116854
rect 259226 116298 259462 116534
rect 259546 116298 259782 116534
rect 259226 80618 259462 80854
rect 259546 80618 259782 80854
rect 259226 80298 259462 80534
rect 259546 80298 259782 80534
rect 259226 44618 259462 44854
rect 259546 44618 259782 44854
rect 259226 44298 259462 44534
rect 259546 44298 259782 44534
rect 259226 8618 259462 8854
rect 259546 8618 259782 8854
rect 259226 8298 259462 8534
rect 259546 8298 259782 8534
rect 259226 -5382 259462 -5146
rect 259546 -5382 259782 -5146
rect 259226 -5702 259462 -5466
rect 259546 -5702 259782 -5466
rect 260466 710362 260702 710598
rect 260786 710362 261022 710598
rect 260466 710042 260702 710278
rect 260786 710042 261022 710278
rect 260466 693858 260702 694094
rect 260786 693858 261022 694094
rect 260466 693538 260702 693774
rect 260786 693538 261022 693774
rect 260466 657858 260702 658094
rect 260786 657858 261022 658094
rect 260466 657538 260702 657774
rect 260786 657538 261022 657774
rect 260466 621858 260702 622094
rect 260786 621858 261022 622094
rect 260466 621538 260702 621774
rect 260786 621538 261022 621774
rect 260466 585858 260702 586094
rect 260786 585858 261022 586094
rect 260466 585538 260702 585774
rect 260786 585538 261022 585774
rect 260466 549858 260702 550094
rect 260786 549858 261022 550094
rect 260466 549538 260702 549774
rect 260786 549538 261022 549774
rect 260466 513858 260702 514094
rect 260786 513858 261022 514094
rect 260466 513538 260702 513774
rect 260786 513538 261022 513774
rect 260466 477858 260702 478094
rect 260786 477858 261022 478094
rect 260466 477538 260702 477774
rect 260786 477538 261022 477774
rect 260466 441858 260702 442094
rect 260786 441858 261022 442094
rect 260466 441538 260702 441774
rect 260786 441538 261022 441774
rect 260466 405858 260702 406094
rect 260786 405858 261022 406094
rect 260466 405538 260702 405774
rect 260786 405538 261022 405774
rect 260466 369858 260702 370094
rect 260786 369858 261022 370094
rect 260466 369538 260702 369774
rect 260786 369538 261022 369774
rect 260466 333858 260702 334094
rect 260786 333858 261022 334094
rect 260466 333538 260702 333774
rect 260786 333538 261022 333774
rect 260466 297858 260702 298094
rect 260786 297858 261022 298094
rect 260466 297538 260702 297774
rect 260786 297538 261022 297774
rect 260466 261858 260702 262094
rect 260786 261858 261022 262094
rect 260466 261538 260702 261774
rect 260786 261538 261022 261774
rect 260466 225858 260702 226094
rect 260786 225858 261022 226094
rect 260466 225538 260702 225774
rect 260786 225538 261022 225774
rect 260466 189858 260702 190094
rect 260786 189858 261022 190094
rect 260466 189538 260702 189774
rect 260786 189538 261022 189774
rect 260466 153858 260702 154094
rect 260786 153858 261022 154094
rect 260466 153538 260702 153774
rect 260786 153538 261022 153774
rect 260466 117858 260702 118094
rect 260786 117858 261022 118094
rect 260466 117538 260702 117774
rect 260786 117538 261022 117774
rect 260466 81858 260702 82094
rect 260786 81858 261022 82094
rect 260466 81538 260702 81774
rect 260786 81538 261022 81774
rect 260466 45858 260702 46094
rect 260786 45858 261022 46094
rect 260466 45538 260702 45774
rect 260786 45538 261022 45774
rect 260466 9858 260702 10094
rect 260786 9858 261022 10094
rect 260466 9538 260702 9774
rect 260786 9538 261022 9774
rect 260466 -6342 260702 -6106
rect 260786 -6342 261022 -6106
rect 260466 -6662 260702 -6426
rect 260786 -6662 261022 -6426
rect 261706 711322 261942 711558
rect 262026 711322 262262 711558
rect 261706 711002 261942 711238
rect 262026 711002 262262 711238
rect 261706 695098 261942 695334
rect 262026 695098 262262 695334
rect 261706 694778 261942 695014
rect 262026 694778 262262 695014
rect 261706 659098 261942 659334
rect 262026 659098 262262 659334
rect 261706 658778 261942 659014
rect 262026 658778 262262 659014
rect 261706 623098 261942 623334
rect 262026 623098 262262 623334
rect 261706 622778 261942 623014
rect 262026 622778 262262 623014
rect 261706 587098 261942 587334
rect 262026 587098 262262 587334
rect 261706 586778 261942 587014
rect 262026 586778 262262 587014
rect 261706 551098 261942 551334
rect 262026 551098 262262 551334
rect 261706 550778 261942 551014
rect 262026 550778 262262 551014
rect 261706 515098 261942 515334
rect 262026 515098 262262 515334
rect 261706 514778 261942 515014
rect 262026 514778 262262 515014
rect 261706 479098 261942 479334
rect 262026 479098 262262 479334
rect 261706 478778 261942 479014
rect 262026 478778 262262 479014
rect 261706 443098 261942 443334
rect 262026 443098 262262 443334
rect 261706 442778 261942 443014
rect 262026 442778 262262 443014
rect 261706 407098 261942 407334
rect 262026 407098 262262 407334
rect 261706 406778 261942 407014
rect 262026 406778 262262 407014
rect 261706 371098 261942 371334
rect 262026 371098 262262 371334
rect 261706 370778 261942 371014
rect 262026 370778 262262 371014
rect 261706 335098 261942 335334
rect 262026 335098 262262 335334
rect 261706 334778 261942 335014
rect 262026 334778 262262 335014
rect 261706 299098 261942 299334
rect 262026 299098 262262 299334
rect 261706 298778 261942 299014
rect 262026 298778 262262 299014
rect 261706 263098 261942 263334
rect 262026 263098 262262 263334
rect 261706 262778 261942 263014
rect 262026 262778 262262 263014
rect 261706 227098 261942 227334
rect 262026 227098 262262 227334
rect 261706 226778 261942 227014
rect 262026 226778 262262 227014
rect 261706 191098 261942 191334
rect 262026 191098 262262 191334
rect 261706 190778 261942 191014
rect 262026 190778 262262 191014
rect 261706 155098 261942 155334
rect 262026 155098 262262 155334
rect 261706 154778 261942 155014
rect 262026 154778 262262 155014
rect 261706 119098 261942 119334
rect 262026 119098 262262 119334
rect 261706 118778 261942 119014
rect 262026 118778 262262 119014
rect 261706 83098 261942 83334
rect 262026 83098 262262 83334
rect 261706 82778 261942 83014
rect 262026 82778 262262 83014
rect 261706 47098 261942 47334
rect 262026 47098 262262 47334
rect 261706 46778 261942 47014
rect 262026 46778 262262 47014
rect 261706 11098 261942 11334
rect 262026 11098 262262 11334
rect 261706 10778 261942 11014
rect 262026 10778 262262 11014
rect 261706 -7302 261942 -7066
rect 262026 -7302 262262 -7066
rect 261706 -7622 261942 -7386
rect 262026 -7622 262262 -7386
rect 289026 704602 289262 704838
rect 289346 704602 289582 704838
rect 289026 704282 289262 704518
rect 289346 704282 289582 704518
rect 289026 686418 289262 686654
rect 289346 686418 289582 686654
rect 289026 686098 289262 686334
rect 289346 686098 289582 686334
rect 289026 650418 289262 650654
rect 289346 650418 289582 650654
rect 289026 650098 289262 650334
rect 289346 650098 289582 650334
rect 289026 614418 289262 614654
rect 289346 614418 289582 614654
rect 289026 614098 289262 614334
rect 289346 614098 289582 614334
rect 289026 578418 289262 578654
rect 289346 578418 289582 578654
rect 289026 578098 289262 578334
rect 289346 578098 289582 578334
rect 289026 542418 289262 542654
rect 289346 542418 289582 542654
rect 289026 542098 289262 542334
rect 289346 542098 289582 542334
rect 289026 506418 289262 506654
rect 289346 506418 289582 506654
rect 289026 506098 289262 506334
rect 289346 506098 289582 506334
rect 289026 470418 289262 470654
rect 289346 470418 289582 470654
rect 289026 470098 289262 470334
rect 289346 470098 289582 470334
rect 289026 434418 289262 434654
rect 289346 434418 289582 434654
rect 289026 434098 289262 434334
rect 289346 434098 289582 434334
rect 289026 398418 289262 398654
rect 289346 398418 289582 398654
rect 289026 398098 289262 398334
rect 289346 398098 289582 398334
rect 289026 362418 289262 362654
rect 289346 362418 289582 362654
rect 289026 362098 289262 362334
rect 289346 362098 289582 362334
rect 289026 326418 289262 326654
rect 289346 326418 289582 326654
rect 289026 326098 289262 326334
rect 289346 326098 289582 326334
rect 289026 290418 289262 290654
rect 289346 290418 289582 290654
rect 289026 290098 289262 290334
rect 289346 290098 289582 290334
rect 289026 254418 289262 254654
rect 289346 254418 289582 254654
rect 289026 254098 289262 254334
rect 289346 254098 289582 254334
rect 289026 218418 289262 218654
rect 289346 218418 289582 218654
rect 289026 218098 289262 218334
rect 289346 218098 289582 218334
rect 289026 182418 289262 182654
rect 289346 182418 289582 182654
rect 289026 182098 289262 182334
rect 289346 182098 289582 182334
rect 289026 146418 289262 146654
rect 289346 146418 289582 146654
rect 289026 146098 289262 146334
rect 289346 146098 289582 146334
rect 289026 110418 289262 110654
rect 289346 110418 289582 110654
rect 289026 110098 289262 110334
rect 289346 110098 289582 110334
rect 289026 74418 289262 74654
rect 289346 74418 289582 74654
rect 289026 74098 289262 74334
rect 289346 74098 289582 74334
rect 289026 38418 289262 38654
rect 289346 38418 289582 38654
rect 289026 38098 289262 38334
rect 289346 38098 289582 38334
rect 289026 2418 289262 2654
rect 289346 2418 289582 2654
rect 289026 2098 289262 2334
rect 289346 2098 289582 2334
rect 289026 -582 289262 -346
rect 289346 -582 289582 -346
rect 289026 -902 289262 -666
rect 289346 -902 289582 -666
rect 290266 705562 290502 705798
rect 290586 705562 290822 705798
rect 290266 705242 290502 705478
rect 290586 705242 290822 705478
rect 290266 687658 290502 687894
rect 290586 687658 290822 687894
rect 290266 687338 290502 687574
rect 290586 687338 290822 687574
rect 290266 651658 290502 651894
rect 290586 651658 290822 651894
rect 290266 651338 290502 651574
rect 290586 651338 290822 651574
rect 290266 615658 290502 615894
rect 290586 615658 290822 615894
rect 290266 615338 290502 615574
rect 290586 615338 290822 615574
rect 290266 579658 290502 579894
rect 290586 579658 290822 579894
rect 290266 579338 290502 579574
rect 290586 579338 290822 579574
rect 290266 543658 290502 543894
rect 290586 543658 290822 543894
rect 290266 543338 290502 543574
rect 290586 543338 290822 543574
rect 290266 507658 290502 507894
rect 290586 507658 290822 507894
rect 290266 507338 290502 507574
rect 290586 507338 290822 507574
rect 290266 471658 290502 471894
rect 290586 471658 290822 471894
rect 290266 471338 290502 471574
rect 290586 471338 290822 471574
rect 290266 435658 290502 435894
rect 290586 435658 290822 435894
rect 290266 435338 290502 435574
rect 290586 435338 290822 435574
rect 290266 399658 290502 399894
rect 290586 399658 290822 399894
rect 290266 399338 290502 399574
rect 290586 399338 290822 399574
rect 290266 363658 290502 363894
rect 290586 363658 290822 363894
rect 290266 363338 290502 363574
rect 290586 363338 290822 363574
rect 290266 327658 290502 327894
rect 290586 327658 290822 327894
rect 290266 327338 290502 327574
rect 290586 327338 290822 327574
rect 290266 291658 290502 291894
rect 290586 291658 290822 291894
rect 290266 291338 290502 291574
rect 290586 291338 290822 291574
rect 290266 255658 290502 255894
rect 290586 255658 290822 255894
rect 290266 255338 290502 255574
rect 290586 255338 290822 255574
rect 290266 219658 290502 219894
rect 290586 219658 290822 219894
rect 290266 219338 290502 219574
rect 290586 219338 290822 219574
rect 290266 183658 290502 183894
rect 290586 183658 290822 183894
rect 290266 183338 290502 183574
rect 290586 183338 290822 183574
rect 290266 147658 290502 147894
rect 290586 147658 290822 147894
rect 290266 147338 290502 147574
rect 290586 147338 290822 147574
rect 290266 111658 290502 111894
rect 290586 111658 290822 111894
rect 290266 111338 290502 111574
rect 290586 111338 290822 111574
rect 290266 75658 290502 75894
rect 290586 75658 290822 75894
rect 290266 75338 290502 75574
rect 290586 75338 290822 75574
rect 290266 39658 290502 39894
rect 290586 39658 290822 39894
rect 290266 39338 290502 39574
rect 290586 39338 290822 39574
rect 290266 3658 290502 3894
rect 290586 3658 290822 3894
rect 290266 3338 290502 3574
rect 290586 3338 290822 3574
rect 290266 -1542 290502 -1306
rect 290586 -1542 290822 -1306
rect 290266 -1862 290502 -1626
rect 290586 -1862 290822 -1626
rect 291506 706522 291742 706758
rect 291826 706522 292062 706758
rect 291506 706202 291742 706438
rect 291826 706202 292062 706438
rect 291506 688898 291742 689134
rect 291826 688898 292062 689134
rect 291506 688578 291742 688814
rect 291826 688578 292062 688814
rect 291506 652898 291742 653134
rect 291826 652898 292062 653134
rect 291506 652578 291742 652814
rect 291826 652578 292062 652814
rect 291506 616898 291742 617134
rect 291826 616898 292062 617134
rect 291506 616578 291742 616814
rect 291826 616578 292062 616814
rect 291506 580898 291742 581134
rect 291826 580898 292062 581134
rect 291506 580578 291742 580814
rect 291826 580578 292062 580814
rect 291506 544898 291742 545134
rect 291826 544898 292062 545134
rect 291506 544578 291742 544814
rect 291826 544578 292062 544814
rect 291506 508898 291742 509134
rect 291826 508898 292062 509134
rect 291506 508578 291742 508814
rect 291826 508578 292062 508814
rect 291506 472898 291742 473134
rect 291826 472898 292062 473134
rect 291506 472578 291742 472814
rect 291826 472578 292062 472814
rect 291506 436898 291742 437134
rect 291826 436898 292062 437134
rect 291506 436578 291742 436814
rect 291826 436578 292062 436814
rect 291506 400898 291742 401134
rect 291826 400898 292062 401134
rect 291506 400578 291742 400814
rect 291826 400578 292062 400814
rect 291506 364898 291742 365134
rect 291826 364898 292062 365134
rect 291506 364578 291742 364814
rect 291826 364578 292062 364814
rect 291506 328898 291742 329134
rect 291826 328898 292062 329134
rect 291506 328578 291742 328814
rect 291826 328578 292062 328814
rect 291506 292898 291742 293134
rect 291826 292898 292062 293134
rect 291506 292578 291742 292814
rect 291826 292578 292062 292814
rect 291506 256898 291742 257134
rect 291826 256898 292062 257134
rect 291506 256578 291742 256814
rect 291826 256578 292062 256814
rect 291506 220898 291742 221134
rect 291826 220898 292062 221134
rect 291506 220578 291742 220814
rect 291826 220578 292062 220814
rect 291506 184898 291742 185134
rect 291826 184898 292062 185134
rect 291506 184578 291742 184814
rect 291826 184578 292062 184814
rect 291506 148898 291742 149134
rect 291826 148898 292062 149134
rect 291506 148578 291742 148814
rect 291826 148578 292062 148814
rect 291506 112898 291742 113134
rect 291826 112898 292062 113134
rect 291506 112578 291742 112814
rect 291826 112578 292062 112814
rect 291506 76898 291742 77134
rect 291826 76898 292062 77134
rect 291506 76578 291742 76814
rect 291826 76578 292062 76814
rect 291506 40898 291742 41134
rect 291826 40898 292062 41134
rect 291506 40578 291742 40814
rect 291826 40578 292062 40814
rect 291506 4898 291742 5134
rect 291826 4898 292062 5134
rect 291506 4578 291742 4814
rect 291826 4578 292062 4814
rect 291506 -2502 291742 -2266
rect 291826 -2502 292062 -2266
rect 291506 -2822 291742 -2586
rect 291826 -2822 292062 -2586
rect 292746 707482 292982 707718
rect 293066 707482 293302 707718
rect 292746 707162 292982 707398
rect 293066 707162 293302 707398
rect 292746 690138 292982 690374
rect 293066 690138 293302 690374
rect 292746 689818 292982 690054
rect 293066 689818 293302 690054
rect 292746 654138 292982 654374
rect 293066 654138 293302 654374
rect 292746 653818 292982 654054
rect 293066 653818 293302 654054
rect 292746 618138 292982 618374
rect 293066 618138 293302 618374
rect 292746 617818 292982 618054
rect 293066 617818 293302 618054
rect 292746 582138 292982 582374
rect 293066 582138 293302 582374
rect 292746 581818 292982 582054
rect 293066 581818 293302 582054
rect 292746 546138 292982 546374
rect 293066 546138 293302 546374
rect 292746 545818 292982 546054
rect 293066 545818 293302 546054
rect 292746 510138 292982 510374
rect 293066 510138 293302 510374
rect 292746 509818 292982 510054
rect 293066 509818 293302 510054
rect 292746 474138 292982 474374
rect 293066 474138 293302 474374
rect 292746 473818 292982 474054
rect 293066 473818 293302 474054
rect 292746 438138 292982 438374
rect 293066 438138 293302 438374
rect 292746 437818 292982 438054
rect 293066 437818 293302 438054
rect 292746 402138 292982 402374
rect 293066 402138 293302 402374
rect 292746 401818 292982 402054
rect 293066 401818 293302 402054
rect 292746 366138 292982 366374
rect 293066 366138 293302 366374
rect 292746 365818 292982 366054
rect 293066 365818 293302 366054
rect 292746 330138 292982 330374
rect 293066 330138 293302 330374
rect 292746 329818 292982 330054
rect 293066 329818 293302 330054
rect 292746 294138 292982 294374
rect 293066 294138 293302 294374
rect 292746 293818 292982 294054
rect 293066 293818 293302 294054
rect 292746 258138 292982 258374
rect 293066 258138 293302 258374
rect 292746 257818 292982 258054
rect 293066 257818 293302 258054
rect 292746 222138 292982 222374
rect 293066 222138 293302 222374
rect 292746 221818 292982 222054
rect 293066 221818 293302 222054
rect 292746 186138 292982 186374
rect 293066 186138 293302 186374
rect 292746 185818 292982 186054
rect 293066 185818 293302 186054
rect 292746 150138 292982 150374
rect 293066 150138 293302 150374
rect 292746 149818 292982 150054
rect 293066 149818 293302 150054
rect 292746 114138 292982 114374
rect 293066 114138 293302 114374
rect 292746 113818 292982 114054
rect 293066 113818 293302 114054
rect 292746 78138 292982 78374
rect 293066 78138 293302 78374
rect 292746 77818 292982 78054
rect 293066 77818 293302 78054
rect 292746 42138 292982 42374
rect 293066 42138 293302 42374
rect 292746 41818 292982 42054
rect 293066 41818 293302 42054
rect 292746 6138 292982 6374
rect 293066 6138 293302 6374
rect 292746 5818 292982 6054
rect 293066 5818 293302 6054
rect 292746 -3462 292982 -3226
rect 293066 -3462 293302 -3226
rect 292746 -3782 292982 -3546
rect 293066 -3782 293302 -3546
rect 293986 708442 294222 708678
rect 294306 708442 294542 708678
rect 293986 708122 294222 708358
rect 294306 708122 294542 708358
rect 293986 691378 294222 691614
rect 294306 691378 294542 691614
rect 293986 691058 294222 691294
rect 294306 691058 294542 691294
rect 293986 655378 294222 655614
rect 294306 655378 294542 655614
rect 293986 655058 294222 655294
rect 294306 655058 294542 655294
rect 293986 619378 294222 619614
rect 294306 619378 294542 619614
rect 293986 619058 294222 619294
rect 294306 619058 294542 619294
rect 293986 583378 294222 583614
rect 294306 583378 294542 583614
rect 293986 583058 294222 583294
rect 294306 583058 294542 583294
rect 293986 547378 294222 547614
rect 294306 547378 294542 547614
rect 293986 547058 294222 547294
rect 294306 547058 294542 547294
rect 293986 511378 294222 511614
rect 294306 511378 294542 511614
rect 293986 511058 294222 511294
rect 294306 511058 294542 511294
rect 293986 475378 294222 475614
rect 294306 475378 294542 475614
rect 293986 475058 294222 475294
rect 294306 475058 294542 475294
rect 293986 439378 294222 439614
rect 294306 439378 294542 439614
rect 293986 439058 294222 439294
rect 294306 439058 294542 439294
rect 293986 403378 294222 403614
rect 294306 403378 294542 403614
rect 293986 403058 294222 403294
rect 294306 403058 294542 403294
rect 293986 367378 294222 367614
rect 294306 367378 294542 367614
rect 293986 367058 294222 367294
rect 294306 367058 294542 367294
rect 293986 331378 294222 331614
rect 294306 331378 294542 331614
rect 293986 331058 294222 331294
rect 294306 331058 294542 331294
rect 293986 295378 294222 295614
rect 294306 295378 294542 295614
rect 293986 295058 294222 295294
rect 294306 295058 294542 295294
rect 293986 259378 294222 259614
rect 294306 259378 294542 259614
rect 293986 259058 294222 259294
rect 294306 259058 294542 259294
rect 293986 223378 294222 223614
rect 294306 223378 294542 223614
rect 293986 223058 294222 223294
rect 294306 223058 294542 223294
rect 293986 187378 294222 187614
rect 294306 187378 294542 187614
rect 293986 187058 294222 187294
rect 294306 187058 294542 187294
rect 293986 151378 294222 151614
rect 294306 151378 294542 151614
rect 293986 151058 294222 151294
rect 294306 151058 294542 151294
rect 293986 115378 294222 115614
rect 294306 115378 294542 115614
rect 293986 115058 294222 115294
rect 294306 115058 294542 115294
rect 293986 79378 294222 79614
rect 294306 79378 294542 79614
rect 293986 79058 294222 79294
rect 294306 79058 294542 79294
rect 293986 43378 294222 43614
rect 294306 43378 294542 43614
rect 293986 43058 294222 43294
rect 294306 43058 294542 43294
rect 293986 7378 294222 7614
rect 294306 7378 294542 7614
rect 293986 7058 294222 7294
rect 294306 7058 294542 7294
rect 293986 -4422 294222 -4186
rect 294306 -4422 294542 -4186
rect 293986 -4742 294222 -4506
rect 294306 -4742 294542 -4506
rect 295226 709402 295462 709638
rect 295546 709402 295782 709638
rect 295226 709082 295462 709318
rect 295546 709082 295782 709318
rect 295226 692618 295462 692854
rect 295546 692618 295782 692854
rect 295226 692298 295462 692534
rect 295546 692298 295782 692534
rect 295226 656618 295462 656854
rect 295546 656618 295782 656854
rect 295226 656298 295462 656534
rect 295546 656298 295782 656534
rect 295226 620618 295462 620854
rect 295546 620618 295782 620854
rect 295226 620298 295462 620534
rect 295546 620298 295782 620534
rect 295226 584618 295462 584854
rect 295546 584618 295782 584854
rect 295226 584298 295462 584534
rect 295546 584298 295782 584534
rect 295226 548618 295462 548854
rect 295546 548618 295782 548854
rect 295226 548298 295462 548534
rect 295546 548298 295782 548534
rect 295226 512618 295462 512854
rect 295546 512618 295782 512854
rect 295226 512298 295462 512534
rect 295546 512298 295782 512534
rect 295226 476618 295462 476854
rect 295546 476618 295782 476854
rect 295226 476298 295462 476534
rect 295546 476298 295782 476534
rect 295226 440618 295462 440854
rect 295546 440618 295782 440854
rect 295226 440298 295462 440534
rect 295546 440298 295782 440534
rect 295226 404618 295462 404854
rect 295546 404618 295782 404854
rect 295226 404298 295462 404534
rect 295546 404298 295782 404534
rect 295226 368618 295462 368854
rect 295546 368618 295782 368854
rect 295226 368298 295462 368534
rect 295546 368298 295782 368534
rect 295226 332618 295462 332854
rect 295546 332618 295782 332854
rect 295226 332298 295462 332534
rect 295546 332298 295782 332534
rect 295226 296618 295462 296854
rect 295546 296618 295782 296854
rect 295226 296298 295462 296534
rect 295546 296298 295782 296534
rect 295226 260618 295462 260854
rect 295546 260618 295782 260854
rect 295226 260298 295462 260534
rect 295546 260298 295782 260534
rect 295226 224618 295462 224854
rect 295546 224618 295782 224854
rect 295226 224298 295462 224534
rect 295546 224298 295782 224534
rect 295226 188618 295462 188854
rect 295546 188618 295782 188854
rect 295226 188298 295462 188534
rect 295546 188298 295782 188534
rect 295226 152618 295462 152854
rect 295546 152618 295782 152854
rect 295226 152298 295462 152534
rect 295546 152298 295782 152534
rect 295226 116618 295462 116854
rect 295546 116618 295782 116854
rect 295226 116298 295462 116534
rect 295546 116298 295782 116534
rect 295226 80618 295462 80854
rect 295546 80618 295782 80854
rect 295226 80298 295462 80534
rect 295546 80298 295782 80534
rect 295226 44618 295462 44854
rect 295546 44618 295782 44854
rect 295226 44298 295462 44534
rect 295546 44298 295782 44534
rect 295226 8618 295462 8854
rect 295546 8618 295782 8854
rect 295226 8298 295462 8534
rect 295546 8298 295782 8534
rect 295226 -5382 295462 -5146
rect 295546 -5382 295782 -5146
rect 295226 -5702 295462 -5466
rect 295546 -5702 295782 -5466
rect 296466 710362 296702 710598
rect 296786 710362 297022 710598
rect 296466 710042 296702 710278
rect 296786 710042 297022 710278
rect 296466 693858 296702 694094
rect 296786 693858 297022 694094
rect 296466 693538 296702 693774
rect 296786 693538 297022 693774
rect 296466 657858 296702 658094
rect 296786 657858 297022 658094
rect 296466 657538 296702 657774
rect 296786 657538 297022 657774
rect 296466 621858 296702 622094
rect 296786 621858 297022 622094
rect 296466 621538 296702 621774
rect 296786 621538 297022 621774
rect 296466 585858 296702 586094
rect 296786 585858 297022 586094
rect 296466 585538 296702 585774
rect 296786 585538 297022 585774
rect 296466 549858 296702 550094
rect 296786 549858 297022 550094
rect 296466 549538 296702 549774
rect 296786 549538 297022 549774
rect 296466 513858 296702 514094
rect 296786 513858 297022 514094
rect 296466 513538 296702 513774
rect 296786 513538 297022 513774
rect 296466 477858 296702 478094
rect 296786 477858 297022 478094
rect 296466 477538 296702 477774
rect 296786 477538 297022 477774
rect 296466 441858 296702 442094
rect 296786 441858 297022 442094
rect 296466 441538 296702 441774
rect 296786 441538 297022 441774
rect 296466 405858 296702 406094
rect 296786 405858 297022 406094
rect 296466 405538 296702 405774
rect 296786 405538 297022 405774
rect 296466 369858 296702 370094
rect 296786 369858 297022 370094
rect 296466 369538 296702 369774
rect 296786 369538 297022 369774
rect 296466 333858 296702 334094
rect 296786 333858 297022 334094
rect 296466 333538 296702 333774
rect 296786 333538 297022 333774
rect 296466 297858 296702 298094
rect 296786 297858 297022 298094
rect 296466 297538 296702 297774
rect 296786 297538 297022 297774
rect 296466 261858 296702 262094
rect 296786 261858 297022 262094
rect 296466 261538 296702 261774
rect 296786 261538 297022 261774
rect 296466 225858 296702 226094
rect 296786 225858 297022 226094
rect 296466 225538 296702 225774
rect 296786 225538 297022 225774
rect 296466 189858 296702 190094
rect 296786 189858 297022 190094
rect 296466 189538 296702 189774
rect 296786 189538 297022 189774
rect 296466 153858 296702 154094
rect 296786 153858 297022 154094
rect 296466 153538 296702 153774
rect 296786 153538 297022 153774
rect 296466 117858 296702 118094
rect 296786 117858 297022 118094
rect 296466 117538 296702 117774
rect 296786 117538 297022 117774
rect 296466 81858 296702 82094
rect 296786 81858 297022 82094
rect 296466 81538 296702 81774
rect 296786 81538 297022 81774
rect 296466 45858 296702 46094
rect 296786 45858 297022 46094
rect 296466 45538 296702 45774
rect 296786 45538 297022 45774
rect 296466 9858 296702 10094
rect 296786 9858 297022 10094
rect 296466 9538 296702 9774
rect 296786 9538 297022 9774
rect 296466 -6342 296702 -6106
rect 296786 -6342 297022 -6106
rect 296466 -6662 296702 -6426
rect 296786 -6662 297022 -6426
rect 297706 711322 297942 711558
rect 298026 711322 298262 711558
rect 297706 711002 297942 711238
rect 298026 711002 298262 711238
rect 297706 695098 297942 695334
rect 298026 695098 298262 695334
rect 297706 694778 297942 695014
rect 298026 694778 298262 695014
rect 297706 659098 297942 659334
rect 298026 659098 298262 659334
rect 297706 658778 297942 659014
rect 298026 658778 298262 659014
rect 297706 623098 297942 623334
rect 298026 623098 298262 623334
rect 297706 622778 297942 623014
rect 298026 622778 298262 623014
rect 297706 587098 297942 587334
rect 298026 587098 298262 587334
rect 297706 586778 297942 587014
rect 298026 586778 298262 587014
rect 297706 551098 297942 551334
rect 298026 551098 298262 551334
rect 297706 550778 297942 551014
rect 298026 550778 298262 551014
rect 297706 515098 297942 515334
rect 298026 515098 298262 515334
rect 297706 514778 297942 515014
rect 298026 514778 298262 515014
rect 297706 479098 297942 479334
rect 298026 479098 298262 479334
rect 297706 478778 297942 479014
rect 298026 478778 298262 479014
rect 297706 443098 297942 443334
rect 298026 443098 298262 443334
rect 297706 442778 297942 443014
rect 298026 442778 298262 443014
rect 297706 407098 297942 407334
rect 298026 407098 298262 407334
rect 297706 406778 297942 407014
rect 298026 406778 298262 407014
rect 297706 371098 297942 371334
rect 298026 371098 298262 371334
rect 297706 370778 297942 371014
rect 298026 370778 298262 371014
rect 297706 335098 297942 335334
rect 298026 335098 298262 335334
rect 297706 334778 297942 335014
rect 298026 334778 298262 335014
rect 297706 299098 297942 299334
rect 298026 299098 298262 299334
rect 297706 298778 297942 299014
rect 298026 298778 298262 299014
rect 297706 263098 297942 263334
rect 298026 263098 298262 263334
rect 297706 262778 297942 263014
rect 298026 262778 298262 263014
rect 297706 227098 297942 227334
rect 298026 227098 298262 227334
rect 297706 226778 297942 227014
rect 298026 226778 298262 227014
rect 297706 191098 297942 191334
rect 298026 191098 298262 191334
rect 297706 190778 297942 191014
rect 298026 190778 298262 191014
rect 297706 155098 297942 155334
rect 298026 155098 298262 155334
rect 297706 154778 297942 155014
rect 298026 154778 298262 155014
rect 297706 119098 297942 119334
rect 298026 119098 298262 119334
rect 297706 118778 297942 119014
rect 298026 118778 298262 119014
rect 297706 83098 297942 83334
rect 298026 83098 298262 83334
rect 297706 82778 297942 83014
rect 298026 82778 298262 83014
rect 297706 47098 297942 47334
rect 298026 47098 298262 47334
rect 297706 46778 297942 47014
rect 298026 46778 298262 47014
rect 297706 11098 297942 11334
rect 298026 11098 298262 11334
rect 297706 10778 297942 11014
rect 298026 10778 298262 11014
rect 297706 -7302 297942 -7066
rect 298026 -7302 298262 -7066
rect 297706 -7622 297942 -7386
rect 298026 -7622 298262 -7386
rect 325026 704602 325262 704838
rect 325346 704602 325582 704838
rect 325026 704282 325262 704518
rect 325346 704282 325582 704518
rect 325026 686418 325262 686654
rect 325346 686418 325582 686654
rect 325026 686098 325262 686334
rect 325346 686098 325582 686334
rect 325026 650418 325262 650654
rect 325346 650418 325582 650654
rect 325026 650098 325262 650334
rect 325346 650098 325582 650334
rect 325026 614418 325262 614654
rect 325346 614418 325582 614654
rect 325026 614098 325262 614334
rect 325346 614098 325582 614334
rect 325026 578418 325262 578654
rect 325346 578418 325582 578654
rect 325026 578098 325262 578334
rect 325346 578098 325582 578334
rect 325026 542418 325262 542654
rect 325346 542418 325582 542654
rect 325026 542098 325262 542334
rect 325346 542098 325582 542334
rect 325026 506418 325262 506654
rect 325346 506418 325582 506654
rect 325026 506098 325262 506334
rect 325346 506098 325582 506334
rect 325026 470418 325262 470654
rect 325346 470418 325582 470654
rect 325026 470098 325262 470334
rect 325346 470098 325582 470334
rect 325026 434418 325262 434654
rect 325346 434418 325582 434654
rect 325026 434098 325262 434334
rect 325346 434098 325582 434334
rect 325026 398418 325262 398654
rect 325346 398418 325582 398654
rect 325026 398098 325262 398334
rect 325346 398098 325582 398334
rect 325026 362418 325262 362654
rect 325346 362418 325582 362654
rect 325026 362098 325262 362334
rect 325346 362098 325582 362334
rect 325026 326418 325262 326654
rect 325346 326418 325582 326654
rect 325026 326098 325262 326334
rect 325346 326098 325582 326334
rect 325026 290418 325262 290654
rect 325346 290418 325582 290654
rect 325026 290098 325262 290334
rect 325346 290098 325582 290334
rect 325026 254418 325262 254654
rect 325346 254418 325582 254654
rect 325026 254098 325262 254334
rect 325346 254098 325582 254334
rect 325026 218418 325262 218654
rect 325346 218418 325582 218654
rect 325026 218098 325262 218334
rect 325346 218098 325582 218334
rect 325026 182418 325262 182654
rect 325346 182418 325582 182654
rect 325026 182098 325262 182334
rect 325346 182098 325582 182334
rect 325026 146418 325262 146654
rect 325346 146418 325582 146654
rect 325026 146098 325262 146334
rect 325346 146098 325582 146334
rect 325026 110418 325262 110654
rect 325346 110418 325582 110654
rect 325026 110098 325262 110334
rect 325346 110098 325582 110334
rect 325026 74418 325262 74654
rect 325346 74418 325582 74654
rect 325026 74098 325262 74334
rect 325346 74098 325582 74334
rect 325026 38418 325262 38654
rect 325346 38418 325582 38654
rect 325026 38098 325262 38334
rect 325346 38098 325582 38334
rect 325026 2418 325262 2654
rect 325346 2418 325582 2654
rect 325026 2098 325262 2334
rect 325346 2098 325582 2334
rect 325026 -582 325262 -346
rect 325346 -582 325582 -346
rect 325026 -902 325262 -666
rect 325346 -902 325582 -666
rect 326266 705562 326502 705798
rect 326586 705562 326822 705798
rect 326266 705242 326502 705478
rect 326586 705242 326822 705478
rect 326266 687658 326502 687894
rect 326586 687658 326822 687894
rect 326266 687338 326502 687574
rect 326586 687338 326822 687574
rect 326266 651658 326502 651894
rect 326586 651658 326822 651894
rect 326266 651338 326502 651574
rect 326586 651338 326822 651574
rect 326266 615658 326502 615894
rect 326586 615658 326822 615894
rect 326266 615338 326502 615574
rect 326586 615338 326822 615574
rect 326266 579658 326502 579894
rect 326586 579658 326822 579894
rect 326266 579338 326502 579574
rect 326586 579338 326822 579574
rect 326266 543658 326502 543894
rect 326586 543658 326822 543894
rect 326266 543338 326502 543574
rect 326586 543338 326822 543574
rect 326266 507658 326502 507894
rect 326586 507658 326822 507894
rect 326266 507338 326502 507574
rect 326586 507338 326822 507574
rect 326266 471658 326502 471894
rect 326586 471658 326822 471894
rect 326266 471338 326502 471574
rect 326586 471338 326822 471574
rect 326266 435658 326502 435894
rect 326586 435658 326822 435894
rect 326266 435338 326502 435574
rect 326586 435338 326822 435574
rect 326266 399658 326502 399894
rect 326586 399658 326822 399894
rect 326266 399338 326502 399574
rect 326586 399338 326822 399574
rect 326266 363658 326502 363894
rect 326586 363658 326822 363894
rect 326266 363338 326502 363574
rect 326586 363338 326822 363574
rect 326266 327658 326502 327894
rect 326586 327658 326822 327894
rect 326266 327338 326502 327574
rect 326586 327338 326822 327574
rect 326266 291658 326502 291894
rect 326586 291658 326822 291894
rect 326266 291338 326502 291574
rect 326586 291338 326822 291574
rect 326266 255658 326502 255894
rect 326586 255658 326822 255894
rect 326266 255338 326502 255574
rect 326586 255338 326822 255574
rect 326266 219658 326502 219894
rect 326586 219658 326822 219894
rect 326266 219338 326502 219574
rect 326586 219338 326822 219574
rect 326266 183658 326502 183894
rect 326586 183658 326822 183894
rect 326266 183338 326502 183574
rect 326586 183338 326822 183574
rect 326266 147658 326502 147894
rect 326586 147658 326822 147894
rect 326266 147338 326502 147574
rect 326586 147338 326822 147574
rect 326266 111658 326502 111894
rect 326586 111658 326822 111894
rect 326266 111338 326502 111574
rect 326586 111338 326822 111574
rect 326266 75658 326502 75894
rect 326586 75658 326822 75894
rect 326266 75338 326502 75574
rect 326586 75338 326822 75574
rect 326266 39658 326502 39894
rect 326586 39658 326822 39894
rect 326266 39338 326502 39574
rect 326586 39338 326822 39574
rect 326266 3658 326502 3894
rect 326586 3658 326822 3894
rect 326266 3338 326502 3574
rect 326586 3338 326822 3574
rect 326266 -1542 326502 -1306
rect 326586 -1542 326822 -1306
rect 326266 -1862 326502 -1626
rect 326586 -1862 326822 -1626
rect 327506 706522 327742 706758
rect 327826 706522 328062 706758
rect 327506 706202 327742 706438
rect 327826 706202 328062 706438
rect 327506 688898 327742 689134
rect 327826 688898 328062 689134
rect 327506 688578 327742 688814
rect 327826 688578 328062 688814
rect 327506 652898 327742 653134
rect 327826 652898 328062 653134
rect 327506 652578 327742 652814
rect 327826 652578 328062 652814
rect 327506 616898 327742 617134
rect 327826 616898 328062 617134
rect 327506 616578 327742 616814
rect 327826 616578 328062 616814
rect 327506 580898 327742 581134
rect 327826 580898 328062 581134
rect 327506 580578 327742 580814
rect 327826 580578 328062 580814
rect 327506 544898 327742 545134
rect 327826 544898 328062 545134
rect 327506 544578 327742 544814
rect 327826 544578 328062 544814
rect 327506 508898 327742 509134
rect 327826 508898 328062 509134
rect 327506 508578 327742 508814
rect 327826 508578 328062 508814
rect 327506 472898 327742 473134
rect 327826 472898 328062 473134
rect 327506 472578 327742 472814
rect 327826 472578 328062 472814
rect 327506 436898 327742 437134
rect 327826 436898 328062 437134
rect 327506 436578 327742 436814
rect 327826 436578 328062 436814
rect 327506 400898 327742 401134
rect 327826 400898 328062 401134
rect 327506 400578 327742 400814
rect 327826 400578 328062 400814
rect 327506 364898 327742 365134
rect 327826 364898 328062 365134
rect 327506 364578 327742 364814
rect 327826 364578 328062 364814
rect 327506 328898 327742 329134
rect 327826 328898 328062 329134
rect 327506 328578 327742 328814
rect 327826 328578 328062 328814
rect 327506 292898 327742 293134
rect 327826 292898 328062 293134
rect 327506 292578 327742 292814
rect 327826 292578 328062 292814
rect 327506 256898 327742 257134
rect 327826 256898 328062 257134
rect 327506 256578 327742 256814
rect 327826 256578 328062 256814
rect 327506 220898 327742 221134
rect 327826 220898 328062 221134
rect 327506 220578 327742 220814
rect 327826 220578 328062 220814
rect 327506 184898 327742 185134
rect 327826 184898 328062 185134
rect 327506 184578 327742 184814
rect 327826 184578 328062 184814
rect 327506 148898 327742 149134
rect 327826 148898 328062 149134
rect 327506 148578 327742 148814
rect 327826 148578 328062 148814
rect 327506 112898 327742 113134
rect 327826 112898 328062 113134
rect 327506 112578 327742 112814
rect 327826 112578 328062 112814
rect 327506 76898 327742 77134
rect 327826 76898 328062 77134
rect 327506 76578 327742 76814
rect 327826 76578 328062 76814
rect 327506 40898 327742 41134
rect 327826 40898 328062 41134
rect 327506 40578 327742 40814
rect 327826 40578 328062 40814
rect 327506 4898 327742 5134
rect 327826 4898 328062 5134
rect 327506 4578 327742 4814
rect 327826 4578 328062 4814
rect 327506 -2502 327742 -2266
rect 327826 -2502 328062 -2266
rect 327506 -2822 327742 -2586
rect 327826 -2822 328062 -2586
rect 328746 707482 328982 707718
rect 329066 707482 329302 707718
rect 328746 707162 328982 707398
rect 329066 707162 329302 707398
rect 328746 690138 328982 690374
rect 329066 690138 329302 690374
rect 328746 689818 328982 690054
rect 329066 689818 329302 690054
rect 328746 654138 328982 654374
rect 329066 654138 329302 654374
rect 328746 653818 328982 654054
rect 329066 653818 329302 654054
rect 328746 618138 328982 618374
rect 329066 618138 329302 618374
rect 328746 617818 328982 618054
rect 329066 617818 329302 618054
rect 328746 582138 328982 582374
rect 329066 582138 329302 582374
rect 328746 581818 328982 582054
rect 329066 581818 329302 582054
rect 328746 546138 328982 546374
rect 329066 546138 329302 546374
rect 328746 545818 328982 546054
rect 329066 545818 329302 546054
rect 328746 510138 328982 510374
rect 329066 510138 329302 510374
rect 328746 509818 328982 510054
rect 329066 509818 329302 510054
rect 328746 474138 328982 474374
rect 329066 474138 329302 474374
rect 328746 473818 328982 474054
rect 329066 473818 329302 474054
rect 328746 438138 328982 438374
rect 329066 438138 329302 438374
rect 328746 437818 328982 438054
rect 329066 437818 329302 438054
rect 328746 402138 328982 402374
rect 329066 402138 329302 402374
rect 328746 401818 328982 402054
rect 329066 401818 329302 402054
rect 328746 366138 328982 366374
rect 329066 366138 329302 366374
rect 328746 365818 328982 366054
rect 329066 365818 329302 366054
rect 328746 330138 328982 330374
rect 329066 330138 329302 330374
rect 328746 329818 328982 330054
rect 329066 329818 329302 330054
rect 328746 294138 328982 294374
rect 329066 294138 329302 294374
rect 328746 293818 328982 294054
rect 329066 293818 329302 294054
rect 328746 258138 328982 258374
rect 329066 258138 329302 258374
rect 328746 257818 328982 258054
rect 329066 257818 329302 258054
rect 328746 222138 328982 222374
rect 329066 222138 329302 222374
rect 328746 221818 328982 222054
rect 329066 221818 329302 222054
rect 328746 186138 328982 186374
rect 329066 186138 329302 186374
rect 328746 185818 328982 186054
rect 329066 185818 329302 186054
rect 328746 150138 328982 150374
rect 329066 150138 329302 150374
rect 328746 149818 328982 150054
rect 329066 149818 329302 150054
rect 328746 114138 328982 114374
rect 329066 114138 329302 114374
rect 328746 113818 328982 114054
rect 329066 113818 329302 114054
rect 328746 78138 328982 78374
rect 329066 78138 329302 78374
rect 328746 77818 328982 78054
rect 329066 77818 329302 78054
rect 328746 42138 328982 42374
rect 329066 42138 329302 42374
rect 328746 41818 328982 42054
rect 329066 41818 329302 42054
rect 328746 6138 328982 6374
rect 329066 6138 329302 6374
rect 328746 5818 328982 6054
rect 329066 5818 329302 6054
rect 328746 -3462 328982 -3226
rect 329066 -3462 329302 -3226
rect 328746 -3782 328982 -3546
rect 329066 -3782 329302 -3546
rect 329986 708442 330222 708678
rect 330306 708442 330542 708678
rect 329986 708122 330222 708358
rect 330306 708122 330542 708358
rect 329986 691378 330222 691614
rect 330306 691378 330542 691614
rect 329986 691058 330222 691294
rect 330306 691058 330542 691294
rect 329986 655378 330222 655614
rect 330306 655378 330542 655614
rect 329986 655058 330222 655294
rect 330306 655058 330542 655294
rect 329986 619378 330222 619614
rect 330306 619378 330542 619614
rect 329986 619058 330222 619294
rect 330306 619058 330542 619294
rect 329986 583378 330222 583614
rect 330306 583378 330542 583614
rect 329986 583058 330222 583294
rect 330306 583058 330542 583294
rect 329986 547378 330222 547614
rect 330306 547378 330542 547614
rect 329986 547058 330222 547294
rect 330306 547058 330542 547294
rect 329986 511378 330222 511614
rect 330306 511378 330542 511614
rect 329986 511058 330222 511294
rect 330306 511058 330542 511294
rect 329986 475378 330222 475614
rect 330306 475378 330542 475614
rect 329986 475058 330222 475294
rect 330306 475058 330542 475294
rect 329986 439378 330222 439614
rect 330306 439378 330542 439614
rect 329986 439058 330222 439294
rect 330306 439058 330542 439294
rect 329986 403378 330222 403614
rect 330306 403378 330542 403614
rect 329986 403058 330222 403294
rect 330306 403058 330542 403294
rect 329986 367378 330222 367614
rect 330306 367378 330542 367614
rect 329986 367058 330222 367294
rect 330306 367058 330542 367294
rect 329986 331378 330222 331614
rect 330306 331378 330542 331614
rect 329986 331058 330222 331294
rect 330306 331058 330542 331294
rect 329986 295378 330222 295614
rect 330306 295378 330542 295614
rect 329986 295058 330222 295294
rect 330306 295058 330542 295294
rect 329986 259378 330222 259614
rect 330306 259378 330542 259614
rect 329986 259058 330222 259294
rect 330306 259058 330542 259294
rect 329986 223378 330222 223614
rect 330306 223378 330542 223614
rect 329986 223058 330222 223294
rect 330306 223058 330542 223294
rect 329986 187378 330222 187614
rect 330306 187378 330542 187614
rect 329986 187058 330222 187294
rect 330306 187058 330542 187294
rect 329986 151378 330222 151614
rect 330306 151378 330542 151614
rect 329986 151058 330222 151294
rect 330306 151058 330542 151294
rect 329986 115378 330222 115614
rect 330306 115378 330542 115614
rect 329986 115058 330222 115294
rect 330306 115058 330542 115294
rect 329986 79378 330222 79614
rect 330306 79378 330542 79614
rect 329986 79058 330222 79294
rect 330306 79058 330542 79294
rect 329986 43378 330222 43614
rect 330306 43378 330542 43614
rect 329986 43058 330222 43294
rect 330306 43058 330542 43294
rect 329986 7378 330222 7614
rect 330306 7378 330542 7614
rect 329986 7058 330222 7294
rect 330306 7058 330542 7294
rect 329986 -4422 330222 -4186
rect 330306 -4422 330542 -4186
rect 329986 -4742 330222 -4506
rect 330306 -4742 330542 -4506
rect 331226 709402 331462 709638
rect 331546 709402 331782 709638
rect 331226 709082 331462 709318
rect 331546 709082 331782 709318
rect 331226 692618 331462 692854
rect 331546 692618 331782 692854
rect 331226 692298 331462 692534
rect 331546 692298 331782 692534
rect 331226 656618 331462 656854
rect 331546 656618 331782 656854
rect 331226 656298 331462 656534
rect 331546 656298 331782 656534
rect 331226 620618 331462 620854
rect 331546 620618 331782 620854
rect 331226 620298 331462 620534
rect 331546 620298 331782 620534
rect 331226 584618 331462 584854
rect 331546 584618 331782 584854
rect 331226 584298 331462 584534
rect 331546 584298 331782 584534
rect 331226 548618 331462 548854
rect 331546 548618 331782 548854
rect 331226 548298 331462 548534
rect 331546 548298 331782 548534
rect 331226 512618 331462 512854
rect 331546 512618 331782 512854
rect 331226 512298 331462 512534
rect 331546 512298 331782 512534
rect 331226 476618 331462 476854
rect 331546 476618 331782 476854
rect 331226 476298 331462 476534
rect 331546 476298 331782 476534
rect 331226 440618 331462 440854
rect 331546 440618 331782 440854
rect 331226 440298 331462 440534
rect 331546 440298 331782 440534
rect 331226 404618 331462 404854
rect 331546 404618 331782 404854
rect 331226 404298 331462 404534
rect 331546 404298 331782 404534
rect 331226 368618 331462 368854
rect 331546 368618 331782 368854
rect 331226 368298 331462 368534
rect 331546 368298 331782 368534
rect 331226 332618 331462 332854
rect 331546 332618 331782 332854
rect 331226 332298 331462 332534
rect 331546 332298 331782 332534
rect 331226 296618 331462 296854
rect 331546 296618 331782 296854
rect 331226 296298 331462 296534
rect 331546 296298 331782 296534
rect 331226 260618 331462 260854
rect 331546 260618 331782 260854
rect 331226 260298 331462 260534
rect 331546 260298 331782 260534
rect 331226 224618 331462 224854
rect 331546 224618 331782 224854
rect 331226 224298 331462 224534
rect 331546 224298 331782 224534
rect 331226 188618 331462 188854
rect 331546 188618 331782 188854
rect 331226 188298 331462 188534
rect 331546 188298 331782 188534
rect 331226 152618 331462 152854
rect 331546 152618 331782 152854
rect 331226 152298 331462 152534
rect 331546 152298 331782 152534
rect 331226 116618 331462 116854
rect 331546 116618 331782 116854
rect 331226 116298 331462 116534
rect 331546 116298 331782 116534
rect 331226 80618 331462 80854
rect 331546 80618 331782 80854
rect 331226 80298 331462 80534
rect 331546 80298 331782 80534
rect 331226 44618 331462 44854
rect 331546 44618 331782 44854
rect 331226 44298 331462 44534
rect 331546 44298 331782 44534
rect 331226 8618 331462 8854
rect 331546 8618 331782 8854
rect 331226 8298 331462 8534
rect 331546 8298 331782 8534
rect 331226 -5382 331462 -5146
rect 331546 -5382 331782 -5146
rect 331226 -5702 331462 -5466
rect 331546 -5702 331782 -5466
rect 332466 710362 332702 710598
rect 332786 710362 333022 710598
rect 332466 710042 332702 710278
rect 332786 710042 333022 710278
rect 332466 693858 332702 694094
rect 332786 693858 333022 694094
rect 332466 693538 332702 693774
rect 332786 693538 333022 693774
rect 332466 657858 332702 658094
rect 332786 657858 333022 658094
rect 332466 657538 332702 657774
rect 332786 657538 333022 657774
rect 332466 621858 332702 622094
rect 332786 621858 333022 622094
rect 332466 621538 332702 621774
rect 332786 621538 333022 621774
rect 332466 585858 332702 586094
rect 332786 585858 333022 586094
rect 332466 585538 332702 585774
rect 332786 585538 333022 585774
rect 332466 549858 332702 550094
rect 332786 549858 333022 550094
rect 332466 549538 332702 549774
rect 332786 549538 333022 549774
rect 332466 513858 332702 514094
rect 332786 513858 333022 514094
rect 332466 513538 332702 513774
rect 332786 513538 333022 513774
rect 332466 477858 332702 478094
rect 332786 477858 333022 478094
rect 332466 477538 332702 477774
rect 332786 477538 333022 477774
rect 332466 441858 332702 442094
rect 332786 441858 333022 442094
rect 332466 441538 332702 441774
rect 332786 441538 333022 441774
rect 332466 405858 332702 406094
rect 332786 405858 333022 406094
rect 332466 405538 332702 405774
rect 332786 405538 333022 405774
rect 332466 369858 332702 370094
rect 332786 369858 333022 370094
rect 332466 369538 332702 369774
rect 332786 369538 333022 369774
rect 332466 333858 332702 334094
rect 332786 333858 333022 334094
rect 332466 333538 332702 333774
rect 332786 333538 333022 333774
rect 332466 297858 332702 298094
rect 332786 297858 333022 298094
rect 332466 297538 332702 297774
rect 332786 297538 333022 297774
rect 332466 261858 332702 262094
rect 332786 261858 333022 262094
rect 332466 261538 332702 261774
rect 332786 261538 333022 261774
rect 332466 225858 332702 226094
rect 332786 225858 333022 226094
rect 332466 225538 332702 225774
rect 332786 225538 333022 225774
rect 332466 189858 332702 190094
rect 332786 189858 333022 190094
rect 332466 189538 332702 189774
rect 332786 189538 333022 189774
rect 332466 153858 332702 154094
rect 332786 153858 333022 154094
rect 332466 153538 332702 153774
rect 332786 153538 333022 153774
rect 332466 117858 332702 118094
rect 332786 117858 333022 118094
rect 332466 117538 332702 117774
rect 332786 117538 333022 117774
rect 332466 81858 332702 82094
rect 332786 81858 333022 82094
rect 332466 81538 332702 81774
rect 332786 81538 333022 81774
rect 332466 45858 332702 46094
rect 332786 45858 333022 46094
rect 332466 45538 332702 45774
rect 332786 45538 333022 45774
rect 332466 9858 332702 10094
rect 332786 9858 333022 10094
rect 332466 9538 332702 9774
rect 332786 9538 333022 9774
rect 332466 -6342 332702 -6106
rect 332786 -6342 333022 -6106
rect 332466 -6662 332702 -6426
rect 332786 -6662 333022 -6426
rect 333706 711322 333942 711558
rect 334026 711322 334262 711558
rect 333706 711002 333942 711238
rect 334026 711002 334262 711238
rect 333706 695098 333942 695334
rect 334026 695098 334262 695334
rect 333706 694778 333942 695014
rect 334026 694778 334262 695014
rect 333706 659098 333942 659334
rect 334026 659098 334262 659334
rect 333706 658778 333942 659014
rect 334026 658778 334262 659014
rect 333706 623098 333942 623334
rect 334026 623098 334262 623334
rect 333706 622778 333942 623014
rect 334026 622778 334262 623014
rect 333706 587098 333942 587334
rect 334026 587098 334262 587334
rect 333706 586778 333942 587014
rect 334026 586778 334262 587014
rect 333706 551098 333942 551334
rect 334026 551098 334262 551334
rect 333706 550778 333942 551014
rect 334026 550778 334262 551014
rect 333706 515098 333942 515334
rect 334026 515098 334262 515334
rect 333706 514778 333942 515014
rect 334026 514778 334262 515014
rect 333706 479098 333942 479334
rect 334026 479098 334262 479334
rect 333706 478778 333942 479014
rect 334026 478778 334262 479014
rect 333706 443098 333942 443334
rect 334026 443098 334262 443334
rect 333706 442778 333942 443014
rect 334026 442778 334262 443014
rect 333706 407098 333942 407334
rect 334026 407098 334262 407334
rect 333706 406778 333942 407014
rect 334026 406778 334262 407014
rect 333706 371098 333942 371334
rect 334026 371098 334262 371334
rect 333706 370778 333942 371014
rect 334026 370778 334262 371014
rect 333706 335098 333942 335334
rect 334026 335098 334262 335334
rect 333706 334778 333942 335014
rect 334026 334778 334262 335014
rect 333706 299098 333942 299334
rect 334026 299098 334262 299334
rect 333706 298778 333942 299014
rect 334026 298778 334262 299014
rect 333706 263098 333942 263334
rect 334026 263098 334262 263334
rect 333706 262778 333942 263014
rect 334026 262778 334262 263014
rect 333706 227098 333942 227334
rect 334026 227098 334262 227334
rect 333706 226778 333942 227014
rect 334026 226778 334262 227014
rect 333706 191098 333942 191334
rect 334026 191098 334262 191334
rect 333706 190778 333942 191014
rect 334026 190778 334262 191014
rect 333706 155098 333942 155334
rect 334026 155098 334262 155334
rect 333706 154778 333942 155014
rect 334026 154778 334262 155014
rect 333706 119098 333942 119334
rect 334026 119098 334262 119334
rect 333706 118778 333942 119014
rect 334026 118778 334262 119014
rect 333706 83098 333942 83334
rect 334026 83098 334262 83334
rect 333706 82778 333942 83014
rect 334026 82778 334262 83014
rect 333706 47098 333942 47334
rect 334026 47098 334262 47334
rect 333706 46778 333942 47014
rect 334026 46778 334262 47014
rect 333706 11098 333942 11334
rect 334026 11098 334262 11334
rect 333706 10778 333942 11014
rect 334026 10778 334262 11014
rect 333706 -7302 333942 -7066
rect 334026 -7302 334262 -7066
rect 333706 -7622 333942 -7386
rect 334026 -7622 334262 -7386
rect 361026 704602 361262 704838
rect 361346 704602 361582 704838
rect 361026 704282 361262 704518
rect 361346 704282 361582 704518
rect 361026 686418 361262 686654
rect 361346 686418 361582 686654
rect 361026 686098 361262 686334
rect 361346 686098 361582 686334
rect 361026 650418 361262 650654
rect 361346 650418 361582 650654
rect 361026 650098 361262 650334
rect 361346 650098 361582 650334
rect 361026 614418 361262 614654
rect 361346 614418 361582 614654
rect 361026 614098 361262 614334
rect 361346 614098 361582 614334
rect 361026 578418 361262 578654
rect 361346 578418 361582 578654
rect 361026 578098 361262 578334
rect 361346 578098 361582 578334
rect 361026 542418 361262 542654
rect 361346 542418 361582 542654
rect 361026 542098 361262 542334
rect 361346 542098 361582 542334
rect 361026 506418 361262 506654
rect 361346 506418 361582 506654
rect 361026 506098 361262 506334
rect 361346 506098 361582 506334
rect 361026 470418 361262 470654
rect 361346 470418 361582 470654
rect 361026 470098 361262 470334
rect 361346 470098 361582 470334
rect 361026 434418 361262 434654
rect 361346 434418 361582 434654
rect 361026 434098 361262 434334
rect 361346 434098 361582 434334
rect 361026 398418 361262 398654
rect 361346 398418 361582 398654
rect 361026 398098 361262 398334
rect 361346 398098 361582 398334
rect 361026 362418 361262 362654
rect 361346 362418 361582 362654
rect 361026 362098 361262 362334
rect 361346 362098 361582 362334
rect 361026 326418 361262 326654
rect 361346 326418 361582 326654
rect 361026 326098 361262 326334
rect 361346 326098 361582 326334
rect 361026 290418 361262 290654
rect 361346 290418 361582 290654
rect 361026 290098 361262 290334
rect 361346 290098 361582 290334
rect 361026 254418 361262 254654
rect 361346 254418 361582 254654
rect 361026 254098 361262 254334
rect 361346 254098 361582 254334
rect 361026 218418 361262 218654
rect 361346 218418 361582 218654
rect 361026 218098 361262 218334
rect 361346 218098 361582 218334
rect 361026 182418 361262 182654
rect 361346 182418 361582 182654
rect 361026 182098 361262 182334
rect 361346 182098 361582 182334
rect 361026 146418 361262 146654
rect 361346 146418 361582 146654
rect 361026 146098 361262 146334
rect 361346 146098 361582 146334
rect 361026 110418 361262 110654
rect 361346 110418 361582 110654
rect 361026 110098 361262 110334
rect 361346 110098 361582 110334
rect 361026 74418 361262 74654
rect 361346 74418 361582 74654
rect 361026 74098 361262 74334
rect 361346 74098 361582 74334
rect 361026 38418 361262 38654
rect 361346 38418 361582 38654
rect 361026 38098 361262 38334
rect 361346 38098 361582 38334
rect 361026 2418 361262 2654
rect 361346 2418 361582 2654
rect 361026 2098 361262 2334
rect 361346 2098 361582 2334
rect 361026 -582 361262 -346
rect 361346 -582 361582 -346
rect 361026 -902 361262 -666
rect 361346 -902 361582 -666
rect 362266 705562 362502 705798
rect 362586 705562 362822 705798
rect 362266 705242 362502 705478
rect 362586 705242 362822 705478
rect 362266 687658 362502 687894
rect 362586 687658 362822 687894
rect 362266 687338 362502 687574
rect 362586 687338 362822 687574
rect 362266 651658 362502 651894
rect 362586 651658 362822 651894
rect 362266 651338 362502 651574
rect 362586 651338 362822 651574
rect 362266 615658 362502 615894
rect 362586 615658 362822 615894
rect 362266 615338 362502 615574
rect 362586 615338 362822 615574
rect 362266 579658 362502 579894
rect 362586 579658 362822 579894
rect 362266 579338 362502 579574
rect 362586 579338 362822 579574
rect 362266 543658 362502 543894
rect 362586 543658 362822 543894
rect 362266 543338 362502 543574
rect 362586 543338 362822 543574
rect 362266 507658 362502 507894
rect 362586 507658 362822 507894
rect 362266 507338 362502 507574
rect 362586 507338 362822 507574
rect 362266 471658 362502 471894
rect 362586 471658 362822 471894
rect 362266 471338 362502 471574
rect 362586 471338 362822 471574
rect 362266 435658 362502 435894
rect 362586 435658 362822 435894
rect 362266 435338 362502 435574
rect 362586 435338 362822 435574
rect 362266 399658 362502 399894
rect 362586 399658 362822 399894
rect 362266 399338 362502 399574
rect 362586 399338 362822 399574
rect 362266 363658 362502 363894
rect 362586 363658 362822 363894
rect 362266 363338 362502 363574
rect 362586 363338 362822 363574
rect 362266 327658 362502 327894
rect 362586 327658 362822 327894
rect 362266 327338 362502 327574
rect 362586 327338 362822 327574
rect 362266 291658 362502 291894
rect 362586 291658 362822 291894
rect 362266 291338 362502 291574
rect 362586 291338 362822 291574
rect 362266 255658 362502 255894
rect 362586 255658 362822 255894
rect 362266 255338 362502 255574
rect 362586 255338 362822 255574
rect 362266 219658 362502 219894
rect 362586 219658 362822 219894
rect 362266 219338 362502 219574
rect 362586 219338 362822 219574
rect 362266 183658 362502 183894
rect 362586 183658 362822 183894
rect 362266 183338 362502 183574
rect 362586 183338 362822 183574
rect 362266 147658 362502 147894
rect 362586 147658 362822 147894
rect 362266 147338 362502 147574
rect 362586 147338 362822 147574
rect 362266 111658 362502 111894
rect 362586 111658 362822 111894
rect 362266 111338 362502 111574
rect 362586 111338 362822 111574
rect 362266 75658 362502 75894
rect 362586 75658 362822 75894
rect 362266 75338 362502 75574
rect 362586 75338 362822 75574
rect 362266 39658 362502 39894
rect 362586 39658 362822 39894
rect 362266 39338 362502 39574
rect 362586 39338 362822 39574
rect 362266 3658 362502 3894
rect 362586 3658 362822 3894
rect 362266 3338 362502 3574
rect 362586 3338 362822 3574
rect 362266 -1542 362502 -1306
rect 362586 -1542 362822 -1306
rect 362266 -1862 362502 -1626
rect 362586 -1862 362822 -1626
rect 363506 706522 363742 706758
rect 363826 706522 364062 706758
rect 363506 706202 363742 706438
rect 363826 706202 364062 706438
rect 363506 688898 363742 689134
rect 363826 688898 364062 689134
rect 363506 688578 363742 688814
rect 363826 688578 364062 688814
rect 363506 652898 363742 653134
rect 363826 652898 364062 653134
rect 363506 652578 363742 652814
rect 363826 652578 364062 652814
rect 363506 616898 363742 617134
rect 363826 616898 364062 617134
rect 363506 616578 363742 616814
rect 363826 616578 364062 616814
rect 363506 580898 363742 581134
rect 363826 580898 364062 581134
rect 363506 580578 363742 580814
rect 363826 580578 364062 580814
rect 363506 544898 363742 545134
rect 363826 544898 364062 545134
rect 363506 544578 363742 544814
rect 363826 544578 364062 544814
rect 363506 508898 363742 509134
rect 363826 508898 364062 509134
rect 363506 508578 363742 508814
rect 363826 508578 364062 508814
rect 363506 472898 363742 473134
rect 363826 472898 364062 473134
rect 363506 472578 363742 472814
rect 363826 472578 364062 472814
rect 363506 436898 363742 437134
rect 363826 436898 364062 437134
rect 363506 436578 363742 436814
rect 363826 436578 364062 436814
rect 363506 400898 363742 401134
rect 363826 400898 364062 401134
rect 363506 400578 363742 400814
rect 363826 400578 364062 400814
rect 363506 364898 363742 365134
rect 363826 364898 364062 365134
rect 363506 364578 363742 364814
rect 363826 364578 364062 364814
rect 363506 328898 363742 329134
rect 363826 328898 364062 329134
rect 363506 328578 363742 328814
rect 363826 328578 364062 328814
rect 363506 292898 363742 293134
rect 363826 292898 364062 293134
rect 363506 292578 363742 292814
rect 363826 292578 364062 292814
rect 363506 256898 363742 257134
rect 363826 256898 364062 257134
rect 363506 256578 363742 256814
rect 363826 256578 364062 256814
rect 363506 220898 363742 221134
rect 363826 220898 364062 221134
rect 363506 220578 363742 220814
rect 363826 220578 364062 220814
rect 363506 184898 363742 185134
rect 363826 184898 364062 185134
rect 363506 184578 363742 184814
rect 363826 184578 364062 184814
rect 363506 148898 363742 149134
rect 363826 148898 364062 149134
rect 363506 148578 363742 148814
rect 363826 148578 364062 148814
rect 363506 112898 363742 113134
rect 363826 112898 364062 113134
rect 363506 112578 363742 112814
rect 363826 112578 364062 112814
rect 363506 76898 363742 77134
rect 363826 76898 364062 77134
rect 363506 76578 363742 76814
rect 363826 76578 364062 76814
rect 363506 40898 363742 41134
rect 363826 40898 364062 41134
rect 363506 40578 363742 40814
rect 363826 40578 364062 40814
rect 363506 4898 363742 5134
rect 363826 4898 364062 5134
rect 363506 4578 363742 4814
rect 363826 4578 364062 4814
rect 363506 -2502 363742 -2266
rect 363826 -2502 364062 -2266
rect 363506 -2822 363742 -2586
rect 363826 -2822 364062 -2586
rect 364746 707482 364982 707718
rect 365066 707482 365302 707718
rect 364746 707162 364982 707398
rect 365066 707162 365302 707398
rect 364746 690138 364982 690374
rect 365066 690138 365302 690374
rect 364746 689818 364982 690054
rect 365066 689818 365302 690054
rect 364746 654138 364982 654374
rect 365066 654138 365302 654374
rect 364746 653818 364982 654054
rect 365066 653818 365302 654054
rect 364746 618138 364982 618374
rect 365066 618138 365302 618374
rect 364746 617818 364982 618054
rect 365066 617818 365302 618054
rect 364746 582138 364982 582374
rect 365066 582138 365302 582374
rect 364746 581818 364982 582054
rect 365066 581818 365302 582054
rect 364746 546138 364982 546374
rect 365066 546138 365302 546374
rect 364746 545818 364982 546054
rect 365066 545818 365302 546054
rect 364746 510138 364982 510374
rect 365066 510138 365302 510374
rect 364746 509818 364982 510054
rect 365066 509818 365302 510054
rect 364746 474138 364982 474374
rect 365066 474138 365302 474374
rect 364746 473818 364982 474054
rect 365066 473818 365302 474054
rect 364746 438138 364982 438374
rect 365066 438138 365302 438374
rect 364746 437818 364982 438054
rect 365066 437818 365302 438054
rect 364746 402138 364982 402374
rect 365066 402138 365302 402374
rect 364746 401818 364982 402054
rect 365066 401818 365302 402054
rect 364746 366138 364982 366374
rect 365066 366138 365302 366374
rect 364746 365818 364982 366054
rect 365066 365818 365302 366054
rect 364746 330138 364982 330374
rect 365066 330138 365302 330374
rect 364746 329818 364982 330054
rect 365066 329818 365302 330054
rect 364746 294138 364982 294374
rect 365066 294138 365302 294374
rect 364746 293818 364982 294054
rect 365066 293818 365302 294054
rect 364746 258138 364982 258374
rect 365066 258138 365302 258374
rect 364746 257818 364982 258054
rect 365066 257818 365302 258054
rect 364746 222138 364982 222374
rect 365066 222138 365302 222374
rect 364746 221818 364982 222054
rect 365066 221818 365302 222054
rect 364746 186138 364982 186374
rect 365066 186138 365302 186374
rect 364746 185818 364982 186054
rect 365066 185818 365302 186054
rect 364746 150138 364982 150374
rect 365066 150138 365302 150374
rect 364746 149818 364982 150054
rect 365066 149818 365302 150054
rect 364746 114138 364982 114374
rect 365066 114138 365302 114374
rect 364746 113818 364982 114054
rect 365066 113818 365302 114054
rect 364746 78138 364982 78374
rect 365066 78138 365302 78374
rect 364746 77818 364982 78054
rect 365066 77818 365302 78054
rect 364746 42138 364982 42374
rect 365066 42138 365302 42374
rect 364746 41818 364982 42054
rect 365066 41818 365302 42054
rect 364746 6138 364982 6374
rect 365066 6138 365302 6374
rect 364746 5818 364982 6054
rect 365066 5818 365302 6054
rect 364746 -3462 364982 -3226
rect 365066 -3462 365302 -3226
rect 364746 -3782 364982 -3546
rect 365066 -3782 365302 -3546
rect 365986 708442 366222 708678
rect 366306 708442 366542 708678
rect 365986 708122 366222 708358
rect 366306 708122 366542 708358
rect 365986 691378 366222 691614
rect 366306 691378 366542 691614
rect 365986 691058 366222 691294
rect 366306 691058 366542 691294
rect 365986 655378 366222 655614
rect 366306 655378 366542 655614
rect 365986 655058 366222 655294
rect 366306 655058 366542 655294
rect 365986 619378 366222 619614
rect 366306 619378 366542 619614
rect 365986 619058 366222 619294
rect 366306 619058 366542 619294
rect 365986 583378 366222 583614
rect 366306 583378 366542 583614
rect 365986 583058 366222 583294
rect 366306 583058 366542 583294
rect 365986 547378 366222 547614
rect 366306 547378 366542 547614
rect 365986 547058 366222 547294
rect 366306 547058 366542 547294
rect 365986 511378 366222 511614
rect 366306 511378 366542 511614
rect 365986 511058 366222 511294
rect 366306 511058 366542 511294
rect 365986 475378 366222 475614
rect 366306 475378 366542 475614
rect 365986 475058 366222 475294
rect 366306 475058 366542 475294
rect 365986 439378 366222 439614
rect 366306 439378 366542 439614
rect 365986 439058 366222 439294
rect 366306 439058 366542 439294
rect 365986 403378 366222 403614
rect 366306 403378 366542 403614
rect 365986 403058 366222 403294
rect 366306 403058 366542 403294
rect 365986 367378 366222 367614
rect 366306 367378 366542 367614
rect 365986 367058 366222 367294
rect 366306 367058 366542 367294
rect 365986 331378 366222 331614
rect 366306 331378 366542 331614
rect 365986 331058 366222 331294
rect 366306 331058 366542 331294
rect 365986 295378 366222 295614
rect 366306 295378 366542 295614
rect 365986 295058 366222 295294
rect 366306 295058 366542 295294
rect 365986 259378 366222 259614
rect 366306 259378 366542 259614
rect 365986 259058 366222 259294
rect 366306 259058 366542 259294
rect 365986 223378 366222 223614
rect 366306 223378 366542 223614
rect 365986 223058 366222 223294
rect 366306 223058 366542 223294
rect 365986 187378 366222 187614
rect 366306 187378 366542 187614
rect 365986 187058 366222 187294
rect 366306 187058 366542 187294
rect 365986 151378 366222 151614
rect 366306 151378 366542 151614
rect 365986 151058 366222 151294
rect 366306 151058 366542 151294
rect 365986 115378 366222 115614
rect 366306 115378 366542 115614
rect 365986 115058 366222 115294
rect 366306 115058 366542 115294
rect 365986 79378 366222 79614
rect 366306 79378 366542 79614
rect 365986 79058 366222 79294
rect 366306 79058 366542 79294
rect 365986 43378 366222 43614
rect 366306 43378 366542 43614
rect 365986 43058 366222 43294
rect 366306 43058 366542 43294
rect 365986 7378 366222 7614
rect 366306 7378 366542 7614
rect 365986 7058 366222 7294
rect 366306 7058 366542 7294
rect 365986 -4422 366222 -4186
rect 366306 -4422 366542 -4186
rect 365986 -4742 366222 -4506
rect 366306 -4742 366542 -4506
rect 367226 709402 367462 709638
rect 367546 709402 367782 709638
rect 367226 709082 367462 709318
rect 367546 709082 367782 709318
rect 367226 692618 367462 692854
rect 367546 692618 367782 692854
rect 367226 692298 367462 692534
rect 367546 692298 367782 692534
rect 367226 656618 367462 656854
rect 367546 656618 367782 656854
rect 367226 656298 367462 656534
rect 367546 656298 367782 656534
rect 367226 620618 367462 620854
rect 367546 620618 367782 620854
rect 367226 620298 367462 620534
rect 367546 620298 367782 620534
rect 367226 584618 367462 584854
rect 367546 584618 367782 584854
rect 367226 584298 367462 584534
rect 367546 584298 367782 584534
rect 367226 548618 367462 548854
rect 367546 548618 367782 548854
rect 367226 548298 367462 548534
rect 367546 548298 367782 548534
rect 367226 512618 367462 512854
rect 367546 512618 367782 512854
rect 367226 512298 367462 512534
rect 367546 512298 367782 512534
rect 367226 476618 367462 476854
rect 367546 476618 367782 476854
rect 367226 476298 367462 476534
rect 367546 476298 367782 476534
rect 367226 440618 367462 440854
rect 367546 440618 367782 440854
rect 367226 440298 367462 440534
rect 367546 440298 367782 440534
rect 367226 404618 367462 404854
rect 367546 404618 367782 404854
rect 367226 404298 367462 404534
rect 367546 404298 367782 404534
rect 367226 368618 367462 368854
rect 367546 368618 367782 368854
rect 367226 368298 367462 368534
rect 367546 368298 367782 368534
rect 367226 332618 367462 332854
rect 367546 332618 367782 332854
rect 367226 332298 367462 332534
rect 367546 332298 367782 332534
rect 367226 296618 367462 296854
rect 367546 296618 367782 296854
rect 367226 296298 367462 296534
rect 367546 296298 367782 296534
rect 367226 260618 367462 260854
rect 367546 260618 367782 260854
rect 367226 260298 367462 260534
rect 367546 260298 367782 260534
rect 367226 224618 367462 224854
rect 367546 224618 367782 224854
rect 367226 224298 367462 224534
rect 367546 224298 367782 224534
rect 367226 188618 367462 188854
rect 367546 188618 367782 188854
rect 367226 188298 367462 188534
rect 367546 188298 367782 188534
rect 367226 152618 367462 152854
rect 367546 152618 367782 152854
rect 367226 152298 367462 152534
rect 367546 152298 367782 152534
rect 367226 116618 367462 116854
rect 367546 116618 367782 116854
rect 367226 116298 367462 116534
rect 367546 116298 367782 116534
rect 367226 80618 367462 80854
rect 367546 80618 367782 80854
rect 367226 80298 367462 80534
rect 367546 80298 367782 80534
rect 367226 44618 367462 44854
rect 367546 44618 367782 44854
rect 367226 44298 367462 44534
rect 367546 44298 367782 44534
rect 367226 8618 367462 8854
rect 367546 8618 367782 8854
rect 367226 8298 367462 8534
rect 367546 8298 367782 8534
rect 367226 -5382 367462 -5146
rect 367546 -5382 367782 -5146
rect 367226 -5702 367462 -5466
rect 367546 -5702 367782 -5466
rect 368466 710362 368702 710598
rect 368786 710362 369022 710598
rect 368466 710042 368702 710278
rect 368786 710042 369022 710278
rect 368466 693858 368702 694094
rect 368786 693858 369022 694094
rect 368466 693538 368702 693774
rect 368786 693538 369022 693774
rect 368466 657858 368702 658094
rect 368786 657858 369022 658094
rect 368466 657538 368702 657774
rect 368786 657538 369022 657774
rect 368466 621858 368702 622094
rect 368786 621858 369022 622094
rect 368466 621538 368702 621774
rect 368786 621538 369022 621774
rect 368466 585858 368702 586094
rect 368786 585858 369022 586094
rect 368466 585538 368702 585774
rect 368786 585538 369022 585774
rect 368466 549858 368702 550094
rect 368786 549858 369022 550094
rect 368466 549538 368702 549774
rect 368786 549538 369022 549774
rect 368466 513858 368702 514094
rect 368786 513858 369022 514094
rect 368466 513538 368702 513774
rect 368786 513538 369022 513774
rect 368466 477858 368702 478094
rect 368786 477858 369022 478094
rect 368466 477538 368702 477774
rect 368786 477538 369022 477774
rect 368466 441858 368702 442094
rect 368786 441858 369022 442094
rect 368466 441538 368702 441774
rect 368786 441538 369022 441774
rect 368466 405858 368702 406094
rect 368786 405858 369022 406094
rect 368466 405538 368702 405774
rect 368786 405538 369022 405774
rect 368466 369858 368702 370094
rect 368786 369858 369022 370094
rect 368466 369538 368702 369774
rect 368786 369538 369022 369774
rect 368466 333858 368702 334094
rect 368786 333858 369022 334094
rect 368466 333538 368702 333774
rect 368786 333538 369022 333774
rect 368466 297858 368702 298094
rect 368786 297858 369022 298094
rect 368466 297538 368702 297774
rect 368786 297538 369022 297774
rect 368466 261858 368702 262094
rect 368786 261858 369022 262094
rect 368466 261538 368702 261774
rect 368786 261538 369022 261774
rect 368466 225858 368702 226094
rect 368786 225858 369022 226094
rect 368466 225538 368702 225774
rect 368786 225538 369022 225774
rect 368466 189858 368702 190094
rect 368786 189858 369022 190094
rect 368466 189538 368702 189774
rect 368786 189538 369022 189774
rect 368466 153858 368702 154094
rect 368786 153858 369022 154094
rect 368466 153538 368702 153774
rect 368786 153538 369022 153774
rect 368466 117858 368702 118094
rect 368786 117858 369022 118094
rect 368466 117538 368702 117774
rect 368786 117538 369022 117774
rect 368466 81858 368702 82094
rect 368786 81858 369022 82094
rect 368466 81538 368702 81774
rect 368786 81538 369022 81774
rect 368466 45858 368702 46094
rect 368786 45858 369022 46094
rect 368466 45538 368702 45774
rect 368786 45538 369022 45774
rect 368466 9858 368702 10094
rect 368786 9858 369022 10094
rect 368466 9538 368702 9774
rect 368786 9538 369022 9774
rect 368466 -6342 368702 -6106
rect 368786 -6342 369022 -6106
rect 368466 -6662 368702 -6426
rect 368786 -6662 369022 -6426
rect 369706 711322 369942 711558
rect 370026 711322 370262 711558
rect 369706 711002 369942 711238
rect 370026 711002 370262 711238
rect 369706 695098 369942 695334
rect 370026 695098 370262 695334
rect 369706 694778 369942 695014
rect 370026 694778 370262 695014
rect 369706 659098 369942 659334
rect 370026 659098 370262 659334
rect 369706 658778 369942 659014
rect 370026 658778 370262 659014
rect 369706 623098 369942 623334
rect 370026 623098 370262 623334
rect 369706 622778 369942 623014
rect 370026 622778 370262 623014
rect 369706 587098 369942 587334
rect 370026 587098 370262 587334
rect 369706 586778 369942 587014
rect 370026 586778 370262 587014
rect 369706 551098 369942 551334
rect 370026 551098 370262 551334
rect 369706 550778 369942 551014
rect 370026 550778 370262 551014
rect 369706 515098 369942 515334
rect 370026 515098 370262 515334
rect 369706 514778 369942 515014
rect 370026 514778 370262 515014
rect 369706 479098 369942 479334
rect 370026 479098 370262 479334
rect 369706 478778 369942 479014
rect 370026 478778 370262 479014
rect 369706 443098 369942 443334
rect 370026 443098 370262 443334
rect 369706 442778 369942 443014
rect 370026 442778 370262 443014
rect 369706 407098 369942 407334
rect 370026 407098 370262 407334
rect 369706 406778 369942 407014
rect 370026 406778 370262 407014
rect 369706 371098 369942 371334
rect 370026 371098 370262 371334
rect 369706 370778 369942 371014
rect 370026 370778 370262 371014
rect 369706 335098 369942 335334
rect 370026 335098 370262 335334
rect 369706 334778 369942 335014
rect 370026 334778 370262 335014
rect 369706 299098 369942 299334
rect 370026 299098 370262 299334
rect 369706 298778 369942 299014
rect 370026 298778 370262 299014
rect 369706 263098 369942 263334
rect 370026 263098 370262 263334
rect 369706 262778 369942 263014
rect 370026 262778 370262 263014
rect 369706 227098 369942 227334
rect 370026 227098 370262 227334
rect 369706 226778 369942 227014
rect 370026 226778 370262 227014
rect 369706 191098 369942 191334
rect 370026 191098 370262 191334
rect 369706 190778 369942 191014
rect 370026 190778 370262 191014
rect 369706 155098 369942 155334
rect 370026 155098 370262 155334
rect 369706 154778 369942 155014
rect 370026 154778 370262 155014
rect 369706 119098 369942 119334
rect 370026 119098 370262 119334
rect 369706 118778 369942 119014
rect 370026 118778 370262 119014
rect 369706 83098 369942 83334
rect 370026 83098 370262 83334
rect 369706 82778 369942 83014
rect 370026 82778 370262 83014
rect 369706 47098 369942 47334
rect 370026 47098 370262 47334
rect 369706 46778 369942 47014
rect 370026 46778 370262 47014
rect 369706 11098 369942 11334
rect 370026 11098 370262 11334
rect 369706 10778 369942 11014
rect 370026 10778 370262 11014
rect 369706 -7302 369942 -7066
rect 370026 -7302 370262 -7066
rect 369706 -7622 369942 -7386
rect 370026 -7622 370262 -7386
rect 397026 704602 397262 704838
rect 397346 704602 397582 704838
rect 397026 704282 397262 704518
rect 397346 704282 397582 704518
rect 397026 686418 397262 686654
rect 397346 686418 397582 686654
rect 397026 686098 397262 686334
rect 397346 686098 397582 686334
rect 397026 650418 397262 650654
rect 397346 650418 397582 650654
rect 397026 650098 397262 650334
rect 397346 650098 397582 650334
rect 397026 614418 397262 614654
rect 397346 614418 397582 614654
rect 397026 614098 397262 614334
rect 397346 614098 397582 614334
rect 397026 578418 397262 578654
rect 397346 578418 397582 578654
rect 397026 578098 397262 578334
rect 397346 578098 397582 578334
rect 397026 542418 397262 542654
rect 397346 542418 397582 542654
rect 397026 542098 397262 542334
rect 397346 542098 397582 542334
rect 397026 506418 397262 506654
rect 397346 506418 397582 506654
rect 397026 506098 397262 506334
rect 397346 506098 397582 506334
rect 397026 470418 397262 470654
rect 397346 470418 397582 470654
rect 397026 470098 397262 470334
rect 397346 470098 397582 470334
rect 397026 434418 397262 434654
rect 397346 434418 397582 434654
rect 397026 434098 397262 434334
rect 397346 434098 397582 434334
rect 397026 398418 397262 398654
rect 397346 398418 397582 398654
rect 397026 398098 397262 398334
rect 397346 398098 397582 398334
rect 397026 362418 397262 362654
rect 397346 362418 397582 362654
rect 397026 362098 397262 362334
rect 397346 362098 397582 362334
rect 397026 326418 397262 326654
rect 397346 326418 397582 326654
rect 397026 326098 397262 326334
rect 397346 326098 397582 326334
rect 397026 290418 397262 290654
rect 397346 290418 397582 290654
rect 397026 290098 397262 290334
rect 397346 290098 397582 290334
rect 397026 254418 397262 254654
rect 397346 254418 397582 254654
rect 397026 254098 397262 254334
rect 397346 254098 397582 254334
rect 397026 218418 397262 218654
rect 397346 218418 397582 218654
rect 397026 218098 397262 218334
rect 397346 218098 397582 218334
rect 397026 182418 397262 182654
rect 397346 182418 397582 182654
rect 397026 182098 397262 182334
rect 397346 182098 397582 182334
rect 397026 146418 397262 146654
rect 397346 146418 397582 146654
rect 397026 146098 397262 146334
rect 397346 146098 397582 146334
rect 397026 110418 397262 110654
rect 397346 110418 397582 110654
rect 397026 110098 397262 110334
rect 397346 110098 397582 110334
rect 397026 74418 397262 74654
rect 397346 74418 397582 74654
rect 397026 74098 397262 74334
rect 397346 74098 397582 74334
rect 397026 38418 397262 38654
rect 397346 38418 397582 38654
rect 397026 38098 397262 38334
rect 397346 38098 397582 38334
rect 397026 2418 397262 2654
rect 397346 2418 397582 2654
rect 397026 2098 397262 2334
rect 397346 2098 397582 2334
rect 397026 -582 397262 -346
rect 397346 -582 397582 -346
rect 397026 -902 397262 -666
rect 397346 -902 397582 -666
rect 398266 705562 398502 705798
rect 398586 705562 398822 705798
rect 398266 705242 398502 705478
rect 398586 705242 398822 705478
rect 398266 687658 398502 687894
rect 398586 687658 398822 687894
rect 398266 687338 398502 687574
rect 398586 687338 398822 687574
rect 398266 651658 398502 651894
rect 398586 651658 398822 651894
rect 398266 651338 398502 651574
rect 398586 651338 398822 651574
rect 398266 615658 398502 615894
rect 398586 615658 398822 615894
rect 398266 615338 398502 615574
rect 398586 615338 398822 615574
rect 398266 579658 398502 579894
rect 398586 579658 398822 579894
rect 398266 579338 398502 579574
rect 398586 579338 398822 579574
rect 398266 543658 398502 543894
rect 398586 543658 398822 543894
rect 398266 543338 398502 543574
rect 398586 543338 398822 543574
rect 398266 507658 398502 507894
rect 398586 507658 398822 507894
rect 398266 507338 398502 507574
rect 398586 507338 398822 507574
rect 398266 471658 398502 471894
rect 398586 471658 398822 471894
rect 398266 471338 398502 471574
rect 398586 471338 398822 471574
rect 398266 435658 398502 435894
rect 398586 435658 398822 435894
rect 398266 435338 398502 435574
rect 398586 435338 398822 435574
rect 398266 399658 398502 399894
rect 398586 399658 398822 399894
rect 398266 399338 398502 399574
rect 398586 399338 398822 399574
rect 398266 363658 398502 363894
rect 398586 363658 398822 363894
rect 398266 363338 398502 363574
rect 398586 363338 398822 363574
rect 398266 327658 398502 327894
rect 398586 327658 398822 327894
rect 398266 327338 398502 327574
rect 398586 327338 398822 327574
rect 398266 291658 398502 291894
rect 398586 291658 398822 291894
rect 398266 291338 398502 291574
rect 398586 291338 398822 291574
rect 398266 255658 398502 255894
rect 398586 255658 398822 255894
rect 398266 255338 398502 255574
rect 398586 255338 398822 255574
rect 398266 219658 398502 219894
rect 398586 219658 398822 219894
rect 398266 219338 398502 219574
rect 398586 219338 398822 219574
rect 398266 183658 398502 183894
rect 398586 183658 398822 183894
rect 398266 183338 398502 183574
rect 398586 183338 398822 183574
rect 398266 147658 398502 147894
rect 398586 147658 398822 147894
rect 398266 147338 398502 147574
rect 398586 147338 398822 147574
rect 398266 111658 398502 111894
rect 398586 111658 398822 111894
rect 398266 111338 398502 111574
rect 398586 111338 398822 111574
rect 398266 75658 398502 75894
rect 398586 75658 398822 75894
rect 398266 75338 398502 75574
rect 398586 75338 398822 75574
rect 398266 39658 398502 39894
rect 398586 39658 398822 39894
rect 398266 39338 398502 39574
rect 398586 39338 398822 39574
rect 398266 3658 398502 3894
rect 398586 3658 398822 3894
rect 398266 3338 398502 3574
rect 398586 3338 398822 3574
rect 398266 -1542 398502 -1306
rect 398586 -1542 398822 -1306
rect 398266 -1862 398502 -1626
rect 398586 -1862 398822 -1626
rect 399506 706522 399742 706758
rect 399826 706522 400062 706758
rect 399506 706202 399742 706438
rect 399826 706202 400062 706438
rect 399506 688898 399742 689134
rect 399826 688898 400062 689134
rect 399506 688578 399742 688814
rect 399826 688578 400062 688814
rect 399506 652898 399742 653134
rect 399826 652898 400062 653134
rect 399506 652578 399742 652814
rect 399826 652578 400062 652814
rect 399506 616898 399742 617134
rect 399826 616898 400062 617134
rect 399506 616578 399742 616814
rect 399826 616578 400062 616814
rect 399506 580898 399742 581134
rect 399826 580898 400062 581134
rect 399506 580578 399742 580814
rect 399826 580578 400062 580814
rect 399506 544898 399742 545134
rect 399826 544898 400062 545134
rect 399506 544578 399742 544814
rect 399826 544578 400062 544814
rect 399506 508898 399742 509134
rect 399826 508898 400062 509134
rect 399506 508578 399742 508814
rect 399826 508578 400062 508814
rect 399506 472898 399742 473134
rect 399826 472898 400062 473134
rect 399506 472578 399742 472814
rect 399826 472578 400062 472814
rect 399506 436898 399742 437134
rect 399826 436898 400062 437134
rect 399506 436578 399742 436814
rect 399826 436578 400062 436814
rect 399506 400898 399742 401134
rect 399826 400898 400062 401134
rect 399506 400578 399742 400814
rect 399826 400578 400062 400814
rect 399506 364898 399742 365134
rect 399826 364898 400062 365134
rect 399506 364578 399742 364814
rect 399826 364578 400062 364814
rect 399506 328898 399742 329134
rect 399826 328898 400062 329134
rect 399506 328578 399742 328814
rect 399826 328578 400062 328814
rect 399506 292898 399742 293134
rect 399826 292898 400062 293134
rect 399506 292578 399742 292814
rect 399826 292578 400062 292814
rect 399506 256898 399742 257134
rect 399826 256898 400062 257134
rect 399506 256578 399742 256814
rect 399826 256578 400062 256814
rect 399506 220898 399742 221134
rect 399826 220898 400062 221134
rect 399506 220578 399742 220814
rect 399826 220578 400062 220814
rect 399506 184898 399742 185134
rect 399826 184898 400062 185134
rect 399506 184578 399742 184814
rect 399826 184578 400062 184814
rect 399506 148898 399742 149134
rect 399826 148898 400062 149134
rect 399506 148578 399742 148814
rect 399826 148578 400062 148814
rect 399506 112898 399742 113134
rect 399826 112898 400062 113134
rect 399506 112578 399742 112814
rect 399826 112578 400062 112814
rect 399506 76898 399742 77134
rect 399826 76898 400062 77134
rect 399506 76578 399742 76814
rect 399826 76578 400062 76814
rect 399506 40898 399742 41134
rect 399826 40898 400062 41134
rect 399506 40578 399742 40814
rect 399826 40578 400062 40814
rect 399506 4898 399742 5134
rect 399826 4898 400062 5134
rect 399506 4578 399742 4814
rect 399826 4578 400062 4814
rect 399506 -2502 399742 -2266
rect 399826 -2502 400062 -2266
rect 399506 -2822 399742 -2586
rect 399826 -2822 400062 -2586
rect 400746 707482 400982 707718
rect 401066 707482 401302 707718
rect 400746 707162 400982 707398
rect 401066 707162 401302 707398
rect 400746 690138 400982 690374
rect 401066 690138 401302 690374
rect 400746 689818 400982 690054
rect 401066 689818 401302 690054
rect 400746 654138 400982 654374
rect 401066 654138 401302 654374
rect 400746 653818 400982 654054
rect 401066 653818 401302 654054
rect 400746 618138 400982 618374
rect 401066 618138 401302 618374
rect 400746 617818 400982 618054
rect 401066 617818 401302 618054
rect 400746 582138 400982 582374
rect 401066 582138 401302 582374
rect 400746 581818 400982 582054
rect 401066 581818 401302 582054
rect 400746 546138 400982 546374
rect 401066 546138 401302 546374
rect 400746 545818 400982 546054
rect 401066 545818 401302 546054
rect 400746 510138 400982 510374
rect 401066 510138 401302 510374
rect 400746 509818 400982 510054
rect 401066 509818 401302 510054
rect 400746 474138 400982 474374
rect 401066 474138 401302 474374
rect 400746 473818 400982 474054
rect 401066 473818 401302 474054
rect 400746 438138 400982 438374
rect 401066 438138 401302 438374
rect 400746 437818 400982 438054
rect 401066 437818 401302 438054
rect 400746 402138 400982 402374
rect 401066 402138 401302 402374
rect 400746 401818 400982 402054
rect 401066 401818 401302 402054
rect 400746 366138 400982 366374
rect 401066 366138 401302 366374
rect 400746 365818 400982 366054
rect 401066 365818 401302 366054
rect 400746 330138 400982 330374
rect 401066 330138 401302 330374
rect 400746 329818 400982 330054
rect 401066 329818 401302 330054
rect 400746 294138 400982 294374
rect 401066 294138 401302 294374
rect 400746 293818 400982 294054
rect 401066 293818 401302 294054
rect 400746 258138 400982 258374
rect 401066 258138 401302 258374
rect 400746 257818 400982 258054
rect 401066 257818 401302 258054
rect 400746 222138 400982 222374
rect 401066 222138 401302 222374
rect 400746 221818 400982 222054
rect 401066 221818 401302 222054
rect 400746 186138 400982 186374
rect 401066 186138 401302 186374
rect 400746 185818 400982 186054
rect 401066 185818 401302 186054
rect 400746 150138 400982 150374
rect 401066 150138 401302 150374
rect 400746 149818 400982 150054
rect 401066 149818 401302 150054
rect 400746 114138 400982 114374
rect 401066 114138 401302 114374
rect 400746 113818 400982 114054
rect 401066 113818 401302 114054
rect 400746 78138 400982 78374
rect 401066 78138 401302 78374
rect 400746 77818 400982 78054
rect 401066 77818 401302 78054
rect 400746 42138 400982 42374
rect 401066 42138 401302 42374
rect 400746 41818 400982 42054
rect 401066 41818 401302 42054
rect 400746 6138 400982 6374
rect 401066 6138 401302 6374
rect 400746 5818 400982 6054
rect 401066 5818 401302 6054
rect 400746 -3462 400982 -3226
rect 401066 -3462 401302 -3226
rect 400746 -3782 400982 -3546
rect 401066 -3782 401302 -3546
rect 401986 708442 402222 708678
rect 402306 708442 402542 708678
rect 401986 708122 402222 708358
rect 402306 708122 402542 708358
rect 401986 691378 402222 691614
rect 402306 691378 402542 691614
rect 401986 691058 402222 691294
rect 402306 691058 402542 691294
rect 401986 655378 402222 655614
rect 402306 655378 402542 655614
rect 401986 655058 402222 655294
rect 402306 655058 402542 655294
rect 401986 619378 402222 619614
rect 402306 619378 402542 619614
rect 401986 619058 402222 619294
rect 402306 619058 402542 619294
rect 401986 583378 402222 583614
rect 402306 583378 402542 583614
rect 401986 583058 402222 583294
rect 402306 583058 402542 583294
rect 401986 547378 402222 547614
rect 402306 547378 402542 547614
rect 401986 547058 402222 547294
rect 402306 547058 402542 547294
rect 401986 511378 402222 511614
rect 402306 511378 402542 511614
rect 401986 511058 402222 511294
rect 402306 511058 402542 511294
rect 401986 475378 402222 475614
rect 402306 475378 402542 475614
rect 401986 475058 402222 475294
rect 402306 475058 402542 475294
rect 401986 439378 402222 439614
rect 402306 439378 402542 439614
rect 401986 439058 402222 439294
rect 402306 439058 402542 439294
rect 401986 403378 402222 403614
rect 402306 403378 402542 403614
rect 401986 403058 402222 403294
rect 402306 403058 402542 403294
rect 401986 367378 402222 367614
rect 402306 367378 402542 367614
rect 401986 367058 402222 367294
rect 402306 367058 402542 367294
rect 401986 331378 402222 331614
rect 402306 331378 402542 331614
rect 401986 331058 402222 331294
rect 402306 331058 402542 331294
rect 401986 295378 402222 295614
rect 402306 295378 402542 295614
rect 401986 295058 402222 295294
rect 402306 295058 402542 295294
rect 401986 259378 402222 259614
rect 402306 259378 402542 259614
rect 401986 259058 402222 259294
rect 402306 259058 402542 259294
rect 401986 223378 402222 223614
rect 402306 223378 402542 223614
rect 401986 223058 402222 223294
rect 402306 223058 402542 223294
rect 401986 187378 402222 187614
rect 402306 187378 402542 187614
rect 401986 187058 402222 187294
rect 402306 187058 402542 187294
rect 401986 151378 402222 151614
rect 402306 151378 402542 151614
rect 401986 151058 402222 151294
rect 402306 151058 402542 151294
rect 401986 115378 402222 115614
rect 402306 115378 402542 115614
rect 401986 115058 402222 115294
rect 402306 115058 402542 115294
rect 401986 79378 402222 79614
rect 402306 79378 402542 79614
rect 401986 79058 402222 79294
rect 402306 79058 402542 79294
rect 401986 43378 402222 43614
rect 402306 43378 402542 43614
rect 401986 43058 402222 43294
rect 402306 43058 402542 43294
rect 401986 7378 402222 7614
rect 402306 7378 402542 7614
rect 401986 7058 402222 7294
rect 402306 7058 402542 7294
rect 401986 -4422 402222 -4186
rect 402306 -4422 402542 -4186
rect 401986 -4742 402222 -4506
rect 402306 -4742 402542 -4506
rect 403226 709402 403462 709638
rect 403546 709402 403782 709638
rect 403226 709082 403462 709318
rect 403546 709082 403782 709318
rect 403226 692618 403462 692854
rect 403546 692618 403782 692854
rect 403226 692298 403462 692534
rect 403546 692298 403782 692534
rect 403226 656618 403462 656854
rect 403546 656618 403782 656854
rect 403226 656298 403462 656534
rect 403546 656298 403782 656534
rect 403226 620618 403462 620854
rect 403546 620618 403782 620854
rect 403226 620298 403462 620534
rect 403546 620298 403782 620534
rect 403226 584618 403462 584854
rect 403546 584618 403782 584854
rect 403226 584298 403462 584534
rect 403546 584298 403782 584534
rect 403226 548618 403462 548854
rect 403546 548618 403782 548854
rect 403226 548298 403462 548534
rect 403546 548298 403782 548534
rect 403226 512618 403462 512854
rect 403546 512618 403782 512854
rect 403226 512298 403462 512534
rect 403546 512298 403782 512534
rect 403226 476618 403462 476854
rect 403546 476618 403782 476854
rect 403226 476298 403462 476534
rect 403546 476298 403782 476534
rect 403226 440618 403462 440854
rect 403546 440618 403782 440854
rect 403226 440298 403462 440534
rect 403546 440298 403782 440534
rect 403226 404618 403462 404854
rect 403546 404618 403782 404854
rect 403226 404298 403462 404534
rect 403546 404298 403782 404534
rect 403226 368618 403462 368854
rect 403546 368618 403782 368854
rect 403226 368298 403462 368534
rect 403546 368298 403782 368534
rect 403226 332618 403462 332854
rect 403546 332618 403782 332854
rect 403226 332298 403462 332534
rect 403546 332298 403782 332534
rect 403226 296618 403462 296854
rect 403546 296618 403782 296854
rect 403226 296298 403462 296534
rect 403546 296298 403782 296534
rect 403226 260618 403462 260854
rect 403546 260618 403782 260854
rect 403226 260298 403462 260534
rect 403546 260298 403782 260534
rect 403226 224618 403462 224854
rect 403546 224618 403782 224854
rect 403226 224298 403462 224534
rect 403546 224298 403782 224534
rect 403226 188618 403462 188854
rect 403546 188618 403782 188854
rect 403226 188298 403462 188534
rect 403546 188298 403782 188534
rect 403226 152618 403462 152854
rect 403546 152618 403782 152854
rect 403226 152298 403462 152534
rect 403546 152298 403782 152534
rect 403226 116618 403462 116854
rect 403546 116618 403782 116854
rect 403226 116298 403462 116534
rect 403546 116298 403782 116534
rect 403226 80618 403462 80854
rect 403546 80618 403782 80854
rect 403226 80298 403462 80534
rect 403546 80298 403782 80534
rect 403226 44618 403462 44854
rect 403546 44618 403782 44854
rect 403226 44298 403462 44534
rect 403546 44298 403782 44534
rect 403226 8618 403462 8854
rect 403546 8618 403782 8854
rect 403226 8298 403462 8534
rect 403546 8298 403782 8534
rect 403226 -5382 403462 -5146
rect 403546 -5382 403782 -5146
rect 403226 -5702 403462 -5466
rect 403546 -5702 403782 -5466
rect 404466 710362 404702 710598
rect 404786 710362 405022 710598
rect 404466 710042 404702 710278
rect 404786 710042 405022 710278
rect 404466 693858 404702 694094
rect 404786 693858 405022 694094
rect 404466 693538 404702 693774
rect 404786 693538 405022 693774
rect 404466 657858 404702 658094
rect 404786 657858 405022 658094
rect 404466 657538 404702 657774
rect 404786 657538 405022 657774
rect 404466 621858 404702 622094
rect 404786 621858 405022 622094
rect 404466 621538 404702 621774
rect 404786 621538 405022 621774
rect 404466 585858 404702 586094
rect 404786 585858 405022 586094
rect 404466 585538 404702 585774
rect 404786 585538 405022 585774
rect 404466 549858 404702 550094
rect 404786 549858 405022 550094
rect 404466 549538 404702 549774
rect 404786 549538 405022 549774
rect 404466 513858 404702 514094
rect 404786 513858 405022 514094
rect 404466 513538 404702 513774
rect 404786 513538 405022 513774
rect 404466 477858 404702 478094
rect 404786 477858 405022 478094
rect 404466 477538 404702 477774
rect 404786 477538 405022 477774
rect 404466 441858 404702 442094
rect 404786 441858 405022 442094
rect 404466 441538 404702 441774
rect 404786 441538 405022 441774
rect 404466 405858 404702 406094
rect 404786 405858 405022 406094
rect 404466 405538 404702 405774
rect 404786 405538 405022 405774
rect 404466 369858 404702 370094
rect 404786 369858 405022 370094
rect 404466 369538 404702 369774
rect 404786 369538 405022 369774
rect 404466 333858 404702 334094
rect 404786 333858 405022 334094
rect 404466 333538 404702 333774
rect 404786 333538 405022 333774
rect 404466 297858 404702 298094
rect 404786 297858 405022 298094
rect 404466 297538 404702 297774
rect 404786 297538 405022 297774
rect 404466 261858 404702 262094
rect 404786 261858 405022 262094
rect 404466 261538 404702 261774
rect 404786 261538 405022 261774
rect 404466 225858 404702 226094
rect 404786 225858 405022 226094
rect 404466 225538 404702 225774
rect 404786 225538 405022 225774
rect 404466 189858 404702 190094
rect 404786 189858 405022 190094
rect 404466 189538 404702 189774
rect 404786 189538 405022 189774
rect 404466 153858 404702 154094
rect 404786 153858 405022 154094
rect 404466 153538 404702 153774
rect 404786 153538 405022 153774
rect 404466 117858 404702 118094
rect 404786 117858 405022 118094
rect 404466 117538 404702 117774
rect 404786 117538 405022 117774
rect 404466 81858 404702 82094
rect 404786 81858 405022 82094
rect 404466 81538 404702 81774
rect 404786 81538 405022 81774
rect 404466 45858 404702 46094
rect 404786 45858 405022 46094
rect 404466 45538 404702 45774
rect 404786 45538 405022 45774
rect 404466 9858 404702 10094
rect 404786 9858 405022 10094
rect 404466 9538 404702 9774
rect 404786 9538 405022 9774
rect 404466 -6342 404702 -6106
rect 404786 -6342 405022 -6106
rect 404466 -6662 404702 -6426
rect 404786 -6662 405022 -6426
rect 405706 711322 405942 711558
rect 406026 711322 406262 711558
rect 405706 711002 405942 711238
rect 406026 711002 406262 711238
rect 405706 695098 405942 695334
rect 406026 695098 406262 695334
rect 405706 694778 405942 695014
rect 406026 694778 406262 695014
rect 405706 659098 405942 659334
rect 406026 659098 406262 659334
rect 405706 658778 405942 659014
rect 406026 658778 406262 659014
rect 405706 623098 405942 623334
rect 406026 623098 406262 623334
rect 405706 622778 405942 623014
rect 406026 622778 406262 623014
rect 405706 587098 405942 587334
rect 406026 587098 406262 587334
rect 405706 586778 405942 587014
rect 406026 586778 406262 587014
rect 405706 551098 405942 551334
rect 406026 551098 406262 551334
rect 405706 550778 405942 551014
rect 406026 550778 406262 551014
rect 405706 515098 405942 515334
rect 406026 515098 406262 515334
rect 405706 514778 405942 515014
rect 406026 514778 406262 515014
rect 405706 479098 405942 479334
rect 406026 479098 406262 479334
rect 405706 478778 405942 479014
rect 406026 478778 406262 479014
rect 405706 443098 405942 443334
rect 406026 443098 406262 443334
rect 405706 442778 405942 443014
rect 406026 442778 406262 443014
rect 405706 407098 405942 407334
rect 406026 407098 406262 407334
rect 405706 406778 405942 407014
rect 406026 406778 406262 407014
rect 405706 371098 405942 371334
rect 406026 371098 406262 371334
rect 405706 370778 405942 371014
rect 406026 370778 406262 371014
rect 405706 335098 405942 335334
rect 406026 335098 406262 335334
rect 405706 334778 405942 335014
rect 406026 334778 406262 335014
rect 405706 299098 405942 299334
rect 406026 299098 406262 299334
rect 405706 298778 405942 299014
rect 406026 298778 406262 299014
rect 405706 263098 405942 263334
rect 406026 263098 406262 263334
rect 405706 262778 405942 263014
rect 406026 262778 406262 263014
rect 405706 227098 405942 227334
rect 406026 227098 406262 227334
rect 405706 226778 405942 227014
rect 406026 226778 406262 227014
rect 405706 191098 405942 191334
rect 406026 191098 406262 191334
rect 405706 190778 405942 191014
rect 406026 190778 406262 191014
rect 405706 155098 405942 155334
rect 406026 155098 406262 155334
rect 405706 154778 405942 155014
rect 406026 154778 406262 155014
rect 405706 119098 405942 119334
rect 406026 119098 406262 119334
rect 405706 118778 405942 119014
rect 406026 118778 406262 119014
rect 405706 83098 405942 83334
rect 406026 83098 406262 83334
rect 405706 82778 405942 83014
rect 406026 82778 406262 83014
rect 405706 47098 405942 47334
rect 406026 47098 406262 47334
rect 405706 46778 405942 47014
rect 406026 46778 406262 47014
rect 405706 11098 405942 11334
rect 406026 11098 406262 11334
rect 405706 10778 405942 11014
rect 406026 10778 406262 11014
rect 405706 -7302 405942 -7066
rect 406026 -7302 406262 -7066
rect 405706 -7622 405942 -7386
rect 406026 -7622 406262 -7386
rect 433026 704602 433262 704838
rect 433346 704602 433582 704838
rect 433026 704282 433262 704518
rect 433346 704282 433582 704518
rect 433026 686418 433262 686654
rect 433346 686418 433582 686654
rect 433026 686098 433262 686334
rect 433346 686098 433582 686334
rect 433026 650418 433262 650654
rect 433346 650418 433582 650654
rect 433026 650098 433262 650334
rect 433346 650098 433582 650334
rect 433026 614418 433262 614654
rect 433346 614418 433582 614654
rect 433026 614098 433262 614334
rect 433346 614098 433582 614334
rect 433026 578418 433262 578654
rect 433346 578418 433582 578654
rect 433026 578098 433262 578334
rect 433346 578098 433582 578334
rect 433026 542418 433262 542654
rect 433346 542418 433582 542654
rect 433026 542098 433262 542334
rect 433346 542098 433582 542334
rect 433026 506418 433262 506654
rect 433346 506418 433582 506654
rect 433026 506098 433262 506334
rect 433346 506098 433582 506334
rect 433026 470418 433262 470654
rect 433346 470418 433582 470654
rect 433026 470098 433262 470334
rect 433346 470098 433582 470334
rect 433026 434418 433262 434654
rect 433346 434418 433582 434654
rect 433026 434098 433262 434334
rect 433346 434098 433582 434334
rect 433026 398418 433262 398654
rect 433346 398418 433582 398654
rect 433026 398098 433262 398334
rect 433346 398098 433582 398334
rect 433026 362418 433262 362654
rect 433346 362418 433582 362654
rect 433026 362098 433262 362334
rect 433346 362098 433582 362334
rect 433026 326418 433262 326654
rect 433346 326418 433582 326654
rect 433026 326098 433262 326334
rect 433346 326098 433582 326334
rect 433026 290418 433262 290654
rect 433346 290418 433582 290654
rect 433026 290098 433262 290334
rect 433346 290098 433582 290334
rect 433026 254418 433262 254654
rect 433346 254418 433582 254654
rect 433026 254098 433262 254334
rect 433346 254098 433582 254334
rect 433026 218418 433262 218654
rect 433346 218418 433582 218654
rect 433026 218098 433262 218334
rect 433346 218098 433582 218334
rect 433026 182418 433262 182654
rect 433346 182418 433582 182654
rect 433026 182098 433262 182334
rect 433346 182098 433582 182334
rect 433026 146418 433262 146654
rect 433346 146418 433582 146654
rect 433026 146098 433262 146334
rect 433346 146098 433582 146334
rect 433026 110418 433262 110654
rect 433346 110418 433582 110654
rect 433026 110098 433262 110334
rect 433346 110098 433582 110334
rect 433026 74418 433262 74654
rect 433346 74418 433582 74654
rect 433026 74098 433262 74334
rect 433346 74098 433582 74334
rect 433026 38418 433262 38654
rect 433346 38418 433582 38654
rect 433026 38098 433262 38334
rect 433346 38098 433582 38334
rect 433026 2418 433262 2654
rect 433346 2418 433582 2654
rect 433026 2098 433262 2334
rect 433346 2098 433582 2334
rect 433026 -582 433262 -346
rect 433346 -582 433582 -346
rect 433026 -902 433262 -666
rect 433346 -902 433582 -666
rect 434266 705562 434502 705798
rect 434586 705562 434822 705798
rect 434266 705242 434502 705478
rect 434586 705242 434822 705478
rect 434266 687658 434502 687894
rect 434586 687658 434822 687894
rect 434266 687338 434502 687574
rect 434586 687338 434822 687574
rect 434266 651658 434502 651894
rect 434586 651658 434822 651894
rect 434266 651338 434502 651574
rect 434586 651338 434822 651574
rect 434266 615658 434502 615894
rect 434586 615658 434822 615894
rect 434266 615338 434502 615574
rect 434586 615338 434822 615574
rect 434266 579658 434502 579894
rect 434586 579658 434822 579894
rect 434266 579338 434502 579574
rect 434586 579338 434822 579574
rect 434266 543658 434502 543894
rect 434586 543658 434822 543894
rect 434266 543338 434502 543574
rect 434586 543338 434822 543574
rect 434266 507658 434502 507894
rect 434586 507658 434822 507894
rect 434266 507338 434502 507574
rect 434586 507338 434822 507574
rect 434266 471658 434502 471894
rect 434586 471658 434822 471894
rect 434266 471338 434502 471574
rect 434586 471338 434822 471574
rect 434266 435658 434502 435894
rect 434586 435658 434822 435894
rect 434266 435338 434502 435574
rect 434586 435338 434822 435574
rect 434266 399658 434502 399894
rect 434586 399658 434822 399894
rect 434266 399338 434502 399574
rect 434586 399338 434822 399574
rect 434266 363658 434502 363894
rect 434586 363658 434822 363894
rect 434266 363338 434502 363574
rect 434586 363338 434822 363574
rect 434266 327658 434502 327894
rect 434586 327658 434822 327894
rect 434266 327338 434502 327574
rect 434586 327338 434822 327574
rect 434266 291658 434502 291894
rect 434586 291658 434822 291894
rect 434266 291338 434502 291574
rect 434586 291338 434822 291574
rect 434266 255658 434502 255894
rect 434586 255658 434822 255894
rect 434266 255338 434502 255574
rect 434586 255338 434822 255574
rect 434266 219658 434502 219894
rect 434586 219658 434822 219894
rect 434266 219338 434502 219574
rect 434586 219338 434822 219574
rect 434266 183658 434502 183894
rect 434586 183658 434822 183894
rect 434266 183338 434502 183574
rect 434586 183338 434822 183574
rect 434266 147658 434502 147894
rect 434586 147658 434822 147894
rect 434266 147338 434502 147574
rect 434586 147338 434822 147574
rect 434266 111658 434502 111894
rect 434586 111658 434822 111894
rect 434266 111338 434502 111574
rect 434586 111338 434822 111574
rect 434266 75658 434502 75894
rect 434586 75658 434822 75894
rect 434266 75338 434502 75574
rect 434586 75338 434822 75574
rect 434266 39658 434502 39894
rect 434586 39658 434822 39894
rect 434266 39338 434502 39574
rect 434586 39338 434822 39574
rect 434266 3658 434502 3894
rect 434586 3658 434822 3894
rect 434266 3338 434502 3574
rect 434586 3338 434822 3574
rect 434266 -1542 434502 -1306
rect 434586 -1542 434822 -1306
rect 434266 -1862 434502 -1626
rect 434586 -1862 434822 -1626
rect 435506 706522 435742 706758
rect 435826 706522 436062 706758
rect 435506 706202 435742 706438
rect 435826 706202 436062 706438
rect 435506 688898 435742 689134
rect 435826 688898 436062 689134
rect 435506 688578 435742 688814
rect 435826 688578 436062 688814
rect 435506 652898 435742 653134
rect 435826 652898 436062 653134
rect 435506 652578 435742 652814
rect 435826 652578 436062 652814
rect 435506 616898 435742 617134
rect 435826 616898 436062 617134
rect 435506 616578 435742 616814
rect 435826 616578 436062 616814
rect 435506 580898 435742 581134
rect 435826 580898 436062 581134
rect 435506 580578 435742 580814
rect 435826 580578 436062 580814
rect 435506 544898 435742 545134
rect 435826 544898 436062 545134
rect 435506 544578 435742 544814
rect 435826 544578 436062 544814
rect 435506 508898 435742 509134
rect 435826 508898 436062 509134
rect 435506 508578 435742 508814
rect 435826 508578 436062 508814
rect 435506 472898 435742 473134
rect 435826 472898 436062 473134
rect 435506 472578 435742 472814
rect 435826 472578 436062 472814
rect 435506 436898 435742 437134
rect 435826 436898 436062 437134
rect 435506 436578 435742 436814
rect 435826 436578 436062 436814
rect 435506 400898 435742 401134
rect 435826 400898 436062 401134
rect 435506 400578 435742 400814
rect 435826 400578 436062 400814
rect 435506 364898 435742 365134
rect 435826 364898 436062 365134
rect 435506 364578 435742 364814
rect 435826 364578 436062 364814
rect 435506 328898 435742 329134
rect 435826 328898 436062 329134
rect 435506 328578 435742 328814
rect 435826 328578 436062 328814
rect 435506 292898 435742 293134
rect 435826 292898 436062 293134
rect 435506 292578 435742 292814
rect 435826 292578 436062 292814
rect 435506 256898 435742 257134
rect 435826 256898 436062 257134
rect 435506 256578 435742 256814
rect 435826 256578 436062 256814
rect 435506 220898 435742 221134
rect 435826 220898 436062 221134
rect 435506 220578 435742 220814
rect 435826 220578 436062 220814
rect 435506 184898 435742 185134
rect 435826 184898 436062 185134
rect 435506 184578 435742 184814
rect 435826 184578 436062 184814
rect 435506 148898 435742 149134
rect 435826 148898 436062 149134
rect 435506 148578 435742 148814
rect 435826 148578 436062 148814
rect 435506 112898 435742 113134
rect 435826 112898 436062 113134
rect 435506 112578 435742 112814
rect 435826 112578 436062 112814
rect 435506 76898 435742 77134
rect 435826 76898 436062 77134
rect 435506 76578 435742 76814
rect 435826 76578 436062 76814
rect 435506 40898 435742 41134
rect 435826 40898 436062 41134
rect 435506 40578 435742 40814
rect 435826 40578 436062 40814
rect 435506 4898 435742 5134
rect 435826 4898 436062 5134
rect 435506 4578 435742 4814
rect 435826 4578 436062 4814
rect 435506 -2502 435742 -2266
rect 435826 -2502 436062 -2266
rect 435506 -2822 435742 -2586
rect 435826 -2822 436062 -2586
rect 436746 707482 436982 707718
rect 437066 707482 437302 707718
rect 436746 707162 436982 707398
rect 437066 707162 437302 707398
rect 436746 690138 436982 690374
rect 437066 690138 437302 690374
rect 436746 689818 436982 690054
rect 437066 689818 437302 690054
rect 436746 654138 436982 654374
rect 437066 654138 437302 654374
rect 436746 653818 436982 654054
rect 437066 653818 437302 654054
rect 436746 618138 436982 618374
rect 437066 618138 437302 618374
rect 436746 617818 436982 618054
rect 437066 617818 437302 618054
rect 436746 582138 436982 582374
rect 437066 582138 437302 582374
rect 436746 581818 436982 582054
rect 437066 581818 437302 582054
rect 436746 546138 436982 546374
rect 437066 546138 437302 546374
rect 436746 545818 436982 546054
rect 437066 545818 437302 546054
rect 436746 510138 436982 510374
rect 437066 510138 437302 510374
rect 436746 509818 436982 510054
rect 437066 509818 437302 510054
rect 436746 474138 436982 474374
rect 437066 474138 437302 474374
rect 436746 473818 436982 474054
rect 437066 473818 437302 474054
rect 436746 438138 436982 438374
rect 437066 438138 437302 438374
rect 436746 437818 436982 438054
rect 437066 437818 437302 438054
rect 436746 402138 436982 402374
rect 437066 402138 437302 402374
rect 436746 401818 436982 402054
rect 437066 401818 437302 402054
rect 436746 366138 436982 366374
rect 437066 366138 437302 366374
rect 436746 365818 436982 366054
rect 437066 365818 437302 366054
rect 436746 330138 436982 330374
rect 437066 330138 437302 330374
rect 436746 329818 436982 330054
rect 437066 329818 437302 330054
rect 436746 294138 436982 294374
rect 437066 294138 437302 294374
rect 436746 293818 436982 294054
rect 437066 293818 437302 294054
rect 436746 258138 436982 258374
rect 437066 258138 437302 258374
rect 436746 257818 436982 258054
rect 437066 257818 437302 258054
rect 436746 222138 436982 222374
rect 437066 222138 437302 222374
rect 436746 221818 436982 222054
rect 437066 221818 437302 222054
rect 436746 186138 436982 186374
rect 437066 186138 437302 186374
rect 436746 185818 436982 186054
rect 437066 185818 437302 186054
rect 436746 150138 436982 150374
rect 437066 150138 437302 150374
rect 436746 149818 436982 150054
rect 437066 149818 437302 150054
rect 436746 114138 436982 114374
rect 437066 114138 437302 114374
rect 436746 113818 436982 114054
rect 437066 113818 437302 114054
rect 436746 78138 436982 78374
rect 437066 78138 437302 78374
rect 436746 77818 436982 78054
rect 437066 77818 437302 78054
rect 436746 42138 436982 42374
rect 437066 42138 437302 42374
rect 436746 41818 436982 42054
rect 437066 41818 437302 42054
rect 436746 6138 436982 6374
rect 437066 6138 437302 6374
rect 436746 5818 436982 6054
rect 437066 5818 437302 6054
rect 436746 -3462 436982 -3226
rect 437066 -3462 437302 -3226
rect 436746 -3782 436982 -3546
rect 437066 -3782 437302 -3546
rect 437986 708442 438222 708678
rect 438306 708442 438542 708678
rect 437986 708122 438222 708358
rect 438306 708122 438542 708358
rect 437986 691378 438222 691614
rect 438306 691378 438542 691614
rect 437986 691058 438222 691294
rect 438306 691058 438542 691294
rect 437986 655378 438222 655614
rect 438306 655378 438542 655614
rect 437986 655058 438222 655294
rect 438306 655058 438542 655294
rect 437986 619378 438222 619614
rect 438306 619378 438542 619614
rect 437986 619058 438222 619294
rect 438306 619058 438542 619294
rect 437986 583378 438222 583614
rect 438306 583378 438542 583614
rect 437986 583058 438222 583294
rect 438306 583058 438542 583294
rect 437986 547378 438222 547614
rect 438306 547378 438542 547614
rect 437986 547058 438222 547294
rect 438306 547058 438542 547294
rect 437986 511378 438222 511614
rect 438306 511378 438542 511614
rect 437986 511058 438222 511294
rect 438306 511058 438542 511294
rect 437986 475378 438222 475614
rect 438306 475378 438542 475614
rect 437986 475058 438222 475294
rect 438306 475058 438542 475294
rect 437986 439378 438222 439614
rect 438306 439378 438542 439614
rect 437986 439058 438222 439294
rect 438306 439058 438542 439294
rect 437986 403378 438222 403614
rect 438306 403378 438542 403614
rect 437986 403058 438222 403294
rect 438306 403058 438542 403294
rect 437986 367378 438222 367614
rect 438306 367378 438542 367614
rect 437986 367058 438222 367294
rect 438306 367058 438542 367294
rect 437986 331378 438222 331614
rect 438306 331378 438542 331614
rect 437986 331058 438222 331294
rect 438306 331058 438542 331294
rect 437986 295378 438222 295614
rect 438306 295378 438542 295614
rect 437986 295058 438222 295294
rect 438306 295058 438542 295294
rect 437986 259378 438222 259614
rect 438306 259378 438542 259614
rect 437986 259058 438222 259294
rect 438306 259058 438542 259294
rect 437986 223378 438222 223614
rect 438306 223378 438542 223614
rect 437986 223058 438222 223294
rect 438306 223058 438542 223294
rect 437986 187378 438222 187614
rect 438306 187378 438542 187614
rect 437986 187058 438222 187294
rect 438306 187058 438542 187294
rect 437986 151378 438222 151614
rect 438306 151378 438542 151614
rect 437986 151058 438222 151294
rect 438306 151058 438542 151294
rect 437986 115378 438222 115614
rect 438306 115378 438542 115614
rect 437986 115058 438222 115294
rect 438306 115058 438542 115294
rect 437986 79378 438222 79614
rect 438306 79378 438542 79614
rect 437986 79058 438222 79294
rect 438306 79058 438542 79294
rect 437986 43378 438222 43614
rect 438306 43378 438542 43614
rect 437986 43058 438222 43294
rect 438306 43058 438542 43294
rect 437986 7378 438222 7614
rect 438306 7378 438542 7614
rect 437986 7058 438222 7294
rect 438306 7058 438542 7294
rect 437986 -4422 438222 -4186
rect 438306 -4422 438542 -4186
rect 437986 -4742 438222 -4506
rect 438306 -4742 438542 -4506
rect 439226 709402 439462 709638
rect 439546 709402 439782 709638
rect 439226 709082 439462 709318
rect 439546 709082 439782 709318
rect 439226 692618 439462 692854
rect 439546 692618 439782 692854
rect 439226 692298 439462 692534
rect 439546 692298 439782 692534
rect 439226 656618 439462 656854
rect 439546 656618 439782 656854
rect 439226 656298 439462 656534
rect 439546 656298 439782 656534
rect 439226 620618 439462 620854
rect 439546 620618 439782 620854
rect 439226 620298 439462 620534
rect 439546 620298 439782 620534
rect 439226 584618 439462 584854
rect 439546 584618 439782 584854
rect 439226 584298 439462 584534
rect 439546 584298 439782 584534
rect 439226 548618 439462 548854
rect 439546 548618 439782 548854
rect 439226 548298 439462 548534
rect 439546 548298 439782 548534
rect 439226 512618 439462 512854
rect 439546 512618 439782 512854
rect 439226 512298 439462 512534
rect 439546 512298 439782 512534
rect 439226 476618 439462 476854
rect 439546 476618 439782 476854
rect 439226 476298 439462 476534
rect 439546 476298 439782 476534
rect 439226 440618 439462 440854
rect 439546 440618 439782 440854
rect 439226 440298 439462 440534
rect 439546 440298 439782 440534
rect 439226 404618 439462 404854
rect 439546 404618 439782 404854
rect 439226 404298 439462 404534
rect 439546 404298 439782 404534
rect 439226 368618 439462 368854
rect 439546 368618 439782 368854
rect 439226 368298 439462 368534
rect 439546 368298 439782 368534
rect 439226 332618 439462 332854
rect 439546 332618 439782 332854
rect 439226 332298 439462 332534
rect 439546 332298 439782 332534
rect 439226 296618 439462 296854
rect 439546 296618 439782 296854
rect 439226 296298 439462 296534
rect 439546 296298 439782 296534
rect 439226 260618 439462 260854
rect 439546 260618 439782 260854
rect 439226 260298 439462 260534
rect 439546 260298 439782 260534
rect 439226 224618 439462 224854
rect 439546 224618 439782 224854
rect 439226 224298 439462 224534
rect 439546 224298 439782 224534
rect 439226 188618 439462 188854
rect 439546 188618 439782 188854
rect 439226 188298 439462 188534
rect 439546 188298 439782 188534
rect 439226 152618 439462 152854
rect 439546 152618 439782 152854
rect 439226 152298 439462 152534
rect 439546 152298 439782 152534
rect 439226 116618 439462 116854
rect 439546 116618 439782 116854
rect 439226 116298 439462 116534
rect 439546 116298 439782 116534
rect 439226 80618 439462 80854
rect 439546 80618 439782 80854
rect 439226 80298 439462 80534
rect 439546 80298 439782 80534
rect 439226 44618 439462 44854
rect 439546 44618 439782 44854
rect 439226 44298 439462 44534
rect 439546 44298 439782 44534
rect 439226 8618 439462 8854
rect 439546 8618 439782 8854
rect 439226 8298 439462 8534
rect 439546 8298 439782 8534
rect 439226 -5382 439462 -5146
rect 439546 -5382 439782 -5146
rect 439226 -5702 439462 -5466
rect 439546 -5702 439782 -5466
rect 440466 710362 440702 710598
rect 440786 710362 441022 710598
rect 440466 710042 440702 710278
rect 440786 710042 441022 710278
rect 440466 693858 440702 694094
rect 440786 693858 441022 694094
rect 440466 693538 440702 693774
rect 440786 693538 441022 693774
rect 440466 657858 440702 658094
rect 440786 657858 441022 658094
rect 440466 657538 440702 657774
rect 440786 657538 441022 657774
rect 440466 621858 440702 622094
rect 440786 621858 441022 622094
rect 440466 621538 440702 621774
rect 440786 621538 441022 621774
rect 440466 585858 440702 586094
rect 440786 585858 441022 586094
rect 440466 585538 440702 585774
rect 440786 585538 441022 585774
rect 440466 549858 440702 550094
rect 440786 549858 441022 550094
rect 440466 549538 440702 549774
rect 440786 549538 441022 549774
rect 440466 513858 440702 514094
rect 440786 513858 441022 514094
rect 440466 513538 440702 513774
rect 440786 513538 441022 513774
rect 440466 477858 440702 478094
rect 440786 477858 441022 478094
rect 440466 477538 440702 477774
rect 440786 477538 441022 477774
rect 440466 441858 440702 442094
rect 440786 441858 441022 442094
rect 440466 441538 440702 441774
rect 440786 441538 441022 441774
rect 440466 405858 440702 406094
rect 440786 405858 441022 406094
rect 440466 405538 440702 405774
rect 440786 405538 441022 405774
rect 440466 369858 440702 370094
rect 440786 369858 441022 370094
rect 440466 369538 440702 369774
rect 440786 369538 441022 369774
rect 440466 333858 440702 334094
rect 440786 333858 441022 334094
rect 440466 333538 440702 333774
rect 440786 333538 441022 333774
rect 440466 297858 440702 298094
rect 440786 297858 441022 298094
rect 440466 297538 440702 297774
rect 440786 297538 441022 297774
rect 440466 261858 440702 262094
rect 440786 261858 441022 262094
rect 440466 261538 440702 261774
rect 440786 261538 441022 261774
rect 440466 225858 440702 226094
rect 440786 225858 441022 226094
rect 440466 225538 440702 225774
rect 440786 225538 441022 225774
rect 440466 189858 440702 190094
rect 440786 189858 441022 190094
rect 440466 189538 440702 189774
rect 440786 189538 441022 189774
rect 440466 153858 440702 154094
rect 440786 153858 441022 154094
rect 440466 153538 440702 153774
rect 440786 153538 441022 153774
rect 440466 117858 440702 118094
rect 440786 117858 441022 118094
rect 440466 117538 440702 117774
rect 440786 117538 441022 117774
rect 440466 81858 440702 82094
rect 440786 81858 441022 82094
rect 440466 81538 440702 81774
rect 440786 81538 441022 81774
rect 440466 45858 440702 46094
rect 440786 45858 441022 46094
rect 440466 45538 440702 45774
rect 440786 45538 441022 45774
rect 440466 9858 440702 10094
rect 440786 9858 441022 10094
rect 440466 9538 440702 9774
rect 440786 9538 441022 9774
rect 440466 -6342 440702 -6106
rect 440786 -6342 441022 -6106
rect 440466 -6662 440702 -6426
rect 440786 -6662 441022 -6426
rect 441706 711322 441942 711558
rect 442026 711322 442262 711558
rect 441706 711002 441942 711238
rect 442026 711002 442262 711238
rect 441706 695098 441942 695334
rect 442026 695098 442262 695334
rect 441706 694778 441942 695014
rect 442026 694778 442262 695014
rect 441706 659098 441942 659334
rect 442026 659098 442262 659334
rect 441706 658778 441942 659014
rect 442026 658778 442262 659014
rect 441706 623098 441942 623334
rect 442026 623098 442262 623334
rect 441706 622778 441942 623014
rect 442026 622778 442262 623014
rect 441706 587098 441942 587334
rect 442026 587098 442262 587334
rect 441706 586778 441942 587014
rect 442026 586778 442262 587014
rect 441706 551098 441942 551334
rect 442026 551098 442262 551334
rect 441706 550778 441942 551014
rect 442026 550778 442262 551014
rect 441706 515098 441942 515334
rect 442026 515098 442262 515334
rect 441706 514778 441942 515014
rect 442026 514778 442262 515014
rect 441706 479098 441942 479334
rect 442026 479098 442262 479334
rect 441706 478778 441942 479014
rect 442026 478778 442262 479014
rect 441706 443098 441942 443334
rect 442026 443098 442262 443334
rect 441706 442778 441942 443014
rect 442026 442778 442262 443014
rect 441706 407098 441942 407334
rect 442026 407098 442262 407334
rect 441706 406778 441942 407014
rect 442026 406778 442262 407014
rect 441706 371098 441942 371334
rect 442026 371098 442262 371334
rect 441706 370778 441942 371014
rect 442026 370778 442262 371014
rect 441706 335098 441942 335334
rect 442026 335098 442262 335334
rect 441706 334778 441942 335014
rect 442026 334778 442262 335014
rect 441706 299098 441942 299334
rect 442026 299098 442262 299334
rect 441706 298778 441942 299014
rect 442026 298778 442262 299014
rect 441706 263098 441942 263334
rect 442026 263098 442262 263334
rect 441706 262778 441942 263014
rect 442026 262778 442262 263014
rect 441706 227098 441942 227334
rect 442026 227098 442262 227334
rect 441706 226778 441942 227014
rect 442026 226778 442262 227014
rect 441706 191098 441942 191334
rect 442026 191098 442262 191334
rect 441706 190778 441942 191014
rect 442026 190778 442262 191014
rect 441706 155098 441942 155334
rect 442026 155098 442262 155334
rect 441706 154778 441942 155014
rect 442026 154778 442262 155014
rect 441706 119098 441942 119334
rect 442026 119098 442262 119334
rect 441706 118778 441942 119014
rect 442026 118778 442262 119014
rect 441706 83098 441942 83334
rect 442026 83098 442262 83334
rect 441706 82778 441942 83014
rect 442026 82778 442262 83014
rect 441706 47098 441942 47334
rect 442026 47098 442262 47334
rect 441706 46778 441942 47014
rect 442026 46778 442262 47014
rect 441706 11098 441942 11334
rect 442026 11098 442262 11334
rect 441706 10778 441942 11014
rect 442026 10778 442262 11014
rect 441706 -7302 441942 -7066
rect 442026 -7302 442262 -7066
rect 441706 -7622 441942 -7386
rect 442026 -7622 442262 -7386
rect 469026 704602 469262 704838
rect 469346 704602 469582 704838
rect 469026 704282 469262 704518
rect 469346 704282 469582 704518
rect 469026 686418 469262 686654
rect 469346 686418 469582 686654
rect 469026 686098 469262 686334
rect 469346 686098 469582 686334
rect 469026 650418 469262 650654
rect 469346 650418 469582 650654
rect 469026 650098 469262 650334
rect 469346 650098 469582 650334
rect 469026 614418 469262 614654
rect 469346 614418 469582 614654
rect 469026 614098 469262 614334
rect 469346 614098 469582 614334
rect 469026 578418 469262 578654
rect 469346 578418 469582 578654
rect 469026 578098 469262 578334
rect 469346 578098 469582 578334
rect 469026 542418 469262 542654
rect 469346 542418 469582 542654
rect 469026 542098 469262 542334
rect 469346 542098 469582 542334
rect 469026 506418 469262 506654
rect 469346 506418 469582 506654
rect 469026 506098 469262 506334
rect 469346 506098 469582 506334
rect 469026 470418 469262 470654
rect 469346 470418 469582 470654
rect 469026 470098 469262 470334
rect 469346 470098 469582 470334
rect 469026 434418 469262 434654
rect 469346 434418 469582 434654
rect 469026 434098 469262 434334
rect 469346 434098 469582 434334
rect 469026 398418 469262 398654
rect 469346 398418 469582 398654
rect 469026 398098 469262 398334
rect 469346 398098 469582 398334
rect 469026 362418 469262 362654
rect 469346 362418 469582 362654
rect 469026 362098 469262 362334
rect 469346 362098 469582 362334
rect 469026 326418 469262 326654
rect 469346 326418 469582 326654
rect 469026 326098 469262 326334
rect 469346 326098 469582 326334
rect 469026 290418 469262 290654
rect 469346 290418 469582 290654
rect 469026 290098 469262 290334
rect 469346 290098 469582 290334
rect 469026 254418 469262 254654
rect 469346 254418 469582 254654
rect 469026 254098 469262 254334
rect 469346 254098 469582 254334
rect 469026 218418 469262 218654
rect 469346 218418 469582 218654
rect 469026 218098 469262 218334
rect 469346 218098 469582 218334
rect 469026 182418 469262 182654
rect 469346 182418 469582 182654
rect 469026 182098 469262 182334
rect 469346 182098 469582 182334
rect 469026 146418 469262 146654
rect 469346 146418 469582 146654
rect 469026 146098 469262 146334
rect 469346 146098 469582 146334
rect 469026 110418 469262 110654
rect 469346 110418 469582 110654
rect 469026 110098 469262 110334
rect 469346 110098 469582 110334
rect 469026 74418 469262 74654
rect 469346 74418 469582 74654
rect 469026 74098 469262 74334
rect 469346 74098 469582 74334
rect 469026 38418 469262 38654
rect 469346 38418 469582 38654
rect 469026 38098 469262 38334
rect 469346 38098 469582 38334
rect 469026 2418 469262 2654
rect 469346 2418 469582 2654
rect 469026 2098 469262 2334
rect 469346 2098 469582 2334
rect 469026 -582 469262 -346
rect 469346 -582 469582 -346
rect 469026 -902 469262 -666
rect 469346 -902 469582 -666
rect 470266 705562 470502 705798
rect 470586 705562 470822 705798
rect 470266 705242 470502 705478
rect 470586 705242 470822 705478
rect 470266 687658 470502 687894
rect 470586 687658 470822 687894
rect 470266 687338 470502 687574
rect 470586 687338 470822 687574
rect 470266 651658 470502 651894
rect 470586 651658 470822 651894
rect 470266 651338 470502 651574
rect 470586 651338 470822 651574
rect 470266 615658 470502 615894
rect 470586 615658 470822 615894
rect 470266 615338 470502 615574
rect 470586 615338 470822 615574
rect 470266 579658 470502 579894
rect 470586 579658 470822 579894
rect 470266 579338 470502 579574
rect 470586 579338 470822 579574
rect 470266 543658 470502 543894
rect 470586 543658 470822 543894
rect 470266 543338 470502 543574
rect 470586 543338 470822 543574
rect 470266 507658 470502 507894
rect 470586 507658 470822 507894
rect 470266 507338 470502 507574
rect 470586 507338 470822 507574
rect 470266 471658 470502 471894
rect 470586 471658 470822 471894
rect 470266 471338 470502 471574
rect 470586 471338 470822 471574
rect 470266 435658 470502 435894
rect 470586 435658 470822 435894
rect 470266 435338 470502 435574
rect 470586 435338 470822 435574
rect 470266 399658 470502 399894
rect 470586 399658 470822 399894
rect 470266 399338 470502 399574
rect 470586 399338 470822 399574
rect 470266 363658 470502 363894
rect 470586 363658 470822 363894
rect 470266 363338 470502 363574
rect 470586 363338 470822 363574
rect 470266 327658 470502 327894
rect 470586 327658 470822 327894
rect 470266 327338 470502 327574
rect 470586 327338 470822 327574
rect 470266 291658 470502 291894
rect 470586 291658 470822 291894
rect 470266 291338 470502 291574
rect 470586 291338 470822 291574
rect 470266 255658 470502 255894
rect 470586 255658 470822 255894
rect 470266 255338 470502 255574
rect 470586 255338 470822 255574
rect 470266 219658 470502 219894
rect 470586 219658 470822 219894
rect 470266 219338 470502 219574
rect 470586 219338 470822 219574
rect 470266 183658 470502 183894
rect 470586 183658 470822 183894
rect 470266 183338 470502 183574
rect 470586 183338 470822 183574
rect 470266 147658 470502 147894
rect 470586 147658 470822 147894
rect 470266 147338 470502 147574
rect 470586 147338 470822 147574
rect 470266 111658 470502 111894
rect 470586 111658 470822 111894
rect 470266 111338 470502 111574
rect 470586 111338 470822 111574
rect 470266 75658 470502 75894
rect 470586 75658 470822 75894
rect 470266 75338 470502 75574
rect 470586 75338 470822 75574
rect 470266 39658 470502 39894
rect 470586 39658 470822 39894
rect 470266 39338 470502 39574
rect 470586 39338 470822 39574
rect 470266 3658 470502 3894
rect 470586 3658 470822 3894
rect 470266 3338 470502 3574
rect 470586 3338 470822 3574
rect 470266 -1542 470502 -1306
rect 470586 -1542 470822 -1306
rect 470266 -1862 470502 -1626
rect 470586 -1862 470822 -1626
rect 471506 706522 471742 706758
rect 471826 706522 472062 706758
rect 471506 706202 471742 706438
rect 471826 706202 472062 706438
rect 471506 688898 471742 689134
rect 471826 688898 472062 689134
rect 471506 688578 471742 688814
rect 471826 688578 472062 688814
rect 471506 652898 471742 653134
rect 471826 652898 472062 653134
rect 471506 652578 471742 652814
rect 471826 652578 472062 652814
rect 471506 616898 471742 617134
rect 471826 616898 472062 617134
rect 471506 616578 471742 616814
rect 471826 616578 472062 616814
rect 471506 580898 471742 581134
rect 471826 580898 472062 581134
rect 471506 580578 471742 580814
rect 471826 580578 472062 580814
rect 471506 544898 471742 545134
rect 471826 544898 472062 545134
rect 471506 544578 471742 544814
rect 471826 544578 472062 544814
rect 471506 508898 471742 509134
rect 471826 508898 472062 509134
rect 471506 508578 471742 508814
rect 471826 508578 472062 508814
rect 471506 472898 471742 473134
rect 471826 472898 472062 473134
rect 471506 472578 471742 472814
rect 471826 472578 472062 472814
rect 471506 436898 471742 437134
rect 471826 436898 472062 437134
rect 471506 436578 471742 436814
rect 471826 436578 472062 436814
rect 471506 400898 471742 401134
rect 471826 400898 472062 401134
rect 471506 400578 471742 400814
rect 471826 400578 472062 400814
rect 471506 364898 471742 365134
rect 471826 364898 472062 365134
rect 471506 364578 471742 364814
rect 471826 364578 472062 364814
rect 472746 707482 472982 707718
rect 473066 707482 473302 707718
rect 472746 707162 472982 707398
rect 473066 707162 473302 707398
rect 472746 690138 472982 690374
rect 473066 690138 473302 690374
rect 472746 689818 472982 690054
rect 473066 689818 473302 690054
rect 472746 654138 472982 654374
rect 473066 654138 473302 654374
rect 472746 653818 472982 654054
rect 473066 653818 473302 654054
rect 472746 618138 472982 618374
rect 473066 618138 473302 618374
rect 472746 617818 472982 618054
rect 473066 617818 473302 618054
rect 472746 582138 472982 582374
rect 473066 582138 473302 582374
rect 472746 581818 472982 582054
rect 473066 581818 473302 582054
rect 472746 546138 472982 546374
rect 473066 546138 473302 546374
rect 472746 545818 472982 546054
rect 473066 545818 473302 546054
rect 472746 510138 472982 510374
rect 473066 510138 473302 510374
rect 472746 509818 472982 510054
rect 473066 509818 473302 510054
rect 472746 474138 472982 474374
rect 473066 474138 473302 474374
rect 472746 473818 472982 474054
rect 473066 473818 473302 474054
rect 473986 708442 474222 708678
rect 474306 708442 474542 708678
rect 473986 708122 474222 708358
rect 474306 708122 474542 708358
rect 473986 691378 474222 691614
rect 474306 691378 474542 691614
rect 473986 691058 474222 691294
rect 474306 691058 474542 691294
rect 473986 655378 474222 655614
rect 474306 655378 474542 655614
rect 473986 655058 474222 655294
rect 474306 655058 474542 655294
rect 473986 619378 474222 619614
rect 474306 619378 474542 619614
rect 473986 619058 474222 619294
rect 474306 619058 474542 619294
rect 473986 583378 474222 583614
rect 474306 583378 474542 583614
rect 473986 583058 474222 583294
rect 474306 583058 474542 583294
rect 473986 547378 474222 547614
rect 474306 547378 474542 547614
rect 473986 547058 474222 547294
rect 474306 547058 474542 547294
rect 473986 511378 474222 511614
rect 474306 511378 474542 511614
rect 473986 511058 474222 511294
rect 474306 511058 474542 511294
rect 473986 475378 474222 475614
rect 474306 475378 474542 475614
rect 473986 475058 474222 475294
rect 474306 475058 474542 475294
rect 472746 438138 472982 438374
rect 473066 438138 473302 438374
rect 472746 437818 472982 438054
rect 473066 437818 473302 438054
rect 473986 439378 474222 439614
rect 474306 439378 474542 439614
rect 473986 439058 474222 439294
rect 474306 439058 474542 439294
rect 472746 402138 472982 402374
rect 473066 402138 473302 402374
rect 472746 401818 472982 402054
rect 473066 401818 473302 402054
rect 473986 403378 474222 403614
rect 474306 403378 474542 403614
rect 473986 403058 474222 403294
rect 474306 403058 474542 403294
rect 472746 366138 472982 366374
rect 473066 366138 473302 366374
rect 472746 365818 472982 366054
rect 473066 365818 473302 366054
rect 475226 709402 475462 709638
rect 475546 709402 475782 709638
rect 475226 709082 475462 709318
rect 475546 709082 475782 709318
rect 475226 692618 475462 692854
rect 475546 692618 475782 692854
rect 475226 692298 475462 692534
rect 475546 692298 475782 692534
rect 475226 656618 475462 656854
rect 475546 656618 475782 656854
rect 475226 656298 475462 656534
rect 475546 656298 475782 656534
rect 475226 620618 475462 620854
rect 475546 620618 475782 620854
rect 475226 620298 475462 620534
rect 475546 620298 475782 620534
rect 475226 584618 475462 584854
rect 475546 584618 475782 584854
rect 475226 584298 475462 584534
rect 475546 584298 475782 584534
rect 475226 548618 475462 548854
rect 475546 548618 475782 548854
rect 475226 548298 475462 548534
rect 475546 548298 475782 548534
rect 475226 512618 475462 512854
rect 475546 512618 475782 512854
rect 475226 512298 475462 512534
rect 475546 512298 475782 512534
rect 475226 476618 475462 476854
rect 475546 476618 475782 476854
rect 475226 476298 475462 476534
rect 475546 476298 475782 476534
rect 475226 440618 475462 440854
rect 475546 440618 475782 440854
rect 475226 440298 475462 440534
rect 475546 440298 475782 440534
rect 475226 404618 475462 404854
rect 475546 404618 475782 404854
rect 475226 404298 475462 404534
rect 475546 404298 475782 404534
rect 473986 367378 474222 367614
rect 474306 367378 474542 367614
rect 473986 367058 474222 367294
rect 474306 367058 474542 367294
rect 475226 368618 475462 368854
rect 475546 368618 475782 368854
rect 475226 368298 475462 368534
rect 475546 368298 475782 368534
rect 476466 710362 476702 710598
rect 476786 710362 477022 710598
rect 476466 710042 476702 710278
rect 476786 710042 477022 710278
rect 476466 693858 476702 694094
rect 476786 693858 477022 694094
rect 476466 693538 476702 693774
rect 476786 693538 477022 693774
rect 476466 657858 476702 658094
rect 476786 657858 477022 658094
rect 476466 657538 476702 657774
rect 476786 657538 477022 657774
rect 476466 621858 476702 622094
rect 476786 621858 477022 622094
rect 476466 621538 476702 621774
rect 476786 621538 477022 621774
rect 476466 585858 476702 586094
rect 476786 585858 477022 586094
rect 476466 585538 476702 585774
rect 476786 585538 477022 585774
rect 476466 549858 476702 550094
rect 476786 549858 477022 550094
rect 476466 549538 476702 549774
rect 476786 549538 477022 549774
rect 476466 513858 476702 514094
rect 476786 513858 477022 514094
rect 476466 513538 476702 513774
rect 476786 513538 477022 513774
rect 476466 477858 476702 478094
rect 476786 477858 477022 478094
rect 476466 477538 476702 477774
rect 476786 477538 477022 477774
rect 476466 441858 476702 442094
rect 476786 441858 477022 442094
rect 476466 441538 476702 441774
rect 476786 441538 477022 441774
rect 476466 405858 476702 406094
rect 476786 405858 477022 406094
rect 476466 405538 476702 405774
rect 476786 405538 477022 405774
rect 476466 369858 476702 370094
rect 476786 369858 477022 370094
rect 476466 369538 476702 369774
rect 476786 369538 477022 369774
rect 477706 711322 477942 711558
rect 478026 711322 478262 711558
rect 477706 711002 477942 711238
rect 478026 711002 478262 711238
rect 477706 695098 477942 695334
rect 478026 695098 478262 695334
rect 477706 694778 477942 695014
rect 478026 694778 478262 695014
rect 477706 659098 477942 659334
rect 478026 659098 478262 659334
rect 477706 658778 477942 659014
rect 478026 658778 478262 659014
rect 477706 623098 477942 623334
rect 478026 623098 478262 623334
rect 477706 622778 477942 623014
rect 478026 622778 478262 623014
rect 477706 587098 477942 587334
rect 478026 587098 478262 587334
rect 477706 586778 477942 587014
rect 478026 586778 478262 587014
rect 477706 551098 477942 551334
rect 478026 551098 478262 551334
rect 477706 550778 477942 551014
rect 478026 550778 478262 551014
rect 477706 515098 477942 515334
rect 478026 515098 478262 515334
rect 477706 514778 477942 515014
rect 478026 514778 478262 515014
rect 477706 479098 477942 479334
rect 478026 479098 478262 479334
rect 477706 478778 477942 479014
rect 478026 478778 478262 479014
rect 505026 704602 505262 704838
rect 505346 704602 505582 704838
rect 505026 704282 505262 704518
rect 505346 704282 505582 704518
rect 505026 686418 505262 686654
rect 505346 686418 505582 686654
rect 505026 686098 505262 686334
rect 505346 686098 505582 686334
rect 505026 650418 505262 650654
rect 505346 650418 505582 650654
rect 505026 650098 505262 650334
rect 505346 650098 505582 650334
rect 505026 614418 505262 614654
rect 505346 614418 505582 614654
rect 505026 614098 505262 614334
rect 505346 614098 505582 614334
rect 505026 578418 505262 578654
rect 505346 578418 505582 578654
rect 505026 578098 505262 578334
rect 505346 578098 505582 578334
rect 505026 542418 505262 542654
rect 505346 542418 505582 542654
rect 505026 542098 505262 542334
rect 505346 542098 505582 542334
rect 505026 506418 505262 506654
rect 505346 506418 505582 506654
rect 505026 506098 505262 506334
rect 505346 506098 505582 506334
rect 505026 470418 505262 470654
rect 505346 470418 505582 470654
rect 505026 470098 505262 470334
rect 505346 470098 505582 470334
rect 477706 443098 477942 443334
rect 478026 443098 478262 443334
rect 477706 442778 477942 443014
rect 478026 442778 478262 443014
rect 477706 407098 477942 407334
rect 478026 407098 478262 407334
rect 477706 406778 477942 407014
rect 478026 406778 478262 407014
rect 505026 434418 505262 434654
rect 505346 434418 505582 434654
rect 505026 434098 505262 434334
rect 505346 434098 505582 434334
rect 477706 371098 477942 371334
rect 478026 371098 478262 371334
rect 477706 370778 477942 371014
rect 478026 370778 478262 371014
rect 471506 328898 471742 329134
rect 471826 328898 472062 329134
rect 471506 328578 471742 328814
rect 471826 328578 472062 328814
rect 471506 292898 471742 293134
rect 471826 292898 472062 293134
rect 471506 292578 471742 292814
rect 471826 292578 472062 292814
rect 472746 330138 472982 330374
rect 473066 330138 473302 330374
rect 472746 329818 472982 330054
rect 473066 329818 473302 330054
rect 473986 331378 474222 331614
rect 474306 331378 474542 331614
rect 473986 331058 474222 331294
rect 474306 331058 474542 331294
rect 472746 294138 472982 294374
rect 473066 294138 473302 294374
rect 472746 293818 472982 294054
rect 473066 293818 473302 294054
rect 473986 295378 474222 295614
rect 474306 295378 474542 295614
rect 473986 295058 474222 295294
rect 474306 295058 474542 295294
rect 475226 332618 475462 332854
rect 475546 332618 475782 332854
rect 475226 332298 475462 332534
rect 475546 332298 475782 332534
rect 475226 296618 475462 296854
rect 475546 296618 475782 296854
rect 475226 296298 475462 296534
rect 475546 296298 475782 296534
rect 476466 333858 476702 334094
rect 476786 333858 477022 334094
rect 476466 333538 476702 333774
rect 476786 333538 477022 333774
rect 476466 297858 476702 298094
rect 476786 297858 477022 298094
rect 476466 297538 476702 297774
rect 476786 297538 477022 297774
rect 477706 335098 477942 335334
rect 478026 335098 478262 335334
rect 477706 334778 477942 335014
rect 478026 334778 478262 335014
rect 505026 398418 505262 398654
rect 505346 398418 505582 398654
rect 505026 398098 505262 398334
rect 505346 398098 505582 398334
rect 505026 362418 505262 362654
rect 505346 362418 505582 362654
rect 505026 362098 505262 362334
rect 505346 362098 505582 362334
rect 477706 299098 477942 299334
rect 478026 299098 478262 299334
rect 477706 298778 477942 299014
rect 478026 298778 478262 299014
rect 505026 326418 505262 326654
rect 505346 326418 505582 326654
rect 505026 326098 505262 326334
rect 505346 326098 505582 326334
rect 505026 290418 505262 290654
rect 505346 290418 505582 290654
rect 505026 290098 505262 290334
rect 505346 290098 505582 290334
rect 471506 256898 471742 257134
rect 471826 256898 472062 257134
rect 471506 256578 471742 256814
rect 471826 256578 472062 256814
rect 471506 220898 471742 221134
rect 471826 220898 472062 221134
rect 471506 220578 471742 220814
rect 471826 220578 472062 220814
rect 471506 184898 471742 185134
rect 471826 184898 472062 185134
rect 471506 184578 471742 184814
rect 471826 184578 472062 184814
rect 471506 148898 471742 149134
rect 471826 148898 472062 149134
rect 471506 148578 471742 148814
rect 471826 148578 472062 148814
rect 471506 112898 471742 113134
rect 471826 112898 472062 113134
rect 471506 112578 471742 112814
rect 471826 112578 472062 112814
rect 471506 76898 471742 77134
rect 471826 76898 472062 77134
rect 471506 76578 471742 76814
rect 471826 76578 472062 76814
rect 471506 40898 471742 41134
rect 471826 40898 472062 41134
rect 471506 40578 471742 40814
rect 471826 40578 472062 40814
rect 471506 4898 471742 5134
rect 471826 4898 472062 5134
rect 471506 4578 471742 4814
rect 471826 4578 472062 4814
rect 471506 -2502 471742 -2266
rect 471826 -2502 472062 -2266
rect 471506 -2822 471742 -2586
rect 471826 -2822 472062 -2586
rect 472746 258138 472982 258374
rect 473066 258138 473302 258374
rect 472746 257818 472982 258054
rect 473066 257818 473302 258054
rect 472746 222138 472982 222374
rect 473066 222138 473302 222374
rect 472746 221818 472982 222054
rect 473066 221818 473302 222054
rect 472746 186138 472982 186374
rect 473066 186138 473302 186374
rect 472746 185818 472982 186054
rect 473066 185818 473302 186054
rect 472746 150138 472982 150374
rect 473066 150138 473302 150374
rect 472746 149818 472982 150054
rect 473066 149818 473302 150054
rect 472746 114138 472982 114374
rect 473066 114138 473302 114374
rect 472746 113818 472982 114054
rect 473066 113818 473302 114054
rect 472746 78138 472982 78374
rect 473066 78138 473302 78374
rect 472746 77818 472982 78054
rect 473066 77818 473302 78054
rect 472746 42138 472982 42374
rect 473066 42138 473302 42374
rect 472746 41818 472982 42054
rect 473066 41818 473302 42054
rect 472746 6138 472982 6374
rect 473066 6138 473302 6374
rect 472746 5818 472982 6054
rect 473066 5818 473302 6054
rect 472746 -3462 472982 -3226
rect 473066 -3462 473302 -3226
rect 472746 -3782 472982 -3546
rect 473066 -3782 473302 -3546
rect 473986 259378 474222 259614
rect 474306 259378 474542 259614
rect 473986 259058 474222 259294
rect 474306 259058 474542 259294
rect 473986 223378 474222 223614
rect 474306 223378 474542 223614
rect 473986 223058 474222 223294
rect 474306 223058 474542 223294
rect 473986 187378 474222 187614
rect 474306 187378 474542 187614
rect 473986 187058 474222 187294
rect 474306 187058 474542 187294
rect 473986 151378 474222 151614
rect 474306 151378 474542 151614
rect 473986 151058 474222 151294
rect 474306 151058 474542 151294
rect 473986 115378 474222 115614
rect 474306 115378 474542 115614
rect 473986 115058 474222 115294
rect 474306 115058 474542 115294
rect 473986 79378 474222 79614
rect 474306 79378 474542 79614
rect 473986 79058 474222 79294
rect 474306 79058 474542 79294
rect 473986 43378 474222 43614
rect 474306 43378 474542 43614
rect 473986 43058 474222 43294
rect 474306 43058 474542 43294
rect 473986 7378 474222 7614
rect 474306 7378 474542 7614
rect 473986 7058 474222 7294
rect 474306 7058 474542 7294
rect 473986 -4422 474222 -4186
rect 474306 -4422 474542 -4186
rect 473986 -4742 474222 -4506
rect 474306 -4742 474542 -4506
rect 475226 260618 475462 260854
rect 475546 260618 475782 260854
rect 475226 260298 475462 260534
rect 475546 260298 475782 260534
rect 475226 224618 475462 224854
rect 475546 224618 475782 224854
rect 475226 224298 475462 224534
rect 475546 224298 475782 224534
rect 475226 188618 475462 188854
rect 475546 188618 475782 188854
rect 475226 188298 475462 188534
rect 475546 188298 475782 188534
rect 475226 152618 475462 152854
rect 475546 152618 475782 152854
rect 475226 152298 475462 152534
rect 475546 152298 475782 152534
rect 475226 116618 475462 116854
rect 475546 116618 475782 116854
rect 475226 116298 475462 116534
rect 475546 116298 475782 116534
rect 475226 80618 475462 80854
rect 475546 80618 475782 80854
rect 475226 80298 475462 80534
rect 475546 80298 475782 80534
rect 475226 44618 475462 44854
rect 475546 44618 475782 44854
rect 475226 44298 475462 44534
rect 475546 44298 475782 44534
rect 475226 8618 475462 8854
rect 475546 8618 475782 8854
rect 475226 8298 475462 8534
rect 475546 8298 475782 8534
rect 475226 -5382 475462 -5146
rect 475546 -5382 475782 -5146
rect 475226 -5702 475462 -5466
rect 475546 -5702 475782 -5466
rect 476466 261858 476702 262094
rect 476786 261858 477022 262094
rect 476466 261538 476702 261774
rect 476786 261538 477022 261774
rect 476466 225858 476702 226094
rect 476786 225858 477022 226094
rect 476466 225538 476702 225774
rect 476786 225538 477022 225774
rect 476466 189858 476702 190094
rect 476786 189858 477022 190094
rect 476466 189538 476702 189774
rect 476786 189538 477022 189774
rect 476466 153858 476702 154094
rect 476786 153858 477022 154094
rect 476466 153538 476702 153774
rect 476786 153538 477022 153774
rect 476466 117858 476702 118094
rect 476786 117858 477022 118094
rect 476466 117538 476702 117774
rect 476786 117538 477022 117774
rect 476466 81858 476702 82094
rect 476786 81858 477022 82094
rect 476466 81538 476702 81774
rect 476786 81538 477022 81774
rect 476466 45858 476702 46094
rect 476786 45858 477022 46094
rect 476466 45538 476702 45774
rect 476786 45538 477022 45774
rect 476466 9858 476702 10094
rect 476786 9858 477022 10094
rect 476466 9538 476702 9774
rect 476786 9538 477022 9774
rect 477706 263098 477942 263334
rect 478026 263098 478262 263334
rect 477706 262778 477942 263014
rect 478026 262778 478262 263014
rect 477706 227098 477942 227334
rect 478026 227098 478262 227334
rect 477706 226778 477942 227014
rect 478026 226778 478262 227014
rect 477706 191098 477942 191334
rect 478026 191098 478262 191334
rect 477706 190778 477942 191014
rect 478026 190778 478262 191014
rect 477706 155098 477942 155334
rect 478026 155098 478262 155334
rect 477706 154778 477942 155014
rect 478026 154778 478262 155014
rect 477706 119098 477942 119334
rect 478026 119098 478262 119334
rect 477706 118778 477942 119014
rect 478026 118778 478262 119014
rect 477706 83098 477942 83334
rect 478026 83098 478262 83334
rect 477706 82778 477942 83014
rect 478026 82778 478262 83014
rect 477706 47098 477942 47334
rect 478026 47098 478262 47334
rect 477706 46778 477942 47014
rect 478026 46778 478262 47014
rect 505026 254418 505262 254654
rect 505346 254418 505582 254654
rect 505026 254098 505262 254334
rect 505346 254098 505582 254334
rect 505026 218418 505262 218654
rect 505346 218418 505582 218654
rect 505026 218098 505262 218334
rect 505346 218098 505582 218334
rect 505026 182418 505262 182654
rect 505346 182418 505582 182654
rect 505026 182098 505262 182334
rect 505346 182098 505582 182334
rect 505026 146418 505262 146654
rect 505346 146418 505582 146654
rect 505026 146098 505262 146334
rect 505346 146098 505582 146334
rect 505026 110418 505262 110654
rect 505346 110418 505582 110654
rect 505026 110098 505262 110334
rect 505346 110098 505582 110334
rect 505026 74418 505262 74654
rect 505346 74418 505582 74654
rect 505026 74098 505262 74334
rect 505346 74098 505582 74334
rect 477706 11098 477942 11334
rect 478026 11098 478262 11334
rect 477706 10778 477942 11014
rect 478026 10778 478262 11014
rect 476466 -6342 476702 -6106
rect 476786 -6342 477022 -6106
rect 476466 -6662 476702 -6426
rect 476786 -6662 477022 -6426
rect 477706 -7302 477942 -7066
rect 478026 -7302 478262 -7066
rect 477706 -7622 477942 -7386
rect 478026 -7622 478262 -7386
rect 505026 38418 505262 38654
rect 505346 38418 505582 38654
rect 505026 38098 505262 38334
rect 505346 38098 505582 38334
rect 505026 2418 505262 2654
rect 505346 2418 505582 2654
rect 505026 2098 505262 2334
rect 505346 2098 505582 2334
rect 505026 -582 505262 -346
rect 505346 -582 505582 -346
rect 505026 -902 505262 -666
rect 505346 -902 505582 -666
rect 506266 705562 506502 705798
rect 506586 705562 506822 705798
rect 506266 705242 506502 705478
rect 506586 705242 506822 705478
rect 506266 687658 506502 687894
rect 506586 687658 506822 687894
rect 506266 687338 506502 687574
rect 506586 687338 506822 687574
rect 506266 651658 506502 651894
rect 506586 651658 506822 651894
rect 506266 651338 506502 651574
rect 506586 651338 506822 651574
rect 506266 615658 506502 615894
rect 506586 615658 506822 615894
rect 506266 615338 506502 615574
rect 506586 615338 506822 615574
rect 506266 579658 506502 579894
rect 506586 579658 506822 579894
rect 506266 579338 506502 579574
rect 506586 579338 506822 579574
rect 506266 543658 506502 543894
rect 506586 543658 506822 543894
rect 506266 543338 506502 543574
rect 506586 543338 506822 543574
rect 506266 507658 506502 507894
rect 506586 507658 506822 507894
rect 506266 507338 506502 507574
rect 506586 507338 506822 507574
rect 506266 471658 506502 471894
rect 506586 471658 506822 471894
rect 506266 471338 506502 471574
rect 506586 471338 506822 471574
rect 506266 435658 506502 435894
rect 506586 435658 506822 435894
rect 506266 435338 506502 435574
rect 506586 435338 506822 435574
rect 506266 399658 506502 399894
rect 506586 399658 506822 399894
rect 506266 399338 506502 399574
rect 506586 399338 506822 399574
rect 506266 363658 506502 363894
rect 506586 363658 506822 363894
rect 506266 363338 506502 363574
rect 506586 363338 506822 363574
rect 506266 327658 506502 327894
rect 506586 327658 506822 327894
rect 506266 327338 506502 327574
rect 506586 327338 506822 327574
rect 506266 291658 506502 291894
rect 506586 291658 506822 291894
rect 506266 291338 506502 291574
rect 506586 291338 506822 291574
rect 506266 255658 506502 255894
rect 506586 255658 506822 255894
rect 506266 255338 506502 255574
rect 506586 255338 506822 255574
rect 506266 219658 506502 219894
rect 506586 219658 506822 219894
rect 506266 219338 506502 219574
rect 506586 219338 506822 219574
rect 506266 183658 506502 183894
rect 506586 183658 506822 183894
rect 506266 183338 506502 183574
rect 506586 183338 506822 183574
rect 506266 147658 506502 147894
rect 506586 147658 506822 147894
rect 506266 147338 506502 147574
rect 506586 147338 506822 147574
rect 506266 111658 506502 111894
rect 506586 111658 506822 111894
rect 506266 111338 506502 111574
rect 506586 111338 506822 111574
rect 506266 75658 506502 75894
rect 506586 75658 506822 75894
rect 506266 75338 506502 75574
rect 506586 75338 506822 75574
rect 506266 39658 506502 39894
rect 506586 39658 506822 39894
rect 506266 39338 506502 39574
rect 506586 39338 506822 39574
rect 506266 3658 506502 3894
rect 506586 3658 506822 3894
rect 506266 3338 506502 3574
rect 506586 3338 506822 3574
rect 506266 -1542 506502 -1306
rect 506586 -1542 506822 -1306
rect 506266 -1862 506502 -1626
rect 506586 -1862 506822 -1626
rect 507506 706522 507742 706758
rect 507826 706522 508062 706758
rect 507506 706202 507742 706438
rect 507826 706202 508062 706438
rect 507506 688898 507742 689134
rect 507826 688898 508062 689134
rect 507506 688578 507742 688814
rect 507826 688578 508062 688814
rect 507506 652898 507742 653134
rect 507826 652898 508062 653134
rect 507506 652578 507742 652814
rect 507826 652578 508062 652814
rect 507506 616898 507742 617134
rect 507826 616898 508062 617134
rect 507506 616578 507742 616814
rect 507826 616578 508062 616814
rect 507506 580898 507742 581134
rect 507826 580898 508062 581134
rect 507506 580578 507742 580814
rect 507826 580578 508062 580814
rect 507506 544898 507742 545134
rect 507826 544898 508062 545134
rect 507506 544578 507742 544814
rect 507826 544578 508062 544814
rect 507506 508898 507742 509134
rect 507826 508898 508062 509134
rect 507506 508578 507742 508814
rect 507826 508578 508062 508814
rect 507506 472898 507742 473134
rect 507826 472898 508062 473134
rect 507506 472578 507742 472814
rect 507826 472578 508062 472814
rect 507506 436898 507742 437134
rect 507826 436898 508062 437134
rect 507506 436578 507742 436814
rect 507826 436578 508062 436814
rect 507506 400898 507742 401134
rect 507826 400898 508062 401134
rect 507506 400578 507742 400814
rect 507826 400578 508062 400814
rect 507506 364898 507742 365134
rect 507826 364898 508062 365134
rect 507506 364578 507742 364814
rect 507826 364578 508062 364814
rect 507506 328898 507742 329134
rect 507826 328898 508062 329134
rect 507506 328578 507742 328814
rect 507826 328578 508062 328814
rect 507506 292898 507742 293134
rect 507826 292898 508062 293134
rect 507506 292578 507742 292814
rect 507826 292578 508062 292814
rect 507506 256898 507742 257134
rect 507826 256898 508062 257134
rect 507506 256578 507742 256814
rect 507826 256578 508062 256814
rect 507506 220898 507742 221134
rect 507826 220898 508062 221134
rect 507506 220578 507742 220814
rect 507826 220578 508062 220814
rect 507506 184898 507742 185134
rect 507826 184898 508062 185134
rect 507506 184578 507742 184814
rect 507826 184578 508062 184814
rect 507506 148898 507742 149134
rect 507826 148898 508062 149134
rect 507506 148578 507742 148814
rect 507826 148578 508062 148814
rect 507506 112898 507742 113134
rect 507826 112898 508062 113134
rect 507506 112578 507742 112814
rect 507826 112578 508062 112814
rect 507506 76898 507742 77134
rect 507826 76898 508062 77134
rect 507506 76578 507742 76814
rect 507826 76578 508062 76814
rect 507506 40898 507742 41134
rect 507826 40898 508062 41134
rect 507506 40578 507742 40814
rect 507826 40578 508062 40814
rect 507506 4898 507742 5134
rect 507826 4898 508062 5134
rect 507506 4578 507742 4814
rect 507826 4578 508062 4814
rect 507506 -2502 507742 -2266
rect 507826 -2502 508062 -2266
rect 507506 -2822 507742 -2586
rect 507826 -2822 508062 -2586
rect 508746 707482 508982 707718
rect 509066 707482 509302 707718
rect 508746 707162 508982 707398
rect 509066 707162 509302 707398
rect 508746 690138 508982 690374
rect 509066 690138 509302 690374
rect 508746 689818 508982 690054
rect 509066 689818 509302 690054
rect 508746 654138 508982 654374
rect 509066 654138 509302 654374
rect 508746 653818 508982 654054
rect 509066 653818 509302 654054
rect 508746 618138 508982 618374
rect 509066 618138 509302 618374
rect 508746 617818 508982 618054
rect 509066 617818 509302 618054
rect 508746 582138 508982 582374
rect 509066 582138 509302 582374
rect 508746 581818 508982 582054
rect 509066 581818 509302 582054
rect 508746 546138 508982 546374
rect 509066 546138 509302 546374
rect 508746 545818 508982 546054
rect 509066 545818 509302 546054
rect 508746 510138 508982 510374
rect 509066 510138 509302 510374
rect 508746 509818 508982 510054
rect 509066 509818 509302 510054
rect 508746 474138 508982 474374
rect 509066 474138 509302 474374
rect 508746 473818 508982 474054
rect 509066 473818 509302 474054
rect 508746 438138 508982 438374
rect 509066 438138 509302 438374
rect 508746 437818 508982 438054
rect 509066 437818 509302 438054
rect 508746 402138 508982 402374
rect 509066 402138 509302 402374
rect 508746 401818 508982 402054
rect 509066 401818 509302 402054
rect 508746 366138 508982 366374
rect 509066 366138 509302 366374
rect 508746 365818 508982 366054
rect 509066 365818 509302 366054
rect 508746 330138 508982 330374
rect 509066 330138 509302 330374
rect 508746 329818 508982 330054
rect 509066 329818 509302 330054
rect 508746 294138 508982 294374
rect 509066 294138 509302 294374
rect 508746 293818 508982 294054
rect 509066 293818 509302 294054
rect 508746 258138 508982 258374
rect 509066 258138 509302 258374
rect 508746 257818 508982 258054
rect 509066 257818 509302 258054
rect 508746 222138 508982 222374
rect 509066 222138 509302 222374
rect 508746 221818 508982 222054
rect 509066 221818 509302 222054
rect 508746 186138 508982 186374
rect 509066 186138 509302 186374
rect 508746 185818 508982 186054
rect 509066 185818 509302 186054
rect 508746 150138 508982 150374
rect 509066 150138 509302 150374
rect 508746 149818 508982 150054
rect 509066 149818 509302 150054
rect 508746 114138 508982 114374
rect 509066 114138 509302 114374
rect 508746 113818 508982 114054
rect 509066 113818 509302 114054
rect 508746 78138 508982 78374
rect 509066 78138 509302 78374
rect 508746 77818 508982 78054
rect 509066 77818 509302 78054
rect 508746 42138 508982 42374
rect 509066 42138 509302 42374
rect 508746 41818 508982 42054
rect 509066 41818 509302 42054
rect 508746 6138 508982 6374
rect 509066 6138 509302 6374
rect 508746 5818 508982 6054
rect 509066 5818 509302 6054
rect 508746 -3462 508982 -3226
rect 509066 -3462 509302 -3226
rect 508746 -3782 508982 -3546
rect 509066 -3782 509302 -3546
rect 509986 708442 510222 708678
rect 510306 708442 510542 708678
rect 509986 708122 510222 708358
rect 510306 708122 510542 708358
rect 509986 691378 510222 691614
rect 510306 691378 510542 691614
rect 509986 691058 510222 691294
rect 510306 691058 510542 691294
rect 509986 655378 510222 655614
rect 510306 655378 510542 655614
rect 509986 655058 510222 655294
rect 510306 655058 510542 655294
rect 509986 619378 510222 619614
rect 510306 619378 510542 619614
rect 509986 619058 510222 619294
rect 510306 619058 510542 619294
rect 509986 583378 510222 583614
rect 510306 583378 510542 583614
rect 509986 583058 510222 583294
rect 510306 583058 510542 583294
rect 509986 547378 510222 547614
rect 510306 547378 510542 547614
rect 509986 547058 510222 547294
rect 510306 547058 510542 547294
rect 509986 511378 510222 511614
rect 510306 511378 510542 511614
rect 509986 511058 510222 511294
rect 510306 511058 510542 511294
rect 509986 475378 510222 475614
rect 510306 475378 510542 475614
rect 509986 475058 510222 475294
rect 510306 475058 510542 475294
rect 509986 439378 510222 439614
rect 510306 439378 510542 439614
rect 509986 439058 510222 439294
rect 510306 439058 510542 439294
rect 509986 403378 510222 403614
rect 510306 403378 510542 403614
rect 509986 403058 510222 403294
rect 510306 403058 510542 403294
rect 509986 367378 510222 367614
rect 510306 367378 510542 367614
rect 509986 367058 510222 367294
rect 510306 367058 510542 367294
rect 509986 331378 510222 331614
rect 510306 331378 510542 331614
rect 509986 331058 510222 331294
rect 510306 331058 510542 331294
rect 509986 295378 510222 295614
rect 510306 295378 510542 295614
rect 509986 295058 510222 295294
rect 510306 295058 510542 295294
rect 509986 259378 510222 259614
rect 510306 259378 510542 259614
rect 509986 259058 510222 259294
rect 510306 259058 510542 259294
rect 509986 223378 510222 223614
rect 510306 223378 510542 223614
rect 509986 223058 510222 223294
rect 510306 223058 510542 223294
rect 509986 187378 510222 187614
rect 510306 187378 510542 187614
rect 509986 187058 510222 187294
rect 510306 187058 510542 187294
rect 509986 151378 510222 151614
rect 510306 151378 510542 151614
rect 509986 151058 510222 151294
rect 510306 151058 510542 151294
rect 509986 115378 510222 115614
rect 510306 115378 510542 115614
rect 509986 115058 510222 115294
rect 510306 115058 510542 115294
rect 509986 79378 510222 79614
rect 510306 79378 510542 79614
rect 509986 79058 510222 79294
rect 510306 79058 510542 79294
rect 509986 43378 510222 43614
rect 510306 43378 510542 43614
rect 509986 43058 510222 43294
rect 510306 43058 510542 43294
rect 509986 7378 510222 7614
rect 510306 7378 510542 7614
rect 509986 7058 510222 7294
rect 510306 7058 510542 7294
rect 509986 -4422 510222 -4186
rect 510306 -4422 510542 -4186
rect 509986 -4742 510222 -4506
rect 510306 -4742 510542 -4506
rect 511226 709402 511462 709638
rect 511546 709402 511782 709638
rect 511226 709082 511462 709318
rect 511546 709082 511782 709318
rect 511226 692618 511462 692854
rect 511546 692618 511782 692854
rect 511226 692298 511462 692534
rect 511546 692298 511782 692534
rect 511226 656618 511462 656854
rect 511546 656618 511782 656854
rect 511226 656298 511462 656534
rect 511546 656298 511782 656534
rect 511226 620618 511462 620854
rect 511546 620618 511782 620854
rect 511226 620298 511462 620534
rect 511546 620298 511782 620534
rect 511226 584618 511462 584854
rect 511546 584618 511782 584854
rect 511226 584298 511462 584534
rect 511546 584298 511782 584534
rect 511226 548618 511462 548854
rect 511546 548618 511782 548854
rect 511226 548298 511462 548534
rect 511546 548298 511782 548534
rect 511226 512618 511462 512854
rect 511546 512618 511782 512854
rect 511226 512298 511462 512534
rect 511546 512298 511782 512534
rect 511226 476618 511462 476854
rect 511546 476618 511782 476854
rect 511226 476298 511462 476534
rect 511546 476298 511782 476534
rect 511226 440618 511462 440854
rect 511546 440618 511782 440854
rect 511226 440298 511462 440534
rect 511546 440298 511782 440534
rect 511226 404618 511462 404854
rect 511546 404618 511782 404854
rect 511226 404298 511462 404534
rect 511546 404298 511782 404534
rect 511226 368618 511462 368854
rect 511546 368618 511782 368854
rect 511226 368298 511462 368534
rect 511546 368298 511782 368534
rect 511226 332618 511462 332854
rect 511546 332618 511782 332854
rect 511226 332298 511462 332534
rect 511546 332298 511782 332534
rect 511226 296618 511462 296854
rect 511546 296618 511782 296854
rect 511226 296298 511462 296534
rect 511546 296298 511782 296534
rect 511226 260618 511462 260854
rect 511546 260618 511782 260854
rect 511226 260298 511462 260534
rect 511546 260298 511782 260534
rect 511226 224618 511462 224854
rect 511546 224618 511782 224854
rect 511226 224298 511462 224534
rect 511546 224298 511782 224534
rect 511226 188618 511462 188854
rect 511546 188618 511782 188854
rect 511226 188298 511462 188534
rect 511546 188298 511782 188534
rect 511226 152618 511462 152854
rect 511546 152618 511782 152854
rect 511226 152298 511462 152534
rect 511546 152298 511782 152534
rect 511226 116618 511462 116854
rect 511546 116618 511782 116854
rect 511226 116298 511462 116534
rect 511546 116298 511782 116534
rect 511226 80618 511462 80854
rect 511546 80618 511782 80854
rect 511226 80298 511462 80534
rect 511546 80298 511782 80534
rect 511226 44618 511462 44854
rect 511546 44618 511782 44854
rect 511226 44298 511462 44534
rect 511546 44298 511782 44534
rect 511226 8618 511462 8854
rect 511546 8618 511782 8854
rect 511226 8298 511462 8534
rect 511546 8298 511782 8534
rect 511226 -5382 511462 -5146
rect 511546 -5382 511782 -5146
rect 511226 -5702 511462 -5466
rect 511546 -5702 511782 -5466
rect 512466 710362 512702 710598
rect 512786 710362 513022 710598
rect 512466 710042 512702 710278
rect 512786 710042 513022 710278
rect 512466 693858 512702 694094
rect 512786 693858 513022 694094
rect 512466 693538 512702 693774
rect 512786 693538 513022 693774
rect 512466 657858 512702 658094
rect 512786 657858 513022 658094
rect 512466 657538 512702 657774
rect 512786 657538 513022 657774
rect 512466 621858 512702 622094
rect 512786 621858 513022 622094
rect 512466 621538 512702 621774
rect 512786 621538 513022 621774
rect 512466 585858 512702 586094
rect 512786 585858 513022 586094
rect 512466 585538 512702 585774
rect 512786 585538 513022 585774
rect 512466 549858 512702 550094
rect 512786 549858 513022 550094
rect 512466 549538 512702 549774
rect 512786 549538 513022 549774
rect 512466 513858 512702 514094
rect 512786 513858 513022 514094
rect 512466 513538 512702 513774
rect 512786 513538 513022 513774
rect 512466 477858 512702 478094
rect 512786 477858 513022 478094
rect 512466 477538 512702 477774
rect 512786 477538 513022 477774
rect 512466 441858 512702 442094
rect 512786 441858 513022 442094
rect 512466 441538 512702 441774
rect 512786 441538 513022 441774
rect 512466 405858 512702 406094
rect 512786 405858 513022 406094
rect 512466 405538 512702 405774
rect 512786 405538 513022 405774
rect 512466 369858 512702 370094
rect 512786 369858 513022 370094
rect 512466 369538 512702 369774
rect 512786 369538 513022 369774
rect 512466 333858 512702 334094
rect 512786 333858 513022 334094
rect 512466 333538 512702 333774
rect 512786 333538 513022 333774
rect 512466 297858 512702 298094
rect 512786 297858 513022 298094
rect 512466 297538 512702 297774
rect 512786 297538 513022 297774
rect 512466 261858 512702 262094
rect 512786 261858 513022 262094
rect 512466 261538 512702 261774
rect 512786 261538 513022 261774
rect 512466 225858 512702 226094
rect 512786 225858 513022 226094
rect 512466 225538 512702 225774
rect 512786 225538 513022 225774
rect 512466 189858 512702 190094
rect 512786 189858 513022 190094
rect 512466 189538 512702 189774
rect 512786 189538 513022 189774
rect 512466 153858 512702 154094
rect 512786 153858 513022 154094
rect 512466 153538 512702 153774
rect 512786 153538 513022 153774
rect 512466 117858 512702 118094
rect 512786 117858 513022 118094
rect 512466 117538 512702 117774
rect 512786 117538 513022 117774
rect 512466 81858 512702 82094
rect 512786 81858 513022 82094
rect 512466 81538 512702 81774
rect 512786 81538 513022 81774
rect 512466 45858 512702 46094
rect 512786 45858 513022 46094
rect 512466 45538 512702 45774
rect 512786 45538 513022 45774
rect 512466 9858 512702 10094
rect 512786 9858 513022 10094
rect 512466 9538 512702 9774
rect 512786 9538 513022 9774
rect 512466 -6342 512702 -6106
rect 512786 -6342 513022 -6106
rect 512466 -6662 512702 -6426
rect 512786 -6662 513022 -6426
rect 513706 711322 513942 711558
rect 514026 711322 514262 711558
rect 513706 711002 513942 711238
rect 514026 711002 514262 711238
rect 513706 695098 513942 695334
rect 514026 695098 514262 695334
rect 513706 694778 513942 695014
rect 514026 694778 514262 695014
rect 513706 659098 513942 659334
rect 514026 659098 514262 659334
rect 513706 658778 513942 659014
rect 514026 658778 514262 659014
rect 513706 623098 513942 623334
rect 514026 623098 514262 623334
rect 513706 622778 513942 623014
rect 514026 622778 514262 623014
rect 513706 587098 513942 587334
rect 514026 587098 514262 587334
rect 513706 586778 513942 587014
rect 514026 586778 514262 587014
rect 513706 551098 513942 551334
rect 514026 551098 514262 551334
rect 513706 550778 513942 551014
rect 514026 550778 514262 551014
rect 513706 515098 513942 515334
rect 514026 515098 514262 515334
rect 513706 514778 513942 515014
rect 514026 514778 514262 515014
rect 513706 479098 513942 479334
rect 514026 479098 514262 479334
rect 513706 478778 513942 479014
rect 514026 478778 514262 479014
rect 541026 704602 541262 704838
rect 541346 704602 541582 704838
rect 541026 704282 541262 704518
rect 541346 704282 541582 704518
rect 541026 686418 541262 686654
rect 541346 686418 541582 686654
rect 541026 686098 541262 686334
rect 541346 686098 541582 686334
rect 541026 650418 541262 650654
rect 541346 650418 541582 650654
rect 541026 650098 541262 650334
rect 541346 650098 541582 650334
rect 541026 614418 541262 614654
rect 541346 614418 541582 614654
rect 541026 614098 541262 614334
rect 541346 614098 541582 614334
rect 541026 578418 541262 578654
rect 541346 578418 541582 578654
rect 541026 578098 541262 578334
rect 541346 578098 541582 578334
rect 541026 542418 541262 542654
rect 541346 542418 541582 542654
rect 541026 542098 541262 542334
rect 541346 542098 541582 542334
rect 541026 506418 541262 506654
rect 541346 506418 541582 506654
rect 541026 506098 541262 506334
rect 541346 506098 541582 506334
rect 541026 470418 541262 470654
rect 541346 470418 541582 470654
rect 541026 470098 541262 470334
rect 541346 470098 541582 470334
rect 542266 705562 542502 705798
rect 542586 705562 542822 705798
rect 542266 705242 542502 705478
rect 542586 705242 542822 705478
rect 542266 687658 542502 687894
rect 542586 687658 542822 687894
rect 542266 687338 542502 687574
rect 542586 687338 542822 687574
rect 542266 651658 542502 651894
rect 542586 651658 542822 651894
rect 542266 651338 542502 651574
rect 542586 651338 542822 651574
rect 542266 615658 542502 615894
rect 542586 615658 542822 615894
rect 542266 615338 542502 615574
rect 542586 615338 542822 615574
rect 542266 579658 542502 579894
rect 542586 579658 542822 579894
rect 542266 579338 542502 579574
rect 542586 579338 542822 579574
rect 542266 543658 542502 543894
rect 542586 543658 542822 543894
rect 542266 543338 542502 543574
rect 542586 543338 542822 543574
rect 542266 507658 542502 507894
rect 542586 507658 542822 507894
rect 542266 507338 542502 507574
rect 542586 507338 542822 507574
rect 542266 471658 542502 471894
rect 542586 471658 542822 471894
rect 542266 471338 542502 471574
rect 542586 471338 542822 471574
rect 543506 706522 543742 706758
rect 543826 706522 544062 706758
rect 543506 706202 543742 706438
rect 543826 706202 544062 706438
rect 543506 688898 543742 689134
rect 543826 688898 544062 689134
rect 543506 688578 543742 688814
rect 543826 688578 544062 688814
rect 543506 652898 543742 653134
rect 543826 652898 544062 653134
rect 543506 652578 543742 652814
rect 543826 652578 544062 652814
rect 543506 616898 543742 617134
rect 543826 616898 544062 617134
rect 543506 616578 543742 616814
rect 543826 616578 544062 616814
rect 543506 580898 543742 581134
rect 543826 580898 544062 581134
rect 543506 580578 543742 580814
rect 543826 580578 544062 580814
rect 543506 544898 543742 545134
rect 543826 544898 544062 545134
rect 543506 544578 543742 544814
rect 543826 544578 544062 544814
rect 543506 508898 543742 509134
rect 543826 508898 544062 509134
rect 543506 508578 543742 508814
rect 543826 508578 544062 508814
rect 543506 472898 543742 473134
rect 543826 472898 544062 473134
rect 543506 472578 543742 472814
rect 543826 472578 544062 472814
rect 544746 707482 544982 707718
rect 545066 707482 545302 707718
rect 544746 707162 544982 707398
rect 545066 707162 545302 707398
rect 544746 690138 544982 690374
rect 545066 690138 545302 690374
rect 544746 689818 544982 690054
rect 545066 689818 545302 690054
rect 544746 654138 544982 654374
rect 545066 654138 545302 654374
rect 544746 653818 544982 654054
rect 545066 653818 545302 654054
rect 544746 618138 544982 618374
rect 545066 618138 545302 618374
rect 544746 617818 544982 618054
rect 545066 617818 545302 618054
rect 544746 582138 544982 582374
rect 545066 582138 545302 582374
rect 544746 581818 544982 582054
rect 545066 581818 545302 582054
rect 544746 546138 544982 546374
rect 545066 546138 545302 546374
rect 544746 545818 544982 546054
rect 545066 545818 545302 546054
rect 544746 510138 544982 510374
rect 545066 510138 545302 510374
rect 544746 509818 544982 510054
rect 545066 509818 545302 510054
rect 544746 474138 544982 474374
rect 545066 474138 545302 474374
rect 544746 473818 544982 474054
rect 545066 473818 545302 474054
rect 545986 708442 546222 708678
rect 546306 708442 546542 708678
rect 545986 708122 546222 708358
rect 546306 708122 546542 708358
rect 545986 691378 546222 691614
rect 546306 691378 546542 691614
rect 545986 691058 546222 691294
rect 546306 691058 546542 691294
rect 545986 655378 546222 655614
rect 546306 655378 546542 655614
rect 545986 655058 546222 655294
rect 546306 655058 546542 655294
rect 545986 619378 546222 619614
rect 546306 619378 546542 619614
rect 545986 619058 546222 619294
rect 546306 619058 546542 619294
rect 545986 583378 546222 583614
rect 546306 583378 546542 583614
rect 545986 583058 546222 583294
rect 546306 583058 546542 583294
rect 545986 547378 546222 547614
rect 546306 547378 546542 547614
rect 545986 547058 546222 547294
rect 546306 547058 546542 547294
rect 545986 511378 546222 511614
rect 546306 511378 546542 511614
rect 545986 511058 546222 511294
rect 546306 511058 546542 511294
rect 545986 475378 546222 475614
rect 546306 475378 546542 475614
rect 545986 475058 546222 475294
rect 546306 475058 546542 475294
rect 547226 709402 547462 709638
rect 547546 709402 547782 709638
rect 547226 709082 547462 709318
rect 547546 709082 547782 709318
rect 547226 692618 547462 692854
rect 547546 692618 547782 692854
rect 547226 692298 547462 692534
rect 547546 692298 547782 692534
rect 547226 656618 547462 656854
rect 547546 656618 547782 656854
rect 547226 656298 547462 656534
rect 547546 656298 547782 656534
rect 547226 620618 547462 620854
rect 547546 620618 547782 620854
rect 547226 620298 547462 620534
rect 547546 620298 547782 620534
rect 547226 584618 547462 584854
rect 547546 584618 547782 584854
rect 547226 584298 547462 584534
rect 547546 584298 547782 584534
rect 547226 548618 547462 548854
rect 547546 548618 547782 548854
rect 547226 548298 547462 548534
rect 547546 548298 547782 548534
rect 547226 512618 547462 512854
rect 547546 512618 547782 512854
rect 547226 512298 547462 512534
rect 547546 512298 547782 512534
rect 547226 476618 547462 476854
rect 547546 476618 547782 476854
rect 547226 476298 547462 476534
rect 547546 476298 547782 476534
rect 513706 443098 513942 443334
rect 514026 443098 514262 443334
rect 513706 442778 513942 443014
rect 514026 442778 514262 443014
rect 540918 435658 541154 435894
rect 540918 435338 541154 435574
rect 539952 434418 540188 434654
rect 539952 434098 540188 434334
rect 542850 435658 543086 435894
rect 542850 435338 543086 435574
rect 541884 434418 542120 434654
rect 541884 434098 542120 434334
rect 543816 434418 544052 434654
rect 543816 434098 544052 434334
rect 547226 440618 547462 440854
rect 547546 440618 547782 440854
rect 547226 440298 547462 440534
rect 547546 440298 547782 440534
rect 544782 435658 545018 435894
rect 544782 435338 545018 435574
rect 546714 435658 546950 435894
rect 546714 435338 546950 435574
rect 545748 434418 545984 434654
rect 545748 434098 545984 434334
rect 513706 407098 513942 407334
rect 514026 407098 514262 407334
rect 513706 406778 513942 407014
rect 514026 406778 514262 407014
rect 540918 399658 541154 399894
rect 540918 399338 541154 399574
rect 539952 398418 540188 398654
rect 539952 398098 540188 398334
rect 542850 399658 543086 399894
rect 542850 399338 543086 399574
rect 541884 398418 542120 398654
rect 541884 398098 542120 398334
rect 543816 398418 544052 398654
rect 543816 398098 544052 398334
rect 547226 404618 547462 404854
rect 547546 404618 547782 404854
rect 547226 404298 547462 404534
rect 547546 404298 547782 404534
rect 544782 399658 545018 399894
rect 544782 399338 545018 399574
rect 546714 399658 546950 399894
rect 546714 399338 546950 399574
rect 545748 398418 545984 398654
rect 545748 398098 545984 398334
rect 513706 371098 513942 371334
rect 514026 371098 514262 371334
rect 513706 370778 513942 371014
rect 514026 370778 514262 371014
rect 540918 363658 541154 363894
rect 540918 363338 541154 363574
rect 539952 362418 540188 362654
rect 539952 362098 540188 362334
rect 542850 363658 543086 363894
rect 542850 363338 543086 363574
rect 541884 362418 542120 362654
rect 541884 362098 542120 362334
rect 543816 362418 544052 362654
rect 543816 362098 544052 362334
rect 547226 368618 547462 368854
rect 547546 368618 547782 368854
rect 547226 368298 547462 368534
rect 547546 368298 547782 368534
rect 544782 363658 545018 363894
rect 544782 363338 545018 363574
rect 546714 363658 546950 363894
rect 546714 363338 546950 363574
rect 545748 362418 545984 362654
rect 545748 362098 545984 362334
rect 513706 335098 513942 335334
rect 514026 335098 514262 335334
rect 513706 334778 513942 335014
rect 514026 334778 514262 335014
rect 540918 327658 541154 327894
rect 540918 327338 541154 327574
rect 539952 326418 540188 326654
rect 539952 326098 540188 326334
rect 542850 327658 543086 327894
rect 542850 327338 543086 327574
rect 541884 326418 542120 326654
rect 541884 326098 542120 326334
rect 543816 326418 544052 326654
rect 543816 326098 544052 326334
rect 547226 332618 547462 332854
rect 547546 332618 547782 332854
rect 547226 332298 547462 332534
rect 547546 332298 547782 332534
rect 544782 327658 545018 327894
rect 544782 327338 545018 327574
rect 546714 327658 546950 327894
rect 546714 327338 546950 327574
rect 545748 326418 545984 326654
rect 545748 326098 545984 326334
rect 513706 299098 513942 299334
rect 514026 299098 514262 299334
rect 513706 298778 513942 299014
rect 514026 298778 514262 299014
rect 547226 296618 547462 296854
rect 547546 296618 547782 296854
rect 547226 296298 547462 296534
rect 547546 296298 547782 296534
rect 540918 291658 541154 291894
rect 540918 291338 541154 291574
rect 542850 291658 543086 291894
rect 542850 291338 543086 291574
rect 544782 291658 545018 291894
rect 544782 291338 545018 291574
rect 546714 291658 546950 291894
rect 546714 291338 546950 291574
rect 539952 290418 540188 290654
rect 539952 290098 540188 290334
rect 541884 290418 542120 290654
rect 541884 290098 542120 290334
rect 543816 290418 544052 290654
rect 543816 290098 544052 290334
rect 545748 290418 545984 290654
rect 545748 290098 545984 290334
rect 513706 263098 513942 263334
rect 514026 263098 514262 263334
rect 513706 262778 513942 263014
rect 514026 262778 514262 263014
rect 513706 227098 513942 227334
rect 514026 227098 514262 227334
rect 513706 226778 513942 227014
rect 514026 226778 514262 227014
rect 513706 191098 513942 191334
rect 514026 191098 514262 191334
rect 513706 190778 513942 191014
rect 514026 190778 514262 191014
rect 513706 155098 513942 155334
rect 514026 155098 514262 155334
rect 513706 154778 513942 155014
rect 514026 154778 514262 155014
rect 513706 119098 513942 119334
rect 514026 119098 514262 119334
rect 513706 118778 513942 119014
rect 514026 118778 514262 119014
rect 513706 83098 513942 83334
rect 514026 83098 514262 83334
rect 513706 82778 513942 83014
rect 514026 82778 514262 83014
rect 513706 47098 513942 47334
rect 514026 47098 514262 47334
rect 513706 46778 513942 47014
rect 514026 46778 514262 47014
rect 513706 11098 513942 11334
rect 514026 11098 514262 11334
rect 513706 10778 513942 11014
rect 514026 10778 514262 11014
rect 513706 -7302 513942 -7066
rect 514026 -7302 514262 -7066
rect 513706 -7622 513942 -7386
rect 514026 -7622 514262 -7386
rect 541026 254418 541262 254654
rect 541346 254418 541582 254654
rect 541026 254098 541262 254334
rect 541346 254098 541582 254334
rect 541026 218418 541262 218654
rect 541346 218418 541582 218654
rect 541026 218098 541262 218334
rect 541346 218098 541582 218334
rect 541026 182418 541262 182654
rect 541346 182418 541582 182654
rect 541026 182098 541262 182334
rect 541346 182098 541582 182334
rect 541026 146418 541262 146654
rect 541346 146418 541582 146654
rect 541026 146098 541262 146334
rect 541346 146098 541582 146334
rect 541026 110418 541262 110654
rect 541346 110418 541582 110654
rect 541026 110098 541262 110334
rect 541346 110098 541582 110334
rect 541026 74418 541262 74654
rect 541346 74418 541582 74654
rect 541026 74098 541262 74334
rect 541346 74098 541582 74334
rect 541026 38418 541262 38654
rect 541346 38418 541582 38654
rect 541026 38098 541262 38334
rect 541346 38098 541582 38334
rect 541026 2418 541262 2654
rect 541346 2418 541582 2654
rect 541026 2098 541262 2334
rect 541346 2098 541582 2334
rect 541026 -582 541262 -346
rect 541346 -582 541582 -346
rect 541026 -902 541262 -666
rect 541346 -902 541582 -666
rect 542266 255658 542502 255894
rect 542586 255658 542822 255894
rect 542266 255338 542502 255574
rect 542586 255338 542822 255574
rect 542266 219658 542502 219894
rect 542586 219658 542822 219894
rect 542266 219338 542502 219574
rect 542586 219338 542822 219574
rect 542266 183658 542502 183894
rect 542586 183658 542822 183894
rect 542266 183338 542502 183574
rect 542586 183338 542822 183574
rect 542266 147658 542502 147894
rect 542586 147658 542822 147894
rect 542266 147338 542502 147574
rect 542586 147338 542822 147574
rect 542266 111658 542502 111894
rect 542586 111658 542822 111894
rect 542266 111338 542502 111574
rect 542586 111338 542822 111574
rect 542266 75658 542502 75894
rect 542586 75658 542822 75894
rect 542266 75338 542502 75574
rect 542586 75338 542822 75574
rect 542266 39658 542502 39894
rect 542586 39658 542822 39894
rect 542266 39338 542502 39574
rect 542586 39338 542822 39574
rect 542266 3658 542502 3894
rect 542586 3658 542822 3894
rect 542266 3338 542502 3574
rect 542586 3338 542822 3574
rect 542266 -1542 542502 -1306
rect 542586 -1542 542822 -1306
rect 542266 -1862 542502 -1626
rect 542586 -1862 542822 -1626
rect 543506 256898 543742 257134
rect 543826 256898 544062 257134
rect 543506 256578 543742 256814
rect 543826 256578 544062 256814
rect 543506 220898 543742 221134
rect 543826 220898 544062 221134
rect 543506 220578 543742 220814
rect 543826 220578 544062 220814
rect 543506 184898 543742 185134
rect 543826 184898 544062 185134
rect 543506 184578 543742 184814
rect 543826 184578 544062 184814
rect 543506 148898 543742 149134
rect 543826 148898 544062 149134
rect 543506 148578 543742 148814
rect 543826 148578 544062 148814
rect 543506 112898 543742 113134
rect 543826 112898 544062 113134
rect 543506 112578 543742 112814
rect 543826 112578 544062 112814
rect 543506 76898 543742 77134
rect 543826 76898 544062 77134
rect 543506 76578 543742 76814
rect 543826 76578 544062 76814
rect 543506 40898 543742 41134
rect 543826 40898 544062 41134
rect 543506 40578 543742 40814
rect 543826 40578 544062 40814
rect 543506 4898 543742 5134
rect 543826 4898 544062 5134
rect 543506 4578 543742 4814
rect 543826 4578 544062 4814
rect 543506 -2502 543742 -2266
rect 543826 -2502 544062 -2266
rect 543506 -2822 543742 -2586
rect 543826 -2822 544062 -2586
rect 544746 258138 544982 258374
rect 545066 258138 545302 258374
rect 544746 257818 544982 258054
rect 545066 257818 545302 258054
rect 544746 222138 544982 222374
rect 545066 222138 545302 222374
rect 544746 221818 544982 222054
rect 545066 221818 545302 222054
rect 544746 186138 544982 186374
rect 545066 186138 545302 186374
rect 544746 185818 544982 186054
rect 545066 185818 545302 186054
rect 544746 150138 544982 150374
rect 545066 150138 545302 150374
rect 544746 149818 544982 150054
rect 545066 149818 545302 150054
rect 544746 114138 544982 114374
rect 545066 114138 545302 114374
rect 544746 113818 544982 114054
rect 545066 113818 545302 114054
rect 544746 78138 544982 78374
rect 545066 78138 545302 78374
rect 544746 77818 544982 78054
rect 545066 77818 545302 78054
rect 544746 42138 544982 42374
rect 545066 42138 545302 42374
rect 544746 41818 544982 42054
rect 545066 41818 545302 42054
rect 544746 6138 544982 6374
rect 545066 6138 545302 6374
rect 544746 5818 544982 6054
rect 545066 5818 545302 6054
rect 544746 -3462 544982 -3226
rect 545066 -3462 545302 -3226
rect 544746 -3782 544982 -3546
rect 545066 -3782 545302 -3546
rect 545986 259378 546222 259614
rect 546306 259378 546542 259614
rect 545986 259058 546222 259294
rect 546306 259058 546542 259294
rect 545986 223378 546222 223614
rect 546306 223378 546542 223614
rect 545986 223058 546222 223294
rect 546306 223058 546542 223294
rect 545986 187378 546222 187614
rect 546306 187378 546542 187614
rect 545986 187058 546222 187294
rect 546306 187058 546542 187294
rect 545986 151378 546222 151614
rect 546306 151378 546542 151614
rect 545986 151058 546222 151294
rect 546306 151058 546542 151294
rect 545986 115378 546222 115614
rect 546306 115378 546542 115614
rect 545986 115058 546222 115294
rect 546306 115058 546542 115294
rect 545986 79378 546222 79614
rect 546306 79378 546542 79614
rect 545986 79058 546222 79294
rect 546306 79058 546542 79294
rect 545986 43378 546222 43614
rect 546306 43378 546542 43614
rect 545986 43058 546222 43294
rect 546306 43058 546542 43294
rect 545986 7378 546222 7614
rect 546306 7378 546542 7614
rect 545986 7058 546222 7294
rect 546306 7058 546542 7294
rect 545986 -4422 546222 -4186
rect 546306 -4422 546542 -4186
rect 545986 -4742 546222 -4506
rect 546306 -4742 546542 -4506
rect 547226 260618 547462 260854
rect 547546 260618 547782 260854
rect 547226 260298 547462 260534
rect 547546 260298 547782 260534
rect 547226 224618 547462 224854
rect 547546 224618 547782 224854
rect 547226 224298 547462 224534
rect 547546 224298 547782 224534
rect 547226 188618 547462 188854
rect 547546 188618 547782 188854
rect 547226 188298 547462 188534
rect 547546 188298 547782 188534
rect 547226 152618 547462 152854
rect 547546 152618 547782 152854
rect 547226 152298 547462 152534
rect 547546 152298 547782 152534
rect 547226 116618 547462 116854
rect 547546 116618 547782 116854
rect 547226 116298 547462 116534
rect 547546 116298 547782 116534
rect 547226 80618 547462 80854
rect 547546 80618 547782 80854
rect 547226 80298 547462 80534
rect 547546 80298 547782 80534
rect 547226 44618 547462 44854
rect 547546 44618 547782 44854
rect 547226 44298 547462 44534
rect 547546 44298 547782 44534
rect 547226 8618 547462 8854
rect 547546 8618 547782 8854
rect 547226 8298 547462 8534
rect 547546 8298 547782 8534
rect 547226 -5382 547462 -5146
rect 547546 -5382 547782 -5146
rect 547226 -5702 547462 -5466
rect 547546 -5702 547782 -5466
rect 548466 710362 548702 710598
rect 548786 710362 549022 710598
rect 548466 710042 548702 710278
rect 548786 710042 549022 710278
rect 548466 693858 548702 694094
rect 548786 693858 549022 694094
rect 548466 693538 548702 693774
rect 548786 693538 549022 693774
rect 548466 657858 548702 658094
rect 548786 657858 549022 658094
rect 548466 657538 548702 657774
rect 548786 657538 549022 657774
rect 548466 621858 548702 622094
rect 548786 621858 549022 622094
rect 548466 621538 548702 621774
rect 548786 621538 549022 621774
rect 548466 585858 548702 586094
rect 548786 585858 549022 586094
rect 548466 585538 548702 585774
rect 548786 585538 549022 585774
rect 548466 549858 548702 550094
rect 548786 549858 549022 550094
rect 548466 549538 548702 549774
rect 548786 549538 549022 549774
rect 548466 513858 548702 514094
rect 548786 513858 549022 514094
rect 548466 513538 548702 513774
rect 548786 513538 549022 513774
rect 548466 477858 548702 478094
rect 548786 477858 549022 478094
rect 548466 477538 548702 477774
rect 548786 477538 549022 477774
rect 548466 441858 548702 442094
rect 548786 441858 549022 442094
rect 548466 441538 548702 441774
rect 548786 441538 549022 441774
rect 549706 711322 549942 711558
rect 550026 711322 550262 711558
rect 549706 711002 549942 711238
rect 550026 711002 550262 711238
rect 549706 695098 549942 695334
rect 550026 695098 550262 695334
rect 549706 694778 549942 695014
rect 550026 694778 550262 695014
rect 549706 659098 549942 659334
rect 550026 659098 550262 659334
rect 549706 658778 549942 659014
rect 550026 658778 550262 659014
rect 549706 623098 549942 623334
rect 550026 623098 550262 623334
rect 549706 622778 549942 623014
rect 550026 622778 550262 623014
rect 549706 587098 549942 587334
rect 550026 587098 550262 587334
rect 549706 586778 549942 587014
rect 550026 586778 550262 587014
rect 549706 551098 549942 551334
rect 550026 551098 550262 551334
rect 549706 550778 549942 551014
rect 550026 550778 550262 551014
rect 549706 515098 549942 515334
rect 550026 515098 550262 515334
rect 549706 514778 549942 515014
rect 550026 514778 550262 515014
rect 549706 479098 549942 479334
rect 550026 479098 550262 479334
rect 549706 478778 549942 479014
rect 550026 478778 550262 479014
rect 549706 443098 549942 443334
rect 550026 443098 550262 443334
rect 549706 442778 549942 443014
rect 550026 442778 550262 443014
rect 548466 405858 548702 406094
rect 548786 405858 549022 406094
rect 548466 405538 548702 405774
rect 548786 405538 549022 405774
rect 549706 407098 549942 407334
rect 550026 407098 550262 407334
rect 549706 406778 549942 407014
rect 550026 406778 550262 407014
rect 548466 369858 548702 370094
rect 548786 369858 549022 370094
rect 548466 369538 548702 369774
rect 548786 369538 549022 369774
rect 549706 371098 549942 371334
rect 550026 371098 550262 371334
rect 549706 370778 549942 371014
rect 550026 370778 550262 371014
rect 548466 333858 548702 334094
rect 548786 333858 549022 334094
rect 548466 333538 548702 333774
rect 548786 333538 549022 333774
rect 549706 335098 549942 335334
rect 550026 335098 550262 335334
rect 549706 334778 549942 335014
rect 550026 334778 550262 335014
rect 548466 297858 548702 298094
rect 548786 297858 549022 298094
rect 548466 297538 548702 297774
rect 548786 297538 549022 297774
rect 549706 299098 549942 299334
rect 550026 299098 550262 299334
rect 549706 298778 549942 299014
rect 550026 298778 550262 299014
rect 548466 261858 548702 262094
rect 548786 261858 549022 262094
rect 548466 261538 548702 261774
rect 548786 261538 549022 261774
rect 548466 225858 548702 226094
rect 548786 225858 549022 226094
rect 548466 225538 548702 225774
rect 548786 225538 549022 225774
rect 548466 189858 548702 190094
rect 548786 189858 549022 190094
rect 548466 189538 548702 189774
rect 548786 189538 549022 189774
rect 548466 153858 548702 154094
rect 548786 153858 549022 154094
rect 548466 153538 548702 153774
rect 548786 153538 549022 153774
rect 548466 117858 548702 118094
rect 548786 117858 549022 118094
rect 548466 117538 548702 117774
rect 548786 117538 549022 117774
rect 548466 81858 548702 82094
rect 548786 81858 549022 82094
rect 548466 81538 548702 81774
rect 548786 81538 549022 81774
rect 548466 45858 548702 46094
rect 548786 45858 549022 46094
rect 548466 45538 548702 45774
rect 548786 45538 549022 45774
rect 549706 263098 549942 263334
rect 550026 263098 550262 263334
rect 549706 262778 549942 263014
rect 550026 262778 550262 263014
rect 549706 227098 549942 227334
rect 550026 227098 550262 227334
rect 549706 226778 549942 227014
rect 550026 226778 550262 227014
rect 549706 191098 549942 191334
rect 550026 191098 550262 191334
rect 549706 190778 549942 191014
rect 550026 190778 550262 191014
rect 549706 155098 549942 155334
rect 550026 155098 550262 155334
rect 549706 154778 549942 155014
rect 550026 154778 550262 155014
rect 549706 119098 549942 119334
rect 550026 119098 550262 119334
rect 549706 118778 549942 119014
rect 550026 118778 550262 119014
rect 549706 83098 549942 83334
rect 550026 83098 550262 83334
rect 549706 82778 549942 83014
rect 550026 82778 550262 83014
rect 549706 47098 549942 47334
rect 550026 47098 550262 47334
rect 549706 46778 549942 47014
rect 550026 46778 550262 47014
rect 548466 9858 548702 10094
rect 548786 9858 549022 10094
rect 548466 9538 548702 9774
rect 548786 9538 549022 9774
rect 548466 -6342 548702 -6106
rect 548786 -6342 549022 -6106
rect 548466 -6662 548702 -6426
rect 548786 -6662 549022 -6426
rect 549706 11098 549942 11334
rect 550026 11098 550262 11334
rect 549706 10778 549942 11014
rect 550026 10778 550262 11014
rect 549706 -7302 549942 -7066
rect 550026 -7302 550262 -7066
rect 549706 -7622 549942 -7386
rect 550026 -7622 550262 -7386
rect 577026 704602 577262 704838
rect 577346 704602 577582 704838
rect 577026 704282 577262 704518
rect 577346 704282 577582 704518
rect 577026 686418 577262 686654
rect 577346 686418 577582 686654
rect 577026 686098 577262 686334
rect 577346 686098 577582 686334
rect 577026 650418 577262 650654
rect 577346 650418 577582 650654
rect 577026 650098 577262 650334
rect 577346 650098 577582 650334
rect 577026 614418 577262 614654
rect 577346 614418 577582 614654
rect 577026 614098 577262 614334
rect 577346 614098 577582 614334
rect 577026 578418 577262 578654
rect 577346 578418 577582 578654
rect 577026 578098 577262 578334
rect 577346 578098 577582 578334
rect 577026 542418 577262 542654
rect 577346 542418 577582 542654
rect 577026 542098 577262 542334
rect 577346 542098 577582 542334
rect 577026 506418 577262 506654
rect 577346 506418 577582 506654
rect 577026 506098 577262 506334
rect 577346 506098 577582 506334
rect 577026 470418 577262 470654
rect 577346 470418 577582 470654
rect 577026 470098 577262 470334
rect 577346 470098 577582 470334
rect 577026 434418 577262 434654
rect 577346 434418 577582 434654
rect 577026 434098 577262 434334
rect 577346 434098 577582 434334
rect 577026 398418 577262 398654
rect 577346 398418 577582 398654
rect 577026 398098 577262 398334
rect 577346 398098 577582 398334
rect 577026 362418 577262 362654
rect 577346 362418 577582 362654
rect 577026 362098 577262 362334
rect 577346 362098 577582 362334
rect 577026 326418 577262 326654
rect 577346 326418 577582 326654
rect 577026 326098 577262 326334
rect 577346 326098 577582 326334
rect 577026 290418 577262 290654
rect 577346 290418 577582 290654
rect 577026 290098 577262 290334
rect 577346 290098 577582 290334
rect 577026 254418 577262 254654
rect 577346 254418 577582 254654
rect 577026 254098 577262 254334
rect 577346 254098 577582 254334
rect 577026 218418 577262 218654
rect 577346 218418 577582 218654
rect 577026 218098 577262 218334
rect 577346 218098 577582 218334
rect 577026 182418 577262 182654
rect 577346 182418 577582 182654
rect 577026 182098 577262 182334
rect 577346 182098 577582 182334
rect 577026 146418 577262 146654
rect 577346 146418 577582 146654
rect 577026 146098 577262 146334
rect 577346 146098 577582 146334
rect 577026 110418 577262 110654
rect 577346 110418 577582 110654
rect 577026 110098 577262 110334
rect 577346 110098 577582 110334
rect 577026 74418 577262 74654
rect 577346 74418 577582 74654
rect 577026 74098 577262 74334
rect 577346 74098 577582 74334
rect 577026 38418 577262 38654
rect 577346 38418 577582 38654
rect 577026 38098 577262 38334
rect 577346 38098 577582 38334
rect 577026 2418 577262 2654
rect 577346 2418 577582 2654
rect 577026 2098 577262 2334
rect 577346 2098 577582 2334
rect 577026 -582 577262 -346
rect 577346 -582 577582 -346
rect 577026 -902 577262 -666
rect 577346 -902 577582 -666
rect 578266 705562 578502 705798
rect 578586 705562 578822 705798
rect 578266 705242 578502 705478
rect 578586 705242 578822 705478
rect 578266 687658 578502 687894
rect 578586 687658 578822 687894
rect 578266 687338 578502 687574
rect 578586 687338 578822 687574
rect 578266 651658 578502 651894
rect 578586 651658 578822 651894
rect 578266 651338 578502 651574
rect 578586 651338 578822 651574
rect 578266 615658 578502 615894
rect 578586 615658 578822 615894
rect 578266 615338 578502 615574
rect 578586 615338 578822 615574
rect 578266 579658 578502 579894
rect 578586 579658 578822 579894
rect 578266 579338 578502 579574
rect 578586 579338 578822 579574
rect 578266 543658 578502 543894
rect 578586 543658 578822 543894
rect 578266 543338 578502 543574
rect 578586 543338 578822 543574
rect 578266 507658 578502 507894
rect 578586 507658 578822 507894
rect 578266 507338 578502 507574
rect 578586 507338 578822 507574
rect 578266 471658 578502 471894
rect 578586 471658 578822 471894
rect 578266 471338 578502 471574
rect 578586 471338 578822 471574
rect 578266 435658 578502 435894
rect 578586 435658 578822 435894
rect 578266 435338 578502 435574
rect 578586 435338 578822 435574
rect 578266 399658 578502 399894
rect 578586 399658 578822 399894
rect 578266 399338 578502 399574
rect 578586 399338 578822 399574
rect 578266 363658 578502 363894
rect 578586 363658 578822 363894
rect 578266 363338 578502 363574
rect 578586 363338 578822 363574
rect 578266 327658 578502 327894
rect 578586 327658 578822 327894
rect 578266 327338 578502 327574
rect 578586 327338 578822 327574
rect 578266 291658 578502 291894
rect 578586 291658 578822 291894
rect 578266 291338 578502 291574
rect 578586 291338 578822 291574
rect 578266 255658 578502 255894
rect 578586 255658 578822 255894
rect 578266 255338 578502 255574
rect 578586 255338 578822 255574
rect 578266 219658 578502 219894
rect 578586 219658 578822 219894
rect 578266 219338 578502 219574
rect 578586 219338 578822 219574
rect 578266 183658 578502 183894
rect 578586 183658 578822 183894
rect 578266 183338 578502 183574
rect 578586 183338 578822 183574
rect 578266 147658 578502 147894
rect 578586 147658 578822 147894
rect 578266 147338 578502 147574
rect 578586 147338 578822 147574
rect 578266 111658 578502 111894
rect 578586 111658 578822 111894
rect 578266 111338 578502 111574
rect 578586 111338 578822 111574
rect 578266 75658 578502 75894
rect 578586 75658 578822 75894
rect 578266 75338 578502 75574
rect 578586 75338 578822 75574
rect 578266 39658 578502 39894
rect 578586 39658 578822 39894
rect 578266 39338 578502 39574
rect 578586 39338 578822 39574
rect 578266 3658 578502 3894
rect 578586 3658 578822 3894
rect 578266 3338 578502 3574
rect 578586 3338 578822 3574
rect 578266 -1542 578502 -1306
rect 578586 -1542 578822 -1306
rect 578266 -1862 578502 -1626
rect 578586 -1862 578822 -1626
rect 579506 706522 579742 706758
rect 579826 706522 580062 706758
rect 579506 706202 579742 706438
rect 579826 706202 580062 706438
rect 579506 688898 579742 689134
rect 579826 688898 580062 689134
rect 579506 688578 579742 688814
rect 579826 688578 580062 688814
rect 579506 652898 579742 653134
rect 579826 652898 580062 653134
rect 579506 652578 579742 652814
rect 579826 652578 580062 652814
rect 579506 616898 579742 617134
rect 579826 616898 580062 617134
rect 579506 616578 579742 616814
rect 579826 616578 580062 616814
rect 579506 580898 579742 581134
rect 579826 580898 580062 581134
rect 579506 580578 579742 580814
rect 579826 580578 580062 580814
rect 579506 544898 579742 545134
rect 579826 544898 580062 545134
rect 579506 544578 579742 544814
rect 579826 544578 580062 544814
rect 579506 508898 579742 509134
rect 579826 508898 580062 509134
rect 579506 508578 579742 508814
rect 579826 508578 580062 508814
rect 579506 472898 579742 473134
rect 579826 472898 580062 473134
rect 579506 472578 579742 472814
rect 579826 472578 580062 472814
rect 579506 436898 579742 437134
rect 579826 436898 580062 437134
rect 579506 436578 579742 436814
rect 579826 436578 580062 436814
rect 579506 400898 579742 401134
rect 579826 400898 580062 401134
rect 579506 400578 579742 400814
rect 579826 400578 580062 400814
rect 579506 364898 579742 365134
rect 579826 364898 580062 365134
rect 579506 364578 579742 364814
rect 579826 364578 580062 364814
rect 579506 328898 579742 329134
rect 579826 328898 580062 329134
rect 579506 328578 579742 328814
rect 579826 328578 580062 328814
rect 579506 292898 579742 293134
rect 579826 292898 580062 293134
rect 579506 292578 579742 292814
rect 579826 292578 580062 292814
rect 579506 256898 579742 257134
rect 579826 256898 580062 257134
rect 579506 256578 579742 256814
rect 579826 256578 580062 256814
rect 579506 220898 579742 221134
rect 579826 220898 580062 221134
rect 579506 220578 579742 220814
rect 579826 220578 580062 220814
rect 579506 184898 579742 185134
rect 579826 184898 580062 185134
rect 579506 184578 579742 184814
rect 579826 184578 580062 184814
rect 579506 148898 579742 149134
rect 579826 148898 580062 149134
rect 579506 148578 579742 148814
rect 579826 148578 580062 148814
rect 579506 112898 579742 113134
rect 579826 112898 580062 113134
rect 579506 112578 579742 112814
rect 579826 112578 580062 112814
rect 579506 76898 579742 77134
rect 579826 76898 580062 77134
rect 579506 76578 579742 76814
rect 579826 76578 580062 76814
rect 579506 40898 579742 41134
rect 579826 40898 580062 41134
rect 579506 40578 579742 40814
rect 579826 40578 580062 40814
rect 579506 4898 579742 5134
rect 579826 4898 580062 5134
rect 579506 4578 579742 4814
rect 579826 4578 580062 4814
rect 579506 -2502 579742 -2266
rect 579826 -2502 580062 -2266
rect 579506 -2822 579742 -2586
rect 579826 -2822 580062 -2586
rect 580746 707482 580982 707718
rect 581066 707482 581302 707718
rect 580746 707162 580982 707398
rect 581066 707162 581302 707398
rect 580746 690138 580982 690374
rect 581066 690138 581302 690374
rect 580746 689818 580982 690054
rect 581066 689818 581302 690054
rect 580746 654138 580982 654374
rect 581066 654138 581302 654374
rect 580746 653818 580982 654054
rect 581066 653818 581302 654054
rect 580746 618138 580982 618374
rect 581066 618138 581302 618374
rect 580746 617818 580982 618054
rect 581066 617818 581302 618054
rect 580746 582138 580982 582374
rect 581066 582138 581302 582374
rect 580746 581818 580982 582054
rect 581066 581818 581302 582054
rect 580746 546138 580982 546374
rect 581066 546138 581302 546374
rect 580746 545818 580982 546054
rect 581066 545818 581302 546054
rect 580746 510138 580982 510374
rect 581066 510138 581302 510374
rect 580746 509818 580982 510054
rect 581066 509818 581302 510054
rect 580746 474138 580982 474374
rect 581066 474138 581302 474374
rect 580746 473818 580982 474054
rect 581066 473818 581302 474054
rect 580746 438138 580982 438374
rect 581066 438138 581302 438374
rect 580746 437818 580982 438054
rect 581066 437818 581302 438054
rect 580746 402138 580982 402374
rect 581066 402138 581302 402374
rect 580746 401818 580982 402054
rect 581066 401818 581302 402054
rect 580746 366138 580982 366374
rect 581066 366138 581302 366374
rect 580746 365818 580982 366054
rect 581066 365818 581302 366054
rect 580746 330138 580982 330374
rect 581066 330138 581302 330374
rect 580746 329818 580982 330054
rect 581066 329818 581302 330054
rect 580746 294138 580982 294374
rect 581066 294138 581302 294374
rect 580746 293818 580982 294054
rect 581066 293818 581302 294054
rect 580746 258138 580982 258374
rect 581066 258138 581302 258374
rect 580746 257818 580982 258054
rect 581066 257818 581302 258054
rect 580746 222138 580982 222374
rect 581066 222138 581302 222374
rect 580746 221818 580982 222054
rect 581066 221818 581302 222054
rect 580746 186138 580982 186374
rect 581066 186138 581302 186374
rect 580746 185818 580982 186054
rect 581066 185818 581302 186054
rect 580746 150138 580982 150374
rect 581066 150138 581302 150374
rect 580746 149818 580982 150054
rect 581066 149818 581302 150054
rect 580746 114138 580982 114374
rect 581066 114138 581302 114374
rect 580746 113818 580982 114054
rect 581066 113818 581302 114054
rect 580746 78138 580982 78374
rect 581066 78138 581302 78374
rect 580746 77818 580982 78054
rect 581066 77818 581302 78054
rect 580746 42138 580982 42374
rect 581066 42138 581302 42374
rect 580746 41818 580982 42054
rect 581066 41818 581302 42054
rect 580746 6138 580982 6374
rect 581066 6138 581302 6374
rect 580746 5818 580982 6054
rect 581066 5818 581302 6054
rect 580746 -3462 580982 -3226
rect 581066 -3462 581302 -3226
rect 580746 -3782 580982 -3546
rect 581066 -3782 581302 -3546
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 581986 708442 582222 708678
rect 582306 708442 582542 708678
rect 581986 708122 582222 708358
rect 582306 708122 582542 708358
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581986 691378 582222 691614
rect 582306 691378 582542 691614
rect 581986 691058 582222 691294
rect 582306 691058 582542 691294
rect 581986 655378 582222 655614
rect 582306 655378 582542 655614
rect 581986 655058 582222 655294
rect 582306 655058 582542 655294
rect 581986 619378 582222 619614
rect 582306 619378 582542 619614
rect 581986 619058 582222 619294
rect 582306 619058 582542 619294
rect 581986 583378 582222 583614
rect 582306 583378 582542 583614
rect 581986 583058 582222 583294
rect 582306 583058 582542 583294
rect 581986 547378 582222 547614
rect 582306 547378 582542 547614
rect 581986 547058 582222 547294
rect 582306 547058 582542 547294
rect 581986 511378 582222 511614
rect 582306 511378 582542 511614
rect 581986 511058 582222 511294
rect 582306 511058 582542 511294
rect 581986 475378 582222 475614
rect 582306 475378 582542 475614
rect 581986 475058 582222 475294
rect 582306 475058 582542 475294
rect 581986 439378 582222 439614
rect 582306 439378 582542 439614
rect 581986 439058 582222 439294
rect 582306 439058 582542 439294
rect 581986 403378 582222 403614
rect 582306 403378 582542 403614
rect 581986 403058 582222 403294
rect 582306 403058 582542 403294
rect 581986 367378 582222 367614
rect 582306 367378 582542 367614
rect 581986 367058 582222 367294
rect 582306 367058 582542 367294
rect 581986 331378 582222 331614
rect 582306 331378 582542 331614
rect 581986 331058 582222 331294
rect 582306 331058 582542 331294
rect 581986 295378 582222 295614
rect 582306 295378 582542 295614
rect 581986 295058 582222 295294
rect 582306 295058 582542 295294
rect 581986 259378 582222 259614
rect 582306 259378 582542 259614
rect 581986 259058 582222 259294
rect 582306 259058 582542 259294
rect 581986 223378 582222 223614
rect 582306 223378 582542 223614
rect 581986 223058 582222 223294
rect 582306 223058 582542 223294
rect 581986 187378 582222 187614
rect 582306 187378 582542 187614
rect 581986 187058 582222 187294
rect 582306 187058 582542 187294
rect 581986 151378 582222 151614
rect 582306 151378 582542 151614
rect 581986 151058 582222 151294
rect 582306 151058 582542 151294
rect 581986 115378 582222 115614
rect 582306 115378 582542 115614
rect 581986 115058 582222 115294
rect 582306 115058 582542 115294
rect 581986 79378 582222 79614
rect 582306 79378 582542 79614
rect 581986 79058 582222 79294
rect 582306 79058 582542 79294
rect 581986 43378 582222 43614
rect 582306 43378 582542 43614
rect 581986 43058 582222 43294
rect 582306 43058 582542 43294
rect 581986 7378 582222 7614
rect 582306 7378 582542 7614
rect 581986 7058 582222 7294
rect 582306 7058 582542 7294
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 686418 585578 686654
rect 585662 686418 585898 686654
rect 585342 686098 585578 686334
rect 585662 686098 585898 686334
rect 585342 650418 585578 650654
rect 585662 650418 585898 650654
rect 585342 650098 585578 650334
rect 585662 650098 585898 650334
rect 585342 614418 585578 614654
rect 585662 614418 585898 614654
rect 585342 614098 585578 614334
rect 585662 614098 585898 614334
rect 585342 578418 585578 578654
rect 585662 578418 585898 578654
rect 585342 578098 585578 578334
rect 585662 578098 585898 578334
rect 585342 542418 585578 542654
rect 585662 542418 585898 542654
rect 585342 542098 585578 542334
rect 585662 542098 585898 542334
rect 585342 506418 585578 506654
rect 585662 506418 585898 506654
rect 585342 506098 585578 506334
rect 585662 506098 585898 506334
rect 585342 470418 585578 470654
rect 585662 470418 585898 470654
rect 585342 470098 585578 470334
rect 585662 470098 585898 470334
rect 585342 434418 585578 434654
rect 585662 434418 585898 434654
rect 585342 434098 585578 434334
rect 585662 434098 585898 434334
rect 585342 398418 585578 398654
rect 585662 398418 585898 398654
rect 585342 398098 585578 398334
rect 585662 398098 585898 398334
rect 585342 362418 585578 362654
rect 585662 362418 585898 362654
rect 585342 362098 585578 362334
rect 585662 362098 585898 362334
rect 585342 326418 585578 326654
rect 585662 326418 585898 326654
rect 585342 326098 585578 326334
rect 585662 326098 585898 326334
rect 585342 290418 585578 290654
rect 585662 290418 585898 290654
rect 585342 290098 585578 290334
rect 585662 290098 585898 290334
rect 585342 254418 585578 254654
rect 585662 254418 585898 254654
rect 585342 254098 585578 254334
rect 585662 254098 585898 254334
rect 585342 218418 585578 218654
rect 585662 218418 585898 218654
rect 585342 218098 585578 218334
rect 585662 218098 585898 218334
rect 585342 182418 585578 182654
rect 585662 182418 585898 182654
rect 585342 182098 585578 182334
rect 585662 182098 585898 182334
rect 585342 146418 585578 146654
rect 585662 146418 585898 146654
rect 585342 146098 585578 146334
rect 585662 146098 585898 146334
rect 585342 110418 585578 110654
rect 585662 110418 585898 110654
rect 585342 110098 585578 110334
rect 585662 110098 585898 110334
rect 585342 74418 585578 74654
rect 585662 74418 585898 74654
rect 585342 74098 585578 74334
rect 585662 74098 585898 74334
rect 585342 38418 585578 38654
rect 585662 38418 585898 38654
rect 585342 38098 585578 38334
rect 585662 38098 585898 38334
rect 585342 2418 585578 2654
rect 585662 2418 585898 2654
rect 585342 2098 585578 2334
rect 585662 2098 585898 2334
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 687658 586538 687894
rect 586622 687658 586858 687894
rect 586302 687338 586538 687574
rect 586622 687338 586858 687574
rect 586302 651658 586538 651894
rect 586622 651658 586858 651894
rect 586302 651338 586538 651574
rect 586622 651338 586858 651574
rect 586302 615658 586538 615894
rect 586622 615658 586858 615894
rect 586302 615338 586538 615574
rect 586622 615338 586858 615574
rect 586302 579658 586538 579894
rect 586622 579658 586858 579894
rect 586302 579338 586538 579574
rect 586622 579338 586858 579574
rect 586302 543658 586538 543894
rect 586622 543658 586858 543894
rect 586302 543338 586538 543574
rect 586622 543338 586858 543574
rect 586302 507658 586538 507894
rect 586622 507658 586858 507894
rect 586302 507338 586538 507574
rect 586622 507338 586858 507574
rect 586302 471658 586538 471894
rect 586622 471658 586858 471894
rect 586302 471338 586538 471574
rect 586622 471338 586858 471574
rect 586302 435658 586538 435894
rect 586622 435658 586858 435894
rect 586302 435338 586538 435574
rect 586622 435338 586858 435574
rect 586302 399658 586538 399894
rect 586622 399658 586858 399894
rect 586302 399338 586538 399574
rect 586622 399338 586858 399574
rect 586302 363658 586538 363894
rect 586622 363658 586858 363894
rect 586302 363338 586538 363574
rect 586622 363338 586858 363574
rect 586302 327658 586538 327894
rect 586622 327658 586858 327894
rect 586302 327338 586538 327574
rect 586622 327338 586858 327574
rect 586302 291658 586538 291894
rect 586622 291658 586858 291894
rect 586302 291338 586538 291574
rect 586622 291338 586858 291574
rect 586302 255658 586538 255894
rect 586622 255658 586858 255894
rect 586302 255338 586538 255574
rect 586622 255338 586858 255574
rect 586302 219658 586538 219894
rect 586622 219658 586858 219894
rect 586302 219338 586538 219574
rect 586622 219338 586858 219574
rect 586302 183658 586538 183894
rect 586622 183658 586858 183894
rect 586302 183338 586538 183574
rect 586622 183338 586858 183574
rect 586302 147658 586538 147894
rect 586622 147658 586858 147894
rect 586302 147338 586538 147574
rect 586622 147338 586858 147574
rect 586302 111658 586538 111894
rect 586622 111658 586858 111894
rect 586302 111338 586538 111574
rect 586622 111338 586858 111574
rect 586302 75658 586538 75894
rect 586622 75658 586858 75894
rect 586302 75338 586538 75574
rect 586622 75338 586858 75574
rect 586302 39658 586538 39894
rect 586622 39658 586858 39894
rect 586302 39338 586538 39574
rect 586622 39338 586858 39574
rect 586302 3658 586538 3894
rect 586622 3658 586858 3894
rect 586302 3338 586538 3574
rect 586622 3338 586858 3574
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 688898 587498 689134
rect 587582 688898 587818 689134
rect 587262 688578 587498 688814
rect 587582 688578 587818 688814
rect 587262 652898 587498 653134
rect 587582 652898 587818 653134
rect 587262 652578 587498 652814
rect 587582 652578 587818 652814
rect 587262 616898 587498 617134
rect 587582 616898 587818 617134
rect 587262 616578 587498 616814
rect 587582 616578 587818 616814
rect 587262 580898 587498 581134
rect 587582 580898 587818 581134
rect 587262 580578 587498 580814
rect 587582 580578 587818 580814
rect 587262 544898 587498 545134
rect 587582 544898 587818 545134
rect 587262 544578 587498 544814
rect 587582 544578 587818 544814
rect 587262 508898 587498 509134
rect 587582 508898 587818 509134
rect 587262 508578 587498 508814
rect 587582 508578 587818 508814
rect 587262 472898 587498 473134
rect 587582 472898 587818 473134
rect 587262 472578 587498 472814
rect 587582 472578 587818 472814
rect 587262 436898 587498 437134
rect 587582 436898 587818 437134
rect 587262 436578 587498 436814
rect 587582 436578 587818 436814
rect 587262 400898 587498 401134
rect 587582 400898 587818 401134
rect 587262 400578 587498 400814
rect 587582 400578 587818 400814
rect 587262 364898 587498 365134
rect 587582 364898 587818 365134
rect 587262 364578 587498 364814
rect 587582 364578 587818 364814
rect 587262 328898 587498 329134
rect 587582 328898 587818 329134
rect 587262 328578 587498 328814
rect 587582 328578 587818 328814
rect 587262 292898 587498 293134
rect 587582 292898 587818 293134
rect 587262 292578 587498 292814
rect 587582 292578 587818 292814
rect 587262 256898 587498 257134
rect 587582 256898 587818 257134
rect 587262 256578 587498 256814
rect 587582 256578 587818 256814
rect 587262 220898 587498 221134
rect 587582 220898 587818 221134
rect 587262 220578 587498 220814
rect 587582 220578 587818 220814
rect 587262 184898 587498 185134
rect 587582 184898 587818 185134
rect 587262 184578 587498 184814
rect 587582 184578 587818 184814
rect 587262 148898 587498 149134
rect 587582 148898 587818 149134
rect 587262 148578 587498 148814
rect 587582 148578 587818 148814
rect 587262 112898 587498 113134
rect 587582 112898 587818 113134
rect 587262 112578 587498 112814
rect 587582 112578 587818 112814
rect 587262 76898 587498 77134
rect 587582 76898 587818 77134
rect 587262 76578 587498 76814
rect 587582 76578 587818 76814
rect 587262 40898 587498 41134
rect 587582 40898 587818 41134
rect 587262 40578 587498 40814
rect 587582 40578 587818 40814
rect 587262 4898 587498 5134
rect 587582 4898 587818 5134
rect 587262 4578 587498 4814
rect 587582 4578 587818 4814
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 690138 588458 690374
rect 588542 690138 588778 690374
rect 588222 689818 588458 690054
rect 588542 689818 588778 690054
rect 588222 654138 588458 654374
rect 588542 654138 588778 654374
rect 588222 653818 588458 654054
rect 588542 653818 588778 654054
rect 588222 618138 588458 618374
rect 588542 618138 588778 618374
rect 588222 617818 588458 618054
rect 588542 617818 588778 618054
rect 588222 582138 588458 582374
rect 588542 582138 588778 582374
rect 588222 581818 588458 582054
rect 588542 581818 588778 582054
rect 588222 546138 588458 546374
rect 588542 546138 588778 546374
rect 588222 545818 588458 546054
rect 588542 545818 588778 546054
rect 588222 510138 588458 510374
rect 588542 510138 588778 510374
rect 588222 509818 588458 510054
rect 588542 509818 588778 510054
rect 588222 474138 588458 474374
rect 588542 474138 588778 474374
rect 588222 473818 588458 474054
rect 588542 473818 588778 474054
rect 588222 438138 588458 438374
rect 588542 438138 588778 438374
rect 588222 437818 588458 438054
rect 588542 437818 588778 438054
rect 588222 402138 588458 402374
rect 588542 402138 588778 402374
rect 588222 401818 588458 402054
rect 588542 401818 588778 402054
rect 588222 366138 588458 366374
rect 588542 366138 588778 366374
rect 588222 365818 588458 366054
rect 588542 365818 588778 366054
rect 588222 330138 588458 330374
rect 588542 330138 588778 330374
rect 588222 329818 588458 330054
rect 588542 329818 588778 330054
rect 588222 294138 588458 294374
rect 588542 294138 588778 294374
rect 588222 293818 588458 294054
rect 588542 293818 588778 294054
rect 588222 258138 588458 258374
rect 588542 258138 588778 258374
rect 588222 257818 588458 258054
rect 588542 257818 588778 258054
rect 588222 222138 588458 222374
rect 588542 222138 588778 222374
rect 588222 221818 588458 222054
rect 588542 221818 588778 222054
rect 588222 186138 588458 186374
rect 588542 186138 588778 186374
rect 588222 185818 588458 186054
rect 588542 185818 588778 186054
rect 588222 150138 588458 150374
rect 588542 150138 588778 150374
rect 588222 149818 588458 150054
rect 588542 149818 588778 150054
rect 588222 114138 588458 114374
rect 588542 114138 588778 114374
rect 588222 113818 588458 114054
rect 588542 113818 588778 114054
rect 588222 78138 588458 78374
rect 588542 78138 588778 78374
rect 588222 77818 588458 78054
rect 588542 77818 588778 78054
rect 588222 42138 588458 42374
rect 588542 42138 588778 42374
rect 588222 41818 588458 42054
rect 588542 41818 588778 42054
rect 588222 6138 588458 6374
rect 588542 6138 588778 6374
rect 588222 5818 588458 6054
rect 588542 5818 588778 6054
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 691378 589418 691614
rect 589502 691378 589738 691614
rect 589182 691058 589418 691294
rect 589502 691058 589738 691294
rect 589182 655378 589418 655614
rect 589502 655378 589738 655614
rect 589182 655058 589418 655294
rect 589502 655058 589738 655294
rect 589182 619378 589418 619614
rect 589502 619378 589738 619614
rect 589182 619058 589418 619294
rect 589502 619058 589738 619294
rect 589182 583378 589418 583614
rect 589502 583378 589738 583614
rect 589182 583058 589418 583294
rect 589502 583058 589738 583294
rect 589182 547378 589418 547614
rect 589502 547378 589738 547614
rect 589182 547058 589418 547294
rect 589502 547058 589738 547294
rect 589182 511378 589418 511614
rect 589502 511378 589738 511614
rect 589182 511058 589418 511294
rect 589502 511058 589738 511294
rect 589182 475378 589418 475614
rect 589502 475378 589738 475614
rect 589182 475058 589418 475294
rect 589502 475058 589738 475294
rect 589182 439378 589418 439614
rect 589502 439378 589738 439614
rect 589182 439058 589418 439294
rect 589502 439058 589738 439294
rect 589182 403378 589418 403614
rect 589502 403378 589738 403614
rect 589182 403058 589418 403294
rect 589502 403058 589738 403294
rect 589182 367378 589418 367614
rect 589502 367378 589738 367614
rect 589182 367058 589418 367294
rect 589502 367058 589738 367294
rect 589182 331378 589418 331614
rect 589502 331378 589738 331614
rect 589182 331058 589418 331294
rect 589502 331058 589738 331294
rect 589182 295378 589418 295614
rect 589502 295378 589738 295614
rect 589182 295058 589418 295294
rect 589502 295058 589738 295294
rect 589182 259378 589418 259614
rect 589502 259378 589738 259614
rect 589182 259058 589418 259294
rect 589502 259058 589738 259294
rect 589182 223378 589418 223614
rect 589502 223378 589738 223614
rect 589182 223058 589418 223294
rect 589502 223058 589738 223294
rect 589182 187378 589418 187614
rect 589502 187378 589738 187614
rect 589182 187058 589418 187294
rect 589502 187058 589738 187294
rect 589182 151378 589418 151614
rect 589502 151378 589738 151614
rect 589182 151058 589418 151294
rect 589502 151058 589738 151294
rect 589182 115378 589418 115614
rect 589502 115378 589738 115614
rect 589182 115058 589418 115294
rect 589502 115058 589738 115294
rect 589182 79378 589418 79614
rect 589502 79378 589738 79614
rect 589182 79058 589418 79294
rect 589502 79058 589738 79294
rect 589182 43378 589418 43614
rect 589502 43378 589738 43614
rect 589182 43058 589418 43294
rect 589502 43058 589738 43294
rect 589182 7378 589418 7614
rect 589502 7378 589738 7614
rect 589182 7058 589418 7294
rect 589502 7058 589738 7294
rect 581986 -4422 582222 -4186
rect 582306 -4422 582542 -4186
rect 581986 -4742 582222 -4506
rect 582306 -4742 582542 -4506
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 692618 590378 692854
rect 590462 692618 590698 692854
rect 590142 692298 590378 692534
rect 590462 692298 590698 692534
rect 590142 656618 590378 656854
rect 590462 656618 590698 656854
rect 590142 656298 590378 656534
rect 590462 656298 590698 656534
rect 590142 620618 590378 620854
rect 590462 620618 590698 620854
rect 590142 620298 590378 620534
rect 590462 620298 590698 620534
rect 590142 584618 590378 584854
rect 590462 584618 590698 584854
rect 590142 584298 590378 584534
rect 590462 584298 590698 584534
rect 590142 548618 590378 548854
rect 590462 548618 590698 548854
rect 590142 548298 590378 548534
rect 590462 548298 590698 548534
rect 590142 512618 590378 512854
rect 590462 512618 590698 512854
rect 590142 512298 590378 512534
rect 590462 512298 590698 512534
rect 590142 476618 590378 476854
rect 590462 476618 590698 476854
rect 590142 476298 590378 476534
rect 590462 476298 590698 476534
rect 590142 440618 590378 440854
rect 590462 440618 590698 440854
rect 590142 440298 590378 440534
rect 590462 440298 590698 440534
rect 590142 404618 590378 404854
rect 590462 404618 590698 404854
rect 590142 404298 590378 404534
rect 590462 404298 590698 404534
rect 590142 368618 590378 368854
rect 590462 368618 590698 368854
rect 590142 368298 590378 368534
rect 590462 368298 590698 368534
rect 590142 332618 590378 332854
rect 590462 332618 590698 332854
rect 590142 332298 590378 332534
rect 590462 332298 590698 332534
rect 590142 296618 590378 296854
rect 590462 296618 590698 296854
rect 590142 296298 590378 296534
rect 590462 296298 590698 296534
rect 590142 260618 590378 260854
rect 590462 260618 590698 260854
rect 590142 260298 590378 260534
rect 590462 260298 590698 260534
rect 590142 224618 590378 224854
rect 590462 224618 590698 224854
rect 590142 224298 590378 224534
rect 590462 224298 590698 224534
rect 590142 188618 590378 188854
rect 590462 188618 590698 188854
rect 590142 188298 590378 188534
rect 590462 188298 590698 188534
rect 590142 152618 590378 152854
rect 590462 152618 590698 152854
rect 590142 152298 590378 152534
rect 590462 152298 590698 152534
rect 590142 116618 590378 116854
rect 590462 116618 590698 116854
rect 590142 116298 590378 116534
rect 590462 116298 590698 116534
rect 590142 80618 590378 80854
rect 590462 80618 590698 80854
rect 590142 80298 590378 80534
rect 590462 80298 590698 80534
rect 590142 44618 590378 44854
rect 590462 44618 590698 44854
rect 590142 44298 590378 44534
rect 590462 44298 590698 44534
rect 590142 8618 590378 8854
rect 590462 8618 590698 8854
rect 590142 8298 590378 8534
rect 590462 8298 590698 8534
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 693858 591338 694094
rect 591422 693858 591658 694094
rect 591102 693538 591338 693774
rect 591422 693538 591658 693774
rect 591102 657858 591338 658094
rect 591422 657858 591658 658094
rect 591102 657538 591338 657774
rect 591422 657538 591658 657774
rect 591102 621858 591338 622094
rect 591422 621858 591658 622094
rect 591102 621538 591338 621774
rect 591422 621538 591658 621774
rect 591102 585858 591338 586094
rect 591422 585858 591658 586094
rect 591102 585538 591338 585774
rect 591422 585538 591658 585774
rect 591102 549858 591338 550094
rect 591422 549858 591658 550094
rect 591102 549538 591338 549774
rect 591422 549538 591658 549774
rect 591102 513858 591338 514094
rect 591422 513858 591658 514094
rect 591102 513538 591338 513774
rect 591422 513538 591658 513774
rect 591102 477858 591338 478094
rect 591422 477858 591658 478094
rect 591102 477538 591338 477774
rect 591422 477538 591658 477774
rect 591102 441858 591338 442094
rect 591422 441858 591658 442094
rect 591102 441538 591338 441774
rect 591422 441538 591658 441774
rect 591102 405858 591338 406094
rect 591422 405858 591658 406094
rect 591102 405538 591338 405774
rect 591422 405538 591658 405774
rect 591102 369858 591338 370094
rect 591422 369858 591658 370094
rect 591102 369538 591338 369774
rect 591422 369538 591658 369774
rect 591102 333858 591338 334094
rect 591422 333858 591658 334094
rect 591102 333538 591338 333774
rect 591422 333538 591658 333774
rect 591102 297858 591338 298094
rect 591422 297858 591658 298094
rect 591102 297538 591338 297774
rect 591422 297538 591658 297774
rect 591102 261858 591338 262094
rect 591422 261858 591658 262094
rect 591102 261538 591338 261774
rect 591422 261538 591658 261774
rect 591102 225858 591338 226094
rect 591422 225858 591658 226094
rect 591102 225538 591338 225774
rect 591422 225538 591658 225774
rect 591102 189858 591338 190094
rect 591422 189858 591658 190094
rect 591102 189538 591338 189774
rect 591422 189538 591658 189774
rect 591102 153858 591338 154094
rect 591422 153858 591658 154094
rect 591102 153538 591338 153774
rect 591422 153538 591658 153774
rect 591102 117858 591338 118094
rect 591422 117858 591658 118094
rect 591102 117538 591338 117774
rect 591422 117538 591658 117774
rect 591102 81858 591338 82094
rect 591422 81858 591658 82094
rect 591102 81538 591338 81774
rect 591422 81538 591658 81774
rect 591102 45858 591338 46094
rect 591422 45858 591658 46094
rect 591102 45538 591338 45774
rect 591422 45538 591658 45774
rect 591102 9858 591338 10094
rect 591422 9858 591658 10094
rect 591102 9538 591338 9774
rect 591422 9538 591658 9774
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 695098 592298 695334
rect 592382 695098 592618 695334
rect 592062 694778 592298 695014
rect 592382 694778 592618 695014
rect 592062 659098 592298 659334
rect 592382 659098 592618 659334
rect 592062 658778 592298 659014
rect 592382 658778 592618 659014
rect 592062 623098 592298 623334
rect 592382 623098 592618 623334
rect 592062 622778 592298 623014
rect 592382 622778 592618 623014
rect 592062 587098 592298 587334
rect 592382 587098 592618 587334
rect 592062 586778 592298 587014
rect 592382 586778 592618 587014
rect 592062 551098 592298 551334
rect 592382 551098 592618 551334
rect 592062 550778 592298 551014
rect 592382 550778 592618 551014
rect 592062 515098 592298 515334
rect 592382 515098 592618 515334
rect 592062 514778 592298 515014
rect 592382 514778 592618 515014
rect 592062 479098 592298 479334
rect 592382 479098 592618 479334
rect 592062 478778 592298 479014
rect 592382 478778 592618 479014
rect 592062 443098 592298 443334
rect 592382 443098 592618 443334
rect 592062 442778 592298 443014
rect 592382 442778 592618 443014
rect 592062 407098 592298 407334
rect 592382 407098 592618 407334
rect 592062 406778 592298 407014
rect 592382 406778 592618 407014
rect 592062 371098 592298 371334
rect 592382 371098 592618 371334
rect 592062 370778 592298 371014
rect 592382 370778 592618 371014
rect 592062 335098 592298 335334
rect 592382 335098 592618 335334
rect 592062 334778 592298 335014
rect 592382 334778 592618 335014
rect 592062 299098 592298 299334
rect 592382 299098 592618 299334
rect 592062 298778 592298 299014
rect 592382 298778 592618 299014
rect 592062 263098 592298 263334
rect 592382 263098 592618 263334
rect 592062 262778 592298 263014
rect 592382 262778 592618 263014
rect 592062 227098 592298 227334
rect 592382 227098 592618 227334
rect 592062 226778 592298 227014
rect 592382 226778 592618 227014
rect 592062 191098 592298 191334
rect 592382 191098 592618 191334
rect 592062 190778 592298 191014
rect 592382 190778 592618 191014
rect 592062 155098 592298 155334
rect 592382 155098 592618 155334
rect 592062 154778 592298 155014
rect 592382 154778 592618 155014
rect 592062 119098 592298 119334
rect 592382 119098 592618 119334
rect 592062 118778 592298 119014
rect 592382 118778 592618 119014
rect 592062 83098 592298 83334
rect 592382 83098 592618 83334
rect 592062 82778 592298 83014
rect 592382 82778 592618 83014
rect 592062 47098 592298 47334
rect 592382 47098 592618 47334
rect 592062 46778 592298 47014
rect 592382 46778 592618 47014
rect 592062 11098 592298 11334
rect 592382 11098 592618 11334
rect 592062 10778 592298 11014
rect 592382 10778 592618 11014
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 9706 711558
rect 9942 711322 10026 711558
rect 10262 711322 45706 711558
rect 45942 711322 46026 711558
rect 46262 711322 81706 711558
rect 81942 711322 82026 711558
rect 82262 711322 117706 711558
rect 117942 711322 118026 711558
rect 118262 711322 153706 711558
rect 153942 711322 154026 711558
rect 154262 711322 189706 711558
rect 189942 711322 190026 711558
rect 190262 711322 225706 711558
rect 225942 711322 226026 711558
rect 226262 711322 261706 711558
rect 261942 711322 262026 711558
rect 262262 711322 297706 711558
rect 297942 711322 298026 711558
rect 298262 711322 333706 711558
rect 333942 711322 334026 711558
rect 334262 711322 369706 711558
rect 369942 711322 370026 711558
rect 370262 711322 405706 711558
rect 405942 711322 406026 711558
rect 406262 711322 441706 711558
rect 441942 711322 442026 711558
rect 442262 711322 477706 711558
rect 477942 711322 478026 711558
rect 478262 711322 513706 711558
rect 513942 711322 514026 711558
rect 514262 711322 549706 711558
rect 549942 711322 550026 711558
rect 550262 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 9706 711238
rect 9942 711002 10026 711238
rect 10262 711002 45706 711238
rect 45942 711002 46026 711238
rect 46262 711002 81706 711238
rect 81942 711002 82026 711238
rect 82262 711002 117706 711238
rect 117942 711002 118026 711238
rect 118262 711002 153706 711238
rect 153942 711002 154026 711238
rect 154262 711002 189706 711238
rect 189942 711002 190026 711238
rect 190262 711002 225706 711238
rect 225942 711002 226026 711238
rect 226262 711002 261706 711238
rect 261942 711002 262026 711238
rect 262262 711002 297706 711238
rect 297942 711002 298026 711238
rect 298262 711002 333706 711238
rect 333942 711002 334026 711238
rect 334262 711002 369706 711238
rect 369942 711002 370026 711238
rect 370262 711002 405706 711238
rect 405942 711002 406026 711238
rect 406262 711002 441706 711238
rect 441942 711002 442026 711238
rect 442262 711002 477706 711238
rect 477942 711002 478026 711238
rect 478262 711002 513706 711238
rect 513942 711002 514026 711238
rect 514262 711002 549706 711238
rect 549942 711002 550026 711238
rect 550262 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 8466 710598
rect 8702 710362 8786 710598
rect 9022 710362 44466 710598
rect 44702 710362 44786 710598
rect 45022 710362 80466 710598
rect 80702 710362 80786 710598
rect 81022 710362 116466 710598
rect 116702 710362 116786 710598
rect 117022 710362 152466 710598
rect 152702 710362 152786 710598
rect 153022 710362 188466 710598
rect 188702 710362 188786 710598
rect 189022 710362 224466 710598
rect 224702 710362 224786 710598
rect 225022 710362 260466 710598
rect 260702 710362 260786 710598
rect 261022 710362 296466 710598
rect 296702 710362 296786 710598
rect 297022 710362 332466 710598
rect 332702 710362 332786 710598
rect 333022 710362 368466 710598
rect 368702 710362 368786 710598
rect 369022 710362 404466 710598
rect 404702 710362 404786 710598
rect 405022 710362 440466 710598
rect 440702 710362 440786 710598
rect 441022 710362 476466 710598
rect 476702 710362 476786 710598
rect 477022 710362 512466 710598
rect 512702 710362 512786 710598
rect 513022 710362 548466 710598
rect 548702 710362 548786 710598
rect 549022 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 8466 710278
rect 8702 710042 8786 710278
rect 9022 710042 44466 710278
rect 44702 710042 44786 710278
rect 45022 710042 80466 710278
rect 80702 710042 80786 710278
rect 81022 710042 116466 710278
rect 116702 710042 116786 710278
rect 117022 710042 152466 710278
rect 152702 710042 152786 710278
rect 153022 710042 188466 710278
rect 188702 710042 188786 710278
rect 189022 710042 224466 710278
rect 224702 710042 224786 710278
rect 225022 710042 260466 710278
rect 260702 710042 260786 710278
rect 261022 710042 296466 710278
rect 296702 710042 296786 710278
rect 297022 710042 332466 710278
rect 332702 710042 332786 710278
rect 333022 710042 368466 710278
rect 368702 710042 368786 710278
rect 369022 710042 404466 710278
rect 404702 710042 404786 710278
rect 405022 710042 440466 710278
rect 440702 710042 440786 710278
rect 441022 710042 476466 710278
rect 476702 710042 476786 710278
rect 477022 710042 512466 710278
rect 512702 710042 512786 710278
rect 513022 710042 548466 710278
rect 548702 710042 548786 710278
rect 549022 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 7226 709638
rect 7462 709402 7546 709638
rect 7782 709402 43226 709638
rect 43462 709402 43546 709638
rect 43782 709402 79226 709638
rect 79462 709402 79546 709638
rect 79782 709402 115226 709638
rect 115462 709402 115546 709638
rect 115782 709402 151226 709638
rect 151462 709402 151546 709638
rect 151782 709402 187226 709638
rect 187462 709402 187546 709638
rect 187782 709402 223226 709638
rect 223462 709402 223546 709638
rect 223782 709402 259226 709638
rect 259462 709402 259546 709638
rect 259782 709402 295226 709638
rect 295462 709402 295546 709638
rect 295782 709402 331226 709638
rect 331462 709402 331546 709638
rect 331782 709402 367226 709638
rect 367462 709402 367546 709638
rect 367782 709402 403226 709638
rect 403462 709402 403546 709638
rect 403782 709402 439226 709638
rect 439462 709402 439546 709638
rect 439782 709402 475226 709638
rect 475462 709402 475546 709638
rect 475782 709402 511226 709638
rect 511462 709402 511546 709638
rect 511782 709402 547226 709638
rect 547462 709402 547546 709638
rect 547782 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 7226 709318
rect 7462 709082 7546 709318
rect 7782 709082 43226 709318
rect 43462 709082 43546 709318
rect 43782 709082 79226 709318
rect 79462 709082 79546 709318
rect 79782 709082 115226 709318
rect 115462 709082 115546 709318
rect 115782 709082 151226 709318
rect 151462 709082 151546 709318
rect 151782 709082 187226 709318
rect 187462 709082 187546 709318
rect 187782 709082 223226 709318
rect 223462 709082 223546 709318
rect 223782 709082 259226 709318
rect 259462 709082 259546 709318
rect 259782 709082 295226 709318
rect 295462 709082 295546 709318
rect 295782 709082 331226 709318
rect 331462 709082 331546 709318
rect 331782 709082 367226 709318
rect 367462 709082 367546 709318
rect 367782 709082 403226 709318
rect 403462 709082 403546 709318
rect 403782 709082 439226 709318
rect 439462 709082 439546 709318
rect 439782 709082 475226 709318
rect 475462 709082 475546 709318
rect 475782 709082 511226 709318
rect 511462 709082 511546 709318
rect 511782 709082 547226 709318
rect 547462 709082 547546 709318
rect 547782 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 5986 708678
rect 6222 708442 6306 708678
rect 6542 708442 41986 708678
rect 42222 708442 42306 708678
rect 42542 708442 77986 708678
rect 78222 708442 78306 708678
rect 78542 708442 113986 708678
rect 114222 708442 114306 708678
rect 114542 708442 149986 708678
rect 150222 708442 150306 708678
rect 150542 708442 185986 708678
rect 186222 708442 186306 708678
rect 186542 708442 221986 708678
rect 222222 708442 222306 708678
rect 222542 708442 257986 708678
rect 258222 708442 258306 708678
rect 258542 708442 293986 708678
rect 294222 708442 294306 708678
rect 294542 708442 329986 708678
rect 330222 708442 330306 708678
rect 330542 708442 365986 708678
rect 366222 708442 366306 708678
rect 366542 708442 401986 708678
rect 402222 708442 402306 708678
rect 402542 708442 437986 708678
rect 438222 708442 438306 708678
rect 438542 708442 473986 708678
rect 474222 708442 474306 708678
rect 474542 708442 509986 708678
rect 510222 708442 510306 708678
rect 510542 708442 545986 708678
rect 546222 708442 546306 708678
rect 546542 708442 581986 708678
rect 582222 708442 582306 708678
rect 582542 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 5986 708358
rect 6222 708122 6306 708358
rect 6542 708122 41986 708358
rect 42222 708122 42306 708358
rect 42542 708122 77986 708358
rect 78222 708122 78306 708358
rect 78542 708122 113986 708358
rect 114222 708122 114306 708358
rect 114542 708122 149986 708358
rect 150222 708122 150306 708358
rect 150542 708122 185986 708358
rect 186222 708122 186306 708358
rect 186542 708122 221986 708358
rect 222222 708122 222306 708358
rect 222542 708122 257986 708358
rect 258222 708122 258306 708358
rect 258542 708122 293986 708358
rect 294222 708122 294306 708358
rect 294542 708122 329986 708358
rect 330222 708122 330306 708358
rect 330542 708122 365986 708358
rect 366222 708122 366306 708358
rect 366542 708122 401986 708358
rect 402222 708122 402306 708358
rect 402542 708122 437986 708358
rect 438222 708122 438306 708358
rect 438542 708122 473986 708358
rect 474222 708122 474306 708358
rect 474542 708122 509986 708358
rect 510222 708122 510306 708358
rect 510542 708122 545986 708358
rect 546222 708122 546306 708358
rect 546542 708122 581986 708358
rect 582222 708122 582306 708358
rect 582542 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 4746 707718
rect 4982 707482 5066 707718
rect 5302 707482 40746 707718
rect 40982 707482 41066 707718
rect 41302 707482 76746 707718
rect 76982 707482 77066 707718
rect 77302 707482 112746 707718
rect 112982 707482 113066 707718
rect 113302 707482 148746 707718
rect 148982 707482 149066 707718
rect 149302 707482 184746 707718
rect 184982 707482 185066 707718
rect 185302 707482 220746 707718
rect 220982 707482 221066 707718
rect 221302 707482 256746 707718
rect 256982 707482 257066 707718
rect 257302 707482 292746 707718
rect 292982 707482 293066 707718
rect 293302 707482 328746 707718
rect 328982 707482 329066 707718
rect 329302 707482 364746 707718
rect 364982 707482 365066 707718
rect 365302 707482 400746 707718
rect 400982 707482 401066 707718
rect 401302 707482 436746 707718
rect 436982 707482 437066 707718
rect 437302 707482 472746 707718
rect 472982 707482 473066 707718
rect 473302 707482 508746 707718
rect 508982 707482 509066 707718
rect 509302 707482 544746 707718
rect 544982 707482 545066 707718
rect 545302 707482 580746 707718
rect 580982 707482 581066 707718
rect 581302 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 4746 707398
rect 4982 707162 5066 707398
rect 5302 707162 40746 707398
rect 40982 707162 41066 707398
rect 41302 707162 76746 707398
rect 76982 707162 77066 707398
rect 77302 707162 112746 707398
rect 112982 707162 113066 707398
rect 113302 707162 148746 707398
rect 148982 707162 149066 707398
rect 149302 707162 184746 707398
rect 184982 707162 185066 707398
rect 185302 707162 220746 707398
rect 220982 707162 221066 707398
rect 221302 707162 256746 707398
rect 256982 707162 257066 707398
rect 257302 707162 292746 707398
rect 292982 707162 293066 707398
rect 293302 707162 328746 707398
rect 328982 707162 329066 707398
rect 329302 707162 364746 707398
rect 364982 707162 365066 707398
rect 365302 707162 400746 707398
rect 400982 707162 401066 707398
rect 401302 707162 436746 707398
rect 436982 707162 437066 707398
rect 437302 707162 472746 707398
rect 472982 707162 473066 707398
rect 473302 707162 508746 707398
rect 508982 707162 509066 707398
rect 509302 707162 544746 707398
rect 544982 707162 545066 707398
rect 545302 707162 580746 707398
rect 580982 707162 581066 707398
rect 581302 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 3506 706758
rect 3742 706522 3826 706758
rect 4062 706522 39506 706758
rect 39742 706522 39826 706758
rect 40062 706522 75506 706758
rect 75742 706522 75826 706758
rect 76062 706522 111506 706758
rect 111742 706522 111826 706758
rect 112062 706522 147506 706758
rect 147742 706522 147826 706758
rect 148062 706522 183506 706758
rect 183742 706522 183826 706758
rect 184062 706522 219506 706758
rect 219742 706522 219826 706758
rect 220062 706522 255506 706758
rect 255742 706522 255826 706758
rect 256062 706522 291506 706758
rect 291742 706522 291826 706758
rect 292062 706522 327506 706758
rect 327742 706522 327826 706758
rect 328062 706522 363506 706758
rect 363742 706522 363826 706758
rect 364062 706522 399506 706758
rect 399742 706522 399826 706758
rect 400062 706522 435506 706758
rect 435742 706522 435826 706758
rect 436062 706522 471506 706758
rect 471742 706522 471826 706758
rect 472062 706522 507506 706758
rect 507742 706522 507826 706758
rect 508062 706522 543506 706758
rect 543742 706522 543826 706758
rect 544062 706522 579506 706758
rect 579742 706522 579826 706758
rect 580062 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 3506 706438
rect 3742 706202 3826 706438
rect 4062 706202 39506 706438
rect 39742 706202 39826 706438
rect 40062 706202 75506 706438
rect 75742 706202 75826 706438
rect 76062 706202 111506 706438
rect 111742 706202 111826 706438
rect 112062 706202 147506 706438
rect 147742 706202 147826 706438
rect 148062 706202 183506 706438
rect 183742 706202 183826 706438
rect 184062 706202 219506 706438
rect 219742 706202 219826 706438
rect 220062 706202 255506 706438
rect 255742 706202 255826 706438
rect 256062 706202 291506 706438
rect 291742 706202 291826 706438
rect 292062 706202 327506 706438
rect 327742 706202 327826 706438
rect 328062 706202 363506 706438
rect 363742 706202 363826 706438
rect 364062 706202 399506 706438
rect 399742 706202 399826 706438
rect 400062 706202 435506 706438
rect 435742 706202 435826 706438
rect 436062 706202 471506 706438
rect 471742 706202 471826 706438
rect 472062 706202 507506 706438
rect 507742 706202 507826 706438
rect 508062 706202 543506 706438
rect 543742 706202 543826 706438
rect 544062 706202 579506 706438
rect 579742 706202 579826 706438
rect 580062 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 2266 705798
rect 2502 705562 2586 705798
rect 2822 705562 38266 705798
rect 38502 705562 38586 705798
rect 38822 705562 74266 705798
rect 74502 705562 74586 705798
rect 74822 705562 110266 705798
rect 110502 705562 110586 705798
rect 110822 705562 146266 705798
rect 146502 705562 146586 705798
rect 146822 705562 182266 705798
rect 182502 705562 182586 705798
rect 182822 705562 218266 705798
rect 218502 705562 218586 705798
rect 218822 705562 254266 705798
rect 254502 705562 254586 705798
rect 254822 705562 290266 705798
rect 290502 705562 290586 705798
rect 290822 705562 326266 705798
rect 326502 705562 326586 705798
rect 326822 705562 362266 705798
rect 362502 705562 362586 705798
rect 362822 705562 398266 705798
rect 398502 705562 398586 705798
rect 398822 705562 434266 705798
rect 434502 705562 434586 705798
rect 434822 705562 470266 705798
rect 470502 705562 470586 705798
rect 470822 705562 506266 705798
rect 506502 705562 506586 705798
rect 506822 705562 542266 705798
rect 542502 705562 542586 705798
rect 542822 705562 578266 705798
rect 578502 705562 578586 705798
rect 578822 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 2266 705478
rect 2502 705242 2586 705478
rect 2822 705242 38266 705478
rect 38502 705242 38586 705478
rect 38822 705242 74266 705478
rect 74502 705242 74586 705478
rect 74822 705242 110266 705478
rect 110502 705242 110586 705478
rect 110822 705242 146266 705478
rect 146502 705242 146586 705478
rect 146822 705242 182266 705478
rect 182502 705242 182586 705478
rect 182822 705242 218266 705478
rect 218502 705242 218586 705478
rect 218822 705242 254266 705478
rect 254502 705242 254586 705478
rect 254822 705242 290266 705478
rect 290502 705242 290586 705478
rect 290822 705242 326266 705478
rect 326502 705242 326586 705478
rect 326822 705242 362266 705478
rect 362502 705242 362586 705478
rect 362822 705242 398266 705478
rect 398502 705242 398586 705478
rect 398822 705242 434266 705478
rect 434502 705242 434586 705478
rect 434822 705242 470266 705478
rect 470502 705242 470586 705478
rect 470822 705242 506266 705478
rect 506502 705242 506586 705478
rect 506822 705242 542266 705478
rect 542502 705242 542586 705478
rect 542822 705242 578266 705478
rect 578502 705242 578586 705478
rect 578822 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1026 704838
rect 1262 704602 1346 704838
rect 1582 704602 37026 704838
rect 37262 704602 37346 704838
rect 37582 704602 73026 704838
rect 73262 704602 73346 704838
rect 73582 704602 109026 704838
rect 109262 704602 109346 704838
rect 109582 704602 145026 704838
rect 145262 704602 145346 704838
rect 145582 704602 181026 704838
rect 181262 704602 181346 704838
rect 181582 704602 217026 704838
rect 217262 704602 217346 704838
rect 217582 704602 253026 704838
rect 253262 704602 253346 704838
rect 253582 704602 289026 704838
rect 289262 704602 289346 704838
rect 289582 704602 325026 704838
rect 325262 704602 325346 704838
rect 325582 704602 361026 704838
rect 361262 704602 361346 704838
rect 361582 704602 397026 704838
rect 397262 704602 397346 704838
rect 397582 704602 433026 704838
rect 433262 704602 433346 704838
rect 433582 704602 469026 704838
rect 469262 704602 469346 704838
rect 469582 704602 505026 704838
rect 505262 704602 505346 704838
rect 505582 704602 541026 704838
rect 541262 704602 541346 704838
rect 541582 704602 577026 704838
rect 577262 704602 577346 704838
rect 577582 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1026 704518
rect 1262 704282 1346 704518
rect 1582 704282 37026 704518
rect 37262 704282 37346 704518
rect 37582 704282 73026 704518
rect 73262 704282 73346 704518
rect 73582 704282 109026 704518
rect 109262 704282 109346 704518
rect 109582 704282 145026 704518
rect 145262 704282 145346 704518
rect 145582 704282 181026 704518
rect 181262 704282 181346 704518
rect 181582 704282 217026 704518
rect 217262 704282 217346 704518
rect 217582 704282 253026 704518
rect 253262 704282 253346 704518
rect 253582 704282 289026 704518
rect 289262 704282 289346 704518
rect 289582 704282 325026 704518
rect 325262 704282 325346 704518
rect 325582 704282 361026 704518
rect 361262 704282 361346 704518
rect 361582 704282 397026 704518
rect 397262 704282 397346 704518
rect 397582 704282 433026 704518
rect 433262 704282 433346 704518
rect 433582 704282 469026 704518
rect 469262 704282 469346 704518
rect 469582 704282 505026 704518
rect 505262 704282 505346 704518
rect 505582 704282 541026 704518
rect 541262 704282 541346 704518
rect 541582 704282 577026 704518
rect 577262 704282 577346 704518
rect 577582 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 695334 592650 695366
rect -8726 695098 -8694 695334
rect -8458 695098 -8374 695334
rect -8138 695098 9706 695334
rect 9942 695098 10026 695334
rect 10262 695098 45706 695334
rect 45942 695098 46026 695334
rect 46262 695098 81706 695334
rect 81942 695098 82026 695334
rect 82262 695098 117706 695334
rect 117942 695098 118026 695334
rect 118262 695098 153706 695334
rect 153942 695098 154026 695334
rect 154262 695098 189706 695334
rect 189942 695098 190026 695334
rect 190262 695098 225706 695334
rect 225942 695098 226026 695334
rect 226262 695098 261706 695334
rect 261942 695098 262026 695334
rect 262262 695098 297706 695334
rect 297942 695098 298026 695334
rect 298262 695098 333706 695334
rect 333942 695098 334026 695334
rect 334262 695098 369706 695334
rect 369942 695098 370026 695334
rect 370262 695098 405706 695334
rect 405942 695098 406026 695334
rect 406262 695098 441706 695334
rect 441942 695098 442026 695334
rect 442262 695098 477706 695334
rect 477942 695098 478026 695334
rect 478262 695098 513706 695334
rect 513942 695098 514026 695334
rect 514262 695098 549706 695334
rect 549942 695098 550026 695334
rect 550262 695098 592062 695334
rect 592298 695098 592382 695334
rect 592618 695098 592650 695334
rect -8726 695014 592650 695098
rect -8726 694778 -8694 695014
rect -8458 694778 -8374 695014
rect -8138 694778 9706 695014
rect 9942 694778 10026 695014
rect 10262 694778 45706 695014
rect 45942 694778 46026 695014
rect 46262 694778 81706 695014
rect 81942 694778 82026 695014
rect 82262 694778 117706 695014
rect 117942 694778 118026 695014
rect 118262 694778 153706 695014
rect 153942 694778 154026 695014
rect 154262 694778 189706 695014
rect 189942 694778 190026 695014
rect 190262 694778 225706 695014
rect 225942 694778 226026 695014
rect 226262 694778 261706 695014
rect 261942 694778 262026 695014
rect 262262 694778 297706 695014
rect 297942 694778 298026 695014
rect 298262 694778 333706 695014
rect 333942 694778 334026 695014
rect 334262 694778 369706 695014
rect 369942 694778 370026 695014
rect 370262 694778 405706 695014
rect 405942 694778 406026 695014
rect 406262 694778 441706 695014
rect 441942 694778 442026 695014
rect 442262 694778 477706 695014
rect 477942 694778 478026 695014
rect 478262 694778 513706 695014
rect 513942 694778 514026 695014
rect 514262 694778 549706 695014
rect 549942 694778 550026 695014
rect 550262 694778 592062 695014
rect 592298 694778 592382 695014
rect 592618 694778 592650 695014
rect -8726 694746 592650 694778
rect -8726 694094 592650 694126
rect -8726 693858 -7734 694094
rect -7498 693858 -7414 694094
rect -7178 693858 8466 694094
rect 8702 693858 8786 694094
rect 9022 693858 44466 694094
rect 44702 693858 44786 694094
rect 45022 693858 80466 694094
rect 80702 693858 80786 694094
rect 81022 693858 116466 694094
rect 116702 693858 116786 694094
rect 117022 693858 152466 694094
rect 152702 693858 152786 694094
rect 153022 693858 188466 694094
rect 188702 693858 188786 694094
rect 189022 693858 224466 694094
rect 224702 693858 224786 694094
rect 225022 693858 260466 694094
rect 260702 693858 260786 694094
rect 261022 693858 296466 694094
rect 296702 693858 296786 694094
rect 297022 693858 332466 694094
rect 332702 693858 332786 694094
rect 333022 693858 368466 694094
rect 368702 693858 368786 694094
rect 369022 693858 404466 694094
rect 404702 693858 404786 694094
rect 405022 693858 440466 694094
rect 440702 693858 440786 694094
rect 441022 693858 476466 694094
rect 476702 693858 476786 694094
rect 477022 693858 512466 694094
rect 512702 693858 512786 694094
rect 513022 693858 548466 694094
rect 548702 693858 548786 694094
rect 549022 693858 591102 694094
rect 591338 693858 591422 694094
rect 591658 693858 592650 694094
rect -8726 693774 592650 693858
rect -8726 693538 -7734 693774
rect -7498 693538 -7414 693774
rect -7178 693538 8466 693774
rect 8702 693538 8786 693774
rect 9022 693538 44466 693774
rect 44702 693538 44786 693774
rect 45022 693538 80466 693774
rect 80702 693538 80786 693774
rect 81022 693538 116466 693774
rect 116702 693538 116786 693774
rect 117022 693538 152466 693774
rect 152702 693538 152786 693774
rect 153022 693538 188466 693774
rect 188702 693538 188786 693774
rect 189022 693538 224466 693774
rect 224702 693538 224786 693774
rect 225022 693538 260466 693774
rect 260702 693538 260786 693774
rect 261022 693538 296466 693774
rect 296702 693538 296786 693774
rect 297022 693538 332466 693774
rect 332702 693538 332786 693774
rect 333022 693538 368466 693774
rect 368702 693538 368786 693774
rect 369022 693538 404466 693774
rect 404702 693538 404786 693774
rect 405022 693538 440466 693774
rect 440702 693538 440786 693774
rect 441022 693538 476466 693774
rect 476702 693538 476786 693774
rect 477022 693538 512466 693774
rect 512702 693538 512786 693774
rect 513022 693538 548466 693774
rect 548702 693538 548786 693774
rect 549022 693538 591102 693774
rect 591338 693538 591422 693774
rect 591658 693538 592650 693774
rect -8726 693506 592650 693538
rect -8726 692854 592650 692886
rect -8726 692618 -6774 692854
rect -6538 692618 -6454 692854
rect -6218 692618 7226 692854
rect 7462 692618 7546 692854
rect 7782 692618 43226 692854
rect 43462 692618 43546 692854
rect 43782 692618 79226 692854
rect 79462 692618 79546 692854
rect 79782 692618 115226 692854
rect 115462 692618 115546 692854
rect 115782 692618 151226 692854
rect 151462 692618 151546 692854
rect 151782 692618 187226 692854
rect 187462 692618 187546 692854
rect 187782 692618 223226 692854
rect 223462 692618 223546 692854
rect 223782 692618 259226 692854
rect 259462 692618 259546 692854
rect 259782 692618 295226 692854
rect 295462 692618 295546 692854
rect 295782 692618 331226 692854
rect 331462 692618 331546 692854
rect 331782 692618 367226 692854
rect 367462 692618 367546 692854
rect 367782 692618 403226 692854
rect 403462 692618 403546 692854
rect 403782 692618 439226 692854
rect 439462 692618 439546 692854
rect 439782 692618 475226 692854
rect 475462 692618 475546 692854
rect 475782 692618 511226 692854
rect 511462 692618 511546 692854
rect 511782 692618 547226 692854
rect 547462 692618 547546 692854
rect 547782 692618 590142 692854
rect 590378 692618 590462 692854
rect 590698 692618 592650 692854
rect -8726 692534 592650 692618
rect -8726 692298 -6774 692534
rect -6538 692298 -6454 692534
rect -6218 692298 7226 692534
rect 7462 692298 7546 692534
rect 7782 692298 43226 692534
rect 43462 692298 43546 692534
rect 43782 692298 79226 692534
rect 79462 692298 79546 692534
rect 79782 692298 115226 692534
rect 115462 692298 115546 692534
rect 115782 692298 151226 692534
rect 151462 692298 151546 692534
rect 151782 692298 187226 692534
rect 187462 692298 187546 692534
rect 187782 692298 223226 692534
rect 223462 692298 223546 692534
rect 223782 692298 259226 692534
rect 259462 692298 259546 692534
rect 259782 692298 295226 692534
rect 295462 692298 295546 692534
rect 295782 692298 331226 692534
rect 331462 692298 331546 692534
rect 331782 692298 367226 692534
rect 367462 692298 367546 692534
rect 367782 692298 403226 692534
rect 403462 692298 403546 692534
rect 403782 692298 439226 692534
rect 439462 692298 439546 692534
rect 439782 692298 475226 692534
rect 475462 692298 475546 692534
rect 475782 692298 511226 692534
rect 511462 692298 511546 692534
rect 511782 692298 547226 692534
rect 547462 692298 547546 692534
rect 547782 692298 590142 692534
rect 590378 692298 590462 692534
rect 590698 692298 592650 692534
rect -8726 692266 592650 692298
rect -8726 691614 592650 691646
rect -8726 691378 -5814 691614
rect -5578 691378 -5494 691614
rect -5258 691378 5986 691614
rect 6222 691378 6306 691614
rect 6542 691378 41986 691614
rect 42222 691378 42306 691614
rect 42542 691378 77986 691614
rect 78222 691378 78306 691614
rect 78542 691378 113986 691614
rect 114222 691378 114306 691614
rect 114542 691378 149986 691614
rect 150222 691378 150306 691614
rect 150542 691378 185986 691614
rect 186222 691378 186306 691614
rect 186542 691378 221986 691614
rect 222222 691378 222306 691614
rect 222542 691378 257986 691614
rect 258222 691378 258306 691614
rect 258542 691378 293986 691614
rect 294222 691378 294306 691614
rect 294542 691378 329986 691614
rect 330222 691378 330306 691614
rect 330542 691378 365986 691614
rect 366222 691378 366306 691614
rect 366542 691378 401986 691614
rect 402222 691378 402306 691614
rect 402542 691378 437986 691614
rect 438222 691378 438306 691614
rect 438542 691378 473986 691614
rect 474222 691378 474306 691614
rect 474542 691378 509986 691614
rect 510222 691378 510306 691614
rect 510542 691378 545986 691614
rect 546222 691378 546306 691614
rect 546542 691378 581986 691614
rect 582222 691378 582306 691614
rect 582542 691378 589182 691614
rect 589418 691378 589502 691614
rect 589738 691378 592650 691614
rect -8726 691294 592650 691378
rect -8726 691058 -5814 691294
rect -5578 691058 -5494 691294
rect -5258 691058 5986 691294
rect 6222 691058 6306 691294
rect 6542 691058 41986 691294
rect 42222 691058 42306 691294
rect 42542 691058 77986 691294
rect 78222 691058 78306 691294
rect 78542 691058 113986 691294
rect 114222 691058 114306 691294
rect 114542 691058 149986 691294
rect 150222 691058 150306 691294
rect 150542 691058 185986 691294
rect 186222 691058 186306 691294
rect 186542 691058 221986 691294
rect 222222 691058 222306 691294
rect 222542 691058 257986 691294
rect 258222 691058 258306 691294
rect 258542 691058 293986 691294
rect 294222 691058 294306 691294
rect 294542 691058 329986 691294
rect 330222 691058 330306 691294
rect 330542 691058 365986 691294
rect 366222 691058 366306 691294
rect 366542 691058 401986 691294
rect 402222 691058 402306 691294
rect 402542 691058 437986 691294
rect 438222 691058 438306 691294
rect 438542 691058 473986 691294
rect 474222 691058 474306 691294
rect 474542 691058 509986 691294
rect 510222 691058 510306 691294
rect 510542 691058 545986 691294
rect 546222 691058 546306 691294
rect 546542 691058 581986 691294
rect 582222 691058 582306 691294
rect 582542 691058 589182 691294
rect 589418 691058 589502 691294
rect 589738 691058 592650 691294
rect -8726 691026 592650 691058
rect -8726 690374 592650 690406
rect -8726 690138 -4854 690374
rect -4618 690138 -4534 690374
rect -4298 690138 4746 690374
rect 4982 690138 5066 690374
rect 5302 690138 40746 690374
rect 40982 690138 41066 690374
rect 41302 690138 76746 690374
rect 76982 690138 77066 690374
rect 77302 690138 112746 690374
rect 112982 690138 113066 690374
rect 113302 690138 148746 690374
rect 148982 690138 149066 690374
rect 149302 690138 184746 690374
rect 184982 690138 185066 690374
rect 185302 690138 220746 690374
rect 220982 690138 221066 690374
rect 221302 690138 256746 690374
rect 256982 690138 257066 690374
rect 257302 690138 292746 690374
rect 292982 690138 293066 690374
rect 293302 690138 328746 690374
rect 328982 690138 329066 690374
rect 329302 690138 364746 690374
rect 364982 690138 365066 690374
rect 365302 690138 400746 690374
rect 400982 690138 401066 690374
rect 401302 690138 436746 690374
rect 436982 690138 437066 690374
rect 437302 690138 472746 690374
rect 472982 690138 473066 690374
rect 473302 690138 508746 690374
rect 508982 690138 509066 690374
rect 509302 690138 544746 690374
rect 544982 690138 545066 690374
rect 545302 690138 580746 690374
rect 580982 690138 581066 690374
rect 581302 690138 588222 690374
rect 588458 690138 588542 690374
rect 588778 690138 592650 690374
rect -8726 690054 592650 690138
rect -8726 689818 -4854 690054
rect -4618 689818 -4534 690054
rect -4298 689818 4746 690054
rect 4982 689818 5066 690054
rect 5302 689818 40746 690054
rect 40982 689818 41066 690054
rect 41302 689818 76746 690054
rect 76982 689818 77066 690054
rect 77302 689818 112746 690054
rect 112982 689818 113066 690054
rect 113302 689818 148746 690054
rect 148982 689818 149066 690054
rect 149302 689818 184746 690054
rect 184982 689818 185066 690054
rect 185302 689818 220746 690054
rect 220982 689818 221066 690054
rect 221302 689818 256746 690054
rect 256982 689818 257066 690054
rect 257302 689818 292746 690054
rect 292982 689818 293066 690054
rect 293302 689818 328746 690054
rect 328982 689818 329066 690054
rect 329302 689818 364746 690054
rect 364982 689818 365066 690054
rect 365302 689818 400746 690054
rect 400982 689818 401066 690054
rect 401302 689818 436746 690054
rect 436982 689818 437066 690054
rect 437302 689818 472746 690054
rect 472982 689818 473066 690054
rect 473302 689818 508746 690054
rect 508982 689818 509066 690054
rect 509302 689818 544746 690054
rect 544982 689818 545066 690054
rect 545302 689818 580746 690054
rect 580982 689818 581066 690054
rect 581302 689818 588222 690054
rect 588458 689818 588542 690054
rect 588778 689818 592650 690054
rect -8726 689786 592650 689818
rect -8726 689134 592650 689166
rect -8726 688898 -3894 689134
rect -3658 688898 -3574 689134
rect -3338 688898 3506 689134
rect 3742 688898 3826 689134
rect 4062 688898 39506 689134
rect 39742 688898 39826 689134
rect 40062 688898 75506 689134
rect 75742 688898 75826 689134
rect 76062 688898 111506 689134
rect 111742 688898 111826 689134
rect 112062 688898 147506 689134
rect 147742 688898 147826 689134
rect 148062 688898 183506 689134
rect 183742 688898 183826 689134
rect 184062 688898 219506 689134
rect 219742 688898 219826 689134
rect 220062 688898 255506 689134
rect 255742 688898 255826 689134
rect 256062 688898 291506 689134
rect 291742 688898 291826 689134
rect 292062 688898 327506 689134
rect 327742 688898 327826 689134
rect 328062 688898 363506 689134
rect 363742 688898 363826 689134
rect 364062 688898 399506 689134
rect 399742 688898 399826 689134
rect 400062 688898 435506 689134
rect 435742 688898 435826 689134
rect 436062 688898 471506 689134
rect 471742 688898 471826 689134
rect 472062 688898 507506 689134
rect 507742 688898 507826 689134
rect 508062 688898 543506 689134
rect 543742 688898 543826 689134
rect 544062 688898 579506 689134
rect 579742 688898 579826 689134
rect 580062 688898 587262 689134
rect 587498 688898 587582 689134
rect 587818 688898 592650 689134
rect -8726 688814 592650 688898
rect -8726 688578 -3894 688814
rect -3658 688578 -3574 688814
rect -3338 688578 3506 688814
rect 3742 688578 3826 688814
rect 4062 688578 39506 688814
rect 39742 688578 39826 688814
rect 40062 688578 75506 688814
rect 75742 688578 75826 688814
rect 76062 688578 111506 688814
rect 111742 688578 111826 688814
rect 112062 688578 147506 688814
rect 147742 688578 147826 688814
rect 148062 688578 183506 688814
rect 183742 688578 183826 688814
rect 184062 688578 219506 688814
rect 219742 688578 219826 688814
rect 220062 688578 255506 688814
rect 255742 688578 255826 688814
rect 256062 688578 291506 688814
rect 291742 688578 291826 688814
rect 292062 688578 327506 688814
rect 327742 688578 327826 688814
rect 328062 688578 363506 688814
rect 363742 688578 363826 688814
rect 364062 688578 399506 688814
rect 399742 688578 399826 688814
rect 400062 688578 435506 688814
rect 435742 688578 435826 688814
rect 436062 688578 471506 688814
rect 471742 688578 471826 688814
rect 472062 688578 507506 688814
rect 507742 688578 507826 688814
rect 508062 688578 543506 688814
rect 543742 688578 543826 688814
rect 544062 688578 579506 688814
rect 579742 688578 579826 688814
rect 580062 688578 587262 688814
rect 587498 688578 587582 688814
rect 587818 688578 592650 688814
rect -8726 688546 592650 688578
rect -8726 687894 592650 687926
rect -8726 687658 -2934 687894
rect -2698 687658 -2614 687894
rect -2378 687658 2266 687894
rect 2502 687658 2586 687894
rect 2822 687658 38266 687894
rect 38502 687658 38586 687894
rect 38822 687658 74266 687894
rect 74502 687658 74586 687894
rect 74822 687658 110266 687894
rect 110502 687658 110586 687894
rect 110822 687658 146266 687894
rect 146502 687658 146586 687894
rect 146822 687658 182266 687894
rect 182502 687658 182586 687894
rect 182822 687658 218266 687894
rect 218502 687658 218586 687894
rect 218822 687658 254266 687894
rect 254502 687658 254586 687894
rect 254822 687658 290266 687894
rect 290502 687658 290586 687894
rect 290822 687658 326266 687894
rect 326502 687658 326586 687894
rect 326822 687658 362266 687894
rect 362502 687658 362586 687894
rect 362822 687658 398266 687894
rect 398502 687658 398586 687894
rect 398822 687658 434266 687894
rect 434502 687658 434586 687894
rect 434822 687658 470266 687894
rect 470502 687658 470586 687894
rect 470822 687658 506266 687894
rect 506502 687658 506586 687894
rect 506822 687658 542266 687894
rect 542502 687658 542586 687894
rect 542822 687658 578266 687894
rect 578502 687658 578586 687894
rect 578822 687658 586302 687894
rect 586538 687658 586622 687894
rect 586858 687658 592650 687894
rect -8726 687574 592650 687658
rect -8726 687338 -2934 687574
rect -2698 687338 -2614 687574
rect -2378 687338 2266 687574
rect 2502 687338 2586 687574
rect 2822 687338 38266 687574
rect 38502 687338 38586 687574
rect 38822 687338 74266 687574
rect 74502 687338 74586 687574
rect 74822 687338 110266 687574
rect 110502 687338 110586 687574
rect 110822 687338 146266 687574
rect 146502 687338 146586 687574
rect 146822 687338 182266 687574
rect 182502 687338 182586 687574
rect 182822 687338 218266 687574
rect 218502 687338 218586 687574
rect 218822 687338 254266 687574
rect 254502 687338 254586 687574
rect 254822 687338 290266 687574
rect 290502 687338 290586 687574
rect 290822 687338 326266 687574
rect 326502 687338 326586 687574
rect 326822 687338 362266 687574
rect 362502 687338 362586 687574
rect 362822 687338 398266 687574
rect 398502 687338 398586 687574
rect 398822 687338 434266 687574
rect 434502 687338 434586 687574
rect 434822 687338 470266 687574
rect 470502 687338 470586 687574
rect 470822 687338 506266 687574
rect 506502 687338 506586 687574
rect 506822 687338 542266 687574
rect 542502 687338 542586 687574
rect 542822 687338 578266 687574
rect 578502 687338 578586 687574
rect 578822 687338 586302 687574
rect 586538 687338 586622 687574
rect 586858 687338 592650 687574
rect -8726 687306 592650 687338
rect -8726 686654 592650 686686
rect -8726 686418 -1974 686654
rect -1738 686418 -1654 686654
rect -1418 686418 1026 686654
rect 1262 686418 1346 686654
rect 1582 686418 37026 686654
rect 37262 686418 37346 686654
rect 37582 686418 73026 686654
rect 73262 686418 73346 686654
rect 73582 686418 109026 686654
rect 109262 686418 109346 686654
rect 109582 686418 145026 686654
rect 145262 686418 145346 686654
rect 145582 686418 181026 686654
rect 181262 686418 181346 686654
rect 181582 686418 217026 686654
rect 217262 686418 217346 686654
rect 217582 686418 253026 686654
rect 253262 686418 253346 686654
rect 253582 686418 289026 686654
rect 289262 686418 289346 686654
rect 289582 686418 325026 686654
rect 325262 686418 325346 686654
rect 325582 686418 361026 686654
rect 361262 686418 361346 686654
rect 361582 686418 397026 686654
rect 397262 686418 397346 686654
rect 397582 686418 433026 686654
rect 433262 686418 433346 686654
rect 433582 686418 469026 686654
rect 469262 686418 469346 686654
rect 469582 686418 505026 686654
rect 505262 686418 505346 686654
rect 505582 686418 541026 686654
rect 541262 686418 541346 686654
rect 541582 686418 577026 686654
rect 577262 686418 577346 686654
rect 577582 686418 585342 686654
rect 585578 686418 585662 686654
rect 585898 686418 592650 686654
rect -8726 686334 592650 686418
rect -8726 686098 -1974 686334
rect -1738 686098 -1654 686334
rect -1418 686098 1026 686334
rect 1262 686098 1346 686334
rect 1582 686098 37026 686334
rect 37262 686098 37346 686334
rect 37582 686098 73026 686334
rect 73262 686098 73346 686334
rect 73582 686098 109026 686334
rect 109262 686098 109346 686334
rect 109582 686098 145026 686334
rect 145262 686098 145346 686334
rect 145582 686098 181026 686334
rect 181262 686098 181346 686334
rect 181582 686098 217026 686334
rect 217262 686098 217346 686334
rect 217582 686098 253026 686334
rect 253262 686098 253346 686334
rect 253582 686098 289026 686334
rect 289262 686098 289346 686334
rect 289582 686098 325026 686334
rect 325262 686098 325346 686334
rect 325582 686098 361026 686334
rect 361262 686098 361346 686334
rect 361582 686098 397026 686334
rect 397262 686098 397346 686334
rect 397582 686098 433026 686334
rect 433262 686098 433346 686334
rect 433582 686098 469026 686334
rect 469262 686098 469346 686334
rect 469582 686098 505026 686334
rect 505262 686098 505346 686334
rect 505582 686098 541026 686334
rect 541262 686098 541346 686334
rect 541582 686098 577026 686334
rect 577262 686098 577346 686334
rect 577582 686098 585342 686334
rect 585578 686098 585662 686334
rect 585898 686098 592650 686334
rect -8726 686066 592650 686098
rect -8726 659334 592650 659366
rect -8726 659098 -8694 659334
rect -8458 659098 -8374 659334
rect -8138 659098 9706 659334
rect 9942 659098 10026 659334
rect 10262 659098 45706 659334
rect 45942 659098 46026 659334
rect 46262 659098 81706 659334
rect 81942 659098 82026 659334
rect 82262 659098 117706 659334
rect 117942 659098 118026 659334
rect 118262 659098 153706 659334
rect 153942 659098 154026 659334
rect 154262 659098 189706 659334
rect 189942 659098 190026 659334
rect 190262 659098 225706 659334
rect 225942 659098 226026 659334
rect 226262 659098 261706 659334
rect 261942 659098 262026 659334
rect 262262 659098 297706 659334
rect 297942 659098 298026 659334
rect 298262 659098 333706 659334
rect 333942 659098 334026 659334
rect 334262 659098 369706 659334
rect 369942 659098 370026 659334
rect 370262 659098 405706 659334
rect 405942 659098 406026 659334
rect 406262 659098 441706 659334
rect 441942 659098 442026 659334
rect 442262 659098 477706 659334
rect 477942 659098 478026 659334
rect 478262 659098 513706 659334
rect 513942 659098 514026 659334
rect 514262 659098 549706 659334
rect 549942 659098 550026 659334
rect 550262 659098 592062 659334
rect 592298 659098 592382 659334
rect 592618 659098 592650 659334
rect -8726 659014 592650 659098
rect -8726 658778 -8694 659014
rect -8458 658778 -8374 659014
rect -8138 658778 9706 659014
rect 9942 658778 10026 659014
rect 10262 658778 45706 659014
rect 45942 658778 46026 659014
rect 46262 658778 81706 659014
rect 81942 658778 82026 659014
rect 82262 658778 117706 659014
rect 117942 658778 118026 659014
rect 118262 658778 153706 659014
rect 153942 658778 154026 659014
rect 154262 658778 189706 659014
rect 189942 658778 190026 659014
rect 190262 658778 225706 659014
rect 225942 658778 226026 659014
rect 226262 658778 261706 659014
rect 261942 658778 262026 659014
rect 262262 658778 297706 659014
rect 297942 658778 298026 659014
rect 298262 658778 333706 659014
rect 333942 658778 334026 659014
rect 334262 658778 369706 659014
rect 369942 658778 370026 659014
rect 370262 658778 405706 659014
rect 405942 658778 406026 659014
rect 406262 658778 441706 659014
rect 441942 658778 442026 659014
rect 442262 658778 477706 659014
rect 477942 658778 478026 659014
rect 478262 658778 513706 659014
rect 513942 658778 514026 659014
rect 514262 658778 549706 659014
rect 549942 658778 550026 659014
rect 550262 658778 592062 659014
rect 592298 658778 592382 659014
rect 592618 658778 592650 659014
rect -8726 658746 592650 658778
rect -8726 658094 592650 658126
rect -8726 657858 -7734 658094
rect -7498 657858 -7414 658094
rect -7178 657858 8466 658094
rect 8702 657858 8786 658094
rect 9022 657858 44466 658094
rect 44702 657858 44786 658094
rect 45022 657858 80466 658094
rect 80702 657858 80786 658094
rect 81022 657858 116466 658094
rect 116702 657858 116786 658094
rect 117022 657858 152466 658094
rect 152702 657858 152786 658094
rect 153022 657858 188466 658094
rect 188702 657858 188786 658094
rect 189022 657858 224466 658094
rect 224702 657858 224786 658094
rect 225022 657858 260466 658094
rect 260702 657858 260786 658094
rect 261022 657858 296466 658094
rect 296702 657858 296786 658094
rect 297022 657858 332466 658094
rect 332702 657858 332786 658094
rect 333022 657858 368466 658094
rect 368702 657858 368786 658094
rect 369022 657858 404466 658094
rect 404702 657858 404786 658094
rect 405022 657858 440466 658094
rect 440702 657858 440786 658094
rect 441022 657858 476466 658094
rect 476702 657858 476786 658094
rect 477022 657858 512466 658094
rect 512702 657858 512786 658094
rect 513022 657858 548466 658094
rect 548702 657858 548786 658094
rect 549022 657858 591102 658094
rect 591338 657858 591422 658094
rect 591658 657858 592650 658094
rect -8726 657774 592650 657858
rect -8726 657538 -7734 657774
rect -7498 657538 -7414 657774
rect -7178 657538 8466 657774
rect 8702 657538 8786 657774
rect 9022 657538 44466 657774
rect 44702 657538 44786 657774
rect 45022 657538 80466 657774
rect 80702 657538 80786 657774
rect 81022 657538 116466 657774
rect 116702 657538 116786 657774
rect 117022 657538 152466 657774
rect 152702 657538 152786 657774
rect 153022 657538 188466 657774
rect 188702 657538 188786 657774
rect 189022 657538 224466 657774
rect 224702 657538 224786 657774
rect 225022 657538 260466 657774
rect 260702 657538 260786 657774
rect 261022 657538 296466 657774
rect 296702 657538 296786 657774
rect 297022 657538 332466 657774
rect 332702 657538 332786 657774
rect 333022 657538 368466 657774
rect 368702 657538 368786 657774
rect 369022 657538 404466 657774
rect 404702 657538 404786 657774
rect 405022 657538 440466 657774
rect 440702 657538 440786 657774
rect 441022 657538 476466 657774
rect 476702 657538 476786 657774
rect 477022 657538 512466 657774
rect 512702 657538 512786 657774
rect 513022 657538 548466 657774
rect 548702 657538 548786 657774
rect 549022 657538 591102 657774
rect 591338 657538 591422 657774
rect 591658 657538 592650 657774
rect -8726 657506 592650 657538
rect -8726 656854 592650 656886
rect -8726 656618 -6774 656854
rect -6538 656618 -6454 656854
rect -6218 656618 7226 656854
rect 7462 656618 7546 656854
rect 7782 656618 43226 656854
rect 43462 656618 43546 656854
rect 43782 656618 79226 656854
rect 79462 656618 79546 656854
rect 79782 656618 115226 656854
rect 115462 656618 115546 656854
rect 115782 656618 151226 656854
rect 151462 656618 151546 656854
rect 151782 656618 187226 656854
rect 187462 656618 187546 656854
rect 187782 656618 223226 656854
rect 223462 656618 223546 656854
rect 223782 656618 259226 656854
rect 259462 656618 259546 656854
rect 259782 656618 295226 656854
rect 295462 656618 295546 656854
rect 295782 656618 331226 656854
rect 331462 656618 331546 656854
rect 331782 656618 367226 656854
rect 367462 656618 367546 656854
rect 367782 656618 403226 656854
rect 403462 656618 403546 656854
rect 403782 656618 439226 656854
rect 439462 656618 439546 656854
rect 439782 656618 475226 656854
rect 475462 656618 475546 656854
rect 475782 656618 511226 656854
rect 511462 656618 511546 656854
rect 511782 656618 547226 656854
rect 547462 656618 547546 656854
rect 547782 656618 590142 656854
rect 590378 656618 590462 656854
rect 590698 656618 592650 656854
rect -8726 656534 592650 656618
rect -8726 656298 -6774 656534
rect -6538 656298 -6454 656534
rect -6218 656298 7226 656534
rect 7462 656298 7546 656534
rect 7782 656298 43226 656534
rect 43462 656298 43546 656534
rect 43782 656298 79226 656534
rect 79462 656298 79546 656534
rect 79782 656298 115226 656534
rect 115462 656298 115546 656534
rect 115782 656298 151226 656534
rect 151462 656298 151546 656534
rect 151782 656298 187226 656534
rect 187462 656298 187546 656534
rect 187782 656298 223226 656534
rect 223462 656298 223546 656534
rect 223782 656298 259226 656534
rect 259462 656298 259546 656534
rect 259782 656298 295226 656534
rect 295462 656298 295546 656534
rect 295782 656298 331226 656534
rect 331462 656298 331546 656534
rect 331782 656298 367226 656534
rect 367462 656298 367546 656534
rect 367782 656298 403226 656534
rect 403462 656298 403546 656534
rect 403782 656298 439226 656534
rect 439462 656298 439546 656534
rect 439782 656298 475226 656534
rect 475462 656298 475546 656534
rect 475782 656298 511226 656534
rect 511462 656298 511546 656534
rect 511782 656298 547226 656534
rect 547462 656298 547546 656534
rect 547782 656298 590142 656534
rect 590378 656298 590462 656534
rect 590698 656298 592650 656534
rect -8726 656266 592650 656298
rect -8726 655614 592650 655646
rect -8726 655378 -5814 655614
rect -5578 655378 -5494 655614
rect -5258 655378 5986 655614
rect 6222 655378 6306 655614
rect 6542 655378 41986 655614
rect 42222 655378 42306 655614
rect 42542 655378 77986 655614
rect 78222 655378 78306 655614
rect 78542 655378 113986 655614
rect 114222 655378 114306 655614
rect 114542 655378 149986 655614
rect 150222 655378 150306 655614
rect 150542 655378 185986 655614
rect 186222 655378 186306 655614
rect 186542 655378 221986 655614
rect 222222 655378 222306 655614
rect 222542 655378 257986 655614
rect 258222 655378 258306 655614
rect 258542 655378 293986 655614
rect 294222 655378 294306 655614
rect 294542 655378 329986 655614
rect 330222 655378 330306 655614
rect 330542 655378 365986 655614
rect 366222 655378 366306 655614
rect 366542 655378 401986 655614
rect 402222 655378 402306 655614
rect 402542 655378 437986 655614
rect 438222 655378 438306 655614
rect 438542 655378 473986 655614
rect 474222 655378 474306 655614
rect 474542 655378 509986 655614
rect 510222 655378 510306 655614
rect 510542 655378 545986 655614
rect 546222 655378 546306 655614
rect 546542 655378 581986 655614
rect 582222 655378 582306 655614
rect 582542 655378 589182 655614
rect 589418 655378 589502 655614
rect 589738 655378 592650 655614
rect -8726 655294 592650 655378
rect -8726 655058 -5814 655294
rect -5578 655058 -5494 655294
rect -5258 655058 5986 655294
rect 6222 655058 6306 655294
rect 6542 655058 41986 655294
rect 42222 655058 42306 655294
rect 42542 655058 77986 655294
rect 78222 655058 78306 655294
rect 78542 655058 113986 655294
rect 114222 655058 114306 655294
rect 114542 655058 149986 655294
rect 150222 655058 150306 655294
rect 150542 655058 185986 655294
rect 186222 655058 186306 655294
rect 186542 655058 221986 655294
rect 222222 655058 222306 655294
rect 222542 655058 257986 655294
rect 258222 655058 258306 655294
rect 258542 655058 293986 655294
rect 294222 655058 294306 655294
rect 294542 655058 329986 655294
rect 330222 655058 330306 655294
rect 330542 655058 365986 655294
rect 366222 655058 366306 655294
rect 366542 655058 401986 655294
rect 402222 655058 402306 655294
rect 402542 655058 437986 655294
rect 438222 655058 438306 655294
rect 438542 655058 473986 655294
rect 474222 655058 474306 655294
rect 474542 655058 509986 655294
rect 510222 655058 510306 655294
rect 510542 655058 545986 655294
rect 546222 655058 546306 655294
rect 546542 655058 581986 655294
rect 582222 655058 582306 655294
rect 582542 655058 589182 655294
rect 589418 655058 589502 655294
rect 589738 655058 592650 655294
rect -8726 655026 592650 655058
rect -8726 654374 592650 654406
rect -8726 654138 -4854 654374
rect -4618 654138 -4534 654374
rect -4298 654138 4746 654374
rect 4982 654138 5066 654374
rect 5302 654138 40746 654374
rect 40982 654138 41066 654374
rect 41302 654138 76746 654374
rect 76982 654138 77066 654374
rect 77302 654138 112746 654374
rect 112982 654138 113066 654374
rect 113302 654138 148746 654374
rect 148982 654138 149066 654374
rect 149302 654138 184746 654374
rect 184982 654138 185066 654374
rect 185302 654138 220746 654374
rect 220982 654138 221066 654374
rect 221302 654138 256746 654374
rect 256982 654138 257066 654374
rect 257302 654138 292746 654374
rect 292982 654138 293066 654374
rect 293302 654138 328746 654374
rect 328982 654138 329066 654374
rect 329302 654138 364746 654374
rect 364982 654138 365066 654374
rect 365302 654138 400746 654374
rect 400982 654138 401066 654374
rect 401302 654138 436746 654374
rect 436982 654138 437066 654374
rect 437302 654138 472746 654374
rect 472982 654138 473066 654374
rect 473302 654138 508746 654374
rect 508982 654138 509066 654374
rect 509302 654138 544746 654374
rect 544982 654138 545066 654374
rect 545302 654138 580746 654374
rect 580982 654138 581066 654374
rect 581302 654138 588222 654374
rect 588458 654138 588542 654374
rect 588778 654138 592650 654374
rect -8726 654054 592650 654138
rect -8726 653818 -4854 654054
rect -4618 653818 -4534 654054
rect -4298 653818 4746 654054
rect 4982 653818 5066 654054
rect 5302 653818 40746 654054
rect 40982 653818 41066 654054
rect 41302 653818 76746 654054
rect 76982 653818 77066 654054
rect 77302 653818 112746 654054
rect 112982 653818 113066 654054
rect 113302 653818 148746 654054
rect 148982 653818 149066 654054
rect 149302 653818 184746 654054
rect 184982 653818 185066 654054
rect 185302 653818 220746 654054
rect 220982 653818 221066 654054
rect 221302 653818 256746 654054
rect 256982 653818 257066 654054
rect 257302 653818 292746 654054
rect 292982 653818 293066 654054
rect 293302 653818 328746 654054
rect 328982 653818 329066 654054
rect 329302 653818 364746 654054
rect 364982 653818 365066 654054
rect 365302 653818 400746 654054
rect 400982 653818 401066 654054
rect 401302 653818 436746 654054
rect 436982 653818 437066 654054
rect 437302 653818 472746 654054
rect 472982 653818 473066 654054
rect 473302 653818 508746 654054
rect 508982 653818 509066 654054
rect 509302 653818 544746 654054
rect 544982 653818 545066 654054
rect 545302 653818 580746 654054
rect 580982 653818 581066 654054
rect 581302 653818 588222 654054
rect 588458 653818 588542 654054
rect 588778 653818 592650 654054
rect -8726 653786 592650 653818
rect -8726 653134 592650 653166
rect -8726 652898 -3894 653134
rect -3658 652898 -3574 653134
rect -3338 652898 3506 653134
rect 3742 652898 3826 653134
rect 4062 652898 39506 653134
rect 39742 652898 39826 653134
rect 40062 652898 75506 653134
rect 75742 652898 75826 653134
rect 76062 652898 111506 653134
rect 111742 652898 111826 653134
rect 112062 652898 147506 653134
rect 147742 652898 147826 653134
rect 148062 652898 183506 653134
rect 183742 652898 183826 653134
rect 184062 652898 219506 653134
rect 219742 652898 219826 653134
rect 220062 652898 255506 653134
rect 255742 652898 255826 653134
rect 256062 652898 291506 653134
rect 291742 652898 291826 653134
rect 292062 652898 327506 653134
rect 327742 652898 327826 653134
rect 328062 652898 363506 653134
rect 363742 652898 363826 653134
rect 364062 652898 399506 653134
rect 399742 652898 399826 653134
rect 400062 652898 435506 653134
rect 435742 652898 435826 653134
rect 436062 652898 471506 653134
rect 471742 652898 471826 653134
rect 472062 652898 507506 653134
rect 507742 652898 507826 653134
rect 508062 652898 543506 653134
rect 543742 652898 543826 653134
rect 544062 652898 579506 653134
rect 579742 652898 579826 653134
rect 580062 652898 587262 653134
rect 587498 652898 587582 653134
rect 587818 652898 592650 653134
rect -8726 652814 592650 652898
rect -8726 652578 -3894 652814
rect -3658 652578 -3574 652814
rect -3338 652578 3506 652814
rect 3742 652578 3826 652814
rect 4062 652578 39506 652814
rect 39742 652578 39826 652814
rect 40062 652578 75506 652814
rect 75742 652578 75826 652814
rect 76062 652578 111506 652814
rect 111742 652578 111826 652814
rect 112062 652578 147506 652814
rect 147742 652578 147826 652814
rect 148062 652578 183506 652814
rect 183742 652578 183826 652814
rect 184062 652578 219506 652814
rect 219742 652578 219826 652814
rect 220062 652578 255506 652814
rect 255742 652578 255826 652814
rect 256062 652578 291506 652814
rect 291742 652578 291826 652814
rect 292062 652578 327506 652814
rect 327742 652578 327826 652814
rect 328062 652578 363506 652814
rect 363742 652578 363826 652814
rect 364062 652578 399506 652814
rect 399742 652578 399826 652814
rect 400062 652578 435506 652814
rect 435742 652578 435826 652814
rect 436062 652578 471506 652814
rect 471742 652578 471826 652814
rect 472062 652578 507506 652814
rect 507742 652578 507826 652814
rect 508062 652578 543506 652814
rect 543742 652578 543826 652814
rect 544062 652578 579506 652814
rect 579742 652578 579826 652814
rect 580062 652578 587262 652814
rect 587498 652578 587582 652814
rect 587818 652578 592650 652814
rect -8726 652546 592650 652578
rect -8726 651894 592650 651926
rect -8726 651658 -2934 651894
rect -2698 651658 -2614 651894
rect -2378 651658 2266 651894
rect 2502 651658 2586 651894
rect 2822 651658 38266 651894
rect 38502 651658 38586 651894
rect 38822 651658 74266 651894
rect 74502 651658 74586 651894
rect 74822 651658 110266 651894
rect 110502 651658 110586 651894
rect 110822 651658 146266 651894
rect 146502 651658 146586 651894
rect 146822 651658 182266 651894
rect 182502 651658 182586 651894
rect 182822 651658 218266 651894
rect 218502 651658 218586 651894
rect 218822 651658 254266 651894
rect 254502 651658 254586 651894
rect 254822 651658 290266 651894
rect 290502 651658 290586 651894
rect 290822 651658 326266 651894
rect 326502 651658 326586 651894
rect 326822 651658 362266 651894
rect 362502 651658 362586 651894
rect 362822 651658 398266 651894
rect 398502 651658 398586 651894
rect 398822 651658 434266 651894
rect 434502 651658 434586 651894
rect 434822 651658 470266 651894
rect 470502 651658 470586 651894
rect 470822 651658 506266 651894
rect 506502 651658 506586 651894
rect 506822 651658 542266 651894
rect 542502 651658 542586 651894
rect 542822 651658 578266 651894
rect 578502 651658 578586 651894
rect 578822 651658 586302 651894
rect 586538 651658 586622 651894
rect 586858 651658 592650 651894
rect -8726 651574 592650 651658
rect -8726 651338 -2934 651574
rect -2698 651338 -2614 651574
rect -2378 651338 2266 651574
rect 2502 651338 2586 651574
rect 2822 651338 38266 651574
rect 38502 651338 38586 651574
rect 38822 651338 74266 651574
rect 74502 651338 74586 651574
rect 74822 651338 110266 651574
rect 110502 651338 110586 651574
rect 110822 651338 146266 651574
rect 146502 651338 146586 651574
rect 146822 651338 182266 651574
rect 182502 651338 182586 651574
rect 182822 651338 218266 651574
rect 218502 651338 218586 651574
rect 218822 651338 254266 651574
rect 254502 651338 254586 651574
rect 254822 651338 290266 651574
rect 290502 651338 290586 651574
rect 290822 651338 326266 651574
rect 326502 651338 326586 651574
rect 326822 651338 362266 651574
rect 362502 651338 362586 651574
rect 362822 651338 398266 651574
rect 398502 651338 398586 651574
rect 398822 651338 434266 651574
rect 434502 651338 434586 651574
rect 434822 651338 470266 651574
rect 470502 651338 470586 651574
rect 470822 651338 506266 651574
rect 506502 651338 506586 651574
rect 506822 651338 542266 651574
rect 542502 651338 542586 651574
rect 542822 651338 578266 651574
rect 578502 651338 578586 651574
rect 578822 651338 586302 651574
rect 586538 651338 586622 651574
rect 586858 651338 592650 651574
rect -8726 651306 592650 651338
rect -8726 650654 592650 650686
rect -8726 650418 -1974 650654
rect -1738 650418 -1654 650654
rect -1418 650418 1026 650654
rect 1262 650418 1346 650654
rect 1582 650418 37026 650654
rect 37262 650418 37346 650654
rect 37582 650418 73026 650654
rect 73262 650418 73346 650654
rect 73582 650418 109026 650654
rect 109262 650418 109346 650654
rect 109582 650418 145026 650654
rect 145262 650418 145346 650654
rect 145582 650418 181026 650654
rect 181262 650418 181346 650654
rect 181582 650418 217026 650654
rect 217262 650418 217346 650654
rect 217582 650418 253026 650654
rect 253262 650418 253346 650654
rect 253582 650418 289026 650654
rect 289262 650418 289346 650654
rect 289582 650418 325026 650654
rect 325262 650418 325346 650654
rect 325582 650418 361026 650654
rect 361262 650418 361346 650654
rect 361582 650418 397026 650654
rect 397262 650418 397346 650654
rect 397582 650418 433026 650654
rect 433262 650418 433346 650654
rect 433582 650418 469026 650654
rect 469262 650418 469346 650654
rect 469582 650418 505026 650654
rect 505262 650418 505346 650654
rect 505582 650418 541026 650654
rect 541262 650418 541346 650654
rect 541582 650418 577026 650654
rect 577262 650418 577346 650654
rect 577582 650418 585342 650654
rect 585578 650418 585662 650654
rect 585898 650418 592650 650654
rect -8726 650334 592650 650418
rect -8726 650098 -1974 650334
rect -1738 650098 -1654 650334
rect -1418 650098 1026 650334
rect 1262 650098 1346 650334
rect 1582 650098 37026 650334
rect 37262 650098 37346 650334
rect 37582 650098 73026 650334
rect 73262 650098 73346 650334
rect 73582 650098 109026 650334
rect 109262 650098 109346 650334
rect 109582 650098 145026 650334
rect 145262 650098 145346 650334
rect 145582 650098 181026 650334
rect 181262 650098 181346 650334
rect 181582 650098 217026 650334
rect 217262 650098 217346 650334
rect 217582 650098 253026 650334
rect 253262 650098 253346 650334
rect 253582 650098 289026 650334
rect 289262 650098 289346 650334
rect 289582 650098 325026 650334
rect 325262 650098 325346 650334
rect 325582 650098 361026 650334
rect 361262 650098 361346 650334
rect 361582 650098 397026 650334
rect 397262 650098 397346 650334
rect 397582 650098 433026 650334
rect 433262 650098 433346 650334
rect 433582 650098 469026 650334
rect 469262 650098 469346 650334
rect 469582 650098 505026 650334
rect 505262 650098 505346 650334
rect 505582 650098 541026 650334
rect 541262 650098 541346 650334
rect 541582 650098 577026 650334
rect 577262 650098 577346 650334
rect 577582 650098 585342 650334
rect 585578 650098 585662 650334
rect 585898 650098 592650 650334
rect -8726 650066 592650 650098
rect -8726 623334 592650 623366
rect -8726 623098 -8694 623334
rect -8458 623098 -8374 623334
rect -8138 623098 9706 623334
rect 9942 623098 10026 623334
rect 10262 623098 45706 623334
rect 45942 623098 46026 623334
rect 46262 623098 81706 623334
rect 81942 623098 82026 623334
rect 82262 623098 117706 623334
rect 117942 623098 118026 623334
rect 118262 623098 153706 623334
rect 153942 623098 154026 623334
rect 154262 623098 189706 623334
rect 189942 623098 190026 623334
rect 190262 623098 225706 623334
rect 225942 623098 226026 623334
rect 226262 623098 261706 623334
rect 261942 623098 262026 623334
rect 262262 623098 297706 623334
rect 297942 623098 298026 623334
rect 298262 623098 333706 623334
rect 333942 623098 334026 623334
rect 334262 623098 369706 623334
rect 369942 623098 370026 623334
rect 370262 623098 405706 623334
rect 405942 623098 406026 623334
rect 406262 623098 441706 623334
rect 441942 623098 442026 623334
rect 442262 623098 477706 623334
rect 477942 623098 478026 623334
rect 478262 623098 513706 623334
rect 513942 623098 514026 623334
rect 514262 623098 549706 623334
rect 549942 623098 550026 623334
rect 550262 623098 592062 623334
rect 592298 623098 592382 623334
rect 592618 623098 592650 623334
rect -8726 623014 592650 623098
rect -8726 622778 -8694 623014
rect -8458 622778 -8374 623014
rect -8138 622778 9706 623014
rect 9942 622778 10026 623014
rect 10262 622778 45706 623014
rect 45942 622778 46026 623014
rect 46262 622778 81706 623014
rect 81942 622778 82026 623014
rect 82262 622778 117706 623014
rect 117942 622778 118026 623014
rect 118262 622778 153706 623014
rect 153942 622778 154026 623014
rect 154262 622778 189706 623014
rect 189942 622778 190026 623014
rect 190262 622778 225706 623014
rect 225942 622778 226026 623014
rect 226262 622778 261706 623014
rect 261942 622778 262026 623014
rect 262262 622778 297706 623014
rect 297942 622778 298026 623014
rect 298262 622778 333706 623014
rect 333942 622778 334026 623014
rect 334262 622778 369706 623014
rect 369942 622778 370026 623014
rect 370262 622778 405706 623014
rect 405942 622778 406026 623014
rect 406262 622778 441706 623014
rect 441942 622778 442026 623014
rect 442262 622778 477706 623014
rect 477942 622778 478026 623014
rect 478262 622778 513706 623014
rect 513942 622778 514026 623014
rect 514262 622778 549706 623014
rect 549942 622778 550026 623014
rect 550262 622778 592062 623014
rect 592298 622778 592382 623014
rect 592618 622778 592650 623014
rect -8726 622746 592650 622778
rect -8726 622094 592650 622126
rect -8726 621858 -7734 622094
rect -7498 621858 -7414 622094
rect -7178 621858 8466 622094
rect 8702 621858 8786 622094
rect 9022 621858 44466 622094
rect 44702 621858 44786 622094
rect 45022 621858 80466 622094
rect 80702 621858 80786 622094
rect 81022 621858 116466 622094
rect 116702 621858 116786 622094
rect 117022 621858 152466 622094
rect 152702 621858 152786 622094
rect 153022 621858 188466 622094
rect 188702 621858 188786 622094
rect 189022 621858 224466 622094
rect 224702 621858 224786 622094
rect 225022 621858 260466 622094
rect 260702 621858 260786 622094
rect 261022 621858 296466 622094
rect 296702 621858 296786 622094
rect 297022 621858 332466 622094
rect 332702 621858 332786 622094
rect 333022 621858 368466 622094
rect 368702 621858 368786 622094
rect 369022 621858 404466 622094
rect 404702 621858 404786 622094
rect 405022 621858 440466 622094
rect 440702 621858 440786 622094
rect 441022 621858 476466 622094
rect 476702 621858 476786 622094
rect 477022 621858 512466 622094
rect 512702 621858 512786 622094
rect 513022 621858 548466 622094
rect 548702 621858 548786 622094
rect 549022 621858 591102 622094
rect 591338 621858 591422 622094
rect 591658 621858 592650 622094
rect -8726 621774 592650 621858
rect -8726 621538 -7734 621774
rect -7498 621538 -7414 621774
rect -7178 621538 8466 621774
rect 8702 621538 8786 621774
rect 9022 621538 44466 621774
rect 44702 621538 44786 621774
rect 45022 621538 80466 621774
rect 80702 621538 80786 621774
rect 81022 621538 116466 621774
rect 116702 621538 116786 621774
rect 117022 621538 152466 621774
rect 152702 621538 152786 621774
rect 153022 621538 188466 621774
rect 188702 621538 188786 621774
rect 189022 621538 224466 621774
rect 224702 621538 224786 621774
rect 225022 621538 260466 621774
rect 260702 621538 260786 621774
rect 261022 621538 296466 621774
rect 296702 621538 296786 621774
rect 297022 621538 332466 621774
rect 332702 621538 332786 621774
rect 333022 621538 368466 621774
rect 368702 621538 368786 621774
rect 369022 621538 404466 621774
rect 404702 621538 404786 621774
rect 405022 621538 440466 621774
rect 440702 621538 440786 621774
rect 441022 621538 476466 621774
rect 476702 621538 476786 621774
rect 477022 621538 512466 621774
rect 512702 621538 512786 621774
rect 513022 621538 548466 621774
rect 548702 621538 548786 621774
rect 549022 621538 591102 621774
rect 591338 621538 591422 621774
rect 591658 621538 592650 621774
rect -8726 621506 592650 621538
rect -8726 620854 592650 620886
rect -8726 620618 -6774 620854
rect -6538 620618 -6454 620854
rect -6218 620618 7226 620854
rect 7462 620618 7546 620854
rect 7782 620618 43226 620854
rect 43462 620618 43546 620854
rect 43782 620618 79226 620854
rect 79462 620618 79546 620854
rect 79782 620618 115226 620854
rect 115462 620618 115546 620854
rect 115782 620618 151226 620854
rect 151462 620618 151546 620854
rect 151782 620618 187226 620854
rect 187462 620618 187546 620854
rect 187782 620618 223226 620854
rect 223462 620618 223546 620854
rect 223782 620618 259226 620854
rect 259462 620618 259546 620854
rect 259782 620618 295226 620854
rect 295462 620618 295546 620854
rect 295782 620618 331226 620854
rect 331462 620618 331546 620854
rect 331782 620618 367226 620854
rect 367462 620618 367546 620854
rect 367782 620618 403226 620854
rect 403462 620618 403546 620854
rect 403782 620618 439226 620854
rect 439462 620618 439546 620854
rect 439782 620618 475226 620854
rect 475462 620618 475546 620854
rect 475782 620618 511226 620854
rect 511462 620618 511546 620854
rect 511782 620618 547226 620854
rect 547462 620618 547546 620854
rect 547782 620618 590142 620854
rect 590378 620618 590462 620854
rect 590698 620618 592650 620854
rect -8726 620534 592650 620618
rect -8726 620298 -6774 620534
rect -6538 620298 -6454 620534
rect -6218 620298 7226 620534
rect 7462 620298 7546 620534
rect 7782 620298 43226 620534
rect 43462 620298 43546 620534
rect 43782 620298 79226 620534
rect 79462 620298 79546 620534
rect 79782 620298 115226 620534
rect 115462 620298 115546 620534
rect 115782 620298 151226 620534
rect 151462 620298 151546 620534
rect 151782 620298 187226 620534
rect 187462 620298 187546 620534
rect 187782 620298 223226 620534
rect 223462 620298 223546 620534
rect 223782 620298 259226 620534
rect 259462 620298 259546 620534
rect 259782 620298 295226 620534
rect 295462 620298 295546 620534
rect 295782 620298 331226 620534
rect 331462 620298 331546 620534
rect 331782 620298 367226 620534
rect 367462 620298 367546 620534
rect 367782 620298 403226 620534
rect 403462 620298 403546 620534
rect 403782 620298 439226 620534
rect 439462 620298 439546 620534
rect 439782 620298 475226 620534
rect 475462 620298 475546 620534
rect 475782 620298 511226 620534
rect 511462 620298 511546 620534
rect 511782 620298 547226 620534
rect 547462 620298 547546 620534
rect 547782 620298 590142 620534
rect 590378 620298 590462 620534
rect 590698 620298 592650 620534
rect -8726 620266 592650 620298
rect -8726 619614 592650 619646
rect -8726 619378 -5814 619614
rect -5578 619378 -5494 619614
rect -5258 619378 5986 619614
rect 6222 619378 6306 619614
rect 6542 619378 41986 619614
rect 42222 619378 42306 619614
rect 42542 619378 77986 619614
rect 78222 619378 78306 619614
rect 78542 619378 113986 619614
rect 114222 619378 114306 619614
rect 114542 619378 149986 619614
rect 150222 619378 150306 619614
rect 150542 619378 185986 619614
rect 186222 619378 186306 619614
rect 186542 619378 221986 619614
rect 222222 619378 222306 619614
rect 222542 619378 257986 619614
rect 258222 619378 258306 619614
rect 258542 619378 293986 619614
rect 294222 619378 294306 619614
rect 294542 619378 329986 619614
rect 330222 619378 330306 619614
rect 330542 619378 365986 619614
rect 366222 619378 366306 619614
rect 366542 619378 401986 619614
rect 402222 619378 402306 619614
rect 402542 619378 437986 619614
rect 438222 619378 438306 619614
rect 438542 619378 473986 619614
rect 474222 619378 474306 619614
rect 474542 619378 509986 619614
rect 510222 619378 510306 619614
rect 510542 619378 545986 619614
rect 546222 619378 546306 619614
rect 546542 619378 581986 619614
rect 582222 619378 582306 619614
rect 582542 619378 589182 619614
rect 589418 619378 589502 619614
rect 589738 619378 592650 619614
rect -8726 619294 592650 619378
rect -8726 619058 -5814 619294
rect -5578 619058 -5494 619294
rect -5258 619058 5986 619294
rect 6222 619058 6306 619294
rect 6542 619058 41986 619294
rect 42222 619058 42306 619294
rect 42542 619058 77986 619294
rect 78222 619058 78306 619294
rect 78542 619058 113986 619294
rect 114222 619058 114306 619294
rect 114542 619058 149986 619294
rect 150222 619058 150306 619294
rect 150542 619058 185986 619294
rect 186222 619058 186306 619294
rect 186542 619058 221986 619294
rect 222222 619058 222306 619294
rect 222542 619058 257986 619294
rect 258222 619058 258306 619294
rect 258542 619058 293986 619294
rect 294222 619058 294306 619294
rect 294542 619058 329986 619294
rect 330222 619058 330306 619294
rect 330542 619058 365986 619294
rect 366222 619058 366306 619294
rect 366542 619058 401986 619294
rect 402222 619058 402306 619294
rect 402542 619058 437986 619294
rect 438222 619058 438306 619294
rect 438542 619058 473986 619294
rect 474222 619058 474306 619294
rect 474542 619058 509986 619294
rect 510222 619058 510306 619294
rect 510542 619058 545986 619294
rect 546222 619058 546306 619294
rect 546542 619058 581986 619294
rect 582222 619058 582306 619294
rect 582542 619058 589182 619294
rect 589418 619058 589502 619294
rect 589738 619058 592650 619294
rect -8726 619026 592650 619058
rect -8726 618374 592650 618406
rect -8726 618138 -4854 618374
rect -4618 618138 -4534 618374
rect -4298 618138 4746 618374
rect 4982 618138 5066 618374
rect 5302 618138 40746 618374
rect 40982 618138 41066 618374
rect 41302 618138 76746 618374
rect 76982 618138 77066 618374
rect 77302 618138 112746 618374
rect 112982 618138 113066 618374
rect 113302 618138 148746 618374
rect 148982 618138 149066 618374
rect 149302 618138 184746 618374
rect 184982 618138 185066 618374
rect 185302 618138 220746 618374
rect 220982 618138 221066 618374
rect 221302 618138 256746 618374
rect 256982 618138 257066 618374
rect 257302 618138 292746 618374
rect 292982 618138 293066 618374
rect 293302 618138 328746 618374
rect 328982 618138 329066 618374
rect 329302 618138 364746 618374
rect 364982 618138 365066 618374
rect 365302 618138 400746 618374
rect 400982 618138 401066 618374
rect 401302 618138 436746 618374
rect 436982 618138 437066 618374
rect 437302 618138 472746 618374
rect 472982 618138 473066 618374
rect 473302 618138 508746 618374
rect 508982 618138 509066 618374
rect 509302 618138 544746 618374
rect 544982 618138 545066 618374
rect 545302 618138 580746 618374
rect 580982 618138 581066 618374
rect 581302 618138 588222 618374
rect 588458 618138 588542 618374
rect 588778 618138 592650 618374
rect -8726 618054 592650 618138
rect -8726 617818 -4854 618054
rect -4618 617818 -4534 618054
rect -4298 617818 4746 618054
rect 4982 617818 5066 618054
rect 5302 617818 40746 618054
rect 40982 617818 41066 618054
rect 41302 617818 76746 618054
rect 76982 617818 77066 618054
rect 77302 617818 112746 618054
rect 112982 617818 113066 618054
rect 113302 617818 148746 618054
rect 148982 617818 149066 618054
rect 149302 617818 184746 618054
rect 184982 617818 185066 618054
rect 185302 617818 220746 618054
rect 220982 617818 221066 618054
rect 221302 617818 256746 618054
rect 256982 617818 257066 618054
rect 257302 617818 292746 618054
rect 292982 617818 293066 618054
rect 293302 617818 328746 618054
rect 328982 617818 329066 618054
rect 329302 617818 364746 618054
rect 364982 617818 365066 618054
rect 365302 617818 400746 618054
rect 400982 617818 401066 618054
rect 401302 617818 436746 618054
rect 436982 617818 437066 618054
rect 437302 617818 472746 618054
rect 472982 617818 473066 618054
rect 473302 617818 508746 618054
rect 508982 617818 509066 618054
rect 509302 617818 544746 618054
rect 544982 617818 545066 618054
rect 545302 617818 580746 618054
rect 580982 617818 581066 618054
rect 581302 617818 588222 618054
rect 588458 617818 588542 618054
rect 588778 617818 592650 618054
rect -8726 617786 592650 617818
rect -8726 617134 592650 617166
rect -8726 616898 -3894 617134
rect -3658 616898 -3574 617134
rect -3338 616898 3506 617134
rect 3742 616898 3826 617134
rect 4062 616898 39506 617134
rect 39742 616898 39826 617134
rect 40062 616898 75506 617134
rect 75742 616898 75826 617134
rect 76062 616898 111506 617134
rect 111742 616898 111826 617134
rect 112062 616898 147506 617134
rect 147742 616898 147826 617134
rect 148062 616898 183506 617134
rect 183742 616898 183826 617134
rect 184062 616898 219506 617134
rect 219742 616898 219826 617134
rect 220062 616898 255506 617134
rect 255742 616898 255826 617134
rect 256062 616898 291506 617134
rect 291742 616898 291826 617134
rect 292062 616898 327506 617134
rect 327742 616898 327826 617134
rect 328062 616898 363506 617134
rect 363742 616898 363826 617134
rect 364062 616898 399506 617134
rect 399742 616898 399826 617134
rect 400062 616898 435506 617134
rect 435742 616898 435826 617134
rect 436062 616898 471506 617134
rect 471742 616898 471826 617134
rect 472062 616898 507506 617134
rect 507742 616898 507826 617134
rect 508062 616898 543506 617134
rect 543742 616898 543826 617134
rect 544062 616898 579506 617134
rect 579742 616898 579826 617134
rect 580062 616898 587262 617134
rect 587498 616898 587582 617134
rect 587818 616898 592650 617134
rect -8726 616814 592650 616898
rect -8726 616578 -3894 616814
rect -3658 616578 -3574 616814
rect -3338 616578 3506 616814
rect 3742 616578 3826 616814
rect 4062 616578 39506 616814
rect 39742 616578 39826 616814
rect 40062 616578 75506 616814
rect 75742 616578 75826 616814
rect 76062 616578 111506 616814
rect 111742 616578 111826 616814
rect 112062 616578 147506 616814
rect 147742 616578 147826 616814
rect 148062 616578 183506 616814
rect 183742 616578 183826 616814
rect 184062 616578 219506 616814
rect 219742 616578 219826 616814
rect 220062 616578 255506 616814
rect 255742 616578 255826 616814
rect 256062 616578 291506 616814
rect 291742 616578 291826 616814
rect 292062 616578 327506 616814
rect 327742 616578 327826 616814
rect 328062 616578 363506 616814
rect 363742 616578 363826 616814
rect 364062 616578 399506 616814
rect 399742 616578 399826 616814
rect 400062 616578 435506 616814
rect 435742 616578 435826 616814
rect 436062 616578 471506 616814
rect 471742 616578 471826 616814
rect 472062 616578 507506 616814
rect 507742 616578 507826 616814
rect 508062 616578 543506 616814
rect 543742 616578 543826 616814
rect 544062 616578 579506 616814
rect 579742 616578 579826 616814
rect 580062 616578 587262 616814
rect 587498 616578 587582 616814
rect 587818 616578 592650 616814
rect -8726 616546 592650 616578
rect -8726 615894 592650 615926
rect -8726 615658 -2934 615894
rect -2698 615658 -2614 615894
rect -2378 615658 2266 615894
rect 2502 615658 2586 615894
rect 2822 615658 38266 615894
rect 38502 615658 38586 615894
rect 38822 615658 74266 615894
rect 74502 615658 74586 615894
rect 74822 615658 110266 615894
rect 110502 615658 110586 615894
rect 110822 615658 146266 615894
rect 146502 615658 146586 615894
rect 146822 615658 182266 615894
rect 182502 615658 182586 615894
rect 182822 615658 218266 615894
rect 218502 615658 218586 615894
rect 218822 615658 254266 615894
rect 254502 615658 254586 615894
rect 254822 615658 290266 615894
rect 290502 615658 290586 615894
rect 290822 615658 326266 615894
rect 326502 615658 326586 615894
rect 326822 615658 362266 615894
rect 362502 615658 362586 615894
rect 362822 615658 398266 615894
rect 398502 615658 398586 615894
rect 398822 615658 434266 615894
rect 434502 615658 434586 615894
rect 434822 615658 470266 615894
rect 470502 615658 470586 615894
rect 470822 615658 506266 615894
rect 506502 615658 506586 615894
rect 506822 615658 542266 615894
rect 542502 615658 542586 615894
rect 542822 615658 578266 615894
rect 578502 615658 578586 615894
rect 578822 615658 586302 615894
rect 586538 615658 586622 615894
rect 586858 615658 592650 615894
rect -8726 615574 592650 615658
rect -8726 615338 -2934 615574
rect -2698 615338 -2614 615574
rect -2378 615338 2266 615574
rect 2502 615338 2586 615574
rect 2822 615338 38266 615574
rect 38502 615338 38586 615574
rect 38822 615338 74266 615574
rect 74502 615338 74586 615574
rect 74822 615338 110266 615574
rect 110502 615338 110586 615574
rect 110822 615338 146266 615574
rect 146502 615338 146586 615574
rect 146822 615338 182266 615574
rect 182502 615338 182586 615574
rect 182822 615338 218266 615574
rect 218502 615338 218586 615574
rect 218822 615338 254266 615574
rect 254502 615338 254586 615574
rect 254822 615338 290266 615574
rect 290502 615338 290586 615574
rect 290822 615338 326266 615574
rect 326502 615338 326586 615574
rect 326822 615338 362266 615574
rect 362502 615338 362586 615574
rect 362822 615338 398266 615574
rect 398502 615338 398586 615574
rect 398822 615338 434266 615574
rect 434502 615338 434586 615574
rect 434822 615338 470266 615574
rect 470502 615338 470586 615574
rect 470822 615338 506266 615574
rect 506502 615338 506586 615574
rect 506822 615338 542266 615574
rect 542502 615338 542586 615574
rect 542822 615338 578266 615574
rect 578502 615338 578586 615574
rect 578822 615338 586302 615574
rect 586538 615338 586622 615574
rect 586858 615338 592650 615574
rect -8726 615306 592650 615338
rect -8726 614654 592650 614686
rect -8726 614418 -1974 614654
rect -1738 614418 -1654 614654
rect -1418 614418 1026 614654
rect 1262 614418 1346 614654
rect 1582 614418 37026 614654
rect 37262 614418 37346 614654
rect 37582 614418 73026 614654
rect 73262 614418 73346 614654
rect 73582 614418 109026 614654
rect 109262 614418 109346 614654
rect 109582 614418 145026 614654
rect 145262 614418 145346 614654
rect 145582 614418 181026 614654
rect 181262 614418 181346 614654
rect 181582 614418 217026 614654
rect 217262 614418 217346 614654
rect 217582 614418 253026 614654
rect 253262 614418 253346 614654
rect 253582 614418 289026 614654
rect 289262 614418 289346 614654
rect 289582 614418 325026 614654
rect 325262 614418 325346 614654
rect 325582 614418 361026 614654
rect 361262 614418 361346 614654
rect 361582 614418 397026 614654
rect 397262 614418 397346 614654
rect 397582 614418 433026 614654
rect 433262 614418 433346 614654
rect 433582 614418 469026 614654
rect 469262 614418 469346 614654
rect 469582 614418 505026 614654
rect 505262 614418 505346 614654
rect 505582 614418 541026 614654
rect 541262 614418 541346 614654
rect 541582 614418 577026 614654
rect 577262 614418 577346 614654
rect 577582 614418 585342 614654
rect 585578 614418 585662 614654
rect 585898 614418 592650 614654
rect -8726 614334 592650 614418
rect -8726 614098 -1974 614334
rect -1738 614098 -1654 614334
rect -1418 614098 1026 614334
rect 1262 614098 1346 614334
rect 1582 614098 37026 614334
rect 37262 614098 37346 614334
rect 37582 614098 73026 614334
rect 73262 614098 73346 614334
rect 73582 614098 109026 614334
rect 109262 614098 109346 614334
rect 109582 614098 145026 614334
rect 145262 614098 145346 614334
rect 145582 614098 181026 614334
rect 181262 614098 181346 614334
rect 181582 614098 217026 614334
rect 217262 614098 217346 614334
rect 217582 614098 253026 614334
rect 253262 614098 253346 614334
rect 253582 614098 289026 614334
rect 289262 614098 289346 614334
rect 289582 614098 325026 614334
rect 325262 614098 325346 614334
rect 325582 614098 361026 614334
rect 361262 614098 361346 614334
rect 361582 614098 397026 614334
rect 397262 614098 397346 614334
rect 397582 614098 433026 614334
rect 433262 614098 433346 614334
rect 433582 614098 469026 614334
rect 469262 614098 469346 614334
rect 469582 614098 505026 614334
rect 505262 614098 505346 614334
rect 505582 614098 541026 614334
rect 541262 614098 541346 614334
rect 541582 614098 577026 614334
rect 577262 614098 577346 614334
rect 577582 614098 585342 614334
rect 585578 614098 585662 614334
rect 585898 614098 592650 614334
rect -8726 614066 592650 614098
rect -8726 587334 592650 587366
rect -8726 587098 -8694 587334
rect -8458 587098 -8374 587334
rect -8138 587098 9706 587334
rect 9942 587098 10026 587334
rect 10262 587098 45706 587334
rect 45942 587098 46026 587334
rect 46262 587098 81706 587334
rect 81942 587098 82026 587334
rect 82262 587098 117706 587334
rect 117942 587098 118026 587334
rect 118262 587098 153706 587334
rect 153942 587098 154026 587334
rect 154262 587098 189706 587334
rect 189942 587098 190026 587334
rect 190262 587098 225706 587334
rect 225942 587098 226026 587334
rect 226262 587098 261706 587334
rect 261942 587098 262026 587334
rect 262262 587098 297706 587334
rect 297942 587098 298026 587334
rect 298262 587098 333706 587334
rect 333942 587098 334026 587334
rect 334262 587098 369706 587334
rect 369942 587098 370026 587334
rect 370262 587098 405706 587334
rect 405942 587098 406026 587334
rect 406262 587098 441706 587334
rect 441942 587098 442026 587334
rect 442262 587098 477706 587334
rect 477942 587098 478026 587334
rect 478262 587098 513706 587334
rect 513942 587098 514026 587334
rect 514262 587098 549706 587334
rect 549942 587098 550026 587334
rect 550262 587098 592062 587334
rect 592298 587098 592382 587334
rect 592618 587098 592650 587334
rect -8726 587014 592650 587098
rect -8726 586778 -8694 587014
rect -8458 586778 -8374 587014
rect -8138 586778 9706 587014
rect 9942 586778 10026 587014
rect 10262 586778 45706 587014
rect 45942 586778 46026 587014
rect 46262 586778 81706 587014
rect 81942 586778 82026 587014
rect 82262 586778 117706 587014
rect 117942 586778 118026 587014
rect 118262 586778 153706 587014
rect 153942 586778 154026 587014
rect 154262 586778 189706 587014
rect 189942 586778 190026 587014
rect 190262 586778 225706 587014
rect 225942 586778 226026 587014
rect 226262 586778 261706 587014
rect 261942 586778 262026 587014
rect 262262 586778 297706 587014
rect 297942 586778 298026 587014
rect 298262 586778 333706 587014
rect 333942 586778 334026 587014
rect 334262 586778 369706 587014
rect 369942 586778 370026 587014
rect 370262 586778 405706 587014
rect 405942 586778 406026 587014
rect 406262 586778 441706 587014
rect 441942 586778 442026 587014
rect 442262 586778 477706 587014
rect 477942 586778 478026 587014
rect 478262 586778 513706 587014
rect 513942 586778 514026 587014
rect 514262 586778 549706 587014
rect 549942 586778 550026 587014
rect 550262 586778 592062 587014
rect 592298 586778 592382 587014
rect 592618 586778 592650 587014
rect -8726 586746 592650 586778
rect -8726 586094 592650 586126
rect -8726 585858 -7734 586094
rect -7498 585858 -7414 586094
rect -7178 585858 8466 586094
rect 8702 585858 8786 586094
rect 9022 585858 44466 586094
rect 44702 585858 44786 586094
rect 45022 585858 80466 586094
rect 80702 585858 80786 586094
rect 81022 585858 116466 586094
rect 116702 585858 116786 586094
rect 117022 585858 152466 586094
rect 152702 585858 152786 586094
rect 153022 585858 188466 586094
rect 188702 585858 188786 586094
rect 189022 585858 224466 586094
rect 224702 585858 224786 586094
rect 225022 585858 260466 586094
rect 260702 585858 260786 586094
rect 261022 585858 296466 586094
rect 296702 585858 296786 586094
rect 297022 585858 332466 586094
rect 332702 585858 332786 586094
rect 333022 585858 368466 586094
rect 368702 585858 368786 586094
rect 369022 585858 404466 586094
rect 404702 585858 404786 586094
rect 405022 585858 440466 586094
rect 440702 585858 440786 586094
rect 441022 585858 476466 586094
rect 476702 585858 476786 586094
rect 477022 585858 512466 586094
rect 512702 585858 512786 586094
rect 513022 585858 548466 586094
rect 548702 585858 548786 586094
rect 549022 585858 591102 586094
rect 591338 585858 591422 586094
rect 591658 585858 592650 586094
rect -8726 585774 592650 585858
rect -8726 585538 -7734 585774
rect -7498 585538 -7414 585774
rect -7178 585538 8466 585774
rect 8702 585538 8786 585774
rect 9022 585538 44466 585774
rect 44702 585538 44786 585774
rect 45022 585538 80466 585774
rect 80702 585538 80786 585774
rect 81022 585538 116466 585774
rect 116702 585538 116786 585774
rect 117022 585538 152466 585774
rect 152702 585538 152786 585774
rect 153022 585538 188466 585774
rect 188702 585538 188786 585774
rect 189022 585538 224466 585774
rect 224702 585538 224786 585774
rect 225022 585538 260466 585774
rect 260702 585538 260786 585774
rect 261022 585538 296466 585774
rect 296702 585538 296786 585774
rect 297022 585538 332466 585774
rect 332702 585538 332786 585774
rect 333022 585538 368466 585774
rect 368702 585538 368786 585774
rect 369022 585538 404466 585774
rect 404702 585538 404786 585774
rect 405022 585538 440466 585774
rect 440702 585538 440786 585774
rect 441022 585538 476466 585774
rect 476702 585538 476786 585774
rect 477022 585538 512466 585774
rect 512702 585538 512786 585774
rect 513022 585538 548466 585774
rect 548702 585538 548786 585774
rect 549022 585538 591102 585774
rect 591338 585538 591422 585774
rect 591658 585538 592650 585774
rect -8726 585506 592650 585538
rect -8726 584854 592650 584886
rect -8726 584618 -6774 584854
rect -6538 584618 -6454 584854
rect -6218 584618 7226 584854
rect 7462 584618 7546 584854
rect 7782 584618 43226 584854
rect 43462 584618 43546 584854
rect 43782 584618 79226 584854
rect 79462 584618 79546 584854
rect 79782 584618 115226 584854
rect 115462 584618 115546 584854
rect 115782 584618 151226 584854
rect 151462 584618 151546 584854
rect 151782 584618 187226 584854
rect 187462 584618 187546 584854
rect 187782 584618 223226 584854
rect 223462 584618 223546 584854
rect 223782 584618 259226 584854
rect 259462 584618 259546 584854
rect 259782 584618 295226 584854
rect 295462 584618 295546 584854
rect 295782 584618 331226 584854
rect 331462 584618 331546 584854
rect 331782 584618 367226 584854
rect 367462 584618 367546 584854
rect 367782 584618 403226 584854
rect 403462 584618 403546 584854
rect 403782 584618 439226 584854
rect 439462 584618 439546 584854
rect 439782 584618 475226 584854
rect 475462 584618 475546 584854
rect 475782 584618 511226 584854
rect 511462 584618 511546 584854
rect 511782 584618 547226 584854
rect 547462 584618 547546 584854
rect 547782 584618 590142 584854
rect 590378 584618 590462 584854
rect 590698 584618 592650 584854
rect -8726 584534 592650 584618
rect -8726 584298 -6774 584534
rect -6538 584298 -6454 584534
rect -6218 584298 7226 584534
rect 7462 584298 7546 584534
rect 7782 584298 43226 584534
rect 43462 584298 43546 584534
rect 43782 584298 79226 584534
rect 79462 584298 79546 584534
rect 79782 584298 115226 584534
rect 115462 584298 115546 584534
rect 115782 584298 151226 584534
rect 151462 584298 151546 584534
rect 151782 584298 187226 584534
rect 187462 584298 187546 584534
rect 187782 584298 223226 584534
rect 223462 584298 223546 584534
rect 223782 584298 259226 584534
rect 259462 584298 259546 584534
rect 259782 584298 295226 584534
rect 295462 584298 295546 584534
rect 295782 584298 331226 584534
rect 331462 584298 331546 584534
rect 331782 584298 367226 584534
rect 367462 584298 367546 584534
rect 367782 584298 403226 584534
rect 403462 584298 403546 584534
rect 403782 584298 439226 584534
rect 439462 584298 439546 584534
rect 439782 584298 475226 584534
rect 475462 584298 475546 584534
rect 475782 584298 511226 584534
rect 511462 584298 511546 584534
rect 511782 584298 547226 584534
rect 547462 584298 547546 584534
rect 547782 584298 590142 584534
rect 590378 584298 590462 584534
rect 590698 584298 592650 584534
rect -8726 584266 592650 584298
rect -8726 583614 592650 583646
rect -8726 583378 -5814 583614
rect -5578 583378 -5494 583614
rect -5258 583378 5986 583614
rect 6222 583378 6306 583614
rect 6542 583378 41986 583614
rect 42222 583378 42306 583614
rect 42542 583378 77986 583614
rect 78222 583378 78306 583614
rect 78542 583378 113986 583614
rect 114222 583378 114306 583614
rect 114542 583378 149986 583614
rect 150222 583378 150306 583614
rect 150542 583378 185986 583614
rect 186222 583378 186306 583614
rect 186542 583378 221986 583614
rect 222222 583378 222306 583614
rect 222542 583378 257986 583614
rect 258222 583378 258306 583614
rect 258542 583378 293986 583614
rect 294222 583378 294306 583614
rect 294542 583378 329986 583614
rect 330222 583378 330306 583614
rect 330542 583378 365986 583614
rect 366222 583378 366306 583614
rect 366542 583378 401986 583614
rect 402222 583378 402306 583614
rect 402542 583378 437986 583614
rect 438222 583378 438306 583614
rect 438542 583378 473986 583614
rect 474222 583378 474306 583614
rect 474542 583378 509986 583614
rect 510222 583378 510306 583614
rect 510542 583378 545986 583614
rect 546222 583378 546306 583614
rect 546542 583378 581986 583614
rect 582222 583378 582306 583614
rect 582542 583378 589182 583614
rect 589418 583378 589502 583614
rect 589738 583378 592650 583614
rect -8726 583294 592650 583378
rect -8726 583058 -5814 583294
rect -5578 583058 -5494 583294
rect -5258 583058 5986 583294
rect 6222 583058 6306 583294
rect 6542 583058 41986 583294
rect 42222 583058 42306 583294
rect 42542 583058 77986 583294
rect 78222 583058 78306 583294
rect 78542 583058 113986 583294
rect 114222 583058 114306 583294
rect 114542 583058 149986 583294
rect 150222 583058 150306 583294
rect 150542 583058 185986 583294
rect 186222 583058 186306 583294
rect 186542 583058 221986 583294
rect 222222 583058 222306 583294
rect 222542 583058 257986 583294
rect 258222 583058 258306 583294
rect 258542 583058 293986 583294
rect 294222 583058 294306 583294
rect 294542 583058 329986 583294
rect 330222 583058 330306 583294
rect 330542 583058 365986 583294
rect 366222 583058 366306 583294
rect 366542 583058 401986 583294
rect 402222 583058 402306 583294
rect 402542 583058 437986 583294
rect 438222 583058 438306 583294
rect 438542 583058 473986 583294
rect 474222 583058 474306 583294
rect 474542 583058 509986 583294
rect 510222 583058 510306 583294
rect 510542 583058 545986 583294
rect 546222 583058 546306 583294
rect 546542 583058 581986 583294
rect 582222 583058 582306 583294
rect 582542 583058 589182 583294
rect 589418 583058 589502 583294
rect 589738 583058 592650 583294
rect -8726 583026 592650 583058
rect -8726 582374 592650 582406
rect -8726 582138 -4854 582374
rect -4618 582138 -4534 582374
rect -4298 582138 4746 582374
rect 4982 582138 5066 582374
rect 5302 582138 40746 582374
rect 40982 582138 41066 582374
rect 41302 582138 76746 582374
rect 76982 582138 77066 582374
rect 77302 582138 112746 582374
rect 112982 582138 113066 582374
rect 113302 582138 148746 582374
rect 148982 582138 149066 582374
rect 149302 582138 184746 582374
rect 184982 582138 185066 582374
rect 185302 582138 220746 582374
rect 220982 582138 221066 582374
rect 221302 582138 256746 582374
rect 256982 582138 257066 582374
rect 257302 582138 292746 582374
rect 292982 582138 293066 582374
rect 293302 582138 328746 582374
rect 328982 582138 329066 582374
rect 329302 582138 364746 582374
rect 364982 582138 365066 582374
rect 365302 582138 400746 582374
rect 400982 582138 401066 582374
rect 401302 582138 436746 582374
rect 436982 582138 437066 582374
rect 437302 582138 472746 582374
rect 472982 582138 473066 582374
rect 473302 582138 508746 582374
rect 508982 582138 509066 582374
rect 509302 582138 544746 582374
rect 544982 582138 545066 582374
rect 545302 582138 580746 582374
rect 580982 582138 581066 582374
rect 581302 582138 588222 582374
rect 588458 582138 588542 582374
rect 588778 582138 592650 582374
rect -8726 582054 592650 582138
rect -8726 581818 -4854 582054
rect -4618 581818 -4534 582054
rect -4298 581818 4746 582054
rect 4982 581818 5066 582054
rect 5302 581818 40746 582054
rect 40982 581818 41066 582054
rect 41302 581818 76746 582054
rect 76982 581818 77066 582054
rect 77302 581818 112746 582054
rect 112982 581818 113066 582054
rect 113302 581818 148746 582054
rect 148982 581818 149066 582054
rect 149302 581818 184746 582054
rect 184982 581818 185066 582054
rect 185302 581818 220746 582054
rect 220982 581818 221066 582054
rect 221302 581818 256746 582054
rect 256982 581818 257066 582054
rect 257302 581818 292746 582054
rect 292982 581818 293066 582054
rect 293302 581818 328746 582054
rect 328982 581818 329066 582054
rect 329302 581818 364746 582054
rect 364982 581818 365066 582054
rect 365302 581818 400746 582054
rect 400982 581818 401066 582054
rect 401302 581818 436746 582054
rect 436982 581818 437066 582054
rect 437302 581818 472746 582054
rect 472982 581818 473066 582054
rect 473302 581818 508746 582054
rect 508982 581818 509066 582054
rect 509302 581818 544746 582054
rect 544982 581818 545066 582054
rect 545302 581818 580746 582054
rect 580982 581818 581066 582054
rect 581302 581818 588222 582054
rect 588458 581818 588542 582054
rect 588778 581818 592650 582054
rect -8726 581786 592650 581818
rect -8726 581134 592650 581166
rect -8726 580898 -3894 581134
rect -3658 580898 -3574 581134
rect -3338 580898 3506 581134
rect 3742 580898 3826 581134
rect 4062 580898 39506 581134
rect 39742 580898 39826 581134
rect 40062 580898 75506 581134
rect 75742 580898 75826 581134
rect 76062 580898 111506 581134
rect 111742 580898 111826 581134
rect 112062 580898 147506 581134
rect 147742 580898 147826 581134
rect 148062 580898 183506 581134
rect 183742 580898 183826 581134
rect 184062 580898 219506 581134
rect 219742 580898 219826 581134
rect 220062 580898 255506 581134
rect 255742 580898 255826 581134
rect 256062 580898 291506 581134
rect 291742 580898 291826 581134
rect 292062 580898 327506 581134
rect 327742 580898 327826 581134
rect 328062 580898 363506 581134
rect 363742 580898 363826 581134
rect 364062 580898 399506 581134
rect 399742 580898 399826 581134
rect 400062 580898 435506 581134
rect 435742 580898 435826 581134
rect 436062 580898 471506 581134
rect 471742 580898 471826 581134
rect 472062 580898 507506 581134
rect 507742 580898 507826 581134
rect 508062 580898 543506 581134
rect 543742 580898 543826 581134
rect 544062 580898 579506 581134
rect 579742 580898 579826 581134
rect 580062 580898 587262 581134
rect 587498 580898 587582 581134
rect 587818 580898 592650 581134
rect -8726 580814 592650 580898
rect -8726 580578 -3894 580814
rect -3658 580578 -3574 580814
rect -3338 580578 3506 580814
rect 3742 580578 3826 580814
rect 4062 580578 39506 580814
rect 39742 580578 39826 580814
rect 40062 580578 75506 580814
rect 75742 580578 75826 580814
rect 76062 580578 111506 580814
rect 111742 580578 111826 580814
rect 112062 580578 147506 580814
rect 147742 580578 147826 580814
rect 148062 580578 183506 580814
rect 183742 580578 183826 580814
rect 184062 580578 219506 580814
rect 219742 580578 219826 580814
rect 220062 580578 255506 580814
rect 255742 580578 255826 580814
rect 256062 580578 291506 580814
rect 291742 580578 291826 580814
rect 292062 580578 327506 580814
rect 327742 580578 327826 580814
rect 328062 580578 363506 580814
rect 363742 580578 363826 580814
rect 364062 580578 399506 580814
rect 399742 580578 399826 580814
rect 400062 580578 435506 580814
rect 435742 580578 435826 580814
rect 436062 580578 471506 580814
rect 471742 580578 471826 580814
rect 472062 580578 507506 580814
rect 507742 580578 507826 580814
rect 508062 580578 543506 580814
rect 543742 580578 543826 580814
rect 544062 580578 579506 580814
rect 579742 580578 579826 580814
rect 580062 580578 587262 580814
rect 587498 580578 587582 580814
rect 587818 580578 592650 580814
rect -8726 580546 592650 580578
rect -8726 579894 592650 579926
rect -8726 579658 -2934 579894
rect -2698 579658 -2614 579894
rect -2378 579658 2266 579894
rect 2502 579658 2586 579894
rect 2822 579658 38266 579894
rect 38502 579658 38586 579894
rect 38822 579658 74266 579894
rect 74502 579658 74586 579894
rect 74822 579658 110266 579894
rect 110502 579658 110586 579894
rect 110822 579658 146266 579894
rect 146502 579658 146586 579894
rect 146822 579658 182266 579894
rect 182502 579658 182586 579894
rect 182822 579658 218266 579894
rect 218502 579658 218586 579894
rect 218822 579658 254266 579894
rect 254502 579658 254586 579894
rect 254822 579658 290266 579894
rect 290502 579658 290586 579894
rect 290822 579658 326266 579894
rect 326502 579658 326586 579894
rect 326822 579658 362266 579894
rect 362502 579658 362586 579894
rect 362822 579658 398266 579894
rect 398502 579658 398586 579894
rect 398822 579658 434266 579894
rect 434502 579658 434586 579894
rect 434822 579658 470266 579894
rect 470502 579658 470586 579894
rect 470822 579658 506266 579894
rect 506502 579658 506586 579894
rect 506822 579658 542266 579894
rect 542502 579658 542586 579894
rect 542822 579658 578266 579894
rect 578502 579658 578586 579894
rect 578822 579658 586302 579894
rect 586538 579658 586622 579894
rect 586858 579658 592650 579894
rect -8726 579574 592650 579658
rect -8726 579338 -2934 579574
rect -2698 579338 -2614 579574
rect -2378 579338 2266 579574
rect 2502 579338 2586 579574
rect 2822 579338 38266 579574
rect 38502 579338 38586 579574
rect 38822 579338 74266 579574
rect 74502 579338 74586 579574
rect 74822 579338 110266 579574
rect 110502 579338 110586 579574
rect 110822 579338 146266 579574
rect 146502 579338 146586 579574
rect 146822 579338 182266 579574
rect 182502 579338 182586 579574
rect 182822 579338 218266 579574
rect 218502 579338 218586 579574
rect 218822 579338 254266 579574
rect 254502 579338 254586 579574
rect 254822 579338 290266 579574
rect 290502 579338 290586 579574
rect 290822 579338 326266 579574
rect 326502 579338 326586 579574
rect 326822 579338 362266 579574
rect 362502 579338 362586 579574
rect 362822 579338 398266 579574
rect 398502 579338 398586 579574
rect 398822 579338 434266 579574
rect 434502 579338 434586 579574
rect 434822 579338 470266 579574
rect 470502 579338 470586 579574
rect 470822 579338 506266 579574
rect 506502 579338 506586 579574
rect 506822 579338 542266 579574
rect 542502 579338 542586 579574
rect 542822 579338 578266 579574
rect 578502 579338 578586 579574
rect 578822 579338 586302 579574
rect 586538 579338 586622 579574
rect 586858 579338 592650 579574
rect -8726 579306 592650 579338
rect -8726 578654 592650 578686
rect -8726 578418 -1974 578654
rect -1738 578418 -1654 578654
rect -1418 578418 1026 578654
rect 1262 578418 1346 578654
rect 1582 578418 37026 578654
rect 37262 578418 37346 578654
rect 37582 578418 73026 578654
rect 73262 578418 73346 578654
rect 73582 578418 109026 578654
rect 109262 578418 109346 578654
rect 109582 578418 145026 578654
rect 145262 578418 145346 578654
rect 145582 578418 181026 578654
rect 181262 578418 181346 578654
rect 181582 578418 217026 578654
rect 217262 578418 217346 578654
rect 217582 578418 253026 578654
rect 253262 578418 253346 578654
rect 253582 578418 289026 578654
rect 289262 578418 289346 578654
rect 289582 578418 325026 578654
rect 325262 578418 325346 578654
rect 325582 578418 361026 578654
rect 361262 578418 361346 578654
rect 361582 578418 397026 578654
rect 397262 578418 397346 578654
rect 397582 578418 433026 578654
rect 433262 578418 433346 578654
rect 433582 578418 469026 578654
rect 469262 578418 469346 578654
rect 469582 578418 505026 578654
rect 505262 578418 505346 578654
rect 505582 578418 541026 578654
rect 541262 578418 541346 578654
rect 541582 578418 577026 578654
rect 577262 578418 577346 578654
rect 577582 578418 585342 578654
rect 585578 578418 585662 578654
rect 585898 578418 592650 578654
rect -8726 578334 592650 578418
rect -8726 578098 -1974 578334
rect -1738 578098 -1654 578334
rect -1418 578098 1026 578334
rect 1262 578098 1346 578334
rect 1582 578098 37026 578334
rect 37262 578098 37346 578334
rect 37582 578098 73026 578334
rect 73262 578098 73346 578334
rect 73582 578098 109026 578334
rect 109262 578098 109346 578334
rect 109582 578098 145026 578334
rect 145262 578098 145346 578334
rect 145582 578098 181026 578334
rect 181262 578098 181346 578334
rect 181582 578098 217026 578334
rect 217262 578098 217346 578334
rect 217582 578098 253026 578334
rect 253262 578098 253346 578334
rect 253582 578098 289026 578334
rect 289262 578098 289346 578334
rect 289582 578098 325026 578334
rect 325262 578098 325346 578334
rect 325582 578098 361026 578334
rect 361262 578098 361346 578334
rect 361582 578098 397026 578334
rect 397262 578098 397346 578334
rect 397582 578098 433026 578334
rect 433262 578098 433346 578334
rect 433582 578098 469026 578334
rect 469262 578098 469346 578334
rect 469582 578098 505026 578334
rect 505262 578098 505346 578334
rect 505582 578098 541026 578334
rect 541262 578098 541346 578334
rect 541582 578098 577026 578334
rect 577262 578098 577346 578334
rect 577582 578098 585342 578334
rect 585578 578098 585662 578334
rect 585898 578098 592650 578334
rect -8726 578066 592650 578098
rect -8726 551334 592650 551366
rect -8726 551098 -8694 551334
rect -8458 551098 -8374 551334
rect -8138 551098 9706 551334
rect 9942 551098 10026 551334
rect 10262 551098 45706 551334
rect 45942 551098 46026 551334
rect 46262 551098 81706 551334
rect 81942 551098 82026 551334
rect 82262 551098 117706 551334
rect 117942 551098 118026 551334
rect 118262 551098 153706 551334
rect 153942 551098 154026 551334
rect 154262 551098 189706 551334
rect 189942 551098 190026 551334
rect 190262 551098 225706 551334
rect 225942 551098 226026 551334
rect 226262 551098 261706 551334
rect 261942 551098 262026 551334
rect 262262 551098 297706 551334
rect 297942 551098 298026 551334
rect 298262 551098 333706 551334
rect 333942 551098 334026 551334
rect 334262 551098 369706 551334
rect 369942 551098 370026 551334
rect 370262 551098 405706 551334
rect 405942 551098 406026 551334
rect 406262 551098 441706 551334
rect 441942 551098 442026 551334
rect 442262 551098 477706 551334
rect 477942 551098 478026 551334
rect 478262 551098 513706 551334
rect 513942 551098 514026 551334
rect 514262 551098 549706 551334
rect 549942 551098 550026 551334
rect 550262 551098 592062 551334
rect 592298 551098 592382 551334
rect 592618 551098 592650 551334
rect -8726 551014 592650 551098
rect -8726 550778 -8694 551014
rect -8458 550778 -8374 551014
rect -8138 550778 9706 551014
rect 9942 550778 10026 551014
rect 10262 550778 45706 551014
rect 45942 550778 46026 551014
rect 46262 550778 81706 551014
rect 81942 550778 82026 551014
rect 82262 550778 117706 551014
rect 117942 550778 118026 551014
rect 118262 550778 153706 551014
rect 153942 550778 154026 551014
rect 154262 550778 189706 551014
rect 189942 550778 190026 551014
rect 190262 550778 225706 551014
rect 225942 550778 226026 551014
rect 226262 550778 261706 551014
rect 261942 550778 262026 551014
rect 262262 550778 297706 551014
rect 297942 550778 298026 551014
rect 298262 550778 333706 551014
rect 333942 550778 334026 551014
rect 334262 550778 369706 551014
rect 369942 550778 370026 551014
rect 370262 550778 405706 551014
rect 405942 550778 406026 551014
rect 406262 550778 441706 551014
rect 441942 550778 442026 551014
rect 442262 550778 477706 551014
rect 477942 550778 478026 551014
rect 478262 550778 513706 551014
rect 513942 550778 514026 551014
rect 514262 550778 549706 551014
rect 549942 550778 550026 551014
rect 550262 550778 592062 551014
rect 592298 550778 592382 551014
rect 592618 550778 592650 551014
rect -8726 550746 592650 550778
rect -8726 550094 592650 550126
rect -8726 549858 -7734 550094
rect -7498 549858 -7414 550094
rect -7178 549858 8466 550094
rect 8702 549858 8786 550094
rect 9022 549858 44466 550094
rect 44702 549858 44786 550094
rect 45022 549858 80466 550094
rect 80702 549858 80786 550094
rect 81022 549858 116466 550094
rect 116702 549858 116786 550094
rect 117022 549858 152466 550094
rect 152702 549858 152786 550094
rect 153022 549858 188466 550094
rect 188702 549858 188786 550094
rect 189022 549858 224466 550094
rect 224702 549858 224786 550094
rect 225022 549858 260466 550094
rect 260702 549858 260786 550094
rect 261022 549858 296466 550094
rect 296702 549858 296786 550094
rect 297022 549858 332466 550094
rect 332702 549858 332786 550094
rect 333022 549858 368466 550094
rect 368702 549858 368786 550094
rect 369022 549858 404466 550094
rect 404702 549858 404786 550094
rect 405022 549858 440466 550094
rect 440702 549858 440786 550094
rect 441022 549858 476466 550094
rect 476702 549858 476786 550094
rect 477022 549858 512466 550094
rect 512702 549858 512786 550094
rect 513022 549858 548466 550094
rect 548702 549858 548786 550094
rect 549022 549858 591102 550094
rect 591338 549858 591422 550094
rect 591658 549858 592650 550094
rect -8726 549774 592650 549858
rect -8726 549538 -7734 549774
rect -7498 549538 -7414 549774
rect -7178 549538 8466 549774
rect 8702 549538 8786 549774
rect 9022 549538 44466 549774
rect 44702 549538 44786 549774
rect 45022 549538 80466 549774
rect 80702 549538 80786 549774
rect 81022 549538 116466 549774
rect 116702 549538 116786 549774
rect 117022 549538 152466 549774
rect 152702 549538 152786 549774
rect 153022 549538 188466 549774
rect 188702 549538 188786 549774
rect 189022 549538 224466 549774
rect 224702 549538 224786 549774
rect 225022 549538 260466 549774
rect 260702 549538 260786 549774
rect 261022 549538 296466 549774
rect 296702 549538 296786 549774
rect 297022 549538 332466 549774
rect 332702 549538 332786 549774
rect 333022 549538 368466 549774
rect 368702 549538 368786 549774
rect 369022 549538 404466 549774
rect 404702 549538 404786 549774
rect 405022 549538 440466 549774
rect 440702 549538 440786 549774
rect 441022 549538 476466 549774
rect 476702 549538 476786 549774
rect 477022 549538 512466 549774
rect 512702 549538 512786 549774
rect 513022 549538 548466 549774
rect 548702 549538 548786 549774
rect 549022 549538 591102 549774
rect 591338 549538 591422 549774
rect 591658 549538 592650 549774
rect -8726 549506 592650 549538
rect -8726 548854 592650 548886
rect -8726 548618 -6774 548854
rect -6538 548618 -6454 548854
rect -6218 548618 7226 548854
rect 7462 548618 7546 548854
rect 7782 548618 43226 548854
rect 43462 548618 43546 548854
rect 43782 548618 79226 548854
rect 79462 548618 79546 548854
rect 79782 548618 115226 548854
rect 115462 548618 115546 548854
rect 115782 548618 151226 548854
rect 151462 548618 151546 548854
rect 151782 548618 187226 548854
rect 187462 548618 187546 548854
rect 187782 548618 223226 548854
rect 223462 548618 223546 548854
rect 223782 548618 259226 548854
rect 259462 548618 259546 548854
rect 259782 548618 295226 548854
rect 295462 548618 295546 548854
rect 295782 548618 331226 548854
rect 331462 548618 331546 548854
rect 331782 548618 367226 548854
rect 367462 548618 367546 548854
rect 367782 548618 403226 548854
rect 403462 548618 403546 548854
rect 403782 548618 439226 548854
rect 439462 548618 439546 548854
rect 439782 548618 475226 548854
rect 475462 548618 475546 548854
rect 475782 548618 511226 548854
rect 511462 548618 511546 548854
rect 511782 548618 547226 548854
rect 547462 548618 547546 548854
rect 547782 548618 590142 548854
rect 590378 548618 590462 548854
rect 590698 548618 592650 548854
rect -8726 548534 592650 548618
rect -8726 548298 -6774 548534
rect -6538 548298 -6454 548534
rect -6218 548298 7226 548534
rect 7462 548298 7546 548534
rect 7782 548298 43226 548534
rect 43462 548298 43546 548534
rect 43782 548298 79226 548534
rect 79462 548298 79546 548534
rect 79782 548298 115226 548534
rect 115462 548298 115546 548534
rect 115782 548298 151226 548534
rect 151462 548298 151546 548534
rect 151782 548298 187226 548534
rect 187462 548298 187546 548534
rect 187782 548298 223226 548534
rect 223462 548298 223546 548534
rect 223782 548298 259226 548534
rect 259462 548298 259546 548534
rect 259782 548298 295226 548534
rect 295462 548298 295546 548534
rect 295782 548298 331226 548534
rect 331462 548298 331546 548534
rect 331782 548298 367226 548534
rect 367462 548298 367546 548534
rect 367782 548298 403226 548534
rect 403462 548298 403546 548534
rect 403782 548298 439226 548534
rect 439462 548298 439546 548534
rect 439782 548298 475226 548534
rect 475462 548298 475546 548534
rect 475782 548298 511226 548534
rect 511462 548298 511546 548534
rect 511782 548298 547226 548534
rect 547462 548298 547546 548534
rect 547782 548298 590142 548534
rect 590378 548298 590462 548534
rect 590698 548298 592650 548534
rect -8726 548266 592650 548298
rect -8726 547614 592650 547646
rect -8726 547378 -5814 547614
rect -5578 547378 -5494 547614
rect -5258 547378 5986 547614
rect 6222 547378 6306 547614
rect 6542 547378 41986 547614
rect 42222 547378 42306 547614
rect 42542 547378 77986 547614
rect 78222 547378 78306 547614
rect 78542 547378 113986 547614
rect 114222 547378 114306 547614
rect 114542 547378 149986 547614
rect 150222 547378 150306 547614
rect 150542 547378 185986 547614
rect 186222 547378 186306 547614
rect 186542 547378 221986 547614
rect 222222 547378 222306 547614
rect 222542 547378 257986 547614
rect 258222 547378 258306 547614
rect 258542 547378 293986 547614
rect 294222 547378 294306 547614
rect 294542 547378 329986 547614
rect 330222 547378 330306 547614
rect 330542 547378 365986 547614
rect 366222 547378 366306 547614
rect 366542 547378 401986 547614
rect 402222 547378 402306 547614
rect 402542 547378 437986 547614
rect 438222 547378 438306 547614
rect 438542 547378 473986 547614
rect 474222 547378 474306 547614
rect 474542 547378 509986 547614
rect 510222 547378 510306 547614
rect 510542 547378 545986 547614
rect 546222 547378 546306 547614
rect 546542 547378 581986 547614
rect 582222 547378 582306 547614
rect 582542 547378 589182 547614
rect 589418 547378 589502 547614
rect 589738 547378 592650 547614
rect -8726 547294 592650 547378
rect -8726 547058 -5814 547294
rect -5578 547058 -5494 547294
rect -5258 547058 5986 547294
rect 6222 547058 6306 547294
rect 6542 547058 41986 547294
rect 42222 547058 42306 547294
rect 42542 547058 77986 547294
rect 78222 547058 78306 547294
rect 78542 547058 113986 547294
rect 114222 547058 114306 547294
rect 114542 547058 149986 547294
rect 150222 547058 150306 547294
rect 150542 547058 185986 547294
rect 186222 547058 186306 547294
rect 186542 547058 221986 547294
rect 222222 547058 222306 547294
rect 222542 547058 257986 547294
rect 258222 547058 258306 547294
rect 258542 547058 293986 547294
rect 294222 547058 294306 547294
rect 294542 547058 329986 547294
rect 330222 547058 330306 547294
rect 330542 547058 365986 547294
rect 366222 547058 366306 547294
rect 366542 547058 401986 547294
rect 402222 547058 402306 547294
rect 402542 547058 437986 547294
rect 438222 547058 438306 547294
rect 438542 547058 473986 547294
rect 474222 547058 474306 547294
rect 474542 547058 509986 547294
rect 510222 547058 510306 547294
rect 510542 547058 545986 547294
rect 546222 547058 546306 547294
rect 546542 547058 581986 547294
rect 582222 547058 582306 547294
rect 582542 547058 589182 547294
rect 589418 547058 589502 547294
rect 589738 547058 592650 547294
rect -8726 547026 592650 547058
rect -8726 546374 592650 546406
rect -8726 546138 -4854 546374
rect -4618 546138 -4534 546374
rect -4298 546138 4746 546374
rect 4982 546138 5066 546374
rect 5302 546138 40746 546374
rect 40982 546138 41066 546374
rect 41302 546138 76746 546374
rect 76982 546138 77066 546374
rect 77302 546138 112746 546374
rect 112982 546138 113066 546374
rect 113302 546138 148746 546374
rect 148982 546138 149066 546374
rect 149302 546138 184746 546374
rect 184982 546138 185066 546374
rect 185302 546138 220746 546374
rect 220982 546138 221066 546374
rect 221302 546138 256746 546374
rect 256982 546138 257066 546374
rect 257302 546138 292746 546374
rect 292982 546138 293066 546374
rect 293302 546138 328746 546374
rect 328982 546138 329066 546374
rect 329302 546138 364746 546374
rect 364982 546138 365066 546374
rect 365302 546138 400746 546374
rect 400982 546138 401066 546374
rect 401302 546138 436746 546374
rect 436982 546138 437066 546374
rect 437302 546138 472746 546374
rect 472982 546138 473066 546374
rect 473302 546138 508746 546374
rect 508982 546138 509066 546374
rect 509302 546138 544746 546374
rect 544982 546138 545066 546374
rect 545302 546138 580746 546374
rect 580982 546138 581066 546374
rect 581302 546138 588222 546374
rect 588458 546138 588542 546374
rect 588778 546138 592650 546374
rect -8726 546054 592650 546138
rect -8726 545818 -4854 546054
rect -4618 545818 -4534 546054
rect -4298 545818 4746 546054
rect 4982 545818 5066 546054
rect 5302 545818 40746 546054
rect 40982 545818 41066 546054
rect 41302 545818 76746 546054
rect 76982 545818 77066 546054
rect 77302 545818 112746 546054
rect 112982 545818 113066 546054
rect 113302 545818 148746 546054
rect 148982 545818 149066 546054
rect 149302 545818 184746 546054
rect 184982 545818 185066 546054
rect 185302 545818 220746 546054
rect 220982 545818 221066 546054
rect 221302 545818 256746 546054
rect 256982 545818 257066 546054
rect 257302 545818 292746 546054
rect 292982 545818 293066 546054
rect 293302 545818 328746 546054
rect 328982 545818 329066 546054
rect 329302 545818 364746 546054
rect 364982 545818 365066 546054
rect 365302 545818 400746 546054
rect 400982 545818 401066 546054
rect 401302 545818 436746 546054
rect 436982 545818 437066 546054
rect 437302 545818 472746 546054
rect 472982 545818 473066 546054
rect 473302 545818 508746 546054
rect 508982 545818 509066 546054
rect 509302 545818 544746 546054
rect 544982 545818 545066 546054
rect 545302 545818 580746 546054
rect 580982 545818 581066 546054
rect 581302 545818 588222 546054
rect 588458 545818 588542 546054
rect 588778 545818 592650 546054
rect -8726 545786 592650 545818
rect -8726 545134 592650 545166
rect -8726 544898 -3894 545134
rect -3658 544898 -3574 545134
rect -3338 544898 3506 545134
rect 3742 544898 3826 545134
rect 4062 544898 39506 545134
rect 39742 544898 39826 545134
rect 40062 544898 75506 545134
rect 75742 544898 75826 545134
rect 76062 544898 111506 545134
rect 111742 544898 111826 545134
rect 112062 544898 147506 545134
rect 147742 544898 147826 545134
rect 148062 544898 183506 545134
rect 183742 544898 183826 545134
rect 184062 544898 219506 545134
rect 219742 544898 219826 545134
rect 220062 544898 255506 545134
rect 255742 544898 255826 545134
rect 256062 544898 291506 545134
rect 291742 544898 291826 545134
rect 292062 544898 327506 545134
rect 327742 544898 327826 545134
rect 328062 544898 363506 545134
rect 363742 544898 363826 545134
rect 364062 544898 399506 545134
rect 399742 544898 399826 545134
rect 400062 544898 435506 545134
rect 435742 544898 435826 545134
rect 436062 544898 471506 545134
rect 471742 544898 471826 545134
rect 472062 544898 507506 545134
rect 507742 544898 507826 545134
rect 508062 544898 543506 545134
rect 543742 544898 543826 545134
rect 544062 544898 579506 545134
rect 579742 544898 579826 545134
rect 580062 544898 587262 545134
rect 587498 544898 587582 545134
rect 587818 544898 592650 545134
rect -8726 544814 592650 544898
rect -8726 544578 -3894 544814
rect -3658 544578 -3574 544814
rect -3338 544578 3506 544814
rect 3742 544578 3826 544814
rect 4062 544578 39506 544814
rect 39742 544578 39826 544814
rect 40062 544578 75506 544814
rect 75742 544578 75826 544814
rect 76062 544578 111506 544814
rect 111742 544578 111826 544814
rect 112062 544578 147506 544814
rect 147742 544578 147826 544814
rect 148062 544578 183506 544814
rect 183742 544578 183826 544814
rect 184062 544578 219506 544814
rect 219742 544578 219826 544814
rect 220062 544578 255506 544814
rect 255742 544578 255826 544814
rect 256062 544578 291506 544814
rect 291742 544578 291826 544814
rect 292062 544578 327506 544814
rect 327742 544578 327826 544814
rect 328062 544578 363506 544814
rect 363742 544578 363826 544814
rect 364062 544578 399506 544814
rect 399742 544578 399826 544814
rect 400062 544578 435506 544814
rect 435742 544578 435826 544814
rect 436062 544578 471506 544814
rect 471742 544578 471826 544814
rect 472062 544578 507506 544814
rect 507742 544578 507826 544814
rect 508062 544578 543506 544814
rect 543742 544578 543826 544814
rect 544062 544578 579506 544814
rect 579742 544578 579826 544814
rect 580062 544578 587262 544814
rect 587498 544578 587582 544814
rect 587818 544578 592650 544814
rect -8726 544546 592650 544578
rect -8726 543894 592650 543926
rect -8726 543658 -2934 543894
rect -2698 543658 -2614 543894
rect -2378 543658 2266 543894
rect 2502 543658 2586 543894
rect 2822 543658 38266 543894
rect 38502 543658 38586 543894
rect 38822 543658 74266 543894
rect 74502 543658 74586 543894
rect 74822 543658 110266 543894
rect 110502 543658 110586 543894
rect 110822 543658 146266 543894
rect 146502 543658 146586 543894
rect 146822 543658 182266 543894
rect 182502 543658 182586 543894
rect 182822 543658 218266 543894
rect 218502 543658 218586 543894
rect 218822 543658 254266 543894
rect 254502 543658 254586 543894
rect 254822 543658 290266 543894
rect 290502 543658 290586 543894
rect 290822 543658 326266 543894
rect 326502 543658 326586 543894
rect 326822 543658 362266 543894
rect 362502 543658 362586 543894
rect 362822 543658 398266 543894
rect 398502 543658 398586 543894
rect 398822 543658 434266 543894
rect 434502 543658 434586 543894
rect 434822 543658 470266 543894
rect 470502 543658 470586 543894
rect 470822 543658 506266 543894
rect 506502 543658 506586 543894
rect 506822 543658 542266 543894
rect 542502 543658 542586 543894
rect 542822 543658 578266 543894
rect 578502 543658 578586 543894
rect 578822 543658 586302 543894
rect 586538 543658 586622 543894
rect 586858 543658 592650 543894
rect -8726 543574 592650 543658
rect -8726 543338 -2934 543574
rect -2698 543338 -2614 543574
rect -2378 543338 2266 543574
rect 2502 543338 2586 543574
rect 2822 543338 38266 543574
rect 38502 543338 38586 543574
rect 38822 543338 74266 543574
rect 74502 543338 74586 543574
rect 74822 543338 110266 543574
rect 110502 543338 110586 543574
rect 110822 543338 146266 543574
rect 146502 543338 146586 543574
rect 146822 543338 182266 543574
rect 182502 543338 182586 543574
rect 182822 543338 218266 543574
rect 218502 543338 218586 543574
rect 218822 543338 254266 543574
rect 254502 543338 254586 543574
rect 254822 543338 290266 543574
rect 290502 543338 290586 543574
rect 290822 543338 326266 543574
rect 326502 543338 326586 543574
rect 326822 543338 362266 543574
rect 362502 543338 362586 543574
rect 362822 543338 398266 543574
rect 398502 543338 398586 543574
rect 398822 543338 434266 543574
rect 434502 543338 434586 543574
rect 434822 543338 470266 543574
rect 470502 543338 470586 543574
rect 470822 543338 506266 543574
rect 506502 543338 506586 543574
rect 506822 543338 542266 543574
rect 542502 543338 542586 543574
rect 542822 543338 578266 543574
rect 578502 543338 578586 543574
rect 578822 543338 586302 543574
rect 586538 543338 586622 543574
rect 586858 543338 592650 543574
rect -8726 543306 592650 543338
rect -8726 542654 592650 542686
rect -8726 542418 -1974 542654
rect -1738 542418 -1654 542654
rect -1418 542418 1026 542654
rect 1262 542418 1346 542654
rect 1582 542418 37026 542654
rect 37262 542418 37346 542654
rect 37582 542418 73026 542654
rect 73262 542418 73346 542654
rect 73582 542418 109026 542654
rect 109262 542418 109346 542654
rect 109582 542418 145026 542654
rect 145262 542418 145346 542654
rect 145582 542418 181026 542654
rect 181262 542418 181346 542654
rect 181582 542418 217026 542654
rect 217262 542418 217346 542654
rect 217582 542418 253026 542654
rect 253262 542418 253346 542654
rect 253582 542418 289026 542654
rect 289262 542418 289346 542654
rect 289582 542418 325026 542654
rect 325262 542418 325346 542654
rect 325582 542418 361026 542654
rect 361262 542418 361346 542654
rect 361582 542418 397026 542654
rect 397262 542418 397346 542654
rect 397582 542418 433026 542654
rect 433262 542418 433346 542654
rect 433582 542418 469026 542654
rect 469262 542418 469346 542654
rect 469582 542418 505026 542654
rect 505262 542418 505346 542654
rect 505582 542418 541026 542654
rect 541262 542418 541346 542654
rect 541582 542418 577026 542654
rect 577262 542418 577346 542654
rect 577582 542418 585342 542654
rect 585578 542418 585662 542654
rect 585898 542418 592650 542654
rect -8726 542334 592650 542418
rect -8726 542098 -1974 542334
rect -1738 542098 -1654 542334
rect -1418 542098 1026 542334
rect 1262 542098 1346 542334
rect 1582 542098 37026 542334
rect 37262 542098 37346 542334
rect 37582 542098 73026 542334
rect 73262 542098 73346 542334
rect 73582 542098 109026 542334
rect 109262 542098 109346 542334
rect 109582 542098 145026 542334
rect 145262 542098 145346 542334
rect 145582 542098 181026 542334
rect 181262 542098 181346 542334
rect 181582 542098 217026 542334
rect 217262 542098 217346 542334
rect 217582 542098 253026 542334
rect 253262 542098 253346 542334
rect 253582 542098 289026 542334
rect 289262 542098 289346 542334
rect 289582 542098 325026 542334
rect 325262 542098 325346 542334
rect 325582 542098 361026 542334
rect 361262 542098 361346 542334
rect 361582 542098 397026 542334
rect 397262 542098 397346 542334
rect 397582 542098 433026 542334
rect 433262 542098 433346 542334
rect 433582 542098 469026 542334
rect 469262 542098 469346 542334
rect 469582 542098 505026 542334
rect 505262 542098 505346 542334
rect 505582 542098 541026 542334
rect 541262 542098 541346 542334
rect 541582 542098 577026 542334
rect 577262 542098 577346 542334
rect 577582 542098 585342 542334
rect 585578 542098 585662 542334
rect 585898 542098 592650 542334
rect -8726 542066 592650 542098
rect -8726 515334 592650 515366
rect -8726 515098 -8694 515334
rect -8458 515098 -8374 515334
rect -8138 515098 9706 515334
rect 9942 515098 10026 515334
rect 10262 515098 45706 515334
rect 45942 515098 46026 515334
rect 46262 515098 81706 515334
rect 81942 515098 82026 515334
rect 82262 515098 117706 515334
rect 117942 515098 118026 515334
rect 118262 515098 153706 515334
rect 153942 515098 154026 515334
rect 154262 515098 189706 515334
rect 189942 515098 190026 515334
rect 190262 515098 225706 515334
rect 225942 515098 226026 515334
rect 226262 515098 261706 515334
rect 261942 515098 262026 515334
rect 262262 515098 297706 515334
rect 297942 515098 298026 515334
rect 298262 515098 333706 515334
rect 333942 515098 334026 515334
rect 334262 515098 369706 515334
rect 369942 515098 370026 515334
rect 370262 515098 405706 515334
rect 405942 515098 406026 515334
rect 406262 515098 441706 515334
rect 441942 515098 442026 515334
rect 442262 515098 477706 515334
rect 477942 515098 478026 515334
rect 478262 515098 513706 515334
rect 513942 515098 514026 515334
rect 514262 515098 549706 515334
rect 549942 515098 550026 515334
rect 550262 515098 592062 515334
rect 592298 515098 592382 515334
rect 592618 515098 592650 515334
rect -8726 515014 592650 515098
rect -8726 514778 -8694 515014
rect -8458 514778 -8374 515014
rect -8138 514778 9706 515014
rect 9942 514778 10026 515014
rect 10262 514778 45706 515014
rect 45942 514778 46026 515014
rect 46262 514778 81706 515014
rect 81942 514778 82026 515014
rect 82262 514778 117706 515014
rect 117942 514778 118026 515014
rect 118262 514778 153706 515014
rect 153942 514778 154026 515014
rect 154262 514778 189706 515014
rect 189942 514778 190026 515014
rect 190262 514778 225706 515014
rect 225942 514778 226026 515014
rect 226262 514778 261706 515014
rect 261942 514778 262026 515014
rect 262262 514778 297706 515014
rect 297942 514778 298026 515014
rect 298262 514778 333706 515014
rect 333942 514778 334026 515014
rect 334262 514778 369706 515014
rect 369942 514778 370026 515014
rect 370262 514778 405706 515014
rect 405942 514778 406026 515014
rect 406262 514778 441706 515014
rect 441942 514778 442026 515014
rect 442262 514778 477706 515014
rect 477942 514778 478026 515014
rect 478262 514778 513706 515014
rect 513942 514778 514026 515014
rect 514262 514778 549706 515014
rect 549942 514778 550026 515014
rect 550262 514778 592062 515014
rect 592298 514778 592382 515014
rect 592618 514778 592650 515014
rect -8726 514746 592650 514778
rect -8726 514094 592650 514126
rect -8726 513858 -7734 514094
rect -7498 513858 -7414 514094
rect -7178 513858 8466 514094
rect 8702 513858 8786 514094
rect 9022 513858 44466 514094
rect 44702 513858 44786 514094
rect 45022 513858 80466 514094
rect 80702 513858 80786 514094
rect 81022 513858 116466 514094
rect 116702 513858 116786 514094
rect 117022 513858 152466 514094
rect 152702 513858 152786 514094
rect 153022 513858 188466 514094
rect 188702 513858 188786 514094
rect 189022 513858 224466 514094
rect 224702 513858 224786 514094
rect 225022 513858 260466 514094
rect 260702 513858 260786 514094
rect 261022 513858 296466 514094
rect 296702 513858 296786 514094
rect 297022 513858 332466 514094
rect 332702 513858 332786 514094
rect 333022 513858 368466 514094
rect 368702 513858 368786 514094
rect 369022 513858 404466 514094
rect 404702 513858 404786 514094
rect 405022 513858 440466 514094
rect 440702 513858 440786 514094
rect 441022 513858 476466 514094
rect 476702 513858 476786 514094
rect 477022 513858 512466 514094
rect 512702 513858 512786 514094
rect 513022 513858 548466 514094
rect 548702 513858 548786 514094
rect 549022 513858 591102 514094
rect 591338 513858 591422 514094
rect 591658 513858 592650 514094
rect -8726 513774 592650 513858
rect -8726 513538 -7734 513774
rect -7498 513538 -7414 513774
rect -7178 513538 8466 513774
rect 8702 513538 8786 513774
rect 9022 513538 44466 513774
rect 44702 513538 44786 513774
rect 45022 513538 80466 513774
rect 80702 513538 80786 513774
rect 81022 513538 116466 513774
rect 116702 513538 116786 513774
rect 117022 513538 152466 513774
rect 152702 513538 152786 513774
rect 153022 513538 188466 513774
rect 188702 513538 188786 513774
rect 189022 513538 224466 513774
rect 224702 513538 224786 513774
rect 225022 513538 260466 513774
rect 260702 513538 260786 513774
rect 261022 513538 296466 513774
rect 296702 513538 296786 513774
rect 297022 513538 332466 513774
rect 332702 513538 332786 513774
rect 333022 513538 368466 513774
rect 368702 513538 368786 513774
rect 369022 513538 404466 513774
rect 404702 513538 404786 513774
rect 405022 513538 440466 513774
rect 440702 513538 440786 513774
rect 441022 513538 476466 513774
rect 476702 513538 476786 513774
rect 477022 513538 512466 513774
rect 512702 513538 512786 513774
rect 513022 513538 548466 513774
rect 548702 513538 548786 513774
rect 549022 513538 591102 513774
rect 591338 513538 591422 513774
rect 591658 513538 592650 513774
rect -8726 513506 592650 513538
rect -8726 512854 592650 512886
rect -8726 512618 -6774 512854
rect -6538 512618 -6454 512854
rect -6218 512618 7226 512854
rect 7462 512618 7546 512854
rect 7782 512618 43226 512854
rect 43462 512618 43546 512854
rect 43782 512618 79226 512854
rect 79462 512618 79546 512854
rect 79782 512618 115226 512854
rect 115462 512618 115546 512854
rect 115782 512618 151226 512854
rect 151462 512618 151546 512854
rect 151782 512618 187226 512854
rect 187462 512618 187546 512854
rect 187782 512618 223226 512854
rect 223462 512618 223546 512854
rect 223782 512618 259226 512854
rect 259462 512618 259546 512854
rect 259782 512618 295226 512854
rect 295462 512618 295546 512854
rect 295782 512618 331226 512854
rect 331462 512618 331546 512854
rect 331782 512618 367226 512854
rect 367462 512618 367546 512854
rect 367782 512618 403226 512854
rect 403462 512618 403546 512854
rect 403782 512618 439226 512854
rect 439462 512618 439546 512854
rect 439782 512618 475226 512854
rect 475462 512618 475546 512854
rect 475782 512618 511226 512854
rect 511462 512618 511546 512854
rect 511782 512618 547226 512854
rect 547462 512618 547546 512854
rect 547782 512618 590142 512854
rect 590378 512618 590462 512854
rect 590698 512618 592650 512854
rect -8726 512534 592650 512618
rect -8726 512298 -6774 512534
rect -6538 512298 -6454 512534
rect -6218 512298 7226 512534
rect 7462 512298 7546 512534
rect 7782 512298 43226 512534
rect 43462 512298 43546 512534
rect 43782 512298 79226 512534
rect 79462 512298 79546 512534
rect 79782 512298 115226 512534
rect 115462 512298 115546 512534
rect 115782 512298 151226 512534
rect 151462 512298 151546 512534
rect 151782 512298 187226 512534
rect 187462 512298 187546 512534
rect 187782 512298 223226 512534
rect 223462 512298 223546 512534
rect 223782 512298 259226 512534
rect 259462 512298 259546 512534
rect 259782 512298 295226 512534
rect 295462 512298 295546 512534
rect 295782 512298 331226 512534
rect 331462 512298 331546 512534
rect 331782 512298 367226 512534
rect 367462 512298 367546 512534
rect 367782 512298 403226 512534
rect 403462 512298 403546 512534
rect 403782 512298 439226 512534
rect 439462 512298 439546 512534
rect 439782 512298 475226 512534
rect 475462 512298 475546 512534
rect 475782 512298 511226 512534
rect 511462 512298 511546 512534
rect 511782 512298 547226 512534
rect 547462 512298 547546 512534
rect 547782 512298 590142 512534
rect 590378 512298 590462 512534
rect 590698 512298 592650 512534
rect -8726 512266 592650 512298
rect -8726 511614 592650 511646
rect -8726 511378 -5814 511614
rect -5578 511378 -5494 511614
rect -5258 511378 5986 511614
rect 6222 511378 6306 511614
rect 6542 511378 41986 511614
rect 42222 511378 42306 511614
rect 42542 511378 77986 511614
rect 78222 511378 78306 511614
rect 78542 511378 113986 511614
rect 114222 511378 114306 511614
rect 114542 511378 149986 511614
rect 150222 511378 150306 511614
rect 150542 511378 185986 511614
rect 186222 511378 186306 511614
rect 186542 511378 221986 511614
rect 222222 511378 222306 511614
rect 222542 511378 257986 511614
rect 258222 511378 258306 511614
rect 258542 511378 293986 511614
rect 294222 511378 294306 511614
rect 294542 511378 329986 511614
rect 330222 511378 330306 511614
rect 330542 511378 365986 511614
rect 366222 511378 366306 511614
rect 366542 511378 401986 511614
rect 402222 511378 402306 511614
rect 402542 511378 437986 511614
rect 438222 511378 438306 511614
rect 438542 511378 473986 511614
rect 474222 511378 474306 511614
rect 474542 511378 509986 511614
rect 510222 511378 510306 511614
rect 510542 511378 545986 511614
rect 546222 511378 546306 511614
rect 546542 511378 581986 511614
rect 582222 511378 582306 511614
rect 582542 511378 589182 511614
rect 589418 511378 589502 511614
rect 589738 511378 592650 511614
rect -8726 511294 592650 511378
rect -8726 511058 -5814 511294
rect -5578 511058 -5494 511294
rect -5258 511058 5986 511294
rect 6222 511058 6306 511294
rect 6542 511058 41986 511294
rect 42222 511058 42306 511294
rect 42542 511058 77986 511294
rect 78222 511058 78306 511294
rect 78542 511058 113986 511294
rect 114222 511058 114306 511294
rect 114542 511058 149986 511294
rect 150222 511058 150306 511294
rect 150542 511058 185986 511294
rect 186222 511058 186306 511294
rect 186542 511058 221986 511294
rect 222222 511058 222306 511294
rect 222542 511058 257986 511294
rect 258222 511058 258306 511294
rect 258542 511058 293986 511294
rect 294222 511058 294306 511294
rect 294542 511058 329986 511294
rect 330222 511058 330306 511294
rect 330542 511058 365986 511294
rect 366222 511058 366306 511294
rect 366542 511058 401986 511294
rect 402222 511058 402306 511294
rect 402542 511058 437986 511294
rect 438222 511058 438306 511294
rect 438542 511058 473986 511294
rect 474222 511058 474306 511294
rect 474542 511058 509986 511294
rect 510222 511058 510306 511294
rect 510542 511058 545986 511294
rect 546222 511058 546306 511294
rect 546542 511058 581986 511294
rect 582222 511058 582306 511294
rect 582542 511058 589182 511294
rect 589418 511058 589502 511294
rect 589738 511058 592650 511294
rect -8726 511026 592650 511058
rect -8726 510374 592650 510406
rect -8726 510138 -4854 510374
rect -4618 510138 -4534 510374
rect -4298 510138 4746 510374
rect 4982 510138 5066 510374
rect 5302 510138 40746 510374
rect 40982 510138 41066 510374
rect 41302 510138 76746 510374
rect 76982 510138 77066 510374
rect 77302 510138 112746 510374
rect 112982 510138 113066 510374
rect 113302 510138 148746 510374
rect 148982 510138 149066 510374
rect 149302 510138 184746 510374
rect 184982 510138 185066 510374
rect 185302 510138 220746 510374
rect 220982 510138 221066 510374
rect 221302 510138 256746 510374
rect 256982 510138 257066 510374
rect 257302 510138 292746 510374
rect 292982 510138 293066 510374
rect 293302 510138 328746 510374
rect 328982 510138 329066 510374
rect 329302 510138 364746 510374
rect 364982 510138 365066 510374
rect 365302 510138 400746 510374
rect 400982 510138 401066 510374
rect 401302 510138 436746 510374
rect 436982 510138 437066 510374
rect 437302 510138 472746 510374
rect 472982 510138 473066 510374
rect 473302 510138 508746 510374
rect 508982 510138 509066 510374
rect 509302 510138 544746 510374
rect 544982 510138 545066 510374
rect 545302 510138 580746 510374
rect 580982 510138 581066 510374
rect 581302 510138 588222 510374
rect 588458 510138 588542 510374
rect 588778 510138 592650 510374
rect -8726 510054 592650 510138
rect -8726 509818 -4854 510054
rect -4618 509818 -4534 510054
rect -4298 509818 4746 510054
rect 4982 509818 5066 510054
rect 5302 509818 40746 510054
rect 40982 509818 41066 510054
rect 41302 509818 76746 510054
rect 76982 509818 77066 510054
rect 77302 509818 112746 510054
rect 112982 509818 113066 510054
rect 113302 509818 148746 510054
rect 148982 509818 149066 510054
rect 149302 509818 184746 510054
rect 184982 509818 185066 510054
rect 185302 509818 220746 510054
rect 220982 509818 221066 510054
rect 221302 509818 256746 510054
rect 256982 509818 257066 510054
rect 257302 509818 292746 510054
rect 292982 509818 293066 510054
rect 293302 509818 328746 510054
rect 328982 509818 329066 510054
rect 329302 509818 364746 510054
rect 364982 509818 365066 510054
rect 365302 509818 400746 510054
rect 400982 509818 401066 510054
rect 401302 509818 436746 510054
rect 436982 509818 437066 510054
rect 437302 509818 472746 510054
rect 472982 509818 473066 510054
rect 473302 509818 508746 510054
rect 508982 509818 509066 510054
rect 509302 509818 544746 510054
rect 544982 509818 545066 510054
rect 545302 509818 580746 510054
rect 580982 509818 581066 510054
rect 581302 509818 588222 510054
rect 588458 509818 588542 510054
rect 588778 509818 592650 510054
rect -8726 509786 592650 509818
rect -8726 509134 592650 509166
rect -8726 508898 -3894 509134
rect -3658 508898 -3574 509134
rect -3338 508898 3506 509134
rect 3742 508898 3826 509134
rect 4062 508898 39506 509134
rect 39742 508898 39826 509134
rect 40062 508898 75506 509134
rect 75742 508898 75826 509134
rect 76062 508898 111506 509134
rect 111742 508898 111826 509134
rect 112062 508898 147506 509134
rect 147742 508898 147826 509134
rect 148062 508898 183506 509134
rect 183742 508898 183826 509134
rect 184062 508898 219506 509134
rect 219742 508898 219826 509134
rect 220062 508898 255506 509134
rect 255742 508898 255826 509134
rect 256062 508898 291506 509134
rect 291742 508898 291826 509134
rect 292062 508898 327506 509134
rect 327742 508898 327826 509134
rect 328062 508898 363506 509134
rect 363742 508898 363826 509134
rect 364062 508898 399506 509134
rect 399742 508898 399826 509134
rect 400062 508898 435506 509134
rect 435742 508898 435826 509134
rect 436062 508898 471506 509134
rect 471742 508898 471826 509134
rect 472062 508898 507506 509134
rect 507742 508898 507826 509134
rect 508062 508898 543506 509134
rect 543742 508898 543826 509134
rect 544062 508898 579506 509134
rect 579742 508898 579826 509134
rect 580062 508898 587262 509134
rect 587498 508898 587582 509134
rect 587818 508898 592650 509134
rect -8726 508814 592650 508898
rect -8726 508578 -3894 508814
rect -3658 508578 -3574 508814
rect -3338 508578 3506 508814
rect 3742 508578 3826 508814
rect 4062 508578 39506 508814
rect 39742 508578 39826 508814
rect 40062 508578 75506 508814
rect 75742 508578 75826 508814
rect 76062 508578 111506 508814
rect 111742 508578 111826 508814
rect 112062 508578 147506 508814
rect 147742 508578 147826 508814
rect 148062 508578 183506 508814
rect 183742 508578 183826 508814
rect 184062 508578 219506 508814
rect 219742 508578 219826 508814
rect 220062 508578 255506 508814
rect 255742 508578 255826 508814
rect 256062 508578 291506 508814
rect 291742 508578 291826 508814
rect 292062 508578 327506 508814
rect 327742 508578 327826 508814
rect 328062 508578 363506 508814
rect 363742 508578 363826 508814
rect 364062 508578 399506 508814
rect 399742 508578 399826 508814
rect 400062 508578 435506 508814
rect 435742 508578 435826 508814
rect 436062 508578 471506 508814
rect 471742 508578 471826 508814
rect 472062 508578 507506 508814
rect 507742 508578 507826 508814
rect 508062 508578 543506 508814
rect 543742 508578 543826 508814
rect 544062 508578 579506 508814
rect 579742 508578 579826 508814
rect 580062 508578 587262 508814
rect 587498 508578 587582 508814
rect 587818 508578 592650 508814
rect -8726 508546 592650 508578
rect -8726 507894 592650 507926
rect -8726 507658 -2934 507894
rect -2698 507658 -2614 507894
rect -2378 507658 2266 507894
rect 2502 507658 2586 507894
rect 2822 507658 38266 507894
rect 38502 507658 38586 507894
rect 38822 507658 74266 507894
rect 74502 507658 74586 507894
rect 74822 507658 110266 507894
rect 110502 507658 110586 507894
rect 110822 507658 146266 507894
rect 146502 507658 146586 507894
rect 146822 507658 182266 507894
rect 182502 507658 182586 507894
rect 182822 507658 218266 507894
rect 218502 507658 218586 507894
rect 218822 507658 254266 507894
rect 254502 507658 254586 507894
rect 254822 507658 290266 507894
rect 290502 507658 290586 507894
rect 290822 507658 326266 507894
rect 326502 507658 326586 507894
rect 326822 507658 362266 507894
rect 362502 507658 362586 507894
rect 362822 507658 398266 507894
rect 398502 507658 398586 507894
rect 398822 507658 434266 507894
rect 434502 507658 434586 507894
rect 434822 507658 470266 507894
rect 470502 507658 470586 507894
rect 470822 507658 506266 507894
rect 506502 507658 506586 507894
rect 506822 507658 542266 507894
rect 542502 507658 542586 507894
rect 542822 507658 578266 507894
rect 578502 507658 578586 507894
rect 578822 507658 586302 507894
rect 586538 507658 586622 507894
rect 586858 507658 592650 507894
rect -8726 507574 592650 507658
rect -8726 507338 -2934 507574
rect -2698 507338 -2614 507574
rect -2378 507338 2266 507574
rect 2502 507338 2586 507574
rect 2822 507338 38266 507574
rect 38502 507338 38586 507574
rect 38822 507338 74266 507574
rect 74502 507338 74586 507574
rect 74822 507338 110266 507574
rect 110502 507338 110586 507574
rect 110822 507338 146266 507574
rect 146502 507338 146586 507574
rect 146822 507338 182266 507574
rect 182502 507338 182586 507574
rect 182822 507338 218266 507574
rect 218502 507338 218586 507574
rect 218822 507338 254266 507574
rect 254502 507338 254586 507574
rect 254822 507338 290266 507574
rect 290502 507338 290586 507574
rect 290822 507338 326266 507574
rect 326502 507338 326586 507574
rect 326822 507338 362266 507574
rect 362502 507338 362586 507574
rect 362822 507338 398266 507574
rect 398502 507338 398586 507574
rect 398822 507338 434266 507574
rect 434502 507338 434586 507574
rect 434822 507338 470266 507574
rect 470502 507338 470586 507574
rect 470822 507338 506266 507574
rect 506502 507338 506586 507574
rect 506822 507338 542266 507574
rect 542502 507338 542586 507574
rect 542822 507338 578266 507574
rect 578502 507338 578586 507574
rect 578822 507338 586302 507574
rect 586538 507338 586622 507574
rect 586858 507338 592650 507574
rect -8726 507306 592650 507338
rect -8726 506654 592650 506686
rect -8726 506418 -1974 506654
rect -1738 506418 -1654 506654
rect -1418 506418 1026 506654
rect 1262 506418 1346 506654
rect 1582 506418 37026 506654
rect 37262 506418 37346 506654
rect 37582 506418 73026 506654
rect 73262 506418 73346 506654
rect 73582 506418 109026 506654
rect 109262 506418 109346 506654
rect 109582 506418 145026 506654
rect 145262 506418 145346 506654
rect 145582 506418 181026 506654
rect 181262 506418 181346 506654
rect 181582 506418 217026 506654
rect 217262 506418 217346 506654
rect 217582 506418 253026 506654
rect 253262 506418 253346 506654
rect 253582 506418 289026 506654
rect 289262 506418 289346 506654
rect 289582 506418 325026 506654
rect 325262 506418 325346 506654
rect 325582 506418 361026 506654
rect 361262 506418 361346 506654
rect 361582 506418 397026 506654
rect 397262 506418 397346 506654
rect 397582 506418 433026 506654
rect 433262 506418 433346 506654
rect 433582 506418 469026 506654
rect 469262 506418 469346 506654
rect 469582 506418 505026 506654
rect 505262 506418 505346 506654
rect 505582 506418 541026 506654
rect 541262 506418 541346 506654
rect 541582 506418 577026 506654
rect 577262 506418 577346 506654
rect 577582 506418 585342 506654
rect 585578 506418 585662 506654
rect 585898 506418 592650 506654
rect -8726 506334 592650 506418
rect -8726 506098 -1974 506334
rect -1738 506098 -1654 506334
rect -1418 506098 1026 506334
rect 1262 506098 1346 506334
rect 1582 506098 37026 506334
rect 37262 506098 37346 506334
rect 37582 506098 73026 506334
rect 73262 506098 73346 506334
rect 73582 506098 109026 506334
rect 109262 506098 109346 506334
rect 109582 506098 145026 506334
rect 145262 506098 145346 506334
rect 145582 506098 181026 506334
rect 181262 506098 181346 506334
rect 181582 506098 217026 506334
rect 217262 506098 217346 506334
rect 217582 506098 253026 506334
rect 253262 506098 253346 506334
rect 253582 506098 289026 506334
rect 289262 506098 289346 506334
rect 289582 506098 325026 506334
rect 325262 506098 325346 506334
rect 325582 506098 361026 506334
rect 361262 506098 361346 506334
rect 361582 506098 397026 506334
rect 397262 506098 397346 506334
rect 397582 506098 433026 506334
rect 433262 506098 433346 506334
rect 433582 506098 469026 506334
rect 469262 506098 469346 506334
rect 469582 506098 505026 506334
rect 505262 506098 505346 506334
rect 505582 506098 541026 506334
rect 541262 506098 541346 506334
rect 541582 506098 577026 506334
rect 577262 506098 577346 506334
rect 577582 506098 585342 506334
rect 585578 506098 585662 506334
rect 585898 506098 592650 506334
rect -8726 506066 592650 506098
rect -8726 479334 592650 479366
rect -8726 479098 -8694 479334
rect -8458 479098 -8374 479334
rect -8138 479098 9706 479334
rect 9942 479098 10026 479334
rect 10262 479098 45706 479334
rect 45942 479098 46026 479334
rect 46262 479098 81706 479334
rect 81942 479098 82026 479334
rect 82262 479098 117706 479334
rect 117942 479098 118026 479334
rect 118262 479098 153706 479334
rect 153942 479098 154026 479334
rect 154262 479098 189706 479334
rect 189942 479098 190026 479334
rect 190262 479098 225706 479334
rect 225942 479098 226026 479334
rect 226262 479098 261706 479334
rect 261942 479098 262026 479334
rect 262262 479098 297706 479334
rect 297942 479098 298026 479334
rect 298262 479098 333706 479334
rect 333942 479098 334026 479334
rect 334262 479098 369706 479334
rect 369942 479098 370026 479334
rect 370262 479098 405706 479334
rect 405942 479098 406026 479334
rect 406262 479098 441706 479334
rect 441942 479098 442026 479334
rect 442262 479098 477706 479334
rect 477942 479098 478026 479334
rect 478262 479098 513706 479334
rect 513942 479098 514026 479334
rect 514262 479098 549706 479334
rect 549942 479098 550026 479334
rect 550262 479098 592062 479334
rect 592298 479098 592382 479334
rect 592618 479098 592650 479334
rect -8726 479014 592650 479098
rect -8726 478778 -8694 479014
rect -8458 478778 -8374 479014
rect -8138 478778 9706 479014
rect 9942 478778 10026 479014
rect 10262 478778 45706 479014
rect 45942 478778 46026 479014
rect 46262 478778 81706 479014
rect 81942 478778 82026 479014
rect 82262 478778 117706 479014
rect 117942 478778 118026 479014
rect 118262 478778 153706 479014
rect 153942 478778 154026 479014
rect 154262 478778 189706 479014
rect 189942 478778 190026 479014
rect 190262 478778 225706 479014
rect 225942 478778 226026 479014
rect 226262 478778 261706 479014
rect 261942 478778 262026 479014
rect 262262 478778 297706 479014
rect 297942 478778 298026 479014
rect 298262 478778 333706 479014
rect 333942 478778 334026 479014
rect 334262 478778 369706 479014
rect 369942 478778 370026 479014
rect 370262 478778 405706 479014
rect 405942 478778 406026 479014
rect 406262 478778 441706 479014
rect 441942 478778 442026 479014
rect 442262 478778 477706 479014
rect 477942 478778 478026 479014
rect 478262 478778 513706 479014
rect 513942 478778 514026 479014
rect 514262 478778 549706 479014
rect 549942 478778 550026 479014
rect 550262 478778 592062 479014
rect 592298 478778 592382 479014
rect 592618 478778 592650 479014
rect -8726 478746 592650 478778
rect -8726 478094 592650 478126
rect -8726 477858 -7734 478094
rect -7498 477858 -7414 478094
rect -7178 477858 8466 478094
rect 8702 477858 8786 478094
rect 9022 477858 44466 478094
rect 44702 477858 44786 478094
rect 45022 477858 80466 478094
rect 80702 477858 80786 478094
rect 81022 477858 116466 478094
rect 116702 477858 116786 478094
rect 117022 477858 152466 478094
rect 152702 477858 152786 478094
rect 153022 477858 188466 478094
rect 188702 477858 188786 478094
rect 189022 477858 224466 478094
rect 224702 477858 224786 478094
rect 225022 477858 260466 478094
rect 260702 477858 260786 478094
rect 261022 477858 296466 478094
rect 296702 477858 296786 478094
rect 297022 477858 332466 478094
rect 332702 477858 332786 478094
rect 333022 477858 368466 478094
rect 368702 477858 368786 478094
rect 369022 477858 404466 478094
rect 404702 477858 404786 478094
rect 405022 477858 440466 478094
rect 440702 477858 440786 478094
rect 441022 477858 476466 478094
rect 476702 477858 476786 478094
rect 477022 477858 512466 478094
rect 512702 477858 512786 478094
rect 513022 477858 548466 478094
rect 548702 477858 548786 478094
rect 549022 477858 591102 478094
rect 591338 477858 591422 478094
rect 591658 477858 592650 478094
rect -8726 477774 592650 477858
rect -8726 477538 -7734 477774
rect -7498 477538 -7414 477774
rect -7178 477538 8466 477774
rect 8702 477538 8786 477774
rect 9022 477538 44466 477774
rect 44702 477538 44786 477774
rect 45022 477538 80466 477774
rect 80702 477538 80786 477774
rect 81022 477538 116466 477774
rect 116702 477538 116786 477774
rect 117022 477538 152466 477774
rect 152702 477538 152786 477774
rect 153022 477538 188466 477774
rect 188702 477538 188786 477774
rect 189022 477538 224466 477774
rect 224702 477538 224786 477774
rect 225022 477538 260466 477774
rect 260702 477538 260786 477774
rect 261022 477538 296466 477774
rect 296702 477538 296786 477774
rect 297022 477538 332466 477774
rect 332702 477538 332786 477774
rect 333022 477538 368466 477774
rect 368702 477538 368786 477774
rect 369022 477538 404466 477774
rect 404702 477538 404786 477774
rect 405022 477538 440466 477774
rect 440702 477538 440786 477774
rect 441022 477538 476466 477774
rect 476702 477538 476786 477774
rect 477022 477538 512466 477774
rect 512702 477538 512786 477774
rect 513022 477538 548466 477774
rect 548702 477538 548786 477774
rect 549022 477538 591102 477774
rect 591338 477538 591422 477774
rect 591658 477538 592650 477774
rect -8726 477506 592650 477538
rect -8726 476854 592650 476886
rect -8726 476618 -6774 476854
rect -6538 476618 -6454 476854
rect -6218 476618 7226 476854
rect 7462 476618 7546 476854
rect 7782 476618 43226 476854
rect 43462 476618 43546 476854
rect 43782 476618 79226 476854
rect 79462 476618 79546 476854
rect 79782 476618 115226 476854
rect 115462 476618 115546 476854
rect 115782 476618 151226 476854
rect 151462 476618 151546 476854
rect 151782 476618 187226 476854
rect 187462 476618 187546 476854
rect 187782 476618 223226 476854
rect 223462 476618 223546 476854
rect 223782 476618 259226 476854
rect 259462 476618 259546 476854
rect 259782 476618 295226 476854
rect 295462 476618 295546 476854
rect 295782 476618 331226 476854
rect 331462 476618 331546 476854
rect 331782 476618 367226 476854
rect 367462 476618 367546 476854
rect 367782 476618 403226 476854
rect 403462 476618 403546 476854
rect 403782 476618 439226 476854
rect 439462 476618 439546 476854
rect 439782 476618 475226 476854
rect 475462 476618 475546 476854
rect 475782 476618 511226 476854
rect 511462 476618 511546 476854
rect 511782 476618 547226 476854
rect 547462 476618 547546 476854
rect 547782 476618 590142 476854
rect 590378 476618 590462 476854
rect 590698 476618 592650 476854
rect -8726 476534 592650 476618
rect -8726 476298 -6774 476534
rect -6538 476298 -6454 476534
rect -6218 476298 7226 476534
rect 7462 476298 7546 476534
rect 7782 476298 43226 476534
rect 43462 476298 43546 476534
rect 43782 476298 79226 476534
rect 79462 476298 79546 476534
rect 79782 476298 115226 476534
rect 115462 476298 115546 476534
rect 115782 476298 151226 476534
rect 151462 476298 151546 476534
rect 151782 476298 187226 476534
rect 187462 476298 187546 476534
rect 187782 476298 223226 476534
rect 223462 476298 223546 476534
rect 223782 476298 259226 476534
rect 259462 476298 259546 476534
rect 259782 476298 295226 476534
rect 295462 476298 295546 476534
rect 295782 476298 331226 476534
rect 331462 476298 331546 476534
rect 331782 476298 367226 476534
rect 367462 476298 367546 476534
rect 367782 476298 403226 476534
rect 403462 476298 403546 476534
rect 403782 476298 439226 476534
rect 439462 476298 439546 476534
rect 439782 476298 475226 476534
rect 475462 476298 475546 476534
rect 475782 476298 511226 476534
rect 511462 476298 511546 476534
rect 511782 476298 547226 476534
rect 547462 476298 547546 476534
rect 547782 476298 590142 476534
rect 590378 476298 590462 476534
rect 590698 476298 592650 476534
rect -8726 476266 592650 476298
rect -8726 475614 592650 475646
rect -8726 475378 -5814 475614
rect -5578 475378 -5494 475614
rect -5258 475378 5986 475614
rect 6222 475378 6306 475614
rect 6542 475378 41986 475614
rect 42222 475378 42306 475614
rect 42542 475378 77986 475614
rect 78222 475378 78306 475614
rect 78542 475378 113986 475614
rect 114222 475378 114306 475614
rect 114542 475378 149986 475614
rect 150222 475378 150306 475614
rect 150542 475378 185986 475614
rect 186222 475378 186306 475614
rect 186542 475378 221986 475614
rect 222222 475378 222306 475614
rect 222542 475378 257986 475614
rect 258222 475378 258306 475614
rect 258542 475378 293986 475614
rect 294222 475378 294306 475614
rect 294542 475378 329986 475614
rect 330222 475378 330306 475614
rect 330542 475378 365986 475614
rect 366222 475378 366306 475614
rect 366542 475378 401986 475614
rect 402222 475378 402306 475614
rect 402542 475378 437986 475614
rect 438222 475378 438306 475614
rect 438542 475378 473986 475614
rect 474222 475378 474306 475614
rect 474542 475378 509986 475614
rect 510222 475378 510306 475614
rect 510542 475378 545986 475614
rect 546222 475378 546306 475614
rect 546542 475378 581986 475614
rect 582222 475378 582306 475614
rect 582542 475378 589182 475614
rect 589418 475378 589502 475614
rect 589738 475378 592650 475614
rect -8726 475294 592650 475378
rect -8726 475058 -5814 475294
rect -5578 475058 -5494 475294
rect -5258 475058 5986 475294
rect 6222 475058 6306 475294
rect 6542 475058 41986 475294
rect 42222 475058 42306 475294
rect 42542 475058 77986 475294
rect 78222 475058 78306 475294
rect 78542 475058 113986 475294
rect 114222 475058 114306 475294
rect 114542 475058 149986 475294
rect 150222 475058 150306 475294
rect 150542 475058 185986 475294
rect 186222 475058 186306 475294
rect 186542 475058 221986 475294
rect 222222 475058 222306 475294
rect 222542 475058 257986 475294
rect 258222 475058 258306 475294
rect 258542 475058 293986 475294
rect 294222 475058 294306 475294
rect 294542 475058 329986 475294
rect 330222 475058 330306 475294
rect 330542 475058 365986 475294
rect 366222 475058 366306 475294
rect 366542 475058 401986 475294
rect 402222 475058 402306 475294
rect 402542 475058 437986 475294
rect 438222 475058 438306 475294
rect 438542 475058 473986 475294
rect 474222 475058 474306 475294
rect 474542 475058 509986 475294
rect 510222 475058 510306 475294
rect 510542 475058 545986 475294
rect 546222 475058 546306 475294
rect 546542 475058 581986 475294
rect 582222 475058 582306 475294
rect 582542 475058 589182 475294
rect 589418 475058 589502 475294
rect 589738 475058 592650 475294
rect -8726 475026 592650 475058
rect -8726 474374 592650 474406
rect -8726 474138 -4854 474374
rect -4618 474138 -4534 474374
rect -4298 474138 4746 474374
rect 4982 474138 5066 474374
rect 5302 474138 40746 474374
rect 40982 474138 41066 474374
rect 41302 474138 76746 474374
rect 76982 474138 77066 474374
rect 77302 474138 112746 474374
rect 112982 474138 113066 474374
rect 113302 474138 148746 474374
rect 148982 474138 149066 474374
rect 149302 474138 184746 474374
rect 184982 474138 185066 474374
rect 185302 474138 220746 474374
rect 220982 474138 221066 474374
rect 221302 474138 256746 474374
rect 256982 474138 257066 474374
rect 257302 474138 292746 474374
rect 292982 474138 293066 474374
rect 293302 474138 328746 474374
rect 328982 474138 329066 474374
rect 329302 474138 364746 474374
rect 364982 474138 365066 474374
rect 365302 474138 400746 474374
rect 400982 474138 401066 474374
rect 401302 474138 436746 474374
rect 436982 474138 437066 474374
rect 437302 474138 472746 474374
rect 472982 474138 473066 474374
rect 473302 474138 508746 474374
rect 508982 474138 509066 474374
rect 509302 474138 544746 474374
rect 544982 474138 545066 474374
rect 545302 474138 580746 474374
rect 580982 474138 581066 474374
rect 581302 474138 588222 474374
rect 588458 474138 588542 474374
rect 588778 474138 592650 474374
rect -8726 474054 592650 474138
rect -8726 473818 -4854 474054
rect -4618 473818 -4534 474054
rect -4298 473818 4746 474054
rect 4982 473818 5066 474054
rect 5302 473818 40746 474054
rect 40982 473818 41066 474054
rect 41302 473818 76746 474054
rect 76982 473818 77066 474054
rect 77302 473818 112746 474054
rect 112982 473818 113066 474054
rect 113302 473818 148746 474054
rect 148982 473818 149066 474054
rect 149302 473818 184746 474054
rect 184982 473818 185066 474054
rect 185302 473818 220746 474054
rect 220982 473818 221066 474054
rect 221302 473818 256746 474054
rect 256982 473818 257066 474054
rect 257302 473818 292746 474054
rect 292982 473818 293066 474054
rect 293302 473818 328746 474054
rect 328982 473818 329066 474054
rect 329302 473818 364746 474054
rect 364982 473818 365066 474054
rect 365302 473818 400746 474054
rect 400982 473818 401066 474054
rect 401302 473818 436746 474054
rect 436982 473818 437066 474054
rect 437302 473818 472746 474054
rect 472982 473818 473066 474054
rect 473302 473818 508746 474054
rect 508982 473818 509066 474054
rect 509302 473818 544746 474054
rect 544982 473818 545066 474054
rect 545302 473818 580746 474054
rect 580982 473818 581066 474054
rect 581302 473818 588222 474054
rect 588458 473818 588542 474054
rect 588778 473818 592650 474054
rect -8726 473786 592650 473818
rect -8726 473134 592650 473166
rect -8726 472898 -3894 473134
rect -3658 472898 -3574 473134
rect -3338 472898 3506 473134
rect 3742 472898 3826 473134
rect 4062 472898 39506 473134
rect 39742 472898 39826 473134
rect 40062 472898 75506 473134
rect 75742 472898 75826 473134
rect 76062 472898 111506 473134
rect 111742 472898 111826 473134
rect 112062 472898 147506 473134
rect 147742 472898 147826 473134
rect 148062 472898 183506 473134
rect 183742 472898 183826 473134
rect 184062 472898 219506 473134
rect 219742 472898 219826 473134
rect 220062 472898 255506 473134
rect 255742 472898 255826 473134
rect 256062 472898 291506 473134
rect 291742 472898 291826 473134
rect 292062 472898 327506 473134
rect 327742 472898 327826 473134
rect 328062 472898 363506 473134
rect 363742 472898 363826 473134
rect 364062 472898 399506 473134
rect 399742 472898 399826 473134
rect 400062 472898 435506 473134
rect 435742 472898 435826 473134
rect 436062 472898 471506 473134
rect 471742 472898 471826 473134
rect 472062 472898 507506 473134
rect 507742 472898 507826 473134
rect 508062 472898 543506 473134
rect 543742 472898 543826 473134
rect 544062 472898 579506 473134
rect 579742 472898 579826 473134
rect 580062 472898 587262 473134
rect 587498 472898 587582 473134
rect 587818 472898 592650 473134
rect -8726 472814 592650 472898
rect -8726 472578 -3894 472814
rect -3658 472578 -3574 472814
rect -3338 472578 3506 472814
rect 3742 472578 3826 472814
rect 4062 472578 39506 472814
rect 39742 472578 39826 472814
rect 40062 472578 75506 472814
rect 75742 472578 75826 472814
rect 76062 472578 111506 472814
rect 111742 472578 111826 472814
rect 112062 472578 147506 472814
rect 147742 472578 147826 472814
rect 148062 472578 183506 472814
rect 183742 472578 183826 472814
rect 184062 472578 219506 472814
rect 219742 472578 219826 472814
rect 220062 472578 255506 472814
rect 255742 472578 255826 472814
rect 256062 472578 291506 472814
rect 291742 472578 291826 472814
rect 292062 472578 327506 472814
rect 327742 472578 327826 472814
rect 328062 472578 363506 472814
rect 363742 472578 363826 472814
rect 364062 472578 399506 472814
rect 399742 472578 399826 472814
rect 400062 472578 435506 472814
rect 435742 472578 435826 472814
rect 436062 472578 471506 472814
rect 471742 472578 471826 472814
rect 472062 472578 507506 472814
rect 507742 472578 507826 472814
rect 508062 472578 543506 472814
rect 543742 472578 543826 472814
rect 544062 472578 579506 472814
rect 579742 472578 579826 472814
rect 580062 472578 587262 472814
rect 587498 472578 587582 472814
rect 587818 472578 592650 472814
rect -8726 472546 592650 472578
rect -8726 471894 592650 471926
rect -8726 471658 -2934 471894
rect -2698 471658 -2614 471894
rect -2378 471658 2266 471894
rect 2502 471658 2586 471894
rect 2822 471658 38266 471894
rect 38502 471658 38586 471894
rect 38822 471658 74266 471894
rect 74502 471658 74586 471894
rect 74822 471658 110266 471894
rect 110502 471658 110586 471894
rect 110822 471658 146266 471894
rect 146502 471658 146586 471894
rect 146822 471658 182266 471894
rect 182502 471658 182586 471894
rect 182822 471658 218266 471894
rect 218502 471658 218586 471894
rect 218822 471658 254266 471894
rect 254502 471658 254586 471894
rect 254822 471658 290266 471894
rect 290502 471658 290586 471894
rect 290822 471658 326266 471894
rect 326502 471658 326586 471894
rect 326822 471658 362266 471894
rect 362502 471658 362586 471894
rect 362822 471658 398266 471894
rect 398502 471658 398586 471894
rect 398822 471658 434266 471894
rect 434502 471658 434586 471894
rect 434822 471658 470266 471894
rect 470502 471658 470586 471894
rect 470822 471658 506266 471894
rect 506502 471658 506586 471894
rect 506822 471658 542266 471894
rect 542502 471658 542586 471894
rect 542822 471658 578266 471894
rect 578502 471658 578586 471894
rect 578822 471658 586302 471894
rect 586538 471658 586622 471894
rect 586858 471658 592650 471894
rect -8726 471574 592650 471658
rect -8726 471338 -2934 471574
rect -2698 471338 -2614 471574
rect -2378 471338 2266 471574
rect 2502 471338 2586 471574
rect 2822 471338 38266 471574
rect 38502 471338 38586 471574
rect 38822 471338 74266 471574
rect 74502 471338 74586 471574
rect 74822 471338 110266 471574
rect 110502 471338 110586 471574
rect 110822 471338 146266 471574
rect 146502 471338 146586 471574
rect 146822 471338 182266 471574
rect 182502 471338 182586 471574
rect 182822 471338 218266 471574
rect 218502 471338 218586 471574
rect 218822 471338 254266 471574
rect 254502 471338 254586 471574
rect 254822 471338 290266 471574
rect 290502 471338 290586 471574
rect 290822 471338 326266 471574
rect 326502 471338 326586 471574
rect 326822 471338 362266 471574
rect 362502 471338 362586 471574
rect 362822 471338 398266 471574
rect 398502 471338 398586 471574
rect 398822 471338 434266 471574
rect 434502 471338 434586 471574
rect 434822 471338 470266 471574
rect 470502 471338 470586 471574
rect 470822 471338 506266 471574
rect 506502 471338 506586 471574
rect 506822 471338 542266 471574
rect 542502 471338 542586 471574
rect 542822 471338 578266 471574
rect 578502 471338 578586 471574
rect 578822 471338 586302 471574
rect 586538 471338 586622 471574
rect 586858 471338 592650 471574
rect -8726 471306 592650 471338
rect -8726 470654 592650 470686
rect -8726 470418 -1974 470654
rect -1738 470418 -1654 470654
rect -1418 470418 1026 470654
rect 1262 470418 1346 470654
rect 1582 470418 37026 470654
rect 37262 470418 37346 470654
rect 37582 470418 73026 470654
rect 73262 470418 73346 470654
rect 73582 470418 109026 470654
rect 109262 470418 109346 470654
rect 109582 470418 145026 470654
rect 145262 470418 145346 470654
rect 145582 470418 181026 470654
rect 181262 470418 181346 470654
rect 181582 470418 217026 470654
rect 217262 470418 217346 470654
rect 217582 470418 253026 470654
rect 253262 470418 253346 470654
rect 253582 470418 289026 470654
rect 289262 470418 289346 470654
rect 289582 470418 325026 470654
rect 325262 470418 325346 470654
rect 325582 470418 361026 470654
rect 361262 470418 361346 470654
rect 361582 470418 397026 470654
rect 397262 470418 397346 470654
rect 397582 470418 433026 470654
rect 433262 470418 433346 470654
rect 433582 470418 469026 470654
rect 469262 470418 469346 470654
rect 469582 470418 505026 470654
rect 505262 470418 505346 470654
rect 505582 470418 541026 470654
rect 541262 470418 541346 470654
rect 541582 470418 577026 470654
rect 577262 470418 577346 470654
rect 577582 470418 585342 470654
rect 585578 470418 585662 470654
rect 585898 470418 592650 470654
rect -8726 470334 592650 470418
rect -8726 470098 -1974 470334
rect -1738 470098 -1654 470334
rect -1418 470098 1026 470334
rect 1262 470098 1346 470334
rect 1582 470098 37026 470334
rect 37262 470098 37346 470334
rect 37582 470098 73026 470334
rect 73262 470098 73346 470334
rect 73582 470098 109026 470334
rect 109262 470098 109346 470334
rect 109582 470098 145026 470334
rect 145262 470098 145346 470334
rect 145582 470098 181026 470334
rect 181262 470098 181346 470334
rect 181582 470098 217026 470334
rect 217262 470098 217346 470334
rect 217582 470098 253026 470334
rect 253262 470098 253346 470334
rect 253582 470098 289026 470334
rect 289262 470098 289346 470334
rect 289582 470098 325026 470334
rect 325262 470098 325346 470334
rect 325582 470098 361026 470334
rect 361262 470098 361346 470334
rect 361582 470098 397026 470334
rect 397262 470098 397346 470334
rect 397582 470098 433026 470334
rect 433262 470098 433346 470334
rect 433582 470098 469026 470334
rect 469262 470098 469346 470334
rect 469582 470098 505026 470334
rect 505262 470098 505346 470334
rect 505582 470098 541026 470334
rect 541262 470098 541346 470334
rect 541582 470098 577026 470334
rect 577262 470098 577346 470334
rect 577582 470098 585342 470334
rect 585578 470098 585662 470334
rect 585898 470098 592650 470334
rect -8726 470066 592650 470098
rect -8726 443334 592650 443366
rect -8726 443098 -8694 443334
rect -8458 443098 -8374 443334
rect -8138 443098 9706 443334
rect 9942 443098 10026 443334
rect 10262 443098 45706 443334
rect 45942 443098 46026 443334
rect 46262 443098 81706 443334
rect 81942 443098 82026 443334
rect 82262 443098 117706 443334
rect 117942 443098 118026 443334
rect 118262 443098 153706 443334
rect 153942 443098 154026 443334
rect 154262 443098 189706 443334
rect 189942 443098 190026 443334
rect 190262 443098 225706 443334
rect 225942 443098 226026 443334
rect 226262 443098 261706 443334
rect 261942 443098 262026 443334
rect 262262 443098 297706 443334
rect 297942 443098 298026 443334
rect 298262 443098 333706 443334
rect 333942 443098 334026 443334
rect 334262 443098 369706 443334
rect 369942 443098 370026 443334
rect 370262 443098 405706 443334
rect 405942 443098 406026 443334
rect 406262 443098 441706 443334
rect 441942 443098 442026 443334
rect 442262 443098 477706 443334
rect 477942 443098 478026 443334
rect 478262 443098 513706 443334
rect 513942 443098 514026 443334
rect 514262 443098 549706 443334
rect 549942 443098 550026 443334
rect 550262 443098 592062 443334
rect 592298 443098 592382 443334
rect 592618 443098 592650 443334
rect -8726 443014 592650 443098
rect -8726 442778 -8694 443014
rect -8458 442778 -8374 443014
rect -8138 442778 9706 443014
rect 9942 442778 10026 443014
rect 10262 442778 45706 443014
rect 45942 442778 46026 443014
rect 46262 442778 81706 443014
rect 81942 442778 82026 443014
rect 82262 442778 117706 443014
rect 117942 442778 118026 443014
rect 118262 442778 153706 443014
rect 153942 442778 154026 443014
rect 154262 442778 189706 443014
rect 189942 442778 190026 443014
rect 190262 442778 225706 443014
rect 225942 442778 226026 443014
rect 226262 442778 261706 443014
rect 261942 442778 262026 443014
rect 262262 442778 297706 443014
rect 297942 442778 298026 443014
rect 298262 442778 333706 443014
rect 333942 442778 334026 443014
rect 334262 442778 369706 443014
rect 369942 442778 370026 443014
rect 370262 442778 405706 443014
rect 405942 442778 406026 443014
rect 406262 442778 441706 443014
rect 441942 442778 442026 443014
rect 442262 442778 477706 443014
rect 477942 442778 478026 443014
rect 478262 442778 513706 443014
rect 513942 442778 514026 443014
rect 514262 442778 549706 443014
rect 549942 442778 550026 443014
rect 550262 442778 592062 443014
rect 592298 442778 592382 443014
rect 592618 442778 592650 443014
rect -8726 442746 592650 442778
rect -8726 442094 592650 442126
rect -8726 441858 -7734 442094
rect -7498 441858 -7414 442094
rect -7178 441858 8466 442094
rect 8702 441858 8786 442094
rect 9022 441858 44466 442094
rect 44702 441858 44786 442094
rect 45022 441858 80466 442094
rect 80702 441858 80786 442094
rect 81022 441858 116466 442094
rect 116702 441858 116786 442094
rect 117022 441858 152466 442094
rect 152702 441858 152786 442094
rect 153022 441858 188466 442094
rect 188702 441858 188786 442094
rect 189022 441858 224466 442094
rect 224702 441858 224786 442094
rect 225022 441858 260466 442094
rect 260702 441858 260786 442094
rect 261022 441858 296466 442094
rect 296702 441858 296786 442094
rect 297022 441858 332466 442094
rect 332702 441858 332786 442094
rect 333022 441858 368466 442094
rect 368702 441858 368786 442094
rect 369022 441858 404466 442094
rect 404702 441858 404786 442094
rect 405022 441858 440466 442094
rect 440702 441858 440786 442094
rect 441022 441858 476466 442094
rect 476702 441858 476786 442094
rect 477022 441858 512466 442094
rect 512702 441858 512786 442094
rect 513022 441858 548466 442094
rect 548702 441858 548786 442094
rect 549022 441858 591102 442094
rect 591338 441858 591422 442094
rect 591658 441858 592650 442094
rect -8726 441774 592650 441858
rect -8726 441538 -7734 441774
rect -7498 441538 -7414 441774
rect -7178 441538 8466 441774
rect 8702 441538 8786 441774
rect 9022 441538 44466 441774
rect 44702 441538 44786 441774
rect 45022 441538 80466 441774
rect 80702 441538 80786 441774
rect 81022 441538 116466 441774
rect 116702 441538 116786 441774
rect 117022 441538 152466 441774
rect 152702 441538 152786 441774
rect 153022 441538 188466 441774
rect 188702 441538 188786 441774
rect 189022 441538 224466 441774
rect 224702 441538 224786 441774
rect 225022 441538 260466 441774
rect 260702 441538 260786 441774
rect 261022 441538 296466 441774
rect 296702 441538 296786 441774
rect 297022 441538 332466 441774
rect 332702 441538 332786 441774
rect 333022 441538 368466 441774
rect 368702 441538 368786 441774
rect 369022 441538 404466 441774
rect 404702 441538 404786 441774
rect 405022 441538 440466 441774
rect 440702 441538 440786 441774
rect 441022 441538 476466 441774
rect 476702 441538 476786 441774
rect 477022 441538 512466 441774
rect 512702 441538 512786 441774
rect 513022 441538 548466 441774
rect 548702 441538 548786 441774
rect 549022 441538 591102 441774
rect 591338 441538 591422 441774
rect 591658 441538 592650 441774
rect -8726 441506 592650 441538
rect -8726 440854 592650 440886
rect -8726 440618 -6774 440854
rect -6538 440618 -6454 440854
rect -6218 440618 7226 440854
rect 7462 440618 7546 440854
rect 7782 440618 43226 440854
rect 43462 440618 43546 440854
rect 43782 440618 79226 440854
rect 79462 440618 79546 440854
rect 79782 440618 115226 440854
rect 115462 440618 115546 440854
rect 115782 440618 151226 440854
rect 151462 440618 151546 440854
rect 151782 440618 187226 440854
rect 187462 440618 187546 440854
rect 187782 440618 223226 440854
rect 223462 440618 223546 440854
rect 223782 440618 259226 440854
rect 259462 440618 259546 440854
rect 259782 440618 295226 440854
rect 295462 440618 295546 440854
rect 295782 440618 331226 440854
rect 331462 440618 331546 440854
rect 331782 440618 367226 440854
rect 367462 440618 367546 440854
rect 367782 440618 403226 440854
rect 403462 440618 403546 440854
rect 403782 440618 439226 440854
rect 439462 440618 439546 440854
rect 439782 440618 475226 440854
rect 475462 440618 475546 440854
rect 475782 440618 511226 440854
rect 511462 440618 511546 440854
rect 511782 440618 547226 440854
rect 547462 440618 547546 440854
rect 547782 440618 590142 440854
rect 590378 440618 590462 440854
rect 590698 440618 592650 440854
rect -8726 440534 592650 440618
rect -8726 440298 -6774 440534
rect -6538 440298 -6454 440534
rect -6218 440298 7226 440534
rect 7462 440298 7546 440534
rect 7782 440298 43226 440534
rect 43462 440298 43546 440534
rect 43782 440298 79226 440534
rect 79462 440298 79546 440534
rect 79782 440298 115226 440534
rect 115462 440298 115546 440534
rect 115782 440298 151226 440534
rect 151462 440298 151546 440534
rect 151782 440298 187226 440534
rect 187462 440298 187546 440534
rect 187782 440298 223226 440534
rect 223462 440298 223546 440534
rect 223782 440298 259226 440534
rect 259462 440298 259546 440534
rect 259782 440298 295226 440534
rect 295462 440298 295546 440534
rect 295782 440298 331226 440534
rect 331462 440298 331546 440534
rect 331782 440298 367226 440534
rect 367462 440298 367546 440534
rect 367782 440298 403226 440534
rect 403462 440298 403546 440534
rect 403782 440298 439226 440534
rect 439462 440298 439546 440534
rect 439782 440298 475226 440534
rect 475462 440298 475546 440534
rect 475782 440298 511226 440534
rect 511462 440298 511546 440534
rect 511782 440298 547226 440534
rect 547462 440298 547546 440534
rect 547782 440298 590142 440534
rect 590378 440298 590462 440534
rect 590698 440298 592650 440534
rect -8726 440266 592650 440298
rect -8726 439614 592650 439646
rect -8726 439378 -5814 439614
rect -5578 439378 -5494 439614
rect -5258 439378 5986 439614
rect 6222 439378 6306 439614
rect 6542 439378 41986 439614
rect 42222 439378 42306 439614
rect 42542 439378 77986 439614
rect 78222 439378 78306 439614
rect 78542 439378 113986 439614
rect 114222 439378 114306 439614
rect 114542 439378 149986 439614
rect 150222 439378 150306 439614
rect 150542 439378 185986 439614
rect 186222 439378 186306 439614
rect 186542 439378 221986 439614
rect 222222 439378 222306 439614
rect 222542 439378 257986 439614
rect 258222 439378 258306 439614
rect 258542 439378 293986 439614
rect 294222 439378 294306 439614
rect 294542 439378 329986 439614
rect 330222 439378 330306 439614
rect 330542 439378 365986 439614
rect 366222 439378 366306 439614
rect 366542 439378 401986 439614
rect 402222 439378 402306 439614
rect 402542 439378 437986 439614
rect 438222 439378 438306 439614
rect 438542 439378 473986 439614
rect 474222 439378 474306 439614
rect 474542 439378 509986 439614
rect 510222 439378 510306 439614
rect 510542 439378 581986 439614
rect 582222 439378 582306 439614
rect 582542 439378 589182 439614
rect 589418 439378 589502 439614
rect 589738 439378 592650 439614
rect -8726 439294 592650 439378
rect -8726 439058 -5814 439294
rect -5578 439058 -5494 439294
rect -5258 439058 5986 439294
rect 6222 439058 6306 439294
rect 6542 439058 41986 439294
rect 42222 439058 42306 439294
rect 42542 439058 77986 439294
rect 78222 439058 78306 439294
rect 78542 439058 113986 439294
rect 114222 439058 114306 439294
rect 114542 439058 149986 439294
rect 150222 439058 150306 439294
rect 150542 439058 185986 439294
rect 186222 439058 186306 439294
rect 186542 439058 221986 439294
rect 222222 439058 222306 439294
rect 222542 439058 257986 439294
rect 258222 439058 258306 439294
rect 258542 439058 293986 439294
rect 294222 439058 294306 439294
rect 294542 439058 329986 439294
rect 330222 439058 330306 439294
rect 330542 439058 365986 439294
rect 366222 439058 366306 439294
rect 366542 439058 401986 439294
rect 402222 439058 402306 439294
rect 402542 439058 437986 439294
rect 438222 439058 438306 439294
rect 438542 439058 473986 439294
rect 474222 439058 474306 439294
rect 474542 439058 509986 439294
rect 510222 439058 510306 439294
rect 510542 439058 581986 439294
rect 582222 439058 582306 439294
rect 582542 439058 589182 439294
rect 589418 439058 589502 439294
rect 589738 439058 592650 439294
rect -8726 439026 592650 439058
rect -8726 438374 592650 438406
rect -8726 438138 -4854 438374
rect -4618 438138 -4534 438374
rect -4298 438138 4746 438374
rect 4982 438138 5066 438374
rect 5302 438138 40746 438374
rect 40982 438138 41066 438374
rect 41302 438138 76746 438374
rect 76982 438138 77066 438374
rect 77302 438138 112746 438374
rect 112982 438138 113066 438374
rect 113302 438138 148746 438374
rect 148982 438138 149066 438374
rect 149302 438138 184746 438374
rect 184982 438138 185066 438374
rect 185302 438138 220746 438374
rect 220982 438138 221066 438374
rect 221302 438138 256746 438374
rect 256982 438138 257066 438374
rect 257302 438138 292746 438374
rect 292982 438138 293066 438374
rect 293302 438138 328746 438374
rect 328982 438138 329066 438374
rect 329302 438138 364746 438374
rect 364982 438138 365066 438374
rect 365302 438138 400746 438374
rect 400982 438138 401066 438374
rect 401302 438138 436746 438374
rect 436982 438138 437066 438374
rect 437302 438138 472746 438374
rect 472982 438138 473066 438374
rect 473302 438138 508746 438374
rect 508982 438138 509066 438374
rect 509302 438138 580746 438374
rect 580982 438138 581066 438374
rect 581302 438138 588222 438374
rect 588458 438138 588542 438374
rect 588778 438138 592650 438374
rect -8726 438054 592650 438138
rect -8726 437818 -4854 438054
rect -4618 437818 -4534 438054
rect -4298 437818 4746 438054
rect 4982 437818 5066 438054
rect 5302 437818 40746 438054
rect 40982 437818 41066 438054
rect 41302 437818 76746 438054
rect 76982 437818 77066 438054
rect 77302 437818 112746 438054
rect 112982 437818 113066 438054
rect 113302 437818 148746 438054
rect 148982 437818 149066 438054
rect 149302 437818 184746 438054
rect 184982 437818 185066 438054
rect 185302 437818 220746 438054
rect 220982 437818 221066 438054
rect 221302 437818 256746 438054
rect 256982 437818 257066 438054
rect 257302 437818 292746 438054
rect 292982 437818 293066 438054
rect 293302 437818 328746 438054
rect 328982 437818 329066 438054
rect 329302 437818 364746 438054
rect 364982 437818 365066 438054
rect 365302 437818 400746 438054
rect 400982 437818 401066 438054
rect 401302 437818 436746 438054
rect 436982 437818 437066 438054
rect 437302 437818 472746 438054
rect 472982 437818 473066 438054
rect 473302 437818 508746 438054
rect 508982 437818 509066 438054
rect 509302 437818 580746 438054
rect 580982 437818 581066 438054
rect 581302 437818 588222 438054
rect 588458 437818 588542 438054
rect 588778 437818 592650 438054
rect -8726 437786 592650 437818
rect -8726 437134 592650 437166
rect -8726 436898 -3894 437134
rect -3658 436898 -3574 437134
rect -3338 436898 3506 437134
rect 3742 436898 3826 437134
rect 4062 436898 39506 437134
rect 39742 436898 39826 437134
rect 40062 436898 75506 437134
rect 75742 436898 75826 437134
rect 76062 436898 111506 437134
rect 111742 436898 111826 437134
rect 112062 436898 147506 437134
rect 147742 436898 147826 437134
rect 148062 436898 183506 437134
rect 183742 436898 183826 437134
rect 184062 436898 219506 437134
rect 219742 436898 219826 437134
rect 220062 436898 255506 437134
rect 255742 436898 255826 437134
rect 256062 436898 291506 437134
rect 291742 436898 291826 437134
rect 292062 436898 327506 437134
rect 327742 436898 327826 437134
rect 328062 436898 363506 437134
rect 363742 436898 363826 437134
rect 364062 436898 399506 437134
rect 399742 436898 399826 437134
rect 400062 436898 435506 437134
rect 435742 436898 435826 437134
rect 436062 436898 471506 437134
rect 471742 436898 471826 437134
rect 472062 436898 507506 437134
rect 507742 436898 507826 437134
rect 508062 436898 579506 437134
rect 579742 436898 579826 437134
rect 580062 436898 587262 437134
rect 587498 436898 587582 437134
rect 587818 436898 592650 437134
rect -8726 436814 592650 436898
rect -8726 436578 -3894 436814
rect -3658 436578 -3574 436814
rect -3338 436578 3506 436814
rect 3742 436578 3826 436814
rect 4062 436578 39506 436814
rect 39742 436578 39826 436814
rect 40062 436578 75506 436814
rect 75742 436578 75826 436814
rect 76062 436578 111506 436814
rect 111742 436578 111826 436814
rect 112062 436578 147506 436814
rect 147742 436578 147826 436814
rect 148062 436578 183506 436814
rect 183742 436578 183826 436814
rect 184062 436578 219506 436814
rect 219742 436578 219826 436814
rect 220062 436578 255506 436814
rect 255742 436578 255826 436814
rect 256062 436578 291506 436814
rect 291742 436578 291826 436814
rect 292062 436578 327506 436814
rect 327742 436578 327826 436814
rect 328062 436578 363506 436814
rect 363742 436578 363826 436814
rect 364062 436578 399506 436814
rect 399742 436578 399826 436814
rect 400062 436578 435506 436814
rect 435742 436578 435826 436814
rect 436062 436578 471506 436814
rect 471742 436578 471826 436814
rect 472062 436578 507506 436814
rect 507742 436578 507826 436814
rect 508062 436578 579506 436814
rect 579742 436578 579826 436814
rect 580062 436578 587262 436814
rect 587498 436578 587582 436814
rect 587818 436578 592650 436814
rect -8726 436546 592650 436578
rect -8726 435894 592650 435926
rect -8726 435658 -2934 435894
rect -2698 435658 -2614 435894
rect -2378 435658 2266 435894
rect 2502 435658 2586 435894
rect 2822 435658 38266 435894
rect 38502 435658 38586 435894
rect 38822 435658 74266 435894
rect 74502 435658 74586 435894
rect 74822 435658 110266 435894
rect 110502 435658 110586 435894
rect 110822 435658 146266 435894
rect 146502 435658 146586 435894
rect 146822 435658 182266 435894
rect 182502 435658 182586 435894
rect 182822 435658 218266 435894
rect 218502 435658 218586 435894
rect 218822 435658 254266 435894
rect 254502 435658 254586 435894
rect 254822 435658 290266 435894
rect 290502 435658 290586 435894
rect 290822 435658 326266 435894
rect 326502 435658 326586 435894
rect 326822 435658 362266 435894
rect 362502 435658 362586 435894
rect 362822 435658 398266 435894
rect 398502 435658 398586 435894
rect 398822 435658 434266 435894
rect 434502 435658 434586 435894
rect 434822 435658 470266 435894
rect 470502 435658 470586 435894
rect 470822 435658 506266 435894
rect 506502 435658 506586 435894
rect 506822 435658 540918 435894
rect 541154 435658 542850 435894
rect 543086 435658 544782 435894
rect 545018 435658 546714 435894
rect 546950 435658 578266 435894
rect 578502 435658 578586 435894
rect 578822 435658 586302 435894
rect 586538 435658 586622 435894
rect 586858 435658 592650 435894
rect -8726 435574 592650 435658
rect -8726 435338 -2934 435574
rect -2698 435338 -2614 435574
rect -2378 435338 2266 435574
rect 2502 435338 2586 435574
rect 2822 435338 38266 435574
rect 38502 435338 38586 435574
rect 38822 435338 74266 435574
rect 74502 435338 74586 435574
rect 74822 435338 110266 435574
rect 110502 435338 110586 435574
rect 110822 435338 146266 435574
rect 146502 435338 146586 435574
rect 146822 435338 182266 435574
rect 182502 435338 182586 435574
rect 182822 435338 218266 435574
rect 218502 435338 218586 435574
rect 218822 435338 254266 435574
rect 254502 435338 254586 435574
rect 254822 435338 290266 435574
rect 290502 435338 290586 435574
rect 290822 435338 326266 435574
rect 326502 435338 326586 435574
rect 326822 435338 362266 435574
rect 362502 435338 362586 435574
rect 362822 435338 398266 435574
rect 398502 435338 398586 435574
rect 398822 435338 434266 435574
rect 434502 435338 434586 435574
rect 434822 435338 470266 435574
rect 470502 435338 470586 435574
rect 470822 435338 506266 435574
rect 506502 435338 506586 435574
rect 506822 435338 540918 435574
rect 541154 435338 542850 435574
rect 543086 435338 544782 435574
rect 545018 435338 546714 435574
rect 546950 435338 578266 435574
rect 578502 435338 578586 435574
rect 578822 435338 586302 435574
rect 586538 435338 586622 435574
rect 586858 435338 592650 435574
rect -8726 435306 592650 435338
rect -8726 434654 592650 434686
rect -8726 434418 -1974 434654
rect -1738 434418 -1654 434654
rect -1418 434418 1026 434654
rect 1262 434418 1346 434654
rect 1582 434418 37026 434654
rect 37262 434418 37346 434654
rect 37582 434418 73026 434654
rect 73262 434418 73346 434654
rect 73582 434418 109026 434654
rect 109262 434418 109346 434654
rect 109582 434418 145026 434654
rect 145262 434418 145346 434654
rect 145582 434418 181026 434654
rect 181262 434418 181346 434654
rect 181582 434418 217026 434654
rect 217262 434418 217346 434654
rect 217582 434418 253026 434654
rect 253262 434418 253346 434654
rect 253582 434418 289026 434654
rect 289262 434418 289346 434654
rect 289582 434418 325026 434654
rect 325262 434418 325346 434654
rect 325582 434418 361026 434654
rect 361262 434418 361346 434654
rect 361582 434418 397026 434654
rect 397262 434418 397346 434654
rect 397582 434418 433026 434654
rect 433262 434418 433346 434654
rect 433582 434418 469026 434654
rect 469262 434418 469346 434654
rect 469582 434418 505026 434654
rect 505262 434418 505346 434654
rect 505582 434418 539952 434654
rect 540188 434418 541884 434654
rect 542120 434418 543816 434654
rect 544052 434418 545748 434654
rect 545984 434418 577026 434654
rect 577262 434418 577346 434654
rect 577582 434418 585342 434654
rect 585578 434418 585662 434654
rect 585898 434418 592650 434654
rect -8726 434334 592650 434418
rect -8726 434098 -1974 434334
rect -1738 434098 -1654 434334
rect -1418 434098 1026 434334
rect 1262 434098 1346 434334
rect 1582 434098 37026 434334
rect 37262 434098 37346 434334
rect 37582 434098 73026 434334
rect 73262 434098 73346 434334
rect 73582 434098 109026 434334
rect 109262 434098 109346 434334
rect 109582 434098 145026 434334
rect 145262 434098 145346 434334
rect 145582 434098 181026 434334
rect 181262 434098 181346 434334
rect 181582 434098 217026 434334
rect 217262 434098 217346 434334
rect 217582 434098 253026 434334
rect 253262 434098 253346 434334
rect 253582 434098 289026 434334
rect 289262 434098 289346 434334
rect 289582 434098 325026 434334
rect 325262 434098 325346 434334
rect 325582 434098 361026 434334
rect 361262 434098 361346 434334
rect 361582 434098 397026 434334
rect 397262 434098 397346 434334
rect 397582 434098 433026 434334
rect 433262 434098 433346 434334
rect 433582 434098 469026 434334
rect 469262 434098 469346 434334
rect 469582 434098 505026 434334
rect 505262 434098 505346 434334
rect 505582 434098 539952 434334
rect 540188 434098 541884 434334
rect 542120 434098 543816 434334
rect 544052 434098 545748 434334
rect 545984 434098 577026 434334
rect 577262 434098 577346 434334
rect 577582 434098 585342 434334
rect 585578 434098 585662 434334
rect 585898 434098 592650 434334
rect -8726 434066 592650 434098
rect -8726 407334 592650 407366
rect -8726 407098 -8694 407334
rect -8458 407098 -8374 407334
rect -8138 407098 9706 407334
rect 9942 407098 10026 407334
rect 10262 407098 45706 407334
rect 45942 407098 46026 407334
rect 46262 407098 81706 407334
rect 81942 407098 82026 407334
rect 82262 407098 117706 407334
rect 117942 407098 118026 407334
rect 118262 407098 153706 407334
rect 153942 407098 154026 407334
rect 154262 407098 189706 407334
rect 189942 407098 190026 407334
rect 190262 407098 225706 407334
rect 225942 407098 226026 407334
rect 226262 407098 261706 407334
rect 261942 407098 262026 407334
rect 262262 407098 297706 407334
rect 297942 407098 298026 407334
rect 298262 407098 333706 407334
rect 333942 407098 334026 407334
rect 334262 407098 369706 407334
rect 369942 407098 370026 407334
rect 370262 407098 405706 407334
rect 405942 407098 406026 407334
rect 406262 407098 441706 407334
rect 441942 407098 442026 407334
rect 442262 407098 477706 407334
rect 477942 407098 478026 407334
rect 478262 407098 513706 407334
rect 513942 407098 514026 407334
rect 514262 407098 549706 407334
rect 549942 407098 550026 407334
rect 550262 407098 592062 407334
rect 592298 407098 592382 407334
rect 592618 407098 592650 407334
rect -8726 407014 592650 407098
rect -8726 406778 -8694 407014
rect -8458 406778 -8374 407014
rect -8138 406778 9706 407014
rect 9942 406778 10026 407014
rect 10262 406778 45706 407014
rect 45942 406778 46026 407014
rect 46262 406778 81706 407014
rect 81942 406778 82026 407014
rect 82262 406778 117706 407014
rect 117942 406778 118026 407014
rect 118262 406778 153706 407014
rect 153942 406778 154026 407014
rect 154262 406778 189706 407014
rect 189942 406778 190026 407014
rect 190262 406778 225706 407014
rect 225942 406778 226026 407014
rect 226262 406778 261706 407014
rect 261942 406778 262026 407014
rect 262262 406778 297706 407014
rect 297942 406778 298026 407014
rect 298262 406778 333706 407014
rect 333942 406778 334026 407014
rect 334262 406778 369706 407014
rect 369942 406778 370026 407014
rect 370262 406778 405706 407014
rect 405942 406778 406026 407014
rect 406262 406778 441706 407014
rect 441942 406778 442026 407014
rect 442262 406778 477706 407014
rect 477942 406778 478026 407014
rect 478262 406778 513706 407014
rect 513942 406778 514026 407014
rect 514262 406778 549706 407014
rect 549942 406778 550026 407014
rect 550262 406778 592062 407014
rect 592298 406778 592382 407014
rect 592618 406778 592650 407014
rect -8726 406746 592650 406778
rect -8726 406094 592650 406126
rect -8726 405858 -7734 406094
rect -7498 405858 -7414 406094
rect -7178 405858 8466 406094
rect 8702 405858 8786 406094
rect 9022 405858 44466 406094
rect 44702 405858 44786 406094
rect 45022 405858 80466 406094
rect 80702 405858 80786 406094
rect 81022 405858 116466 406094
rect 116702 405858 116786 406094
rect 117022 405858 152466 406094
rect 152702 405858 152786 406094
rect 153022 405858 188466 406094
rect 188702 405858 188786 406094
rect 189022 405858 224466 406094
rect 224702 405858 224786 406094
rect 225022 405858 260466 406094
rect 260702 405858 260786 406094
rect 261022 405858 296466 406094
rect 296702 405858 296786 406094
rect 297022 405858 332466 406094
rect 332702 405858 332786 406094
rect 333022 405858 368466 406094
rect 368702 405858 368786 406094
rect 369022 405858 404466 406094
rect 404702 405858 404786 406094
rect 405022 405858 440466 406094
rect 440702 405858 440786 406094
rect 441022 405858 476466 406094
rect 476702 405858 476786 406094
rect 477022 405858 512466 406094
rect 512702 405858 512786 406094
rect 513022 405858 548466 406094
rect 548702 405858 548786 406094
rect 549022 405858 591102 406094
rect 591338 405858 591422 406094
rect 591658 405858 592650 406094
rect -8726 405774 592650 405858
rect -8726 405538 -7734 405774
rect -7498 405538 -7414 405774
rect -7178 405538 8466 405774
rect 8702 405538 8786 405774
rect 9022 405538 44466 405774
rect 44702 405538 44786 405774
rect 45022 405538 80466 405774
rect 80702 405538 80786 405774
rect 81022 405538 116466 405774
rect 116702 405538 116786 405774
rect 117022 405538 152466 405774
rect 152702 405538 152786 405774
rect 153022 405538 188466 405774
rect 188702 405538 188786 405774
rect 189022 405538 224466 405774
rect 224702 405538 224786 405774
rect 225022 405538 260466 405774
rect 260702 405538 260786 405774
rect 261022 405538 296466 405774
rect 296702 405538 296786 405774
rect 297022 405538 332466 405774
rect 332702 405538 332786 405774
rect 333022 405538 368466 405774
rect 368702 405538 368786 405774
rect 369022 405538 404466 405774
rect 404702 405538 404786 405774
rect 405022 405538 440466 405774
rect 440702 405538 440786 405774
rect 441022 405538 476466 405774
rect 476702 405538 476786 405774
rect 477022 405538 512466 405774
rect 512702 405538 512786 405774
rect 513022 405538 548466 405774
rect 548702 405538 548786 405774
rect 549022 405538 591102 405774
rect 591338 405538 591422 405774
rect 591658 405538 592650 405774
rect -8726 405506 592650 405538
rect -8726 404854 592650 404886
rect -8726 404618 -6774 404854
rect -6538 404618 -6454 404854
rect -6218 404618 7226 404854
rect 7462 404618 7546 404854
rect 7782 404618 43226 404854
rect 43462 404618 43546 404854
rect 43782 404618 79226 404854
rect 79462 404618 79546 404854
rect 79782 404618 115226 404854
rect 115462 404618 115546 404854
rect 115782 404618 151226 404854
rect 151462 404618 151546 404854
rect 151782 404618 187226 404854
rect 187462 404618 187546 404854
rect 187782 404618 223226 404854
rect 223462 404618 223546 404854
rect 223782 404618 259226 404854
rect 259462 404618 259546 404854
rect 259782 404618 295226 404854
rect 295462 404618 295546 404854
rect 295782 404618 331226 404854
rect 331462 404618 331546 404854
rect 331782 404618 367226 404854
rect 367462 404618 367546 404854
rect 367782 404618 403226 404854
rect 403462 404618 403546 404854
rect 403782 404618 439226 404854
rect 439462 404618 439546 404854
rect 439782 404618 475226 404854
rect 475462 404618 475546 404854
rect 475782 404618 511226 404854
rect 511462 404618 511546 404854
rect 511782 404618 547226 404854
rect 547462 404618 547546 404854
rect 547782 404618 590142 404854
rect 590378 404618 590462 404854
rect 590698 404618 592650 404854
rect -8726 404534 592650 404618
rect -8726 404298 -6774 404534
rect -6538 404298 -6454 404534
rect -6218 404298 7226 404534
rect 7462 404298 7546 404534
rect 7782 404298 43226 404534
rect 43462 404298 43546 404534
rect 43782 404298 79226 404534
rect 79462 404298 79546 404534
rect 79782 404298 115226 404534
rect 115462 404298 115546 404534
rect 115782 404298 151226 404534
rect 151462 404298 151546 404534
rect 151782 404298 187226 404534
rect 187462 404298 187546 404534
rect 187782 404298 223226 404534
rect 223462 404298 223546 404534
rect 223782 404298 259226 404534
rect 259462 404298 259546 404534
rect 259782 404298 295226 404534
rect 295462 404298 295546 404534
rect 295782 404298 331226 404534
rect 331462 404298 331546 404534
rect 331782 404298 367226 404534
rect 367462 404298 367546 404534
rect 367782 404298 403226 404534
rect 403462 404298 403546 404534
rect 403782 404298 439226 404534
rect 439462 404298 439546 404534
rect 439782 404298 475226 404534
rect 475462 404298 475546 404534
rect 475782 404298 511226 404534
rect 511462 404298 511546 404534
rect 511782 404298 547226 404534
rect 547462 404298 547546 404534
rect 547782 404298 590142 404534
rect 590378 404298 590462 404534
rect 590698 404298 592650 404534
rect -8726 404266 592650 404298
rect -8726 403614 592650 403646
rect -8726 403378 -5814 403614
rect -5578 403378 -5494 403614
rect -5258 403378 5986 403614
rect 6222 403378 6306 403614
rect 6542 403378 41986 403614
rect 42222 403378 42306 403614
rect 42542 403378 77986 403614
rect 78222 403378 78306 403614
rect 78542 403378 113986 403614
rect 114222 403378 114306 403614
rect 114542 403378 149986 403614
rect 150222 403378 150306 403614
rect 150542 403378 185986 403614
rect 186222 403378 186306 403614
rect 186542 403378 221986 403614
rect 222222 403378 222306 403614
rect 222542 403378 257986 403614
rect 258222 403378 258306 403614
rect 258542 403378 293986 403614
rect 294222 403378 294306 403614
rect 294542 403378 329986 403614
rect 330222 403378 330306 403614
rect 330542 403378 365986 403614
rect 366222 403378 366306 403614
rect 366542 403378 401986 403614
rect 402222 403378 402306 403614
rect 402542 403378 437986 403614
rect 438222 403378 438306 403614
rect 438542 403378 473986 403614
rect 474222 403378 474306 403614
rect 474542 403378 509986 403614
rect 510222 403378 510306 403614
rect 510542 403378 581986 403614
rect 582222 403378 582306 403614
rect 582542 403378 589182 403614
rect 589418 403378 589502 403614
rect 589738 403378 592650 403614
rect -8726 403294 592650 403378
rect -8726 403058 -5814 403294
rect -5578 403058 -5494 403294
rect -5258 403058 5986 403294
rect 6222 403058 6306 403294
rect 6542 403058 41986 403294
rect 42222 403058 42306 403294
rect 42542 403058 77986 403294
rect 78222 403058 78306 403294
rect 78542 403058 113986 403294
rect 114222 403058 114306 403294
rect 114542 403058 149986 403294
rect 150222 403058 150306 403294
rect 150542 403058 185986 403294
rect 186222 403058 186306 403294
rect 186542 403058 221986 403294
rect 222222 403058 222306 403294
rect 222542 403058 257986 403294
rect 258222 403058 258306 403294
rect 258542 403058 293986 403294
rect 294222 403058 294306 403294
rect 294542 403058 329986 403294
rect 330222 403058 330306 403294
rect 330542 403058 365986 403294
rect 366222 403058 366306 403294
rect 366542 403058 401986 403294
rect 402222 403058 402306 403294
rect 402542 403058 437986 403294
rect 438222 403058 438306 403294
rect 438542 403058 473986 403294
rect 474222 403058 474306 403294
rect 474542 403058 509986 403294
rect 510222 403058 510306 403294
rect 510542 403058 581986 403294
rect 582222 403058 582306 403294
rect 582542 403058 589182 403294
rect 589418 403058 589502 403294
rect 589738 403058 592650 403294
rect -8726 403026 592650 403058
rect -8726 402374 592650 402406
rect -8726 402138 -4854 402374
rect -4618 402138 -4534 402374
rect -4298 402138 4746 402374
rect 4982 402138 5066 402374
rect 5302 402138 40746 402374
rect 40982 402138 41066 402374
rect 41302 402138 76746 402374
rect 76982 402138 77066 402374
rect 77302 402138 112746 402374
rect 112982 402138 113066 402374
rect 113302 402138 148746 402374
rect 148982 402138 149066 402374
rect 149302 402138 184746 402374
rect 184982 402138 185066 402374
rect 185302 402138 220746 402374
rect 220982 402138 221066 402374
rect 221302 402138 256746 402374
rect 256982 402138 257066 402374
rect 257302 402138 292746 402374
rect 292982 402138 293066 402374
rect 293302 402138 328746 402374
rect 328982 402138 329066 402374
rect 329302 402138 364746 402374
rect 364982 402138 365066 402374
rect 365302 402138 400746 402374
rect 400982 402138 401066 402374
rect 401302 402138 436746 402374
rect 436982 402138 437066 402374
rect 437302 402138 472746 402374
rect 472982 402138 473066 402374
rect 473302 402138 508746 402374
rect 508982 402138 509066 402374
rect 509302 402138 580746 402374
rect 580982 402138 581066 402374
rect 581302 402138 588222 402374
rect 588458 402138 588542 402374
rect 588778 402138 592650 402374
rect -8726 402054 592650 402138
rect -8726 401818 -4854 402054
rect -4618 401818 -4534 402054
rect -4298 401818 4746 402054
rect 4982 401818 5066 402054
rect 5302 401818 40746 402054
rect 40982 401818 41066 402054
rect 41302 401818 76746 402054
rect 76982 401818 77066 402054
rect 77302 401818 112746 402054
rect 112982 401818 113066 402054
rect 113302 401818 148746 402054
rect 148982 401818 149066 402054
rect 149302 401818 184746 402054
rect 184982 401818 185066 402054
rect 185302 401818 220746 402054
rect 220982 401818 221066 402054
rect 221302 401818 256746 402054
rect 256982 401818 257066 402054
rect 257302 401818 292746 402054
rect 292982 401818 293066 402054
rect 293302 401818 328746 402054
rect 328982 401818 329066 402054
rect 329302 401818 364746 402054
rect 364982 401818 365066 402054
rect 365302 401818 400746 402054
rect 400982 401818 401066 402054
rect 401302 401818 436746 402054
rect 436982 401818 437066 402054
rect 437302 401818 472746 402054
rect 472982 401818 473066 402054
rect 473302 401818 508746 402054
rect 508982 401818 509066 402054
rect 509302 401818 580746 402054
rect 580982 401818 581066 402054
rect 581302 401818 588222 402054
rect 588458 401818 588542 402054
rect 588778 401818 592650 402054
rect -8726 401786 592650 401818
rect -8726 401134 592650 401166
rect -8726 400898 -3894 401134
rect -3658 400898 -3574 401134
rect -3338 400898 3506 401134
rect 3742 400898 3826 401134
rect 4062 400898 39506 401134
rect 39742 400898 39826 401134
rect 40062 400898 75506 401134
rect 75742 400898 75826 401134
rect 76062 400898 111506 401134
rect 111742 400898 111826 401134
rect 112062 400898 147506 401134
rect 147742 400898 147826 401134
rect 148062 400898 183506 401134
rect 183742 400898 183826 401134
rect 184062 400898 219506 401134
rect 219742 400898 219826 401134
rect 220062 400898 255506 401134
rect 255742 400898 255826 401134
rect 256062 400898 291506 401134
rect 291742 400898 291826 401134
rect 292062 400898 327506 401134
rect 327742 400898 327826 401134
rect 328062 400898 363506 401134
rect 363742 400898 363826 401134
rect 364062 400898 399506 401134
rect 399742 400898 399826 401134
rect 400062 400898 435506 401134
rect 435742 400898 435826 401134
rect 436062 400898 471506 401134
rect 471742 400898 471826 401134
rect 472062 400898 507506 401134
rect 507742 400898 507826 401134
rect 508062 400898 579506 401134
rect 579742 400898 579826 401134
rect 580062 400898 587262 401134
rect 587498 400898 587582 401134
rect 587818 400898 592650 401134
rect -8726 400814 592650 400898
rect -8726 400578 -3894 400814
rect -3658 400578 -3574 400814
rect -3338 400578 3506 400814
rect 3742 400578 3826 400814
rect 4062 400578 39506 400814
rect 39742 400578 39826 400814
rect 40062 400578 75506 400814
rect 75742 400578 75826 400814
rect 76062 400578 111506 400814
rect 111742 400578 111826 400814
rect 112062 400578 147506 400814
rect 147742 400578 147826 400814
rect 148062 400578 183506 400814
rect 183742 400578 183826 400814
rect 184062 400578 219506 400814
rect 219742 400578 219826 400814
rect 220062 400578 255506 400814
rect 255742 400578 255826 400814
rect 256062 400578 291506 400814
rect 291742 400578 291826 400814
rect 292062 400578 327506 400814
rect 327742 400578 327826 400814
rect 328062 400578 363506 400814
rect 363742 400578 363826 400814
rect 364062 400578 399506 400814
rect 399742 400578 399826 400814
rect 400062 400578 435506 400814
rect 435742 400578 435826 400814
rect 436062 400578 471506 400814
rect 471742 400578 471826 400814
rect 472062 400578 507506 400814
rect 507742 400578 507826 400814
rect 508062 400578 579506 400814
rect 579742 400578 579826 400814
rect 580062 400578 587262 400814
rect 587498 400578 587582 400814
rect 587818 400578 592650 400814
rect -8726 400546 592650 400578
rect -8726 399894 592650 399926
rect -8726 399658 -2934 399894
rect -2698 399658 -2614 399894
rect -2378 399658 2266 399894
rect 2502 399658 2586 399894
rect 2822 399658 38266 399894
rect 38502 399658 38586 399894
rect 38822 399658 74266 399894
rect 74502 399658 74586 399894
rect 74822 399658 110266 399894
rect 110502 399658 110586 399894
rect 110822 399658 146266 399894
rect 146502 399658 146586 399894
rect 146822 399658 182266 399894
rect 182502 399658 182586 399894
rect 182822 399658 218266 399894
rect 218502 399658 218586 399894
rect 218822 399658 254266 399894
rect 254502 399658 254586 399894
rect 254822 399658 290266 399894
rect 290502 399658 290586 399894
rect 290822 399658 326266 399894
rect 326502 399658 326586 399894
rect 326822 399658 362266 399894
rect 362502 399658 362586 399894
rect 362822 399658 398266 399894
rect 398502 399658 398586 399894
rect 398822 399658 434266 399894
rect 434502 399658 434586 399894
rect 434822 399658 470266 399894
rect 470502 399658 470586 399894
rect 470822 399658 506266 399894
rect 506502 399658 506586 399894
rect 506822 399658 540918 399894
rect 541154 399658 542850 399894
rect 543086 399658 544782 399894
rect 545018 399658 546714 399894
rect 546950 399658 578266 399894
rect 578502 399658 578586 399894
rect 578822 399658 586302 399894
rect 586538 399658 586622 399894
rect 586858 399658 592650 399894
rect -8726 399574 592650 399658
rect -8726 399338 -2934 399574
rect -2698 399338 -2614 399574
rect -2378 399338 2266 399574
rect 2502 399338 2586 399574
rect 2822 399338 38266 399574
rect 38502 399338 38586 399574
rect 38822 399338 74266 399574
rect 74502 399338 74586 399574
rect 74822 399338 110266 399574
rect 110502 399338 110586 399574
rect 110822 399338 146266 399574
rect 146502 399338 146586 399574
rect 146822 399338 182266 399574
rect 182502 399338 182586 399574
rect 182822 399338 218266 399574
rect 218502 399338 218586 399574
rect 218822 399338 254266 399574
rect 254502 399338 254586 399574
rect 254822 399338 290266 399574
rect 290502 399338 290586 399574
rect 290822 399338 326266 399574
rect 326502 399338 326586 399574
rect 326822 399338 362266 399574
rect 362502 399338 362586 399574
rect 362822 399338 398266 399574
rect 398502 399338 398586 399574
rect 398822 399338 434266 399574
rect 434502 399338 434586 399574
rect 434822 399338 470266 399574
rect 470502 399338 470586 399574
rect 470822 399338 506266 399574
rect 506502 399338 506586 399574
rect 506822 399338 540918 399574
rect 541154 399338 542850 399574
rect 543086 399338 544782 399574
rect 545018 399338 546714 399574
rect 546950 399338 578266 399574
rect 578502 399338 578586 399574
rect 578822 399338 586302 399574
rect 586538 399338 586622 399574
rect 586858 399338 592650 399574
rect -8726 399306 592650 399338
rect -8726 398654 592650 398686
rect -8726 398418 -1974 398654
rect -1738 398418 -1654 398654
rect -1418 398418 1026 398654
rect 1262 398418 1346 398654
rect 1582 398418 37026 398654
rect 37262 398418 37346 398654
rect 37582 398418 73026 398654
rect 73262 398418 73346 398654
rect 73582 398418 109026 398654
rect 109262 398418 109346 398654
rect 109582 398418 145026 398654
rect 145262 398418 145346 398654
rect 145582 398418 181026 398654
rect 181262 398418 181346 398654
rect 181582 398418 217026 398654
rect 217262 398418 217346 398654
rect 217582 398418 253026 398654
rect 253262 398418 253346 398654
rect 253582 398418 289026 398654
rect 289262 398418 289346 398654
rect 289582 398418 325026 398654
rect 325262 398418 325346 398654
rect 325582 398418 361026 398654
rect 361262 398418 361346 398654
rect 361582 398418 397026 398654
rect 397262 398418 397346 398654
rect 397582 398418 433026 398654
rect 433262 398418 433346 398654
rect 433582 398418 469026 398654
rect 469262 398418 469346 398654
rect 469582 398418 505026 398654
rect 505262 398418 505346 398654
rect 505582 398418 539952 398654
rect 540188 398418 541884 398654
rect 542120 398418 543816 398654
rect 544052 398418 545748 398654
rect 545984 398418 577026 398654
rect 577262 398418 577346 398654
rect 577582 398418 585342 398654
rect 585578 398418 585662 398654
rect 585898 398418 592650 398654
rect -8726 398334 592650 398418
rect -8726 398098 -1974 398334
rect -1738 398098 -1654 398334
rect -1418 398098 1026 398334
rect 1262 398098 1346 398334
rect 1582 398098 37026 398334
rect 37262 398098 37346 398334
rect 37582 398098 73026 398334
rect 73262 398098 73346 398334
rect 73582 398098 109026 398334
rect 109262 398098 109346 398334
rect 109582 398098 145026 398334
rect 145262 398098 145346 398334
rect 145582 398098 181026 398334
rect 181262 398098 181346 398334
rect 181582 398098 217026 398334
rect 217262 398098 217346 398334
rect 217582 398098 253026 398334
rect 253262 398098 253346 398334
rect 253582 398098 289026 398334
rect 289262 398098 289346 398334
rect 289582 398098 325026 398334
rect 325262 398098 325346 398334
rect 325582 398098 361026 398334
rect 361262 398098 361346 398334
rect 361582 398098 397026 398334
rect 397262 398098 397346 398334
rect 397582 398098 433026 398334
rect 433262 398098 433346 398334
rect 433582 398098 469026 398334
rect 469262 398098 469346 398334
rect 469582 398098 505026 398334
rect 505262 398098 505346 398334
rect 505582 398098 539952 398334
rect 540188 398098 541884 398334
rect 542120 398098 543816 398334
rect 544052 398098 545748 398334
rect 545984 398098 577026 398334
rect 577262 398098 577346 398334
rect 577582 398098 585342 398334
rect 585578 398098 585662 398334
rect 585898 398098 592650 398334
rect -8726 398066 592650 398098
rect -8726 371334 592650 371366
rect -8726 371098 -8694 371334
rect -8458 371098 -8374 371334
rect -8138 371098 9706 371334
rect 9942 371098 10026 371334
rect 10262 371098 45706 371334
rect 45942 371098 46026 371334
rect 46262 371098 81706 371334
rect 81942 371098 82026 371334
rect 82262 371098 117706 371334
rect 117942 371098 118026 371334
rect 118262 371098 153706 371334
rect 153942 371098 154026 371334
rect 154262 371098 189706 371334
rect 189942 371098 190026 371334
rect 190262 371098 225706 371334
rect 225942 371098 226026 371334
rect 226262 371098 261706 371334
rect 261942 371098 262026 371334
rect 262262 371098 297706 371334
rect 297942 371098 298026 371334
rect 298262 371098 333706 371334
rect 333942 371098 334026 371334
rect 334262 371098 369706 371334
rect 369942 371098 370026 371334
rect 370262 371098 405706 371334
rect 405942 371098 406026 371334
rect 406262 371098 441706 371334
rect 441942 371098 442026 371334
rect 442262 371098 477706 371334
rect 477942 371098 478026 371334
rect 478262 371098 513706 371334
rect 513942 371098 514026 371334
rect 514262 371098 549706 371334
rect 549942 371098 550026 371334
rect 550262 371098 592062 371334
rect 592298 371098 592382 371334
rect 592618 371098 592650 371334
rect -8726 371014 592650 371098
rect -8726 370778 -8694 371014
rect -8458 370778 -8374 371014
rect -8138 370778 9706 371014
rect 9942 370778 10026 371014
rect 10262 370778 45706 371014
rect 45942 370778 46026 371014
rect 46262 370778 81706 371014
rect 81942 370778 82026 371014
rect 82262 370778 117706 371014
rect 117942 370778 118026 371014
rect 118262 370778 153706 371014
rect 153942 370778 154026 371014
rect 154262 370778 189706 371014
rect 189942 370778 190026 371014
rect 190262 370778 225706 371014
rect 225942 370778 226026 371014
rect 226262 370778 261706 371014
rect 261942 370778 262026 371014
rect 262262 370778 297706 371014
rect 297942 370778 298026 371014
rect 298262 370778 333706 371014
rect 333942 370778 334026 371014
rect 334262 370778 369706 371014
rect 369942 370778 370026 371014
rect 370262 370778 405706 371014
rect 405942 370778 406026 371014
rect 406262 370778 441706 371014
rect 441942 370778 442026 371014
rect 442262 370778 477706 371014
rect 477942 370778 478026 371014
rect 478262 370778 513706 371014
rect 513942 370778 514026 371014
rect 514262 370778 549706 371014
rect 549942 370778 550026 371014
rect 550262 370778 592062 371014
rect 592298 370778 592382 371014
rect 592618 370778 592650 371014
rect -8726 370746 592650 370778
rect -8726 370094 592650 370126
rect -8726 369858 -7734 370094
rect -7498 369858 -7414 370094
rect -7178 369858 8466 370094
rect 8702 369858 8786 370094
rect 9022 369858 44466 370094
rect 44702 369858 44786 370094
rect 45022 369858 80466 370094
rect 80702 369858 80786 370094
rect 81022 369858 116466 370094
rect 116702 369858 116786 370094
rect 117022 369858 152466 370094
rect 152702 369858 152786 370094
rect 153022 369858 188466 370094
rect 188702 369858 188786 370094
rect 189022 369858 224466 370094
rect 224702 369858 224786 370094
rect 225022 369858 260466 370094
rect 260702 369858 260786 370094
rect 261022 369858 296466 370094
rect 296702 369858 296786 370094
rect 297022 369858 332466 370094
rect 332702 369858 332786 370094
rect 333022 369858 368466 370094
rect 368702 369858 368786 370094
rect 369022 369858 404466 370094
rect 404702 369858 404786 370094
rect 405022 369858 440466 370094
rect 440702 369858 440786 370094
rect 441022 369858 476466 370094
rect 476702 369858 476786 370094
rect 477022 369858 512466 370094
rect 512702 369858 512786 370094
rect 513022 369858 548466 370094
rect 548702 369858 548786 370094
rect 549022 369858 591102 370094
rect 591338 369858 591422 370094
rect 591658 369858 592650 370094
rect -8726 369774 592650 369858
rect -8726 369538 -7734 369774
rect -7498 369538 -7414 369774
rect -7178 369538 8466 369774
rect 8702 369538 8786 369774
rect 9022 369538 44466 369774
rect 44702 369538 44786 369774
rect 45022 369538 80466 369774
rect 80702 369538 80786 369774
rect 81022 369538 116466 369774
rect 116702 369538 116786 369774
rect 117022 369538 152466 369774
rect 152702 369538 152786 369774
rect 153022 369538 188466 369774
rect 188702 369538 188786 369774
rect 189022 369538 224466 369774
rect 224702 369538 224786 369774
rect 225022 369538 260466 369774
rect 260702 369538 260786 369774
rect 261022 369538 296466 369774
rect 296702 369538 296786 369774
rect 297022 369538 332466 369774
rect 332702 369538 332786 369774
rect 333022 369538 368466 369774
rect 368702 369538 368786 369774
rect 369022 369538 404466 369774
rect 404702 369538 404786 369774
rect 405022 369538 440466 369774
rect 440702 369538 440786 369774
rect 441022 369538 476466 369774
rect 476702 369538 476786 369774
rect 477022 369538 512466 369774
rect 512702 369538 512786 369774
rect 513022 369538 548466 369774
rect 548702 369538 548786 369774
rect 549022 369538 591102 369774
rect 591338 369538 591422 369774
rect 591658 369538 592650 369774
rect -8726 369506 592650 369538
rect -8726 368854 592650 368886
rect -8726 368618 -6774 368854
rect -6538 368618 -6454 368854
rect -6218 368618 7226 368854
rect 7462 368618 7546 368854
rect 7782 368618 43226 368854
rect 43462 368618 43546 368854
rect 43782 368618 79226 368854
rect 79462 368618 79546 368854
rect 79782 368618 115226 368854
rect 115462 368618 115546 368854
rect 115782 368618 151226 368854
rect 151462 368618 151546 368854
rect 151782 368618 187226 368854
rect 187462 368618 187546 368854
rect 187782 368618 223226 368854
rect 223462 368618 223546 368854
rect 223782 368618 259226 368854
rect 259462 368618 259546 368854
rect 259782 368618 295226 368854
rect 295462 368618 295546 368854
rect 295782 368618 331226 368854
rect 331462 368618 331546 368854
rect 331782 368618 367226 368854
rect 367462 368618 367546 368854
rect 367782 368618 403226 368854
rect 403462 368618 403546 368854
rect 403782 368618 439226 368854
rect 439462 368618 439546 368854
rect 439782 368618 475226 368854
rect 475462 368618 475546 368854
rect 475782 368618 511226 368854
rect 511462 368618 511546 368854
rect 511782 368618 547226 368854
rect 547462 368618 547546 368854
rect 547782 368618 590142 368854
rect 590378 368618 590462 368854
rect 590698 368618 592650 368854
rect -8726 368534 592650 368618
rect -8726 368298 -6774 368534
rect -6538 368298 -6454 368534
rect -6218 368298 7226 368534
rect 7462 368298 7546 368534
rect 7782 368298 43226 368534
rect 43462 368298 43546 368534
rect 43782 368298 79226 368534
rect 79462 368298 79546 368534
rect 79782 368298 115226 368534
rect 115462 368298 115546 368534
rect 115782 368298 151226 368534
rect 151462 368298 151546 368534
rect 151782 368298 187226 368534
rect 187462 368298 187546 368534
rect 187782 368298 223226 368534
rect 223462 368298 223546 368534
rect 223782 368298 259226 368534
rect 259462 368298 259546 368534
rect 259782 368298 295226 368534
rect 295462 368298 295546 368534
rect 295782 368298 331226 368534
rect 331462 368298 331546 368534
rect 331782 368298 367226 368534
rect 367462 368298 367546 368534
rect 367782 368298 403226 368534
rect 403462 368298 403546 368534
rect 403782 368298 439226 368534
rect 439462 368298 439546 368534
rect 439782 368298 475226 368534
rect 475462 368298 475546 368534
rect 475782 368298 511226 368534
rect 511462 368298 511546 368534
rect 511782 368298 547226 368534
rect 547462 368298 547546 368534
rect 547782 368298 590142 368534
rect 590378 368298 590462 368534
rect 590698 368298 592650 368534
rect -8726 368266 592650 368298
rect -8726 367614 592650 367646
rect -8726 367378 -5814 367614
rect -5578 367378 -5494 367614
rect -5258 367378 5986 367614
rect 6222 367378 6306 367614
rect 6542 367378 41986 367614
rect 42222 367378 42306 367614
rect 42542 367378 77986 367614
rect 78222 367378 78306 367614
rect 78542 367378 113986 367614
rect 114222 367378 114306 367614
rect 114542 367378 149986 367614
rect 150222 367378 150306 367614
rect 150542 367378 185986 367614
rect 186222 367378 186306 367614
rect 186542 367378 221986 367614
rect 222222 367378 222306 367614
rect 222542 367378 257986 367614
rect 258222 367378 258306 367614
rect 258542 367378 293986 367614
rect 294222 367378 294306 367614
rect 294542 367378 329986 367614
rect 330222 367378 330306 367614
rect 330542 367378 365986 367614
rect 366222 367378 366306 367614
rect 366542 367378 401986 367614
rect 402222 367378 402306 367614
rect 402542 367378 437986 367614
rect 438222 367378 438306 367614
rect 438542 367378 473986 367614
rect 474222 367378 474306 367614
rect 474542 367378 509986 367614
rect 510222 367378 510306 367614
rect 510542 367378 581986 367614
rect 582222 367378 582306 367614
rect 582542 367378 589182 367614
rect 589418 367378 589502 367614
rect 589738 367378 592650 367614
rect -8726 367294 592650 367378
rect -8726 367058 -5814 367294
rect -5578 367058 -5494 367294
rect -5258 367058 5986 367294
rect 6222 367058 6306 367294
rect 6542 367058 41986 367294
rect 42222 367058 42306 367294
rect 42542 367058 77986 367294
rect 78222 367058 78306 367294
rect 78542 367058 113986 367294
rect 114222 367058 114306 367294
rect 114542 367058 149986 367294
rect 150222 367058 150306 367294
rect 150542 367058 185986 367294
rect 186222 367058 186306 367294
rect 186542 367058 221986 367294
rect 222222 367058 222306 367294
rect 222542 367058 257986 367294
rect 258222 367058 258306 367294
rect 258542 367058 293986 367294
rect 294222 367058 294306 367294
rect 294542 367058 329986 367294
rect 330222 367058 330306 367294
rect 330542 367058 365986 367294
rect 366222 367058 366306 367294
rect 366542 367058 401986 367294
rect 402222 367058 402306 367294
rect 402542 367058 437986 367294
rect 438222 367058 438306 367294
rect 438542 367058 473986 367294
rect 474222 367058 474306 367294
rect 474542 367058 509986 367294
rect 510222 367058 510306 367294
rect 510542 367058 581986 367294
rect 582222 367058 582306 367294
rect 582542 367058 589182 367294
rect 589418 367058 589502 367294
rect 589738 367058 592650 367294
rect -8726 367026 592650 367058
rect -8726 366374 592650 366406
rect -8726 366138 -4854 366374
rect -4618 366138 -4534 366374
rect -4298 366138 4746 366374
rect 4982 366138 5066 366374
rect 5302 366138 40746 366374
rect 40982 366138 41066 366374
rect 41302 366138 76746 366374
rect 76982 366138 77066 366374
rect 77302 366138 112746 366374
rect 112982 366138 113066 366374
rect 113302 366138 148746 366374
rect 148982 366138 149066 366374
rect 149302 366138 184746 366374
rect 184982 366138 185066 366374
rect 185302 366138 220746 366374
rect 220982 366138 221066 366374
rect 221302 366138 256746 366374
rect 256982 366138 257066 366374
rect 257302 366138 292746 366374
rect 292982 366138 293066 366374
rect 293302 366138 328746 366374
rect 328982 366138 329066 366374
rect 329302 366138 364746 366374
rect 364982 366138 365066 366374
rect 365302 366138 400746 366374
rect 400982 366138 401066 366374
rect 401302 366138 436746 366374
rect 436982 366138 437066 366374
rect 437302 366138 472746 366374
rect 472982 366138 473066 366374
rect 473302 366138 508746 366374
rect 508982 366138 509066 366374
rect 509302 366138 580746 366374
rect 580982 366138 581066 366374
rect 581302 366138 588222 366374
rect 588458 366138 588542 366374
rect 588778 366138 592650 366374
rect -8726 366054 592650 366138
rect -8726 365818 -4854 366054
rect -4618 365818 -4534 366054
rect -4298 365818 4746 366054
rect 4982 365818 5066 366054
rect 5302 365818 40746 366054
rect 40982 365818 41066 366054
rect 41302 365818 76746 366054
rect 76982 365818 77066 366054
rect 77302 365818 112746 366054
rect 112982 365818 113066 366054
rect 113302 365818 148746 366054
rect 148982 365818 149066 366054
rect 149302 365818 184746 366054
rect 184982 365818 185066 366054
rect 185302 365818 220746 366054
rect 220982 365818 221066 366054
rect 221302 365818 256746 366054
rect 256982 365818 257066 366054
rect 257302 365818 292746 366054
rect 292982 365818 293066 366054
rect 293302 365818 328746 366054
rect 328982 365818 329066 366054
rect 329302 365818 364746 366054
rect 364982 365818 365066 366054
rect 365302 365818 400746 366054
rect 400982 365818 401066 366054
rect 401302 365818 436746 366054
rect 436982 365818 437066 366054
rect 437302 365818 472746 366054
rect 472982 365818 473066 366054
rect 473302 365818 508746 366054
rect 508982 365818 509066 366054
rect 509302 365818 580746 366054
rect 580982 365818 581066 366054
rect 581302 365818 588222 366054
rect 588458 365818 588542 366054
rect 588778 365818 592650 366054
rect -8726 365786 592650 365818
rect -8726 365134 592650 365166
rect -8726 364898 -3894 365134
rect -3658 364898 -3574 365134
rect -3338 364898 3506 365134
rect 3742 364898 3826 365134
rect 4062 364898 39506 365134
rect 39742 364898 39826 365134
rect 40062 364898 75506 365134
rect 75742 364898 75826 365134
rect 76062 364898 111506 365134
rect 111742 364898 111826 365134
rect 112062 364898 147506 365134
rect 147742 364898 147826 365134
rect 148062 364898 183506 365134
rect 183742 364898 183826 365134
rect 184062 364898 219506 365134
rect 219742 364898 219826 365134
rect 220062 364898 255506 365134
rect 255742 364898 255826 365134
rect 256062 364898 291506 365134
rect 291742 364898 291826 365134
rect 292062 364898 327506 365134
rect 327742 364898 327826 365134
rect 328062 364898 363506 365134
rect 363742 364898 363826 365134
rect 364062 364898 399506 365134
rect 399742 364898 399826 365134
rect 400062 364898 435506 365134
rect 435742 364898 435826 365134
rect 436062 364898 471506 365134
rect 471742 364898 471826 365134
rect 472062 364898 507506 365134
rect 507742 364898 507826 365134
rect 508062 364898 579506 365134
rect 579742 364898 579826 365134
rect 580062 364898 587262 365134
rect 587498 364898 587582 365134
rect 587818 364898 592650 365134
rect -8726 364814 592650 364898
rect -8726 364578 -3894 364814
rect -3658 364578 -3574 364814
rect -3338 364578 3506 364814
rect 3742 364578 3826 364814
rect 4062 364578 39506 364814
rect 39742 364578 39826 364814
rect 40062 364578 75506 364814
rect 75742 364578 75826 364814
rect 76062 364578 111506 364814
rect 111742 364578 111826 364814
rect 112062 364578 147506 364814
rect 147742 364578 147826 364814
rect 148062 364578 183506 364814
rect 183742 364578 183826 364814
rect 184062 364578 219506 364814
rect 219742 364578 219826 364814
rect 220062 364578 255506 364814
rect 255742 364578 255826 364814
rect 256062 364578 291506 364814
rect 291742 364578 291826 364814
rect 292062 364578 327506 364814
rect 327742 364578 327826 364814
rect 328062 364578 363506 364814
rect 363742 364578 363826 364814
rect 364062 364578 399506 364814
rect 399742 364578 399826 364814
rect 400062 364578 435506 364814
rect 435742 364578 435826 364814
rect 436062 364578 471506 364814
rect 471742 364578 471826 364814
rect 472062 364578 507506 364814
rect 507742 364578 507826 364814
rect 508062 364578 579506 364814
rect 579742 364578 579826 364814
rect 580062 364578 587262 364814
rect 587498 364578 587582 364814
rect 587818 364578 592650 364814
rect -8726 364546 592650 364578
rect -8726 363894 592650 363926
rect -8726 363658 -2934 363894
rect -2698 363658 -2614 363894
rect -2378 363658 2266 363894
rect 2502 363658 2586 363894
rect 2822 363658 38266 363894
rect 38502 363658 38586 363894
rect 38822 363658 74266 363894
rect 74502 363658 74586 363894
rect 74822 363658 110266 363894
rect 110502 363658 110586 363894
rect 110822 363658 146266 363894
rect 146502 363658 146586 363894
rect 146822 363658 182266 363894
rect 182502 363658 182586 363894
rect 182822 363658 218266 363894
rect 218502 363658 218586 363894
rect 218822 363658 254266 363894
rect 254502 363658 254586 363894
rect 254822 363658 290266 363894
rect 290502 363658 290586 363894
rect 290822 363658 326266 363894
rect 326502 363658 326586 363894
rect 326822 363658 362266 363894
rect 362502 363658 362586 363894
rect 362822 363658 398266 363894
rect 398502 363658 398586 363894
rect 398822 363658 434266 363894
rect 434502 363658 434586 363894
rect 434822 363658 470266 363894
rect 470502 363658 470586 363894
rect 470822 363658 506266 363894
rect 506502 363658 506586 363894
rect 506822 363658 540918 363894
rect 541154 363658 542850 363894
rect 543086 363658 544782 363894
rect 545018 363658 546714 363894
rect 546950 363658 578266 363894
rect 578502 363658 578586 363894
rect 578822 363658 586302 363894
rect 586538 363658 586622 363894
rect 586858 363658 592650 363894
rect -8726 363574 592650 363658
rect -8726 363338 -2934 363574
rect -2698 363338 -2614 363574
rect -2378 363338 2266 363574
rect 2502 363338 2586 363574
rect 2822 363338 38266 363574
rect 38502 363338 38586 363574
rect 38822 363338 74266 363574
rect 74502 363338 74586 363574
rect 74822 363338 110266 363574
rect 110502 363338 110586 363574
rect 110822 363338 146266 363574
rect 146502 363338 146586 363574
rect 146822 363338 182266 363574
rect 182502 363338 182586 363574
rect 182822 363338 218266 363574
rect 218502 363338 218586 363574
rect 218822 363338 254266 363574
rect 254502 363338 254586 363574
rect 254822 363338 290266 363574
rect 290502 363338 290586 363574
rect 290822 363338 326266 363574
rect 326502 363338 326586 363574
rect 326822 363338 362266 363574
rect 362502 363338 362586 363574
rect 362822 363338 398266 363574
rect 398502 363338 398586 363574
rect 398822 363338 434266 363574
rect 434502 363338 434586 363574
rect 434822 363338 470266 363574
rect 470502 363338 470586 363574
rect 470822 363338 506266 363574
rect 506502 363338 506586 363574
rect 506822 363338 540918 363574
rect 541154 363338 542850 363574
rect 543086 363338 544782 363574
rect 545018 363338 546714 363574
rect 546950 363338 578266 363574
rect 578502 363338 578586 363574
rect 578822 363338 586302 363574
rect 586538 363338 586622 363574
rect 586858 363338 592650 363574
rect -8726 363306 592650 363338
rect -8726 362654 592650 362686
rect -8726 362418 -1974 362654
rect -1738 362418 -1654 362654
rect -1418 362418 1026 362654
rect 1262 362418 1346 362654
rect 1582 362418 37026 362654
rect 37262 362418 37346 362654
rect 37582 362418 73026 362654
rect 73262 362418 73346 362654
rect 73582 362418 109026 362654
rect 109262 362418 109346 362654
rect 109582 362418 145026 362654
rect 145262 362418 145346 362654
rect 145582 362418 181026 362654
rect 181262 362418 181346 362654
rect 181582 362418 217026 362654
rect 217262 362418 217346 362654
rect 217582 362418 253026 362654
rect 253262 362418 253346 362654
rect 253582 362418 289026 362654
rect 289262 362418 289346 362654
rect 289582 362418 325026 362654
rect 325262 362418 325346 362654
rect 325582 362418 361026 362654
rect 361262 362418 361346 362654
rect 361582 362418 397026 362654
rect 397262 362418 397346 362654
rect 397582 362418 433026 362654
rect 433262 362418 433346 362654
rect 433582 362418 469026 362654
rect 469262 362418 469346 362654
rect 469582 362418 505026 362654
rect 505262 362418 505346 362654
rect 505582 362418 539952 362654
rect 540188 362418 541884 362654
rect 542120 362418 543816 362654
rect 544052 362418 545748 362654
rect 545984 362418 577026 362654
rect 577262 362418 577346 362654
rect 577582 362418 585342 362654
rect 585578 362418 585662 362654
rect 585898 362418 592650 362654
rect -8726 362334 592650 362418
rect -8726 362098 -1974 362334
rect -1738 362098 -1654 362334
rect -1418 362098 1026 362334
rect 1262 362098 1346 362334
rect 1582 362098 37026 362334
rect 37262 362098 37346 362334
rect 37582 362098 73026 362334
rect 73262 362098 73346 362334
rect 73582 362098 109026 362334
rect 109262 362098 109346 362334
rect 109582 362098 145026 362334
rect 145262 362098 145346 362334
rect 145582 362098 181026 362334
rect 181262 362098 181346 362334
rect 181582 362098 217026 362334
rect 217262 362098 217346 362334
rect 217582 362098 253026 362334
rect 253262 362098 253346 362334
rect 253582 362098 289026 362334
rect 289262 362098 289346 362334
rect 289582 362098 325026 362334
rect 325262 362098 325346 362334
rect 325582 362098 361026 362334
rect 361262 362098 361346 362334
rect 361582 362098 397026 362334
rect 397262 362098 397346 362334
rect 397582 362098 433026 362334
rect 433262 362098 433346 362334
rect 433582 362098 469026 362334
rect 469262 362098 469346 362334
rect 469582 362098 505026 362334
rect 505262 362098 505346 362334
rect 505582 362098 539952 362334
rect 540188 362098 541884 362334
rect 542120 362098 543816 362334
rect 544052 362098 545748 362334
rect 545984 362098 577026 362334
rect 577262 362098 577346 362334
rect 577582 362098 585342 362334
rect 585578 362098 585662 362334
rect 585898 362098 592650 362334
rect -8726 362066 592650 362098
rect -8726 335334 592650 335366
rect -8726 335098 -8694 335334
rect -8458 335098 -8374 335334
rect -8138 335098 9706 335334
rect 9942 335098 10026 335334
rect 10262 335098 45706 335334
rect 45942 335098 46026 335334
rect 46262 335098 81706 335334
rect 81942 335098 82026 335334
rect 82262 335098 117706 335334
rect 117942 335098 118026 335334
rect 118262 335098 153706 335334
rect 153942 335098 154026 335334
rect 154262 335098 189706 335334
rect 189942 335098 190026 335334
rect 190262 335098 225706 335334
rect 225942 335098 226026 335334
rect 226262 335098 261706 335334
rect 261942 335098 262026 335334
rect 262262 335098 297706 335334
rect 297942 335098 298026 335334
rect 298262 335098 333706 335334
rect 333942 335098 334026 335334
rect 334262 335098 369706 335334
rect 369942 335098 370026 335334
rect 370262 335098 405706 335334
rect 405942 335098 406026 335334
rect 406262 335098 441706 335334
rect 441942 335098 442026 335334
rect 442262 335098 477706 335334
rect 477942 335098 478026 335334
rect 478262 335098 513706 335334
rect 513942 335098 514026 335334
rect 514262 335098 549706 335334
rect 549942 335098 550026 335334
rect 550262 335098 592062 335334
rect 592298 335098 592382 335334
rect 592618 335098 592650 335334
rect -8726 335014 592650 335098
rect -8726 334778 -8694 335014
rect -8458 334778 -8374 335014
rect -8138 334778 9706 335014
rect 9942 334778 10026 335014
rect 10262 334778 45706 335014
rect 45942 334778 46026 335014
rect 46262 334778 81706 335014
rect 81942 334778 82026 335014
rect 82262 334778 117706 335014
rect 117942 334778 118026 335014
rect 118262 334778 153706 335014
rect 153942 334778 154026 335014
rect 154262 334778 189706 335014
rect 189942 334778 190026 335014
rect 190262 334778 225706 335014
rect 225942 334778 226026 335014
rect 226262 334778 261706 335014
rect 261942 334778 262026 335014
rect 262262 334778 297706 335014
rect 297942 334778 298026 335014
rect 298262 334778 333706 335014
rect 333942 334778 334026 335014
rect 334262 334778 369706 335014
rect 369942 334778 370026 335014
rect 370262 334778 405706 335014
rect 405942 334778 406026 335014
rect 406262 334778 441706 335014
rect 441942 334778 442026 335014
rect 442262 334778 477706 335014
rect 477942 334778 478026 335014
rect 478262 334778 513706 335014
rect 513942 334778 514026 335014
rect 514262 334778 549706 335014
rect 549942 334778 550026 335014
rect 550262 334778 592062 335014
rect 592298 334778 592382 335014
rect 592618 334778 592650 335014
rect -8726 334746 592650 334778
rect -8726 334094 592650 334126
rect -8726 333858 -7734 334094
rect -7498 333858 -7414 334094
rect -7178 333858 8466 334094
rect 8702 333858 8786 334094
rect 9022 333858 44466 334094
rect 44702 333858 44786 334094
rect 45022 333858 80466 334094
rect 80702 333858 80786 334094
rect 81022 333858 116466 334094
rect 116702 333858 116786 334094
rect 117022 333858 152466 334094
rect 152702 333858 152786 334094
rect 153022 333858 188466 334094
rect 188702 333858 188786 334094
rect 189022 333858 224466 334094
rect 224702 333858 224786 334094
rect 225022 333858 260466 334094
rect 260702 333858 260786 334094
rect 261022 333858 296466 334094
rect 296702 333858 296786 334094
rect 297022 333858 332466 334094
rect 332702 333858 332786 334094
rect 333022 333858 368466 334094
rect 368702 333858 368786 334094
rect 369022 333858 404466 334094
rect 404702 333858 404786 334094
rect 405022 333858 440466 334094
rect 440702 333858 440786 334094
rect 441022 333858 476466 334094
rect 476702 333858 476786 334094
rect 477022 333858 512466 334094
rect 512702 333858 512786 334094
rect 513022 333858 548466 334094
rect 548702 333858 548786 334094
rect 549022 333858 591102 334094
rect 591338 333858 591422 334094
rect 591658 333858 592650 334094
rect -8726 333774 592650 333858
rect -8726 333538 -7734 333774
rect -7498 333538 -7414 333774
rect -7178 333538 8466 333774
rect 8702 333538 8786 333774
rect 9022 333538 44466 333774
rect 44702 333538 44786 333774
rect 45022 333538 80466 333774
rect 80702 333538 80786 333774
rect 81022 333538 116466 333774
rect 116702 333538 116786 333774
rect 117022 333538 152466 333774
rect 152702 333538 152786 333774
rect 153022 333538 188466 333774
rect 188702 333538 188786 333774
rect 189022 333538 224466 333774
rect 224702 333538 224786 333774
rect 225022 333538 260466 333774
rect 260702 333538 260786 333774
rect 261022 333538 296466 333774
rect 296702 333538 296786 333774
rect 297022 333538 332466 333774
rect 332702 333538 332786 333774
rect 333022 333538 368466 333774
rect 368702 333538 368786 333774
rect 369022 333538 404466 333774
rect 404702 333538 404786 333774
rect 405022 333538 440466 333774
rect 440702 333538 440786 333774
rect 441022 333538 476466 333774
rect 476702 333538 476786 333774
rect 477022 333538 512466 333774
rect 512702 333538 512786 333774
rect 513022 333538 548466 333774
rect 548702 333538 548786 333774
rect 549022 333538 591102 333774
rect 591338 333538 591422 333774
rect 591658 333538 592650 333774
rect -8726 333506 592650 333538
rect -8726 332854 592650 332886
rect -8726 332618 -6774 332854
rect -6538 332618 -6454 332854
rect -6218 332618 7226 332854
rect 7462 332618 7546 332854
rect 7782 332618 43226 332854
rect 43462 332618 43546 332854
rect 43782 332618 79226 332854
rect 79462 332618 79546 332854
rect 79782 332618 115226 332854
rect 115462 332618 115546 332854
rect 115782 332618 151226 332854
rect 151462 332618 151546 332854
rect 151782 332618 187226 332854
rect 187462 332618 187546 332854
rect 187782 332618 223226 332854
rect 223462 332618 223546 332854
rect 223782 332618 259226 332854
rect 259462 332618 259546 332854
rect 259782 332618 295226 332854
rect 295462 332618 295546 332854
rect 295782 332618 331226 332854
rect 331462 332618 331546 332854
rect 331782 332618 367226 332854
rect 367462 332618 367546 332854
rect 367782 332618 403226 332854
rect 403462 332618 403546 332854
rect 403782 332618 439226 332854
rect 439462 332618 439546 332854
rect 439782 332618 475226 332854
rect 475462 332618 475546 332854
rect 475782 332618 511226 332854
rect 511462 332618 511546 332854
rect 511782 332618 547226 332854
rect 547462 332618 547546 332854
rect 547782 332618 590142 332854
rect 590378 332618 590462 332854
rect 590698 332618 592650 332854
rect -8726 332534 592650 332618
rect -8726 332298 -6774 332534
rect -6538 332298 -6454 332534
rect -6218 332298 7226 332534
rect 7462 332298 7546 332534
rect 7782 332298 43226 332534
rect 43462 332298 43546 332534
rect 43782 332298 79226 332534
rect 79462 332298 79546 332534
rect 79782 332298 115226 332534
rect 115462 332298 115546 332534
rect 115782 332298 151226 332534
rect 151462 332298 151546 332534
rect 151782 332298 187226 332534
rect 187462 332298 187546 332534
rect 187782 332298 223226 332534
rect 223462 332298 223546 332534
rect 223782 332298 259226 332534
rect 259462 332298 259546 332534
rect 259782 332298 295226 332534
rect 295462 332298 295546 332534
rect 295782 332298 331226 332534
rect 331462 332298 331546 332534
rect 331782 332298 367226 332534
rect 367462 332298 367546 332534
rect 367782 332298 403226 332534
rect 403462 332298 403546 332534
rect 403782 332298 439226 332534
rect 439462 332298 439546 332534
rect 439782 332298 475226 332534
rect 475462 332298 475546 332534
rect 475782 332298 511226 332534
rect 511462 332298 511546 332534
rect 511782 332298 547226 332534
rect 547462 332298 547546 332534
rect 547782 332298 590142 332534
rect 590378 332298 590462 332534
rect 590698 332298 592650 332534
rect -8726 332266 592650 332298
rect -8726 331614 592650 331646
rect -8726 331378 -5814 331614
rect -5578 331378 -5494 331614
rect -5258 331378 5986 331614
rect 6222 331378 6306 331614
rect 6542 331378 41986 331614
rect 42222 331378 42306 331614
rect 42542 331378 77986 331614
rect 78222 331378 78306 331614
rect 78542 331378 113986 331614
rect 114222 331378 114306 331614
rect 114542 331378 149986 331614
rect 150222 331378 150306 331614
rect 150542 331378 185986 331614
rect 186222 331378 186306 331614
rect 186542 331378 221986 331614
rect 222222 331378 222306 331614
rect 222542 331378 257986 331614
rect 258222 331378 258306 331614
rect 258542 331378 293986 331614
rect 294222 331378 294306 331614
rect 294542 331378 329986 331614
rect 330222 331378 330306 331614
rect 330542 331378 365986 331614
rect 366222 331378 366306 331614
rect 366542 331378 401986 331614
rect 402222 331378 402306 331614
rect 402542 331378 437986 331614
rect 438222 331378 438306 331614
rect 438542 331378 473986 331614
rect 474222 331378 474306 331614
rect 474542 331378 509986 331614
rect 510222 331378 510306 331614
rect 510542 331378 581986 331614
rect 582222 331378 582306 331614
rect 582542 331378 589182 331614
rect 589418 331378 589502 331614
rect 589738 331378 592650 331614
rect -8726 331294 592650 331378
rect -8726 331058 -5814 331294
rect -5578 331058 -5494 331294
rect -5258 331058 5986 331294
rect 6222 331058 6306 331294
rect 6542 331058 41986 331294
rect 42222 331058 42306 331294
rect 42542 331058 77986 331294
rect 78222 331058 78306 331294
rect 78542 331058 113986 331294
rect 114222 331058 114306 331294
rect 114542 331058 149986 331294
rect 150222 331058 150306 331294
rect 150542 331058 185986 331294
rect 186222 331058 186306 331294
rect 186542 331058 221986 331294
rect 222222 331058 222306 331294
rect 222542 331058 257986 331294
rect 258222 331058 258306 331294
rect 258542 331058 293986 331294
rect 294222 331058 294306 331294
rect 294542 331058 329986 331294
rect 330222 331058 330306 331294
rect 330542 331058 365986 331294
rect 366222 331058 366306 331294
rect 366542 331058 401986 331294
rect 402222 331058 402306 331294
rect 402542 331058 437986 331294
rect 438222 331058 438306 331294
rect 438542 331058 473986 331294
rect 474222 331058 474306 331294
rect 474542 331058 509986 331294
rect 510222 331058 510306 331294
rect 510542 331058 581986 331294
rect 582222 331058 582306 331294
rect 582542 331058 589182 331294
rect 589418 331058 589502 331294
rect 589738 331058 592650 331294
rect -8726 331026 592650 331058
rect -8726 330374 592650 330406
rect -8726 330138 -4854 330374
rect -4618 330138 -4534 330374
rect -4298 330138 4746 330374
rect 4982 330138 5066 330374
rect 5302 330138 40746 330374
rect 40982 330138 41066 330374
rect 41302 330138 76746 330374
rect 76982 330138 77066 330374
rect 77302 330138 112746 330374
rect 112982 330138 113066 330374
rect 113302 330138 148746 330374
rect 148982 330138 149066 330374
rect 149302 330138 184746 330374
rect 184982 330138 185066 330374
rect 185302 330138 220746 330374
rect 220982 330138 221066 330374
rect 221302 330138 256746 330374
rect 256982 330138 257066 330374
rect 257302 330138 292746 330374
rect 292982 330138 293066 330374
rect 293302 330138 328746 330374
rect 328982 330138 329066 330374
rect 329302 330138 364746 330374
rect 364982 330138 365066 330374
rect 365302 330138 400746 330374
rect 400982 330138 401066 330374
rect 401302 330138 436746 330374
rect 436982 330138 437066 330374
rect 437302 330138 472746 330374
rect 472982 330138 473066 330374
rect 473302 330138 508746 330374
rect 508982 330138 509066 330374
rect 509302 330138 580746 330374
rect 580982 330138 581066 330374
rect 581302 330138 588222 330374
rect 588458 330138 588542 330374
rect 588778 330138 592650 330374
rect -8726 330054 592650 330138
rect -8726 329818 -4854 330054
rect -4618 329818 -4534 330054
rect -4298 329818 4746 330054
rect 4982 329818 5066 330054
rect 5302 329818 40746 330054
rect 40982 329818 41066 330054
rect 41302 329818 76746 330054
rect 76982 329818 77066 330054
rect 77302 329818 112746 330054
rect 112982 329818 113066 330054
rect 113302 329818 148746 330054
rect 148982 329818 149066 330054
rect 149302 329818 184746 330054
rect 184982 329818 185066 330054
rect 185302 329818 220746 330054
rect 220982 329818 221066 330054
rect 221302 329818 256746 330054
rect 256982 329818 257066 330054
rect 257302 329818 292746 330054
rect 292982 329818 293066 330054
rect 293302 329818 328746 330054
rect 328982 329818 329066 330054
rect 329302 329818 364746 330054
rect 364982 329818 365066 330054
rect 365302 329818 400746 330054
rect 400982 329818 401066 330054
rect 401302 329818 436746 330054
rect 436982 329818 437066 330054
rect 437302 329818 472746 330054
rect 472982 329818 473066 330054
rect 473302 329818 508746 330054
rect 508982 329818 509066 330054
rect 509302 329818 580746 330054
rect 580982 329818 581066 330054
rect 581302 329818 588222 330054
rect 588458 329818 588542 330054
rect 588778 329818 592650 330054
rect -8726 329786 592650 329818
rect -8726 329134 592650 329166
rect -8726 328898 -3894 329134
rect -3658 328898 -3574 329134
rect -3338 328898 3506 329134
rect 3742 328898 3826 329134
rect 4062 328898 39506 329134
rect 39742 328898 39826 329134
rect 40062 328898 75506 329134
rect 75742 328898 75826 329134
rect 76062 328898 111506 329134
rect 111742 328898 111826 329134
rect 112062 328898 147506 329134
rect 147742 328898 147826 329134
rect 148062 328898 183506 329134
rect 183742 328898 183826 329134
rect 184062 328898 219506 329134
rect 219742 328898 219826 329134
rect 220062 328898 255506 329134
rect 255742 328898 255826 329134
rect 256062 328898 291506 329134
rect 291742 328898 291826 329134
rect 292062 328898 327506 329134
rect 327742 328898 327826 329134
rect 328062 328898 363506 329134
rect 363742 328898 363826 329134
rect 364062 328898 399506 329134
rect 399742 328898 399826 329134
rect 400062 328898 435506 329134
rect 435742 328898 435826 329134
rect 436062 328898 471506 329134
rect 471742 328898 471826 329134
rect 472062 328898 507506 329134
rect 507742 328898 507826 329134
rect 508062 328898 579506 329134
rect 579742 328898 579826 329134
rect 580062 328898 587262 329134
rect 587498 328898 587582 329134
rect 587818 328898 592650 329134
rect -8726 328814 592650 328898
rect -8726 328578 -3894 328814
rect -3658 328578 -3574 328814
rect -3338 328578 3506 328814
rect 3742 328578 3826 328814
rect 4062 328578 39506 328814
rect 39742 328578 39826 328814
rect 40062 328578 75506 328814
rect 75742 328578 75826 328814
rect 76062 328578 111506 328814
rect 111742 328578 111826 328814
rect 112062 328578 147506 328814
rect 147742 328578 147826 328814
rect 148062 328578 183506 328814
rect 183742 328578 183826 328814
rect 184062 328578 219506 328814
rect 219742 328578 219826 328814
rect 220062 328578 255506 328814
rect 255742 328578 255826 328814
rect 256062 328578 291506 328814
rect 291742 328578 291826 328814
rect 292062 328578 327506 328814
rect 327742 328578 327826 328814
rect 328062 328578 363506 328814
rect 363742 328578 363826 328814
rect 364062 328578 399506 328814
rect 399742 328578 399826 328814
rect 400062 328578 435506 328814
rect 435742 328578 435826 328814
rect 436062 328578 471506 328814
rect 471742 328578 471826 328814
rect 472062 328578 507506 328814
rect 507742 328578 507826 328814
rect 508062 328578 579506 328814
rect 579742 328578 579826 328814
rect 580062 328578 587262 328814
rect 587498 328578 587582 328814
rect 587818 328578 592650 328814
rect -8726 328546 592650 328578
rect -8726 327894 592650 327926
rect -8726 327658 -2934 327894
rect -2698 327658 -2614 327894
rect -2378 327658 2266 327894
rect 2502 327658 2586 327894
rect 2822 327658 38266 327894
rect 38502 327658 38586 327894
rect 38822 327658 74266 327894
rect 74502 327658 74586 327894
rect 74822 327658 110266 327894
rect 110502 327658 110586 327894
rect 110822 327658 146266 327894
rect 146502 327658 146586 327894
rect 146822 327658 182266 327894
rect 182502 327658 182586 327894
rect 182822 327658 218266 327894
rect 218502 327658 218586 327894
rect 218822 327658 254266 327894
rect 254502 327658 254586 327894
rect 254822 327658 290266 327894
rect 290502 327658 290586 327894
rect 290822 327658 326266 327894
rect 326502 327658 326586 327894
rect 326822 327658 362266 327894
rect 362502 327658 362586 327894
rect 362822 327658 398266 327894
rect 398502 327658 398586 327894
rect 398822 327658 434266 327894
rect 434502 327658 434586 327894
rect 434822 327658 470266 327894
rect 470502 327658 470586 327894
rect 470822 327658 506266 327894
rect 506502 327658 506586 327894
rect 506822 327658 540918 327894
rect 541154 327658 542850 327894
rect 543086 327658 544782 327894
rect 545018 327658 546714 327894
rect 546950 327658 578266 327894
rect 578502 327658 578586 327894
rect 578822 327658 586302 327894
rect 586538 327658 586622 327894
rect 586858 327658 592650 327894
rect -8726 327574 592650 327658
rect -8726 327338 -2934 327574
rect -2698 327338 -2614 327574
rect -2378 327338 2266 327574
rect 2502 327338 2586 327574
rect 2822 327338 38266 327574
rect 38502 327338 38586 327574
rect 38822 327338 74266 327574
rect 74502 327338 74586 327574
rect 74822 327338 110266 327574
rect 110502 327338 110586 327574
rect 110822 327338 146266 327574
rect 146502 327338 146586 327574
rect 146822 327338 182266 327574
rect 182502 327338 182586 327574
rect 182822 327338 218266 327574
rect 218502 327338 218586 327574
rect 218822 327338 254266 327574
rect 254502 327338 254586 327574
rect 254822 327338 290266 327574
rect 290502 327338 290586 327574
rect 290822 327338 326266 327574
rect 326502 327338 326586 327574
rect 326822 327338 362266 327574
rect 362502 327338 362586 327574
rect 362822 327338 398266 327574
rect 398502 327338 398586 327574
rect 398822 327338 434266 327574
rect 434502 327338 434586 327574
rect 434822 327338 470266 327574
rect 470502 327338 470586 327574
rect 470822 327338 506266 327574
rect 506502 327338 506586 327574
rect 506822 327338 540918 327574
rect 541154 327338 542850 327574
rect 543086 327338 544782 327574
rect 545018 327338 546714 327574
rect 546950 327338 578266 327574
rect 578502 327338 578586 327574
rect 578822 327338 586302 327574
rect 586538 327338 586622 327574
rect 586858 327338 592650 327574
rect -8726 327306 592650 327338
rect -8726 326654 592650 326686
rect -8726 326418 -1974 326654
rect -1738 326418 -1654 326654
rect -1418 326418 1026 326654
rect 1262 326418 1346 326654
rect 1582 326418 37026 326654
rect 37262 326418 37346 326654
rect 37582 326418 73026 326654
rect 73262 326418 73346 326654
rect 73582 326418 109026 326654
rect 109262 326418 109346 326654
rect 109582 326418 145026 326654
rect 145262 326418 145346 326654
rect 145582 326418 181026 326654
rect 181262 326418 181346 326654
rect 181582 326418 217026 326654
rect 217262 326418 217346 326654
rect 217582 326418 253026 326654
rect 253262 326418 253346 326654
rect 253582 326418 289026 326654
rect 289262 326418 289346 326654
rect 289582 326418 325026 326654
rect 325262 326418 325346 326654
rect 325582 326418 361026 326654
rect 361262 326418 361346 326654
rect 361582 326418 397026 326654
rect 397262 326418 397346 326654
rect 397582 326418 433026 326654
rect 433262 326418 433346 326654
rect 433582 326418 469026 326654
rect 469262 326418 469346 326654
rect 469582 326418 505026 326654
rect 505262 326418 505346 326654
rect 505582 326418 539952 326654
rect 540188 326418 541884 326654
rect 542120 326418 543816 326654
rect 544052 326418 545748 326654
rect 545984 326418 577026 326654
rect 577262 326418 577346 326654
rect 577582 326418 585342 326654
rect 585578 326418 585662 326654
rect 585898 326418 592650 326654
rect -8726 326334 592650 326418
rect -8726 326098 -1974 326334
rect -1738 326098 -1654 326334
rect -1418 326098 1026 326334
rect 1262 326098 1346 326334
rect 1582 326098 37026 326334
rect 37262 326098 37346 326334
rect 37582 326098 73026 326334
rect 73262 326098 73346 326334
rect 73582 326098 109026 326334
rect 109262 326098 109346 326334
rect 109582 326098 145026 326334
rect 145262 326098 145346 326334
rect 145582 326098 181026 326334
rect 181262 326098 181346 326334
rect 181582 326098 217026 326334
rect 217262 326098 217346 326334
rect 217582 326098 253026 326334
rect 253262 326098 253346 326334
rect 253582 326098 289026 326334
rect 289262 326098 289346 326334
rect 289582 326098 325026 326334
rect 325262 326098 325346 326334
rect 325582 326098 361026 326334
rect 361262 326098 361346 326334
rect 361582 326098 397026 326334
rect 397262 326098 397346 326334
rect 397582 326098 433026 326334
rect 433262 326098 433346 326334
rect 433582 326098 469026 326334
rect 469262 326098 469346 326334
rect 469582 326098 505026 326334
rect 505262 326098 505346 326334
rect 505582 326098 539952 326334
rect 540188 326098 541884 326334
rect 542120 326098 543816 326334
rect 544052 326098 545748 326334
rect 545984 326098 577026 326334
rect 577262 326098 577346 326334
rect 577582 326098 585342 326334
rect 585578 326098 585662 326334
rect 585898 326098 592650 326334
rect -8726 326066 592650 326098
rect -8726 299334 592650 299366
rect -8726 299098 -8694 299334
rect -8458 299098 -8374 299334
rect -8138 299098 9706 299334
rect 9942 299098 10026 299334
rect 10262 299098 45706 299334
rect 45942 299098 46026 299334
rect 46262 299098 81706 299334
rect 81942 299098 82026 299334
rect 82262 299098 117706 299334
rect 117942 299098 118026 299334
rect 118262 299098 153706 299334
rect 153942 299098 154026 299334
rect 154262 299098 189706 299334
rect 189942 299098 190026 299334
rect 190262 299098 225706 299334
rect 225942 299098 226026 299334
rect 226262 299098 261706 299334
rect 261942 299098 262026 299334
rect 262262 299098 297706 299334
rect 297942 299098 298026 299334
rect 298262 299098 333706 299334
rect 333942 299098 334026 299334
rect 334262 299098 369706 299334
rect 369942 299098 370026 299334
rect 370262 299098 405706 299334
rect 405942 299098 406026 299334
rect 406262 299098 441706 299334
rect 441942 299098 442026 299334
rect 442262 299098 477706 299334
rect 477942 299098 478026 299334
rect 478262 299098 513706 299334
rect 513942 299098 514026 299334
rect 514262 299098 549706 299334
rect 549942 299098 550026 299334
rect 550262 299098 592062 299334
rect 592298 299098 592382 299334
rect 592618 299098 592650 299334
rect -8726 299014 592650 299098
rect -8726 298778 -8694 299014
rect -8458 298778 -8374 299014
rect -8138 298778 9706 299014
rect 9942 298778 10026 299014
rect 10262 298778 45706 299014
rect 45942 298778 46026 299014
rect 46262 298778 81706 299014
rect 81942 298778 82026 299014
rect 82262 298778 117706 299014
rect 117942 298778 118026 299014
rect 118262 298778 153706 299014
rect 153942 298778 154026 299014
rect 154262 298778 189706 299014
rect 189942 298778 190026 299014
rect 190262 298778 225706 299014
rect 225942 298778 226026 299014
rect 226262 298778 261706 299014
rect 261942 298778 262026 299014
rect 262262 298778 297706 299014
rect 297942 298778 298026 299014
rect 298262 298778 333706 299014
rect 333942 298778 334026 299014
rect 334262 298778 369706 299014
rect 369942 298778 370026 299014
rect 370262 298778 405706 299014
rect 405942 298778 406026 299014
rect 406262 298778 441706 299014
rect 441942 298778 442026 299014
rect 442262 298778 477706 299014
rect 477942 298778 478026 299014
rect 478262 298778 513706 299014
rect 513942 298778 514026 299014
rect 514262 298778 549706 299014
rect 549942 298778 550026 299014
rect 550262 298778 592062 299014
rect 592298 298778 592382 299014
rect 592618 298778 592650 299014
rect -8726 298746 592650 298778
rect -8726 298094 592650 298126
rect -8726 297858 -7734 298094
rect -7498 297858 -7414 298094
rect -7178 297858 8466 298094
rect 8702 297858 8786 298094
rect 9022 297858 44466 298094
rect 44702 297858 44786 298094
rect 45022 297858 80466 298094
rect 80702 297858 80786 298094
rect 81022 297858 116466 298094
rect 116702 297858 116786 298094
rect 117022 297858 152466 298094
rect 152702 297858 152786 298094
rect 153022 297858 188466 298094
rect 188702 297858 188786 298094
rect 189022 297858 224466 298094
rect 224702 297858 224786 298094
rect 225022 297858 260466 298094
rect 260702 297858 260786 298094
rect 261022 297858 296466 298094
rect 296702 297858 296786 298094
rect 297022 297858 332466 298094
rect 332702 297858 332786 298094
rect 333022 297858 368466 298094
rect 368702 297858 368786 298094
rect 369022 297858 404466 298094
rect 404702 297858 404786 298094
rect 405022 297858 440466 298094
rect 440702 297858 440786 298094
rect 441022 297858 476466 298094
rect 476702 297858 476786 298094
rect 477022 297858 512466 298094
rect 512702 297858 512786 298094
rect 513022 297858 548466 298094
rect 548702 297858 548786 298094
rect 549022 297858 591102 298094
rect 591338 297858 591422 298094
rect 591658 297858 592650 298094
rect -8726 297774 592650 297858
rect -8726 297538 -7734 297774
rect -7498 297538 -7414 297774
rect -7178 297538 8466 297774
rect 8702 297538 8786 297774
rect 9022 297538 44466 297774
rect 44702 297538 44786 297774
rect 45022 297538 80466 297774
rect 80702 297538 80786 297774
rect 81022 297538 116466 297774
rect 116702 297538 116786 297774
rect 117022 297538 152466 297774
rect 152702 297538 152786 297774
rect 153022 297538 188466 297774
rect 188702 297538 188786 297774
rect 189022 297538 224466 297774
rect 224702 297538 224786 297774
rect 225022 297538 260466 297774
rect 260702 297538 260786 297774
rect 261022 297538 296466 297774
rect 296702 297538 296786 297774
rect 297022 297538 332466 297774
rect 332702 297538 332786 297774
rect 333022 297538 368466 297774
rect 368702 297538 368786 297774
rect 369022 297538 404466 297774
rect 404702 297538 404786 297774
rect 405022 297538 440466 297774
rect 440702 297538 440786 297774
rect 441022 297538 476466 297774
rect 476702 297538 476786 297774
rect 477022 297538 512466 297774
rect 512702 297538 512786 297774
rect 513022 297538 548466 297774
rect 548702 297538 548786 297774
rect 549022 297538 591102 297774
rect 591338 297538 591422 297774
rect 591658 297538 592650 297774
rect -8726 297506 592650 297538
rect -8726 296854 592650 296886
rect -8726 296618 -6774 296854
rect -6538 296618 -6454 296854
rect -6218 296618 7226 296854
rect 7462 296618 7546 296854
rect 7782 296618 43226 296854
rect 43462 296618 43546 296854
rect 43782 296618 79226 296854
rect 79462 296618 79546 296854
rect 79782 296618 115226 296854
rect 115462 296618 115546 296854
rect 115782 296618 151226 296854
rect 151462 296618 151546 296854
rect 151782 296618 187226 296854
rect 187462 296618 187546 296854
rect 187782 296618 223226 296854
rect 223462 296618 223546 296854
rect 223782 296618 259226 296854
rect 259462 296618 259546 296854
rect 259782 296618 295226 296854
rect 295462 296618 295546 296854
rect 295782 296618 331226 296854
rect 331462 296618 331546 296854
rect 331782 296618 367226 296854
rect 367462 296618 367546 296854
rect 367782 296618 403226 296854
rect 403462 296618 403546 296854
rect 403782 296618 439226 296854
rect 439462 296618 439546 296854
rect 439782 296618 475226 296854
rect 475462 296618 475546 296854
rect 475782 296618 511226 296854
rect 511462 296618 511546 296854
rect 511782 296618 547226 296854
rect 547462 296618 547546 296854
rect 547782 296618 590142 296854
rect 590378 296618 590462 296854
rect 590698 296618 592650 296854
rect -8726 296534 592650 296618
rect -8726 296298 -6774 296534
rect -6538 296298 -6454 296534
rect -6218 296298 7226 296534
rect 7462 296298 7546 296534
rect 7782 296298 43226 296534
rect 43462 296298 43546 296534
rect 43782 296298 79226 296534
rect 79462 296298 79546 296534
rect 79782 296298 115226 296534
rect 115462 296298 115546 296534
rect 115782 296298 151226 296534
rect 151462 296298 151546 296534
rect 151782 296298 187226 296534
rect 187462 296298 187546 296534
rect 187782 296298 223226 296534
rect 223462 296298 223546 296534
rect 223782 296298 259226 296534
rect 259462 296298 259546 296534
rect 259782 296298 295226 296534
rect 295462 296298 295546 296534
rect 295782 296298 331226 296534
rect 331462 296298 331546 296534
rect 331782 296298 367226 296534
rect 367462 296298 367546 296534
rect 367782 296298 403226 296534
rect 403462 296298 403546 296534
rect 403782 296298 439226 296534
rect 439462 296298 439546 296534
rect 439782 296298 475226 296534
rect 475462 296298 475546 296534
rect 475782 296298 511226 296534
rect 511462 296298 511546 296534
rect 511782 296298 547226 296534
rect 547462 296298 547546 296534
rect 547782 296298 590142 296534
rect 590378 296298 590462 296534
rect 590698 296298 592650 296534
rect -8726 296266 592650 296298
rect -8726 295614 592650 295646
rect -8726 295378 -5814 295614
rect -5578 295378 -5494 295614
rect -5258 295378 5986 295614
rect 6222 295378 6306 295614
rect 6542 295378 41986 295614
rect 42222 295378 42306 295614
rect 42542 295378 77986 295614
rect 78222 295378 78306 295614
rect 78542 295378 113986 295614
rect 114222 295378 114306 295614
rect 114542 295378 149986 295614
rect 150222 295378 150306 295614
rect 150542 295378 185986 295614
rect 186222 295378 186306 295614
rect 186542 295378 221986 295614
rect 222222 295378 222306 295614
rect 222542 295378 257986 295614
rect 258222 295378 258306 295614
rect 258542 295378 293986 295614
rect 294222 295378 294306 295614
rect 294542 295378 329986 295614
rect 330222 295378 330306 295614
rect 330542 295378 365986 295614
rect 366222 295378 366306 295614
rect 366542 295378 401986 295614
rect 402222 295378 402306 295614
rect 402542 295378 437986 295614
rect 438222 295378 438306 295614
rect 438542 295378 473986 295614
rect 474222 295378 474306 295614
rect 474542 295378 509986 295614
rect 510222 295378 510306 295614
rect 510542 295378 581986 295614
rect 582222 295378 582306 295614
rect 582542 295378 589182 295614
rect 589418 295378 589502 295614
rect 589738 295378 592650 295614
rect -8726 295294 592650 295378
rect -8726 295058 -5814 295294
rect -5578 295058 -5494 295294
rect -5258 295058 5986 295294
rect 6222 295058 6306 295294
rect 6542 295058 41986 295294
rect 42222 295058 42306 295294
rect 42542 295058 77986 295294
rect 78222 295058 78306 295294
rect 78542 295058 113986 295294
rect 114222 295058 114306 295294
rect 114542 295058 149986 295294
rect 150222 295058 150306 295294
rect 150542 295058 185986 295294
rect 186222 295058 186306 295294
rect 186542 295058 221986 295294
rect 222222 295058 222306 295294
rect 222542 295058 257986 295294
rect 258222 295058 258306 295294
rect 258542 295058 293986 295294
rect 294222 295058 294306 295294
rect 294542 295058 329986 295294
rect 330222 295058 330306 295294
rect 330542 295058 365986 295294
rect 366222 295058 366306 295294
rect 366542 295058 401986 295294
rect 402222 295058 402306 295294
rect 402542 295058 437986 295294
rect 438222 295058 438306 295294
rect 438542 295058 473986 295294
rect 474222 295058 474306 295294
rect 474542 295058 509986 295294
rect 510222 295058 510306 295294
rect 510542 295058 581986 295294
rect 582222 295058 582306 295294
rect 582542 295058 589182 295294
rect 589418 295058 589502 295294
rect 589738 295058 592650 295294
rect -8726 295026 592650 295058
rect -8726 294374 592650 294406
rect -8726 294138 -4854 294374
rect -4618 294138 -4534 294374
rect -4298 294138 4746 294374
rect 4982 294138 5066 294374
rect 5302 294138 40746 294374
rect 40982 294138 41066 294374
rect 41302 294138 76746 294374
rect 76982 294138 77066 294374
rect 77302 294138 112746 294374
rect 112982 294138 113066 294374
rect 113302 294138 148746 294374
rect 148982 294138 149066 294374
rect 149302 294138 184746 294374
rect 184982 294138 185066 294374
rect 185302 294138 220746 294374
rect 220982 294138 221066 294374
rect 221302 294138 256746 294374
rect 256982 294138 257066 294374
rect 257302 294138 292746 294374
rect 292982 294138 293066 294374
rect 293302 294138 328746 294374
rect 328982 294138 329066 294374
rect 329302 294138 364746 294374
rect 364982 294138 365066 294374
rect 365302 294138 400746 294374
rect 400982 294138 401066 294374
rect 401302 294138 436746 294374
rect 436982 294138 437066 294374
rect 437302 294138 472746 294374
rect 472982 294138 473066 294374
rect 473302 294138 508746 294374
rect 508982 294138 509066 294374
rect 509302 294138 580746 294374
rect 580982 294138 581066 294374
rect 581302 294138 588222 294374
rect 588458 294138 588542 294374
rect 588778 294138 592650 294374
rect -8726 294054 592650 294138
rect -8726 293818 -4854 294054
rect -4618 293818 -4534 294054
rect -4298 293818 4746 294054
rect 4982 293818 5066 294054
rect 5302 293818 40746 294054
rect 40982 293818 41066 294054
rect 41302 293818 76746 294054
rect 76982 293818 77066 294054
rect 77302 293818 112746 294054
rect 112982 293818 113066 294054
rect 113302 293818 148746 294054
rect 148982 293818 149066 294054
rect 149302 293818 184746 294054
rect 184982 293818 185066 294054
rect 185302 293818 220746 294054
rect 220982 293818 221066 294054
rect 221302 293818 256746 294054
rect 256982 293818 257066 294054
rect 257302 293818 292746 294054
rect 292982 293818 293066 294054
rect 293302 293818 328746 294054
rect 328982 293818 329066 294054
rect 329302 293818 364746 294054
rect 364982 293818 365066 294054
rect 365302 293818 400746 294054
rect 400982 293818 401066 294054
rect 401302 293818 436746 294054
rect 436982 293818 437066 294054
rect 437302 293818 472746 294054
rect 472982 293818 473066 294054
rect 473302 293818 508746 294054
rect 508982 293818 509066 294054
rect 509302 293818 580746 294054
rect 580982 293818 581066 294054
rect 581302 293818 588222 294054
rect 588458 293818 588542 294054
rect 588778 293818 592650 294054
rect -8726 293786 592650 293818
rect -8726 293134 592650 293166
rect -8726 292898 -3894 293134
rect -3658 292898 -3574 293134
rect -3338 292898 3506 293134
rect 3742 292898 3826 293134
rect 4062 292898 39506 293134
rect 39742 292898 39826 293134
rect 40062 292898 75506 293134
rect 75742 292898 75826 293134
rect 76062 292898 111506 293134
rect 111742 292898 111826 293134
rect 112062 292898 147506 293134
rect 147742 292898 147826 293134
rect 148062 292898 183506 293134
rect 183742 292898 183826 293134
rect 184062 292898 219506 293134
rect 219742 292898 219826 293134
rect 220062 292898 255506 293134
rect 255742 292898 255826 293134
rect 256062 292898 291506 293134
rect 291742 292898 291826 293134
rect 292062 292898 327506 293134
rect 327742 292898 327826 293134
rect 328062 292898 363506 293134
rect 363742 292898 363826 293134
rect 364062 292898 399506 293134
rect 399742 292898 399826 293134
rect 400062 292898 435506 293134
rect 435742 292898 435826 293134
rect 436062 292898 471506 293134
rect 471742 292898 471826 293134
rect 472062 292898 507506 293134
rect 507742 292898 507826 293134
rect 508062 292898 579506 293134
rect 579742 292898 579826 293134
rect 580062 292898 587262 293134
rect 587498 292898 587582 293134
rect 587818 292898 592650 293134
rect -8726 292814 592650 292898
rect -8726 292578 -3894 292814
rect -3658 292578 -3574 292814
rect -3338 292578 3506 292814
rect 3742 292578 3826 292814
rect 4062 292578 39506 292814
rect 39742 292578 39826 292814
rect 40062 292578 75506 292814
rect 75742 292578 75826 292814
rect 76062 292578 111506 292814
rect 111742 292578 111826 292814
rect 112062 292578 147506 292814
rect 147742 292578 147826 292814
rect 148062 292578 183506 292814
rect 183742 292578 183826 292814
rect 184062 292578 219506 292814
rect 219742 292578 219826 292814
rect 220062 292578 255506 292814
rect 255742 292578 255826 292814
rect 256062 292578 291506 292814
rect 291742 292578 291826 292814
rect 292062 292578 327506 292814
rect 327742 292578 327826 292814
rect 328062 292578 363506 292814
rect 363742 292578 363826 292814
rect 364062 292578 399506 292814
rect 399742 292578 399826 292814
rect 400062 292578 435506 292814
rect 435742 292578 435826 292814
rect 436062 292578 471506 292814
rect 471742 292578 471826 292814
rect 472062 292578 507506 292814
rect 507742 292578 507826 292814
rect 508062 292578 579506 292814
rect 579742 292578 579826 292814
rect 580062 292578 587262 292814
rect 587498 292578 587582 292814
rect 587818 292578 592650 292814
rect -8726 292546 592650 292578
rect -8726 291894 592650 291926
rect -8726 291658 -2934 291894
rect -2698 291658 -2614 291894
rect -2378 291658 2266 291894
rect 2502 291658 2586 291894
rect 2822 291658 38266 291894
rect 38502 291658 38586 291894
rect 38822 291658 74266 291894
rect 74502 291658 74586 291894
rect 74822 291658 110266 291894
rect 110502 291658 110586 291894
rect 110822 291658 146266 291894
rect 146502 291658 146586 291894
rect 146822 291658 182266 291894
rect 182502 291658 182586 291894
rect 182822 291658 218266 291894
rect 218502 291658 218586 291894
rect 218822 291658 254266 291894
rect 254502 291658 254586 291894
rect 254822 291658 290266 291894
rect 290502 291658 290586 291894
rect 290822 291658 326266 291894
rect 326502 291658 326586 291894
rect 326822 291658 362266 291894
rect 362502 291658 362586 291894
rect 362822 291658 398266 291894
rect 398502 291658 398586 291894
rect 398822 291658 434266 291894
rect 434502 291658 434586 291894
rect 434822 291658 470266 291894
rect 470502 291658 470586 291894
rect 470822 291658 506266 291894
rect 506502 291658 506586 291894
rect 506822 291658 540918 291894
rect 541154 291658 542850 291894
rect 543086 291658 544782 291894
rect 545018 291658 546714 291894
rect 546950 291658 578266 291894
rect 578502 291658 578586 291894
rect 578822 291658 586302 291894
rect 586538 291658 586622 291894
rect 586858 291658 592650 291894
rect -8726 291574 592650 291658
rect -8726 291338 -2934 291574
rect -2698 291338 -2614 291574
rect -2378 291338 2266 291574
rect 2502 291338 2586 291574
rect 2822 291338 38266 291574
rect 38502 291338 38586 291574
rect 38822 291338 74266 291574
rect 74502 291338 74586 291574
rect 74822 291338 110266 291574
rect 110502 291338 110586 291574
rect 110822 291338 146266 291574
rect 146502 291338 146586 291574
rect 146822 291338 182266 291574
rect 182502 291338 182586 291574
rect 182822 291338 218266 291574
rect 218502 291338 218586 291574
rect 218822 291338 254266 291574
rect 254502 291338 254586 291574
rect 254822 291338 290266 291574
rect 290502 291338 290586 291574
rect 290822 291338 326266 291574
rect 326502 291338 326586 291574
rect 326822 291338 362266 291574
rect 362502 291338 362586 291574
rect 362822 291338 398266 291574
rect 398502 291338 398586 291574
rect 398822 291338 434266 291574
rect 434502 291338 434586 291574
rect 434822 291338 470266 291574
rect 470502 291338 470586 291574
rect 470822 291338 506266 291574
rect 506502 291338 506586 291574
rect 506822 291338 540918 291574
rect 541154 291338 542850 291574
rect 543086 291338 544782 291574
rect 545018 291338 546714 291574
rect 546950 291338 578266 291574
rect 578502 291338 578586 291574
rect 578822 291338 586302 291574
rect 586538 291338 586622 291574
rect 586858 291338 592650 291574
rect -8726 291306 592650 291338
rect -8726 290654 592650 290686
rect -8726 290418 -1974 290654
rect -1738 290418 -1654 290654
rect -1418 290418 1026 290654
rect 1262 290418 1346 290654
rect 1582 290418 37026 290654
rect 37262 290418 37346 290654
rect 37582 290418 73026 290654
rect 73262 290418 73346 290654
rect 73582 290418 109026 290654
rect 109262 290418 109346 290654
rect 109582 290418 145026 290654
rect 145262 290418 145346 290654
rect 145582 290418 181026 290654
rect 181262 290418 181346 290654
rect 181582 290418 217026 290654
rect 217262 290418 217346 290654
rect 217582 290418 253026 290654
rect 253262 290418 253346 290654
rect 253582 290418 289026 290654
rect 289262 290418 289346 290654
rect 289582 290418 325026 290654
rect 325262 290418 325346 290654
rect 325582 290418 361026 290654
rect 361262 290418 361346 290654
rect 361582 290418 397026 290654
rect 397262 290418 397346 290654
rect 397582 290418 433026 290654
rect 433262 290418 433346 290654
rect 433582 290418 469026 290654
rect 469262 290418 469346 290654
rect 469582 290418 505026 290654
rect 505262 290418 505346 290654
rect 505582 290418 539952 290654
rect 540188 290418 541884 290654
rect 542120 290418 543816 290654
rect 544052 290418 545748 290654
rect 545984 290418 577026 290654
rect 577262 290418 577346 290654
rect 577582 290418 585342 290654
rect 585578 290418 585662 290654
rect 585898 290418 592650 290654
rect -8726 290334 592650 290418
rect -8726 290098 -1974 290334
rect -1738 290098 -1654 290334
rect -1418 290098 1026 290334
rect 1262 290098 1346 290334
rect 1582 290098 37026 290334
rect 37262 290098 37346 290334
rect 37582 290098 73026 290334
rect 73262 290098 73346 290334
rect 73582 290098 109026 290334
rect 109262 290098 109346 290334
rect 109582 290098 145026 290334
rect 145262 290098 145346 290334
rect 145582 290098 181026 290334
rect 181262 290098 181346 290334
rect 181582 290098 217026 290334
rect 217262 290098 217346 290334
rect 217582 290098 253026 290334
rect 253262 290098 253346 290334
rect 253582 290098 289026 290334
rect 289262 290098 289346 290334
rect 289582 290098 325026 290334
rect 325262 290098 325346 290334
rect 325582 290098 361026 290334
rect 361262 290098 361346 290334
rect 361582 290098 397026 290334
rect 397262 290098 397346 290334
rect 397582 290098 433026 290334
rect 433262 290098 433346 290334
rect 433582 290098 469026 290334
rect 469262 290098 469346 290334
rect 469582 290098 505026 290334
rect 505262 290098 505346 290334
rect 505582 290098 539952 290334
rect 540188 290098 541884 290334
rect 542120 290098 543816 290334
rect 544052 290098 545748 290334
rect 545984 290098 577026 290334
rect 577262 290098 577346 290334
rect 577582 290098 585342 290334
rect 585578 290098 585662 290334
rect 585898 290098 592650 290334
rect -8726 290066 592650 290098
rect -8726 263334 592650 263366
rect -8726 263098 -8694 263334
rect -8458 263098 -8374 263334
rect -8138 263098 9706 263334
rect 9942 263098 10026 263334
rect 10262 263098 45706 263334
rect 45942 263098 46026 263334
rect 46262 263098 81706 263334
rect 81942 263098 82026 263334
rect 82262 263098 117706 263334
rect 117942 263098 118026 263334
rect 118262 263098 153706 263334
rect 153942 263098 154026 263334
rect 154262 263098 189706 263334
rect 189942 263098 190026 263334
rect 190262 263098 225706 263334
rect 225942 263098 226026 263334
rect 226262 263098 261706 263334
rect 261942 263098 262026 263334
rect 262262 263098 297706 263334
rect 297942 263098 298026 263334
rect 298262 263098 333706 263334
rect 333942 263098 334026 263334
rect 334262 263098 369706 263334
rect 369942 263098 370026 263334
rect 370262 263098 405706 263334
rect 405942 263098 406026 263334
rect 406262 263098 441706 263334
rect 441942 263098 442026 263334
rect 442262 263098 477706 263334
rect 477942 263098 478026 263334
rect 478262 263098 513706 263334
rect 513942 263098 514026 263334
rect 514262 263098 549706 263334
rect 549942 263098 550026 263334
rect 550262 263098 592062 263334
rect 592298 263098 592382 263334
rect 592618 263098 592650 263334
rect -8726 263014 592650 263098
rect -8726 262778 -8694 263014
rect -8458 262778 -8374 263014
rect -8138 262778 9706 263014
rect 9942 262778 10026 263014
rect 10262 262778 45706 263014
rect 45942 262778 46026 263014
rect 46262 262778 81706 263014
rect 81942 262778 82026 263014
rect 82262 262778 117706 263014
rect 117942 262778 118026 263014
rect 118262 262778 153706 263014
rect 153942 262778 154026 263014
rect 154262 262778 189706 263014
rect 189942 262778 190026 263014
rect 190262 262778 225706 263014
rect 225942 262778 226026 263014
rect 226262 262778 261706 263014
rect 261942 262778 262026 263014
rect 262262 262778 297706 263014
rect 297942 262778 298026 263014
rect 298262 262778 333706 263014
rect 333942 262778 334026 263014
rect 334262 262778 369706 263014
rect 369942 262778 370026 263014
rect 370262 262778 405706 263014
rect 405942 262778 406026 263014
rect 406262 262778 441706 263014
rect 441942 262778 442026 263014
rect 442262 262778 477706 263014
rect 477942 262778 478026 263014
rect 478262 262778 513706 263014
rect 513942 262778 514026 263014
rect 514262 262778 549706 263014
rect 549942 262778 550026 263014
rect 550262 262778 592062 263014
rect 592298 262778 592382 263014
rect 592618 262778 592650 263014
rect -8726 262746 592650 262778
rect -8726 262094 592650 262126
rect -8726 261858 -7734 262094
rect -7498 261858 -7414 262094
rect -7178 261858 8466 262094
rect 8702 261858 8786 262094
rect 9022 261858 44466 262094
rect 44702 261858 44786 262094
rect 45022 261858 80466 262094
rect 80702 261858 80786 262094
rect 81022 261858 116466 262094
rect 116702 261858 116786 262094
rect 117022 261858 152466 262094
rect 152702 261858 152786 262094
rect 153022 261858 188466 262094
rect 188702 261858 188786 262094
rect 189022 261858 224466 262094
rect 224702 261858 224786 262094
rect 225022 261858 260466 262094
rect 260702 261858 260786 262094
rect 261022 261858 296466 262094
rect 296702 261858 296786 262094
rect 297022 261858 332466 262094
rect 332702 261858 332786 262094
rect 333022 261858 368466 262094
rect 368702 261858 368786 262094
rect 369022 261858 404466 262094
rect 404702 261858 404786 262094
rect 405022 261858 440466 262094
rect 440702 261858 440786 262094
rect 441022 261858 476466 262094
rect 476702 261858 476786 262094
rect 477022 261858 512466 262094
rect 512702 261858 512786 262094
rect 513022 261858 548466 262094
rect 548702 261858 548786 262094
rect 549022 261858 591102 262094
rect 591338 261858 591422 262094
rect 591658 261858 592650 262094
rect -8726 261774 592650 261858
rect -8726 261538 -7734 261774
rect -7498 261538 -7414 261774
rect -7178 261538 8466 261774
rect 8702 261538 8786 261774
rect 9022 261538 44466 261774
rect 44702 261538 44786 261774
rect 45022 261538 80466 261774
rect 80702 261538 80786 261774
rect 81022 261538 116466 261774
rect 116702 261538 116786 261774
rect 117022 261538 152466 261774
rect 152702 261538 152786 261774
rect 153022 261538 188466 261774
rect 188702 261538 188786 261774
rect 189022 261538 224466 261774
rect 224702 261538 224786 261774
rect 225022 261538 260466 261774
rect 260702 261538 260786 261774
rect 261022 261538 296466 261774
rect 296702 261538 296786 261774
rect 297022 261538 332466 261774
rect 332702 261538 332786 261774
rect 333022 261538 368466 261774
rect 368702 261538 368786 261774
rect 369022 261538 404466 261774
rect 404702 261538 404786 261774
rect 405022 261538 440466 261774
rect 440702 261538 440786 261774
rect 441022 261538 476466 261774
rect 476702 261538 476786 261774
rect 477022 261538 512466 261774
rect 512702 261538 512786 261774
rect 513022 261538 548466 261774
rect 548702 261538 548786 261774
rect 549022 261538 591102 261774
rect 591338 261538 591422 261774
rect 591658 261538 592650 261774
rect -8726 261506 592650 261538
rect -8726 260854 592650 260886
rect -8726 260618 -6774 260854
rect -6538 260618 -6454 260854
rect -6218 260618 7226 260854
rect 7462 260618 7546 260854
rect 7782 260618 43226 260854
rect 43462 260618 43546 260854
rect 43782 260618 79226 260854
rect 79462 260618 79546 260854
rect 79782 260618 115226 260854
rect 115462 260618 115546 260854
rect 115782 260618 151226 260854
rect 151462 260618 151546 260854
rect 151782 260618 187226 260854
rect 187462 260618 187546 260854
rect 187782 260618 223226 260854
rect 223462 260618 223546 260854
rect 223782 260618 259226 260854
rect 259462 260618 259546 260854
rect 259782 260618 295226 260854
rect 295462 260618 295546 260854
rect 295782 260618 331226 260854
rect 331462 260618 331546 260854
rect 331782 260618 367226 260854
rect 367462 260618 367546 260854
rect 367782 260618 403226 260854
rect 403462 260618 403546 260854
rect 403782 260618 439226 260854
rect 439462 260618 439546 260854
rect 439782 260618 475226 260854
rect 475462 260618 475546 260854
rect 475782 260618 511226 260854
rect 511462 260618 511546 260854
rect 511782 260618 547226 260854
rect 547462 260618 547546 260854
rect 547782 260618 590142 260854
rect 590378 260618 590462 260854
rect 590698 260618 592650 260854
rect -8726 260534 592650 260618
rect -8726 260298 -6774 260534
rect -6538 260298 -6454 260534
rect -6218 260298 7226 260534
rect 7462 260298 7546 260534
rect 7782 260298 43226 260534
rect 43462 260298 43546 260534
rect 43782 260298 79226 260534
rect 79462 260298 79546 260534
rect 79782 260298 115226 260534
rect 115462 260298 115546 260534
rect 115782 260298 151226 260534
rect 151462 260298 151546 260534
rect 151782 260298 187226 260534
rect 187462 260298 187546 260534
rect 187782 260298 223226 260534
rect 223462 260298 223546 260534
rect 223782 260298 259226 260534
rect 259462 260298 259546 260534
rect 259782 260298 295226 260534
rect 295462 260298 295546 260534
rect 295782 260298 331226 260534
rect 331462 260298 331546 260534
rect 331782 260298 367226 260534
rect 367462 260298 367546 260534
rect 367782 260298 403226 260534
rect 403462 260298 403546 260534
rect 403782 260298 439226 260534
rect 439462 260298 439546 260534
rect 439782 260298 475226 260534
rect 475462 260298 475546 260534
rect 475782 260298 511226 260534
rect 511462 260298 511546 260534
rect 511782 260298 547226 260534
rect 547462 260298 547546 260534
rect 547782 260298 590142 260534
rect 590378 260298 590462 260534
rect 590698 260298 592650 260534
rect -8726 260266 592650 260298
rect -8726 259614 592650 259646
rect -8726 259378 -5814 259614
rect -5578 259378 -5494 259614
rect -5258 259378 5986 259614
rect 6222 259378 6306 259614
rect 6542 259378 41986 259614
rect 42222 259378 42306 259614
rect 42542 259378 77986 259614
rect 78222 259378 78306 259614
rect 78542 259378 113986 259614
rect 114222 259378 114306 259614
rect 114542 259378 149986 259614
rect 150222 259378 150306 259614
rect 150542 259378 185986 259614
rect 186222 259378 186306 259614
rect 186542 259378 221986 259614
rect 222222 259378 222306 259614
rect 222542 259378 257986 259614
rect 258222 259378 258306 259614
rect 258542 259378 293986 259614
rect 294222 259378 294306 259614
rect 294542 259378 329986 259614
rect 330222 259378 330306 259614
rect 330542 259378 365986 259614
rect 366222 259378 366306 259614
rect 366542 259378 401986 259614
rect 402222 259378 402306 259614
rect 402542 259378 437986 259614
rect 438222 259378 438306 259614
rect 438542 259378 473986 259614
rect 474222 259378 474306 259614
rect 474542 259378 509986 259614
rect 510222 259378 510306 259614
rect 510542 259378 545986 259614
rect 546222 259378 546306 259614
rect 546542 259378 581986 259614
rect 582222 259378 582306 259614
rect 582542 259378 589182 259614
rect 589418 259378 589502 259614
rect 589738 259378 592650 259614
rect -8726 259294 592650 259378
rect -8726 259058 -5814 259294
rect -5578 259058 -5494 259294
rect -5258 259058 5986 259294
rect 6222 259058 6306 259294
rect 6542 259058 41986 259294
rect 42222 259058 42306 259294
rect 42542 259058 77986 259294
rect 78222 259058 78306 259294
rect 78542 259058 113986 259294
rect 114222 259058 114306 259294
rect 114542 259058 149986 259294
rect 150222 259058 150306 259294
rect 150542 259058 185986 259294
rect 186222 259058 186306 259294
rect 186542 259058 221986 259294
rect 222222 259058 222306 259294
rect 222542 259058 257986 259294
rect 258222 259058 258306 259294
rect 258542 259058 293986 259294
rect 294222 259058 294306 259294
rect 294542 259058 329986 259294
rect 330222 259058 330306 259294
rect 330542 259058 365986 259294
rect 366222 259058 366306 259294
rect 366542 259058 401986 259294
rect 402222 259058 402306 259294
rect 402542 259058 437986 259294
rect 438222 259058 438306 259294
rect 438542 259058 473986 259294
rect 474222 259058 474306 259294
rect 474542 259058 509986 259294
rect 510222 259058 510306 259294
rect 510542 259058 545986 259294
rect 546222 259058 546306 259294
rect 546542 259058 581986 259294
rect 582222 259058 582306 259294
rect 582542 259058 589182 259294
rect 589418 259058 589502 259294
rect 589738 259058 592650 259294
rect -8726 259026 592650 259058
rect -8726 258374 592650 258406
rect -8726 258138 -4854 258374
rect -4618 258138 -4534 258374
rect -4298 258138 4746 258374
rect 4982 258138 5066 258374
rect 5302 258138 40746 258374
rect 40982 258138 41066 258374
rect 41302 258138 76746 258374
rect 76982 258138 77066 258374
rect 77302 258138 112746 258374
rect 112982 258138 113066 258374
rect 113302 258138 148746 258374
rect 148982 258138 149066 258374
rect 149302 258138 184746 258374
rect 184982 258138 185066 258374
rect 185302 258138 220746 258374
rect 220982 258138 221066 258374
rect 221302 258138 256746 258374
rect 256982 258138 257066 258374
rect 257302 258138 292746 258374
rect 292982 258138 293066 258374
rect 293302 258138 328746 258374
rect 328982 258138 329066 258374
rect 329302 258138 364746 258374
rect 364982 258138 365066 258374
rect 365302 258138 400746 258374
rect 400982 258138 401066 258374
rect 401302 258138 436746 258374
rect 436982 258138 437066 258374
rect 437302 258138 472746 258374
rect 472982 258138 473066 258374
rect 473302 258138 508746 258374
rect 508982 258138 509066 258374
rect 509302 258138 544746 258374
rect 544982 258138 545066 258374
rect 545302 258138 580746 258374
rect 580982 258138 581066 258374
rect 581302 258138 588222 258374
rect 588458 258138 588542 258374
rect 588778 258138 592650 258374
rect -8726 258054 592650 258138
rect -8726 257818 -4854 258054
rect -4618 257818 -4534 258054
rect -4298 257818 4746 258054
rect 4982 257818 5066 258054
rect 5302 257818 40746 258054
rect 40982 257818 41066 258054
rect 41302 257818 76746 258054
rect 76982 257818 77066 258054
rect 77302 257818 112746 258054
rect 112982 257818 113066 258054
rect 113302 257818 148746 258054
rect 148982 257818 149066 258054
rect 149302 257818 184746 258054
rect 184982 257818 185066 258054
rect 185302 257818 220746 258054
rect 220982 257818 221066 258054
rect 221302 257818 256746 258054
rect 256982 257818 257066 258054
rect 257302 257818 292746 258054
rect 292982 257818 293066 258054
rect 293302 257818 328746 258054
rect 328982 257818 329066 258054
rect 329302 257818 364746 258054
rect 364982 257818 365066 258054
rect 365302 257818 400746 258054
rect 400982 257818 401066 258054
rect 401302 257818 436746 258054
rect 436982 257818 437066 258054
rect 437302 257818 472746 258054
rect 472982 257818 473066 258054
rect 473302 257818 508746 258054
rect 508982 257818 509066 258054
rect 509302 257818 544746 258054
rect 544982 257818 545066 258054
rect 545302 257818 580746 258054
rect 580982 257818 581066 258054
rect 581302 257818 588222 258054
rect 588458 257818 588542 258054
rect 588778 257818 592650 258054
rect -8726 257786 592650 257818
rect -8726 257134 592650 257166
rect -8726 256898 -3894 257134
rect -3658 256898 -3574 257134
rect -3338 256898 3506 257134
rect 3742 256898 3826 257134
rect 4062 256898 39506 257134
rect 39742 256898 39826 257134
rect 40062 256898 75506 257134
rect 75742 256898 75826 257134
rect 76062 256898 111506 257134
rect 111742 256898 111826 257134
rect 112062 256898 147506 257134
rect 147742 256898 147826 257134
rect 148062 256898 183506 257134
rect 183742 256898 183826 257134
rect 184062 256898 219506 257134
rect 219742 256898 219826 257134
rect 220062 256898 255506 257134
rect 255742 256898 255826 257134
rect 256062 256898 291506 257134
rect 291742 256898 291826 257134
rect 292062 256898 327506 257134
rect 327742 256898 327826 257134
rect 328062 256898 363506 257134
rect 363742 256898 363826 257134
rect 364062 256898 399506 257134
rect 399742 256898 399826 257134
rect 400062 256898 435506 257134
rect 435742 256898 435826 257134
rect 436062 256898 471506 257134
rect 471742 256898 471826 257134
rect 472062 256898 507506 257134
rect 507742 256898 507826 257134
rect 508062 256898 543506 257134
rect 543742 256898 543826 257134
rect 544062 256898 579506 257134
rect 579742 256898 579826 257134
rect 580062 256898 587262 257134
rect 587498 256898 587582 257134
rect 587818 256898 592650 257134
rect -8726 256814 592650 256898
rect -8726 256578 -3894 256814
rect -3658 256578 -3574 256814
rect -3338 256578 3506 256814
rect 3742 256578 3826 256814
rect 4062 256578 39506 256814
rect 39742 256578 39826 256814
rect 40062 256578 75506 256814
rect 75742 256578 75826 256814
rect 76062 256578 111506 256814
rect 111742 256578 111826 256814
rect 112062 256578 147506 256814
rect 147742 256578 147826 256814
rect 148062 256578 183506 256814
rect 183742 256578 183826 256814
rect 184062 256578 219506 256814
rect 219742 256578 219826 256814
rect 220062 256578 255506 256814
rect 255742 256578 255826 256814
rect 256062 256578 291506 256814
rect 291742 256578 291826 256814
rect 292062 256578 327506 256814
rect 327742 256578 327826 256814
rect 328062 256578 363506 256814
rect 363742 256578 363826 256814
rect 364062 256578 399506 256814
rect 399742 256578 399826 256814
rect 400062 256578 435506 256814
rect 435742 256578 435826 256814
rect 436062 256578 471506 256814
rect 471742 256578 471826 256814
rect 472062 256578 507506 256814
rect 507742 256578 507826 256814
rect 508062 256578 543506 256814
rect 543742 256578 543826 256814
rect 544062 256578 579506 256814
rect 579742 256578 579826 256814
rect 580062 256578 587262 256814
rect 587498 256578 587582 256814
rect 587818 256578 592650 256814
rect -8726 256546 592650 256578
rect -8726 255894 592650 255926
rect -8726 255658 -2934 255894
rect -2698 255658 -2614 255894
rect -2378 255658 2266 255894
rect 2502 255658 2586 255894
rect 2822 255658 38266 255894
rect 38502 255658 38586 255894
rect 38822 255658 74266 255894
rect 74502 255658 74586 255894
rect 74822 255658 110266 255894
rect 110502 255658 110586 255894
rect 110822 255658 146266 255894
rect 146502 255658 146586 255894
rect 146822 255658 182266 255894
rect 182502 255658 182586 255894
rect 182822 255658 218266 255894
rect 218502 255658 218586 255894
rect 218822 255658 254266 255894
rect 254502 255658 254586 255894
rect 254822 255658 290266 255894
rect 290502 255658 290586 255894
rect 290822 255658 326266 255894
rect 326502 255658 326586 255894
rect 326822 255658 362266 255894
rect 362502 255658 362586 255894
rect 362822 255658 398266 255894
rect 398502 255658 398586 255894
rect 398822 255658 434266 255894
rect 434502 255658 434586 255894
rect 434822 255658 470266 255894
rect 470502 255658 470586 255894
rect 470822 255658 506266 255894
rect 506502 255658 506586 255894
rect 506822 255658 542266 255894
rect 542502 255658 542586 255894
rect 542822 255658 578266 255894
rect 578502 255658 578586 255894
rect 578822 255658 586302 255894
rect 586538 255658 586622 255894
rect 586858 255658 592650 255894
rect -8726 255574 592650 255658
rect -8726 255338 -2934 255574
rect -2698 255338 -2614 255574
rect -2378 255338 2266 255574
rect 2502 255338 2586 255574
rect 2822 255338 38266 255574
rect 38502 255338 38586 255574
rect 38822 255338 74266 255574
rect 74502 255338 74586 255574
rect 74822 255338 110266 255574
rect 110502 255338 110586 255574
rect 110822 255338 146266 255574
rect 146502 255338 146586 255574
rect 146822 255338 182266 255574
rect 182502 255338 182586 255574
rect 182822 255338 218266 255574
rect 218502 255338 218586 255574
rect 218822 255338 254266 255574
rect 254502 255338 254586 255574
rect 254822 255338 290266 255574
rect 290502 255338 290586 255574
rect 290822 255338 326266 255574
rect 326502 255338 326586 255574
rect 326822 255338 362266 255574
rect 362502 255338 362586 255574
rect 362822 255338 398266 255574
rect 398502 255338 398586 255574
rect 398822 255338 434266 255574
rect 434502 255338 434586 255574
rect 434822 255338 470266 255574
rect 470502 255338 470586 255574
rect 470822 255338 506266 255574
rect 506502 255338 506586 255574
rect 506822 255338 542266 255574
rect 542502 255338 542586 255574
rect 542822 255338 578266 255574
rect 578502 255338 578586 255574
rect 578822 255338 586302 255574
rect 586538 255338 586622 255574
rect 586858 255338 592650 255574
rect -8726 255306 592650 255338
rect -8726 254654 592650 254686
rect -8726 254418 -1974 254654
rect -1738 254418 -1654 254654
rect -1418 254418 1026 254654
rect 1262 254418 1346 254654
rect 1582 254418 37026 254654
rect 37262 254418 37346 254654
rect 37582 254418 73026 254654
rect 73262 254418 73346 254654
rect 73582 254418 109026 254654
rect 109262 254418 109346 254654
rect 109582 254418 145026 254654
rect 145262 254418 145346 254654
rect 145582 254418 181026 254654
rect 181262 254418 181346 254654
rect 181582 254418 217026 254654
rect 217262 254418 217346 254654
rect 217582 254418 253026 254654
rect 253262 254418 253346 254654
rect 253582 254418 289026 254654
rect 289262 254418 289346 254654
rect 289582 254418 325026 254654
rect 325262 254418 325346 254654
rect 325582 254418 361026 254654
rect 361262 254418 361346 254654
rect 361582 254418 397026 254654
rect 397262 254418 397346 254654
rect 397582 254418 433026 254654
rect 433262 254418 433346 254654
rect 433582 254418 469026 254654
rect 469262 254418 469346 254654
rect 469582 254418 505026 254654
rect 505262 254418 505346 254654
rect 505582 254418 541026 254654
rect 541262 254418 541346 254654
rect 541582 254418 577026 254654
rect 577262 254418 577346 254654
rect 577582 254418 585342 254654
rect 585578 254418 585662 254654
rect 585898 254418 592650 254654
rect -8726 254334 592650 254418
rect -8726 254098 -1974 254334
rect -1738 254098 -1654 254334
rect -1418 254098 1026 254334
rect 1262 254098 1346 254334
rect 1582 254098 37026 254334
rect 37262 254098 37346 254334
rect 37582 254098 73026 254334
rect 73262 254098 73346 254334
rect 73582 254098 109026 254334
rect 109262 254098 109346 254334
rect 109582 254098 145026 254334
rect 145262 254098 145346 254334
rect 145582 254098 181026 254334
rect 181262 254098 181346 254334
rect 181582 254098 217026 254334
rect 217262 254098 217346 254334
rect 217582 254098 253026 254334
rect 253262 254098 253346 254334
rect 253582 254098 289026 254334
rect 289262 254098 289346 254334
rect 289582 254098 325026 254334
rect 325262 254098 325346 254334
rect 325582 254098 361026 254334
rect 361262 254098 361346 254334
rect 361582 254098 397026 254334
rect 397262 254098 397346 254334
rect 397582 254098 433026 254334
rect 433262 254098 433346 254334
rect 433582 254098 469026 254334
rect 469262 254098 469346 254334
rect 469582 254098 505026 254334
rect 505262 254098 505346 254334
rect 505582 254098 541026 254334
rect 541262 254098 541346 254334
rect 541582 254098 577026 254334
rect 577262 254098 577346 254334
rect 577582 254098 585342 254334
rect 585578 254098 585662 254334
rect 585898 254098 592650 254334
rect -8726 254066 592650 254098
rect -8726 227334 592650 227366
rect -8726 227098 -8694 227334
rect -8458 227098 -8374 227334
rect -8138 227098 9706 227334
rect 9942 227098 10026 227334
rect 10262 227098 45706 227334
rect 45942 227098 46026 227334
rect 46262 227098 81706 227334
rect 81942 227098 82026 227334
rect 82262 227098 117706 227334
rect 117942 227098 118026 227334
rect 118262 227098 153706 227334
rect 153942 227098 154026 227334
rect 154262 227098 189706 227334
rect 189942 227098 190026 227334
rect 190262 227098 225706 227334
rect 225942 227098 226026 227334
rect 226262 227098 261706 227334
rect 261942 227098 262026 227334
rect 262262 227098 297706 227334
rect 297942 227098 298026 227334
rect 298262 227098 333706 227334
rect 333942 227098 334026 227334
rect 334262 227098 369706 227334
rect 369942 227098 370026 227334
rect 370262 227098 405706 227334
rect 405942 227098 406026 227334
rect 406262 227098 441706 227334
rect 441942 227098 442026 227334
rect 442262 227098 477706 227334
rect 477942 227098 478026 227334
rect 478262 227098 513706 227334
rect 513942 227098 514026 227334
rect 514262 227098 549706 227334
rect 549942 227098 550026 227334
rect 550262 227098 592062 227334
rect 592298 227098 592382 227334
rect 592618 227098 592650 227334
rect -8726 227014 592650 227098
rect -8726 226778 -8694 227014
rect -8458 226778 -8374 227014
rect -8138 226778 9706 227014
rect 9942 226778 10026 227014
rect 10262 226778 45706 227014
rect 45942 226778 46026 227014
rect 46262 226778 81706 227014
rect 81942 226778 82026 227014
rect 82262 226778 117706 227014
rect 117942 226778 118026 227014
rect 118262 226778 153706 227014
rect 153942 226778 154026 227014
rect 154262 226778 189706 227014
rect 189942 226778 190026 227014
rect 190262 226778 225706 227014
rect 225942 226778 226026 227014
rect 226262 226778 261706 227014
rect 261942 226778 262026 227014
rect 262262 226778 297706 227014
rect 297942 226778 298026 227014
rect 298262 226778 333706 227014
rect 333942 226778 334026 227014
rect 334262 226778 369706 227014
rect 369942 226778 370026 227014
rect 370262 226778 405706 227014
rect 405942 226778 406026 227014
rect 406262 226778 441706 227014
rect 441942 226778 442026 227014
rect 442262 226778 477706 227014
rect 477942 226778 478026 227014
rect 478262 226778 513706 227014
rect 513942 226778 514026 227014
rect 514262 226778 549706 227014
rect 549942 226778 550026 227014
rect 550262 226778 592062 227014
rect 592298 226778 592382 227014
rect 592618 226778 592650 227014
rect -8726 226746 592650 226778
rect -8726 226094 592650 226126
rect -8726 225858 -7734 226094
rect -7498 225858 -7414 226094
rect -7178 225858 8466 226094
rect 8702 225858 8786 226094
rect 9022 225858 44466 226094
rect 44702 225858 44786 226094
rect 45022 225858 80466 226094
rect 80702 225858 80786 226094
rect 81022 225858 116466 226094
rect 116702 225858 116786 226094
rect 117022 225858 152466 226094
rect 152702 225858 152786 226094
rect 153022 225858 188466 226094
rect 188702 225858 188786 226094
rect 189022 225858 224466 226094
rect 224702 225858 224786 226094
rect 225022 225858 260466 226094
rect 260702 225858 260786 226094
rect 261022 225858 296466 226094
rect 296702 225858 296786 226094
rect 297022 225858 332466 226094
rect 332702 225858 332786 226094
rect 333022 225858 368466 226094
rect 368702 225858 368786 226094
rect 369022 225858 404466 226094
rect 404702 225858 404786 226094
rect 405022 225858 440466 226094
rect 440702 225858 440786 226094
rect 441022 225858 476466 226094
rect 476702 225858 476786 226094
rect 477022 225858 512466 226094
rect 512702 225858 512786 226094
rect 513022 225858 548466 226094
rect 548702 225858 548786 226094
rect 549022 225858 591102 226094
rect 591338 225858 591422 226094
rect 591658 225858 592650 226094
rect -8726 225774 592650 225858
rect -8726 225538 -7734 225774
rect -7498 225538 -7414 225774
rect -7178 225538 8466 225774
rect 8702 225538 8786 225774
rect 9022 225538 44466 225774
rect 44702 225538 44786 225774
rect 45022 225538 80466 225774
rect 80702 225538 80786 225774
rect 81022 225538 116466 225774
rect 116702 225538 116786 225774
rect 117022 225538 152466 225774
rect 152702 225538 152786 225774
rect 153022 225538 188466 225774
rect 188702 225538 188786 225774
rect 189022 225538 224466 225774
rect 224702 225538 224786 225774
rect 225022 225538 260466 225774
rect 260702 225538 260786 225774
rect 261022 225538 296466 225774
rect 296702 225538 296786 225774
rect 297022 225538 332466 225774
rect 332702 225538 332786 225774
rect 333022 225538 368466 225774
rect 368702 225538 368786 225774
rect 369022 225538 404466 225774
rect 404702 225538 404786 225774
rect 405022 225538 440466 225774
rect 440702 225538 440786 225774
rect 441022 225538 476466 225774
rect 476702 225538 476786 225774
rect 477022 225538 512466 225774
rect 512702 225538 512786 225774
rect 513022 225538 548466 225774
rect 548702 225538 548786 225774
rect 549022 225538 591102 225774
rect 591338 225538 591422 225774
rect 591658 225538 592650 225774
rect -8726 225506 592650 225538
rect -8726 224854 592650 224886
rect -8726 224618 -6774 224854
rect -6538 224618 -6454 224854
rect -6218 224618 7226 224854
rect 7462 224618 7546 224854
rect 7782 224618 43226 224854
rect 43462 224618 43546 224854
rect 43782 224618 79226 224854
rect 79462 224618 79546 224854
rect 79782 224618 115226 224854
rect 115462 224618 115546 224854
rect 115782 224618 151226 224854
rect 151462 224618 151546 224854
rect 151782 224618 187226 224854
rect 187462 224618 187546 224854
rect 187782 224618 223226 224854
rect 223462 224618 223546 224854
rect 223782 224618 259226 224854
rect 259462 224618 259546 224854
rect 259782 224618 295226 224854
rect 295462 224618 295546 224854
rect 295782 224618 331226 224854
rect 331462 224618 331546 224854
rect 331782 224618 367226 224854
rect 367462 224618 367546 224854
rect 367782 224618 403226 224854
rect 403462 224618 403546 224854
rect 403782 224618 439226 224854
rect 439462 224618 439546 224854
rect 439782 224618 475226 224854
rect 475462 224618 475546 224854
rect 475782 224618 511226 224854
rect 511462 224618 511546 224854
rect 511782 224618 547226 224854
rect 547462 224618 547546 224854
rect 547782 224618 590142 224854
rect 590378 224618 590462 224854
rect 590698 224618 592650 224854
rect -8726 224534 592650 224618
rect -8726 224298 -6774 224534
rect -6538 224298 -6454 224534
rect -6218 224298 7226 224534
rect 7462 224298 7546 224534
rect 7782 224298 43226 224534
rect 43462 224298 43546 224534
rect 43782 224298 79226 224534
rect 79462 224298 79546 224534
rect 79782 224298 115226 224534
rect 115462 224298 115546 224534
rect 115782 224298 151226 224534
rect 151462 224298 151546 224534
rect 151782 224298 187226 224534
rect 187462 224298 187546 224534
rect 187782 224298 223226 224534
rect 223462 224298 223546 224534
rect 223782 224298 259226 224534
rect 259462 224298 259546 224534
rect 259782 224298 295226 224534
rect 295462 224298 295546 224534
rect 295782 224298 331226 224534
rect 331462 224298 331546 224534
rect 331782 224298 367226 224534
rect 367462 224298 367546 224534
rect 367782 224298 403226 224534
rect 403462 224298 403546 224534
rect 403782 224298 439226 224534
rect 439462 224298 439546 224534
rect 439782 224298 475226 224534
rect 475462 224298 475546 224534
rect 475782 224298 511226 224534
rect 511462 224298 511546 224534
rect 511782 224298 547226 224534
rect 547462 224298 547546 224534
rect 547782 224298 590142 224534
rect 590378 224298 590462 224534
rect 590698 224298 592650 224534
rect -8726 224266 592650 224298
rect -8726 223614 592650 223646
rect -8726 223378 -5814 223614
rect -5578 223378 -5494 223614
rect -5258 223378 5986 223614
rect 6222 223378 6306 223614
rect 6542 223378 41986 223614
rect 42222 223378 42306 223614
rect 42542 223378 77986 223614
rect 78222 223378 78306 223614
rect 78542 223378 113986 223614
rect 114222 223378 114306 223614
rect 114542 223378 149986 223614
rect 150222 223378 150306 223614
rect 150542 223378 185986 223614
rect 186222 223378 186306 223614
rect 186542 223378 221986 223614
rect 222222 223378 222306 223614
rect 222542 223378 257986 223614
rect 258222 223378 258306 223614
rect 258542 223378 293986 223614
rect 294222 223378 294306 223614
rect 294542 223378 329986 223614
rect 330222 223378 330306 223614
rect 330542 223378 365986 223614
rect 366222 223378 366306 223614
rect 366542 223378 401986 223614
rect 402222 223378 402306 223614
rect 402542 223378 437986 223614
rect 438222 223378 438306 223614
rect 438542 223378 473986 223614
rect 474222 223378 474306 223614
rect 474542 223378 509986 223614
rect 510222 223378 510306 223614
rect 510542 223378 545986 223614
rect 546222 223378 546306 223614
rect 546542 223378 581986 223614
rect 582222 223378 582306 223614
rect 582542 223378 589182 223614
rect 589418 223378 589502 223614
rect 589738 223378 592650 223614
rect -8726 223294 592650 223378
rect -8726 223058 -5814 223294
rect -5578 223058 -5494 223294
rect -5258 223058 5986 223294
rect 6222 223058 6306 223294
rect 6542 223058 41986 223294
rect 42222 223058 42306 223294
rect 42542 223058 77986 223294
rect 78222 223058 78306 223294
rect 78542 223058 113986 223294
rect 114222 223058 114306 223294
rect 114542 223058 149986 223294
rect 150222 223058 150306 223294
rect 150542 223058 185986 223294
rect 186222 223058 186306 223294
rect 186542 223058 221986 223294
rect 222222 223058 222306 223294
rect 222542 223058 257986 223294
rect 258222 223058 258306 223294
rect 258542 223058 293986 223294
rect 294222 223058 294306 223294
rect 294542 223058 329986 223294
rect 330222 223058 330306 223294
rect 330542 223058 365986 223294
rect 366222 223058 366306 223294
rect 366542 223058 401986 223294
rect 402222 223058 402306 223294
rect 402542 223058 437986 223294
rect 438222 223058 438306 223294
rect 438542 223058 473986 223294
rect 474222 223058 474306 223294
rect 474542 223058 509986 223294
rect 510222 223058 510306 223294
rect 510542 223058 545986 223294
rect 546222 223058 546306 223294
rect 546542 223058 581986 223294
rect 582222 223058 582306 223294
rect 582542 223058 589182 223294
rect 589418 223058 589502 223294
rect 589738 223058 592650 223294
rect -8726 223026 592650 223058
rect -8726 222374 592650 222406
rect -8726 222138 -4854 222374
rect -4618 222138 -4534 222374
rect -4298 222138 4746 222374
rect 4982 222138 5066 222374
rect 5302 222138 40746 222374
rect 40982 222138 41066 222374
rect 41302 222138 76746 222374
rect 76982 222138 77066 222374
rect 77302 222138 112746 222374
rect 112982 222138 113066 222374
rect 113302 222138 148746 222374
rect 148982 222138 149066 222374
rect 149302 222138 184746 222374
rect 184982 222138 185066 222374
rect 185302 222138 220746 222374
rect 220982 222138 221066 222374
rect 221302 222138 256746 222374
rect 256982 222138 257066 222374
rect 257302 222138 292746 222374
rect 292982 222138 293066 222374
rect 293302 222138 328746 222374
rect 328982 222138 329066 222374
rect 329302 222138 364746 222374
rect 364982 222138 365066 222374
rect 365302 222138 400746 222374
rect 400982 222138 401066 222374
rect 401302 222138 436746 222374
rect 436982 222138 437066 222374
rect 437302 222138 472746 222374
rect 472982 222138 473066 222374
rect 473302 222138 508746 222374
rect 508982 222138 509066 222374
rect 509302 222138 544746 222374
rect 544982 222138 545066 222374
rect 545302 222138 580746 222374
rect 580982 222138 581066 222374
rect 581302 222138 588222 222374
rect 588458 222138 588542 222374
rect 588778 222138 592650 222374
rect -8726 222054 592650 222138
rect -8726 221818 -4854 222054
rect -4618 221818 -4534 222054
rect -4298 221818 4746 222054
rect 4982 221818 5066 222054
rect 5302 221818 40746 222054
rect 40982 221818 41066 222054
rect 41302 221818 76746 222054
rect 76982 221818 77066 222054
rect 77302 221818 112746 222054
rect 112982 221818 113066 222054
rect 113302 221818 148746 222054
rect 148982 221818 149066 222054
rect 149302 221818 184746 222054
rect 184982 221818 185066 222054
rect 185302 221818 220746 222054
rect 220982 221818 221066 222054
rect 221302 221818 256746 222054
rect 256982 221818 257066 222054
rect 257302 221818 292746 222054
rect 292982 221818 293066 222054
rect 293302 221818 328746 222054
rect 328982 221818 329066 222054
rect 329302 221818 364746 222054
rect 364982 221818 365066 222054
rect 365302 221818 400746 222054
rect 400982 221818 401066 222054
rect 401302 221818 436746 222054
rect 436982 221818 437066 222054
rect 437302 221818 472746 222054
rect 472982 221818 473066 222054
rect 473302 221818 508746 222054
rect 508982 221818 509066 222054
rect 509302 221818 544746 222054
rect 544982 221818 545066 222054
rect 545302 221818 580746 222054
rect 580982 221818 581066 222054
rect 581302 221818 588222 222054
rect 588458 221818 588542 222054
rect 588778 221818 592650 222054
rect -8726 221786 592650 221818
rect -8726 221134 592650 221166
rect -8726 220898 -3894 221134
rect -3658 220898 -3574 221134
rect -3338 220898 3506 221134
rect 3742 220898 3826 221134
rect 4062 220898 39506 221134
rect 39742 220898 39826 221134
rect 40062 220898 75506 221134
rect 75742 220898 75826 221134
rect 76062 220898 111506 221134
rect 111742 220898 111826 221134
rect 112062 220898 147506 221134
rect 147742 220898 147826 221134
rect 148062 220898 183506 221134
rect 183742 220898 183826 221134
rect 184062 220898 219506 221134
rect 219742 220898 219826 221134
rect 220062 220898 255506 221134
rect 255742 220898 255826 221134
rect 256062 220898 291506 221134
rect 291742 220898 291826 221134
rect 292062 220898 327506 221134
rect 327742 220898 327826 221134
rect 328062 220898 363506 221134
rect 363742 220898 363826 221134
rect 364062 220898 399506 221134
rect 399742 220898 399826 221134
rect 400062 220898 435506 221134
rect 435742 220898 435826 221134
rect 436062 220898 471506 221134
rect 471742 220898 471826 221134
rect 472062 220898 507506 221134
rect 507742 220898 507826 221134
rect 508062 220898 543506 221134
rect 543742 220898 543826 221134
rect 544062 220898 579506 221134
rect 579742 220898 579826 221134
rect 580062 220898 587262 221134
rect 587498 220898 587582 221134
rect 587818 220898 592650 221134
rect -8726 220814 592650 220898
rect -8726 220578 -3894 220814
rect -3658 220578 -3574 220814
rect -3338 220578 3506 220814
rect 3742 220578 3826 220814
rect 4062 220578 39506 220814
rect 39742 220578 39826 220814
rect 40062 220578 75506 220814
rect 75742 220578 75826 220814
rect 76062 220578 111506 220814
rect 111742 220578 111826 220814
rect 112062 220578 147506 220814
rect 147742 220578 147826 220814
rect 148062 220578 183506 220814
rect 183742 220578 183826 220814
rect 184062 220578 219506 220814
rect 219742 220578 219826 220814
rect 220062 220578 255506 220814
rect 255742 220578 255826 220814
rect 256062 220578 291506 220814
rect 291742 220578 291826 220814
rect 292062 220578 327506 220814
rect 327742 220578 327826 220814
rect 328062 220578 363506 220814
rect 363742 220578 363826 220814
rect 364062 220578 399506 220814
rect 399742 220578 399826 220814
rect 400062 220578 435506 220814
rect 435742 220578 435826 220814
rect 436062 220578 471506 220814
rect 471742 220578 471826 220814
rect 472062 220578 507506 220814
rect 507742 220578 507826 220814
rect 508062 220578 543506 220814
rect 543742 220578 543826 220814
rect 544062 220578 579506 220814
rect 579742 220578 579826 220814
rect 580062 220578 587262 220814
rect 587498 220578 587582 220814
rect 587818 220578 592650 220814
rect -8726 220546 592650 220578
rect -8726 219894 592650 219926
rect -8726 219658 -2934 219894
rect -2698 219658 -2614 219894
rect -2378 219658 2266 219894
rect 2502 219658 2586 219894
rect 2822 219658 38266 219894
rect 38502 219658 38586 219894
rect 38822 219658 74266 219894
rect 74502 219658 74586 219894
rect 74822 219658 110266 219894
rect 110502 219658 110586 219894
rect 110822 219658 146266 219894
rect 146502 219658 146586 219894
rect 146822 219658 182266 219894
rect 182502 219658 182586 219894
rect 182822 219658 218266 219894
rect 218502 219658 218586 219894
rect 218822 219658 254266 219894
rect 254502 219658 254586 219894
rect 254822 219658 290266 219894
rect 290502 219658 290586 219894
rect 290822 219658 326266 219894
rect 326502 219658 326586 219894
rect 326822 219658 362266 219894
rect 362502 219658 362586 219894
rect 362822 219658 398266 219894
rect 398502 219658 398586 219894
rect 398822 219658 434266 219894
rect 434502 219658 434586 219894
rect 434822 219658 470266 219894
rect 470502 219658 470586 219894
rect 470822 219658 506266 219894
rect 506502 219658 506586 219894
rect 506822 219658 542266 219894
rect 542502 219658 542586 219894
rect 542822 219658 578266 219894
rect 578502 219658 578586 219894
rect 578822 219658 586302 219894
rect 586538 219658 586622 219894
rect 586858 219658 592650 219894
rect -8726 219574 592650 219658
rect -8726 219338 -2934 219574
rect -2698 219338 -2614 219574
rect -2378 219338 2266 219574
rect 2502 219338 2586 219574
rect 2822 219338 38266 219574
rect 38502 219338 38586 219574
rect 38822 219338 74266 219574
rect 74502 219338 74586 219574
rect 74822 219338 110266 219574
rect 110502 219338 110586 219574
rect 110822 219338 146266 219574
rect 146502 219338 146586 219574
rect 146822 219338 182266 219574
rect 182502 219338 182586 219574
rect 182822 219338 218266 219574
rect 218502 219338 218586 219574
rect 218822 219338 254266 219574
rect 254502 219338 254586 219574
rect 254822 219338 290266 219574
rect 290502 219338 290586 219574
rect 290822 219338 326266 219574
rect 326502 219338 326586 219574
rect 326822 219338 362266 219574
rect 362502 219338 362586 219574
rect 362822 219338 398266 219574
rect 398502 219338 398586 219574
rect 398822 219338 434266 219574
rect 434502 219338 434586 219574
rect 434822 219338 470266 219574
rect 470502 219338 470586 219574
rect 470822 219338 506266 219574
rect 506502 219338 506586 219574
rect 506822 219338 542266 219574
rect 542502 219338 542586 219574
rect 542822 219338 578266 219574
rect 578502 219338 578586 219574
rect 578822 219338 586302 219574
rect 586538 219338 586622 219574
rect 586858 219338 592650 219574
rect -8726 219306 592650 219338
rect -8726 218654 592650 218686
rect -8726 218418 -1974 218654
rect -1738 218418 -1654 218654
rect -1418 218418 1026 218654
rect 1262 218418 1346 218654
rect 1582 218418 37026 218654
rect 37262 218418 37346 218654
rect 37582 218418 73026 218654
rect 73262 218418 73346 218654
rect 73582 218418 109026 218654
rect 109262 218418 109346 218654
rect 109582 218418 145026 218654
rect 145262 218418 145346 218654
rect 145582 218418 181026 218654
rect 181262 218418 181346 218654
rect 181582 218418 217026 218654
rect 217262 218418 217346 218654
rect 217582 218418 253026 218654
rect 253262 218418 253346 218654
rect 253582 218418 289026 218654
rect 289262 218418 289346 218654
rect 289582 218418 325026 218654
rect 325262 218418 325346 218654
rect 325582 218418 361026 218654
rect 361262 218418 361346 218654
rect 361582 218418 397026 218654
rect 397262 218418 397346 218654
rect 397582 218418 433026 218654
rect 433262 218418 433346 218654
rect 433582 218418 469026 218654
rect 469262 218418 469346 218654
rect 469582 218418 505026 218654
rect 505262 218418 505346 218654
rect 505582 218418 541026 218654
rect 541262 218418 541346 218654
rect 541582 218418 577026 218654
rect 577262 218418 577346 218654
rect 577582 218418 585342 218654
rect 585578 218418 585662 218654
rect 585898 218418 592650 218654
rect -8726 218334 592650 218418
rect -8726 218098 -1974 218334
rect -1738 218098 -1654 218334
rect -1418 218098 1026 218334
rect 1262 218098 1346 218334
rect 1582 218098 37026 218334
rect 37262 218098 37346 218334
rect 37582 218098 73026 218334
rect 73262 218098 73346 218334
rect 73582 218098 109026 218334
rect 109262 218098 109346 218334
rect 109582 218098 145026 218334
rect 145262 218098 145346 218334
rect 145582 218098 181026 218334
rect 181262 218098 181346 218334
rect 181582 218098 217026 218334
rect 217262 218098 217346 218334
rect 217582 218098 253026 218334
rect 253262 218098 253346 218334
rect 253582 218098 289026 218334
rect 289262 218098 289346 218334
rect 289582 218098 325026 218334
rect 325262 218098 325346 218334
rect 325582 218098 361026 218334
rect 361262 218098 361346 218334
rect 361582 218098 397026 218334
rect 397262 218098 397346 218334
rect 397582 218098 433026 218334
rect 433262 218098 433346 218334
rect 433582 218098 469026 218334
rect 469262 218098 469346 218334
rect 469582 218098 505026 218334
rect 505262 218098 505346 218334
rect 505582 218098 541026 218334
rect 541262 218098 541346 218334
rect 541582 218098 577026 218334
rect 577262 218098 577346 218334
rect 577582 218098 585342 218334
rect 585578 218098 585662 218334
rect 585898 218098 592650 218334
rect -8726 218066 592650 218098
rect -8726 191334 592650 191366
rect -8726 191098 -8694 191334
rect -8458 191098 -8374 191334
rect -8138 191098 9706 191334
rect 9942 191098 10026 191334
rect 10262 191098 45706 191334
rect 45942 191098 46026 191334
rect 46262 191098 81706 191334
rect 81942 191098 82026 191334
rect 82262 191098 117706 191334
rect 117942 191098 118026 191334
rect 118262 191098 153706 191334
rect 153942 191098 154026 191334
rect 154262 191098 189706 191334
rect 189942 191098 190026 191334
rect 190262 191098 225706 191334
rect 225942 191098 226026 191334
rect 226262 191098 261706 191334
rect 261942 191098 262026 191334
rect 262262 191098 297706 191334
rect 297942 191098 298026 191334
rect 298262 191098 333706 191334
rect 333942 191098 334026 191334
rect 334262 191098 369706 191334
rect 369942 191098 370026 191334
rect 370262 191098 405706 191334
rect 405942 191098 406026 191334
rect 406262 191098 441706 191334
rect 441942 191098 442026 191334
rect 442262 191098 477706 191334
rect 477942 191098 478026 191334
rect 478262 191098 513706 191334
rect 513942 191098 514026 191334
rect 514262 191098 549706 191334
rect 549942 191098 550026 191334
rect 550262 191098 592062 191334
rect 592298 191098 592382 191334
rect 592618 191098 592650 191334
rect -8726 191014 592650 191098
rect -8726 190778 -8694 191014
rect -8458 190778 -8374 191014
rect -8138 190778 9706 191014
rect 9942 190778 10026 191014
rect 10262 190778 45706 191014
rect 45942 190778 46026 191014
rect 46262 190778 81706 191014
rect 81942 190778 82026 191014
rect 82262 190778 117706 191014
rect 117942 190778 118026 191014
rect 118262 190778 153706 191014
rect 153942 190778 154026 191014
rect 154262 190778 189706 191014
rect 189942 190778 190026 191014
rect 190262 190778 225706 191014
rect 225942 190778 226026 191014
rect 226262 190778 261706 191014
rect 261942 190778 262026 191014
rect 262262 190778 297706 191014
rect 297942 190778 298026 191014
rect 298262 190778 333706 191014
rect 333942 190778 334026 191014
rect 334262 190778 369706 191014
rect 369942 190778 370026 191014
rect 370262 190778 405706 191014
rect 405942 190778 406026 191014
rect 406262 190778 441706 191014
rect 441942 190778 442026 191014
rect 442262 190778 477706 191014
rect 477942 190778 478026 191014
rect 478262 190778 513706 191014
rect 513942 190778 514026 191014
rect 514262 190778 549706 191014
rect 549942 190778 550026 191014
rect 550262 190778 592062 191014
rect 592298 190778 592382 191014
rect 592618 190778 592650 191014
rect -8726 190746 592650 190778
rect -8726 190094 592650 190126
rect -8726 189858 -7734 190094
rect -7498 189858 -7414 190094
rect -7178 189858 8466 190094
rect 8702 189858 8786 190094
rect 9022 189858 44466 190094
rect 44702 189858 44786 190094
rect 45022 189858 80466 190094
rect 80702 189858 80786 190094
rect 81022 189858 116466 190094
rect 116702 189858 116786 190094
rect 117022 189858 152466 190094
rect 152702 189858 152786 190094
rect 153022 189858 188466 190094
rect 188702 189858 188786 190094
rect 189022 189858 224466 190094
rect 224702 189858 224786 190094
rect 225022 189858 260466 190094
rect 260702 189858 260786 190094
rect 261022 189858 296466 190094
rect 296702 189858 296786 190094
rect 297022 189858 332466 190094
rect 332702 189858 332786 190094
rect 333022 189858 368466 190094
rect 368702 189858 368786 190094
rect 369022 189858 404466 190094
rect 404702 189858 404786 190094
rect 405022 189858 440466 190094
rect 440702 189858 440786 190094
rect 441022 189858 476466 190094
rect 476702 189858 476786 190094
rect 477022 189858 512466 190094
rect 512702 189858 512786 190094
rect 513022 189858 548466 190094
rect 548702 189858 548786 190094
rect 549022 189858 591102 190094
rect 591338 189858 591422 190094
rect 591658 189858 592650 190094
rect -8726 189774 592650 189858
rect -8726 189538 -7734 189774
rect -7498 189538 -7414 189774
rect -7178 189538 8466 189774
rect 8702 189538 8786 189774
rect 9022 189538 44466 189774
rect 44702 189538 44786 189774
rect 45022 189538 80466 189774
rect 80702 189538 80786 189774
rect 81022 189538 116466 189774
rect 116702 189538 116786 189774
rect 117022 189538 152466 189774
rect 152702 189538 152786 189774
rect 153022 189538 188466 189774
rect 188702 189538 188786 189774
rect 189022 189538 224466 189774
rect 224702 189538 224786 189774
rect 225022 189538 260466 189774
rect 260702 189538 260786 189774
rect 261022 189538 296466 189774
rect 296702 189538 296786 189774
rect 297022 189538 332466 189774
rect 332702 189538 332786 189774
rect 333022 189538 368466 189774
rect 368702 189538 368786 189774
rect 369022 189538 404466 189774
rect 404702 189538 404786 189774
rect 405022 189538 440466 189774
rect 440702 189538 440786 189774
rect 441022 189538 476466 189774
rect 476702 189538 476786 189774
rect 477022 189538 512466 189774
rect 512702 189538 512786 189774
rect 513022 189538 548466 189774
rect 548702 189538 548786 189774
rect 549022 189538 591102 189774
rect 591338 189538 591422 189774
rect 591658 189538 592650 189774
rect -8726 189506 592650 189538
rect -8726 188854 592650 188886
rect -8726 188618 -6774 188854
rect -6538 188618 -6454 188854
rect -6218 188618 7226 188854
rect 7462 188618 7546 188854
rect 7782 188618 43226 188854
rect 43462 188618 43546 188854
rect 43782 188618 79226 188854
rect 79462 188618 79546 188854
rect 79782 188618 115226 188854
rect 115462 188618 115546 188854
rect 115782 188618 151226 188854
rect 151462 188618 151546 188854
rect 151782 188618 187226 188854
rect 187462 188618 187546 188854
rect 187782 188618 223226 188854
rect 223462 188618 223546 188854
rect 223782 188618 259226 188854
rect 259462 188618 259546 188854
rect 259782 188618 295226 188854
rect 295462 188618 295546 188854
rect 295782 188618 331226 188854
rect 331462 188618 331546 188854
rect 331782 188618 367226 188854
rect 367462 188618 367546 188854
rect 367782 188618 403226 188854
rect 403462 188618 403546 188854
rect 403782 188618 439226 188854
rect 439462 188618 439546 188854
rect 439782 188618 475226 188854
rect 475462 188618 475546 188854
rect 475782 188618 511226 188854
rect 511462 188618 511546 188854
rect 511782 188618 547226 188854
rect 547462 188618 547546 188854
rect 547782 188618 590142 188854
rect 590378 188618 590462 188854
rect 590698 188618 592650 188854
rect -8726 188534 592650 188618
rect -8726 188298 -6774 188534
rect -6538 188298 -6454 188534
rect -6218 188298 7226 188534
rect 7462 188298 7546 188534
rect 7782 188298 43226 188534
rect 43462 188298 43546 188534
rect 43782 188298 79226 188534
rect 79462 188298 79546 188534
rect 79782 188298 115226 188534
rect 115462 188298 115546 188534
rect 115782 188298 151226 188534
rect 151462 188298 151546 188534
rect 151782 188298 187226 188534
rect 187462 188298 187546 188534
rect 187782 188298 223226 188534
rect 223462 188298 223546 188534
rect 223782 188298 259226 188534
rect 259462 188298 259546 188534
rect 259782 188298 295226 188534
rect 295462 188298 295546 188534
rect 295782 188298 331226 188534
rect 331462 188298 331546 188534
rect 331782 188298 367226 188534
rect 367462 188298 367546 188534
rect 367782 188298 403226 188534
rect 403462 188298 403546 188534
rect 403782 188298 439226 188534
rect 439462 188298 439546 188534
rect 439782 188298 475226 188534
rect 475462 188298 475546 188534
rect 475782 188298 511226 188534
rect 511462 188298 511546 188534
rect 511782 188298 547226 188534
rect 547462 188298 547546 188534
rect 547782 188298 590142 188534
rect 590378 188298 590462 188534
rect 590698 188298 592650 188534
rect -8726 188266 592650 188298
rect -8726 187614 592650 187646
rect -8726 187378 -5814 187614
rect -5578 187378 -5494 187614
rect -5258 187378 5986 187614
rect 6222 187378 6306 187614
rect 6542 187378 41986 187614
rect 42222 187378 42306 187614
rect 42542 187378 77986 187614
rect 78222 187378 78306 187614
rect 78542 187378 113986 187614
rect 114222 187378 114306 187614
rect 114542 187378 149986 187614
rect 150222 187378 150306 187614
rect 150542 187378 185986 187614
rect 186222 187378 186306 187614
rect 186542 187378 221986 187614
rect 222222 187378 222306 187614
rect 222542 187378 257986 187614
rect 258222 187378 258306 187614
rect 258542 187378 293986 187614
rect 294222 187378 294306 187614
rect 294542 187378 329986 187614
rect 330222 187378 330306 187614
rect 330542 187378 365986 187614
rect 366222 187378 366306 187614
rect 366542 187378 401986 187614
rect 402222 187378 402306 187614
rect 402542 187378 437986 187614
rect 438222 187378 438306 187614
rect 438542 187378 473986 187614
rect 474222 187378 474306 187614
rect 474542 187378 509986 187614
rect 510222 187378 510306 187614
rect 510542 187378 545986 187614
rect 546222 187378 546306 187614
rect 546542 187378 581986 187614
rect 582222 187378 582306 187614
rect 582542 187378 589182 187614
rect 589418 187378 589502 187614
rect 589738 187378 592650 187614
rect -8726 187294 592650 187378
rect -8726 187058 -5814 187294
rect -5578 187058 -5494 187294
rect -5258 187058 5986 187294
rect 6222 187058 6306 187294
rect 6542 187058 41986 187294
rect 42222 187058 42306 187294
rect 42542 187058 77986 187294
rect 78222 187058 78306 187294
rect 78542 187058 113986 187294
rect 114222 187058 114306 187294
rect 114542 187058 149986 187294
rect 150222 187058 150306 187294
rect 150542 187058 185986 187294
rect 186222 187058 186306 187294
rect 186542 187058 221986 187294
rect 222222 187058 222306 187294
rect 222542 187058 257986 187294
rect 258222 187058 258306 187294
rect 258542 187058 293986 187294
rect 294222 187058 294306 187294
rect 294542 187058 329986 187294
rect 330222 187058 330306 187294
rect 330542 187058 365986 187294
rect 366222 187058 366306 187294
rect 366542 187058 401986 187294
rect 402222 187058 402306 187294
rect 402542 187058 437986 187294
rect 438222 187058 438306 187294
rect 438542 187058 473986 187294
rect 474222 187058 474306 187294
rect 474542 187058 509986 187294
rect 510222 187058 510306 187294
rect 510542 187058 545986 187294
rect 546222 187058 546306 187294
rect 546542 187058 581986 187294
rect 582222 187058 582306 187294
rect 582542 187058 589182 187294
rect 589418 187058 589502 187294
rect 589738 187058 592650 187294
rect -8726 187026 592650 187058
rect -8726 186374 592650 186406
rect -8726 186138 -4854 186374
rect -4618 186138 -4534 186374
rect -4298 186138 4746 186374
rect 4982 186138 5066 186374
rect 5302 186138 40746 186374
rect 40982 186138 41066 186374
rect 41302 186138 76746 186374
rect 76982 186138 77066 186374
rect 77302 186138 112746 186374
rect 112982 186138 113066 186374
rect 113302 186138 148746 186374
rect 148982 186138 149066 186374
rect 149302 186138 184746 186374
rect 184982 186138 185066 186374
rect 185302 186138 220746 186374
rect 220982 186138 221066 186374
rect 221302 186138 256746 186374
rect 256982 186138 257066 186374
rect 257302 186138 292746 186374
rect 292982 186138 293066 186374
rect 293302 186138 328746 186374
rect 328982 186138 329066 186374
rect 329302 186138 364746 186374
rect 364982 186138 365066 186374
rect 365302 186138 400746 186374
rect 400982 186138 401066 186374
rect 401302 186138 436746 186374
rect 436982 186138 437066 186374
rect 437302 186138 472746 186374
rect 472982 186138 473066 186374
rect 473302 186138 508746 186374
rect 508982 186138 509066 186374
rect 509302 186138 544746 186374
rect 544982 186138 545066 186374
rect 545302 186138 580746 186374
rect 580982 186138 581066 186374
rect 581302 186138 588222 186374
rect 588458 186138 588542 186374
rect 588778 186138 592650 186374
rect -8726 186054 592650 186138
rect -8726 185818 -4854 186054
rect -4618 185818 -4534 186054
rect -4298 185818 4746 186054
rect 4982 185818 5066 186054
rect 5302 185818 40746 186054
rect 40982 185818 41066 186054
rect 41302 185818 76746 186054
rect 76982 185818 77066 186054
rect 77302 185818 112746 186054
rect 112982 185818 113066 186054
rect 113302 185818 148746 186054
rect 148982 185818 149066 186054
rect 149302 185818 184746 186054
rect 184982 185818 185066 186054
rect 185302 185818 220746 186054
rect 220982 185818 221066 186054
rect 221302 185818 256746 186054
rect 256982 185818 257066 186054
rect 257302 185818 292746 186054
rect 292982 185818 293066 186054
rect 293302 185818 328746 186054
rect 328982 185818 329066 186054
rect 329302 185818 364746 186054
rect 364982 185818 365066 186054
rect 365302 185818 400746 186054
rect 400982 185818 401066 186054
rect 401302 185818 436746 186054
rect 436982 185818 437066 186054
rect 437302 185818 472746 186054
rect 472982 185818 473066 186054
rect 473302 185818 508746 186054
rect 508982 185818 509066 186054
rect 509302 185818 544746 186054
rect 544982 185818 545066 186054
rect 545302 185818 580746 186054
rect 580982 185818 581066 186054
rect 581302 185818 588222 186054
rect 588458 185818 588542 186054
rect 588778 185818 592650 186054
rect -8726 185786 592650 185818
rect -8726 185134 592650 185166
rect -8726 184898 -3894 185134
rect -3658 184898 -3574 185134
rect -3338 184898 3506 185134
rect 3742 184898 3826 185134
rect 4062 184898 39506 185134
rect 39742 184898 39826 185134
rect 40062 184898 75506 185134
rect 75742 184898 75826 185134
rect 76062 184898 111506 185134
rect 111742 184898 111826 185134
rect 112062 184898 147506 185134
rect 147742 184898 147826 185134
rect 148062 184898 183506 185134
rect 183742 184898 183826 185134
rect 184062 184898 219506 185134
rect 219742 184898 219826 185134
rect 220062 184898 255506 185134
rect 255742 184898 255826 185134
rect 256062 184898 291506 185134
rect 291742 184898 291826 185134
rect 292062 184898 327506 185134
rect 327742 184898 327826 185134
rect 328062 184898 363506 185134
rect 363742 184898 363826 185134
rect 364062 184898 399506 185134
rect 399742 184898 399826 185134
rect 400062 184898 435506 185134
rect 435742 184898 435826 185134
rect 436062 184898 471506 185134
rect 471742 184898 471826 185134
rect 472062 184898 507506 185134
rect 507742 184898 507826 185134
rect 508062 184898 543506 185134
rect 543742 184898 543826 185134
rect 544062 184898 579506 185134
rect 579742 184898 579826 185134
rect 580062 184898 587262 185134
rect 587498 184898 587582 185134
rect 587818 184898 592650 185134
rect -8726 184814 592650 184898
rect -8726 184578 -3894 184814
rect -3658 184578 -3574 184814
rect -3338 184578 3506 184814
rect 3742 184578 3826 184814
rect 4062 184578 39506 184814
rect 39742 184578 39826 184814
rect 40062 184578 75506 184814
rect 75742 184578 75826 184814
rect 76062 184578 111506 184814
rect 111742 184578 111826 184814
rect 112062 184578 147506 184814
rect 147742 184578 147826 184814
rect 148062 184578 183506 184814
rect 183742 184578 183826 184814
rect 184062 184578 219506 184814
rect 219742 184578 219826 184814
rect 220062 184578 255506 184814
rect 255742 184578 255826 184814
rect 256062 184578 291506 184814
rect 291742 184578 291826 184814
rect 292062 184578 327506 184814
rect 327742 184578 327826 184814
rect 328062 184578 363506 184814
rect 363742 184578 363826 184814
rect 364062 184578 399506 184814
rect 399742 184578 399826 184814
rect 400062 184578 435506 184814
rect 435742 184578 435826 184814
rect 436062 184578 471506 184814
rect 471742 184578 471826 184814
rect 472062 184578 507506 184814
rect 507742 184578 507826 184814
rect 508062 184578 543506 184814
rect 543742 184578 543826 184814
rect 544062 184578 579506 184814
rect 579742 184578 579826 184814
rect 580062 184578 587262 184814
rect 587498 184578 587582 184814
rect 587818 184578 592650 184814
rect -8726 184546 592650 184578
rect -8726 183894 592650 183926
rect -8726 183658 -2934 183894
rect -2698 183658 -2614 183894
rect -2378 183658 2266 183894
rect 2502 183658 2586 183894
rect 2822 183658 38266 183894
rect 38502 183658 38586 183894
rect 38822 183658 74266 183894
rect 74502 183658 74586 183894
rect 74822 183658 110266 183894
rect 110502 183658 110586 183894
rect 110822 183658 146266 183894
rect 146502 183658 146586 183894
rect 146822 183658 182266 183894
rect 182502 183658 182586 183894
rect 182822 183658 218266 183894
rect 218502 183658 218586 183894
rect 218822 183658 254266 183894
rect 254502 183658 254586 183894
rect 254822 183658 290266 183894
rect 290502 183658 290586 183894
rect 290822 183658 326266 183894
rect 326502 183658 326586 183894
rect 326822 183658 362266 183894
rect 362502 183658 362586 183894
rect 362822 183658 398266 183894
rect 398502 183658 398586 183894
rect 398822 183658 434266 183894
rect 434502 183658 434586 183894
rect 434822 183658 470266 183894
rect 470502 183658 470586 183894
rect 470822 183658 506266 183894
rect 506502 183658 506586 183894
rect 506822 183658 542266 183894
rect 542502 183658 542586 183894
rect 542822 183658 578266 183894
rect 578502 183658 578586 183894
rect 578822 183658 586302 183894
rect 586538 183658 586622 183894
rect 586858 183658 592650 183894
rect -8726 183574 592650 183658
rect -8726 183338 -2934 183574
rect -2698 183338 -2614 183574
rect -2378 183338 2266 183574
rect 2502 183338 2586 183574
rect 2822 183338 38266 183574
rect 38502 183338 38586 183574
rect 38822 183338 74266 183574
rect 74502 183338 74586 183574
rect 74822 183338 110266 183574
rect 110502 183338 110586 183574
rect 110822 183338 146266 183574
rect 146502 183338 146586 183574
rect 146822 183338 182266 183574
rect 182502 183338 182586 183574
rect 182822 183338 218266 183574
rect 218502 183338 218586 183574
rect 218822 183338 254266 183574
rect 254502 183338 254586 183574
rect 254822 183338 290266 183574
rect 290502 183338 290586 183574
rect 290822 183338 326266 183574
rect 326502 183338 326586 183574
rect 326822 183338 362266 183574
rect 362502 183338 362586 183574
rect 362822 183338 398266 183574
rect 398502 183338 398586 183574
rect 398822 183338 434266 183574
rect 434502 183338 434586 183574
rect 434822 183338 470266 183574
rect 470502 183338 470586 183574
rect 470822 183338 506266 183574
rect 506502 183338 506586 183574
rect 506822 183338 542266 183574
rect 542502 183338 542586 183574
rect 542822 183338 578266 183574
rect 578502 183338 578586 183574
rect 578822 183338 586302 183574
rect 586538 183338 586622 183574
rect 586858 183338 592650 183574
rect -8726 183306 592650 183338
rect -8726 182654 592650 182686
rect -8726 182418 -1974 182654
rect -1738 182418 -1654 182654
rect -1418 182418 1026 182654
rect 1262 182418 1346 182654
rect 1582 182418 37026 182654
rect 37262 182418 37346 182654
rect 37582 182418 73026 182654
rect 73262 182418 73346 182654
rect 73582 182418 109026 182654
rect 109262 182418 109346 182654
rect 109582 182418 145026 182654
rect 145262 182418 145346 182654
rect 145582 182418 181026 182654
rect 181262 182418 181346 182654
rect 181582 182418 217026 182654
rect 217262 182418 217346 182654
rect 217582 182418 253026 182654
rect 253262 182418 253346 182654
rect 253582 182418 289026 182654
rect 289262 182418 289346 182654
rect 289582 182418 325026 182654
rect 325262 182418 325346 182654
rect 325582 182418 361026 182654
rect 361262 182418 361346 182654
rect 361582 182418 397026 182654
rect 397262 182418 397346 182654
rect 397582 182418 433026 182654
rect 433262 182418 433346 182654
rect 433582 182418 469026 182654
rect 469262 182418 469346 182654
rect 469582 182418 505026 182654
rect 505262 182418 505346 182654
rect 505582 182418 541026 182654
rect 541262 182418 541346 182654
rect 541582 182418 577026 182654
rect 577262 182418 577346 182654
rect 577582 182418 585342 182654
rect 585578 182418 585662 182654
rect 585898 182418 592650 182654
rect -8726 182334 592650 182418
rect -8726 182098 -1974 182334
rect -1738 182098 -1654 182334
rect -1418 182098 1026 182334
rect 1262 182098 1346 182334
rect 1582 182098 37026 182334
rect 37262 182098 37346 182334
rect 37582 182098 73026 182334
rect 73262 182098 73346 182334
rect 73582 182098 109026 182334
rect 109262 182098 109346 182334
rect 109582 182098 145026 182334
rect 145262 182098 145346 182334
rect 145582 182098 181026 182334
rect 181262 182098 181346 182334
rect 181582 182098 217026 182334
rect 217262 182098 217346 182334
rect 217582 182098 253026 182334
rect 253262 182098 253346 182334
rect 253582 182098 289026 182334
rect 289262 182098 289346 182334
rect 289582 182098 325026 182334
rect 325262 182098 325346 182334
rect 325582 182098 361026 182334
rect 361262 182098 361346 182334
rect 361582 182098 397026 182334
rect 397262 182098 397346 182334
rect 397582 182098 433026 182334
rect 433262 182098 433346 182334
rect 433582 182098 469026 182334
rect 469262 182098 469346 182334
rect 469582 182098 505026 182334
rect 505262 182098 505346 182334
rect 505582 182098 541026 182334
rect 541262 182098 541346 182334
rect 541582 182098 577026 182334
rect 577262 182098 577346 182334
rect 577582 182098 585342 182334
rect 585578 182098 585662 182334
rect 585898 182098 592650 182334
rect -8726 182066 592650 182098
rect -8726 155334 592650 155366
rect -8726 155098 -8694 155334
rect -8458 155098 -8374 155334
rect -8138 155098 9706 155334
rect 9942 155098 10026 155334
rect 10262 155098 45706 155334
rect 45942 155098 46026 155334
rect 46262 155098 81706 155334
rect 81942 155098 82026 155334
rect 82262 155098 117706 155334
rect 117942 155098 118026 155334
rect 118262 155098 153706 155334
rect 153942 155098 154026 155334
rect 154262 155098 189706 155334
rect 189942 155098 190026 155334
rect 190262 155098 225706 155334
rect 225942 155098 226026 155334
rect 226262 155098 261706 155334
rect 261942 155098 262026 155334
rect 262262 155098 297706 155334
rect 297942 155098 298026 155334
rect 298262 155098 333706 155334
rect 333942 155098 334026 155334
rect 334262 155098 369706 155334
rect 369942 155098 370026 155334
rect 370262 155098 405706 155334
rect 405942 155098 406026 155334
rect 406262 155098 441706 155334
rect 441942 155098 442026 155334
rect 442262 155098 477706 155334
rect 477942 155098 478026 155334
rect 478262 155098 513706 155334
rect 513942 155098 514026 155334
rect 514262 155098 549706 155334
rect 549942 155098 550026 155334
rect 550262 155098 592062 155334
rect 592298 155098 592382 155334
rect 592618 155098 592650 155334
rect -8726 155014 592650 155098
rect -8726 154778 -8694 155014
rect -8458 154778 -8374 155014
rect -8138 154778 9706 155014
rect 9942 154778 10026 155014
rect 10262 154778 45706 155014
rect 45942 154778 46026 155014
rect 46262 154778 81706 155014
rect 81942 154778 82026 155014
rect 82262 154778 117706 155014
rect 117942 154778 118026 155014
rect 118262 154778 153706 155014
rect 153942 154778 154026 155014
rect 154262 154778 189706 155014
rect 189942 154778 190026 155014
rect 190262 154778 225706 155014
rect 225942 154778 226026 155014
rect 226262 154778 261706 155014
rect 261942 154778 262026 155014
rect 262262 154778 297706 155014
rect 297942 154778 298026 155014
rect 298262 154778 333706 155014
rect 333942 154778 334026 155014
rect 334262 154778 369706 155014
rect 369942 154778 370026 155014
rect 370262 154778 405706 155014
rect 405942 154778 406026 155014
rect 406262 154778 441706 155014
rect 441942 154778 442026 155014
rect 442262 154778 477706 155014
rect 477942 154778 478026 155014
rect 478262 154778 513706 155014
rect 513942 154778 514026 155014
rect 514262 154778 549706 155014
rect 549942 154778 550026 155014
rect 550262 154778 592062 155014
rect 592298 154778 592382 155014
rect 592618 154778 592650 155014
rect -8726 154746 592650 154778
rect -8726 154094 592650 154126
rect -8726 153858 -7734 154094
rect -7498 153858 -7414 154094
rect -7178 153858 8466 154094
rect 8702 153858 8786 154094
rect 9022 153858 44466 154094
rect 44702 153858 44786 154094
rect 45022 153858 80466 154094
rect 80702 153858 80786 154094
rect 81022 153858 116466 154094
rect 116702 153858 116786 154094
rect 117022 153858 152466 154094
rect 152702 153858 152786 154094
rect 153022 153858 188466 154094
rect 188702 153858 188786 154094
rect 189022 153858 224466 154094
rect 224702 153858 224786 154094
rect 225022 153858 260466 154094
rect 260702 153858 260786 154094
rect 261022 153858 296466 154094
rect 296702 153858 296786 154094
rect 297022 153858 332466 154094
rect 332702 153858 332786 154094
rect 333022 153858 368466 154094
rect 368702 153858 368786 154094
rect 369022 153858 404466 154094
rect 404702 153858 404786 154094
rect 405022 153858 440466 154094
rect 440702 153858 440786 154094
rect 441022 153858 476466 154094
rect 476702 153858 476786 154094
rect 477022 153858 512466 154094
rect 512702 153858 512786 154094
rect 513022 153858 548466 154094
rect 548702 153858 548786 154094
rect 549022 153858 591102 154094
rect 591338 153858 591422 154094
rect 591658 153858 592650 154094
rect -8726 153774 592650 153858
rect -8726 153538 -7734 153774
rect -7498 153538 -7414 153774
rect -7178 153538 8466 153774
rect 8702 153538 8786 153774
rect 9022 153538 44466 153774
rect 44702 153538 44786 153774
rect 45022 153538 80466 153774
rect 80702 153538 80786 153774
rect 81022 153538 116466 153774
rect 116702 153538 116786 153774
rect 117022 153538 152466 153774
rect 152702 153538 152786 153774
rect 153022 153538 188466 153774
rect 188702 153538 188786 153774
rect 189022 153538 224466 153774
rect 224702 153538 224786 153774
rect 225022 153538 260466 153774
rect 260702 153538 260786 153774
rect 261022 153538 296466 153774
rect 296702 153538 296786 153774
rect 297022 153538 332466 153774
rect 332702 153538 332786 153774
rect 333022 153538 368466 153774
rect 368702 153538 368786 153774
rect 369022 153538 404466 153774
rect 404702 153538 404786 153774
rect 405022 153538 440466 153774
rect 440702 153538 440786 153774
rect 441022 153538 476466 153774
rect 476702 153538 476786 153774
rect 477022 153538 512466 153774
rect 512702 153538 512786 153774
rect 513022 153538 548466 153774
rect 548702 153538 548786 153774
rect 549022 153538 591102 153774
rect 591338 153538 591422 153774
rect 591658 153538 592650 153774
rect -8726 153506 592650 153538
rect -8726 152854 592650 152886
rect -8726 152618 -6774 152854
rect -6538 152618 -6454 152854
rect -6218 152618 7226 152854
rect 7462 152618 7546 152854
rect 7782 152618 43226 152854
rect 43462 152618 43546 152854
rect 43782 152618 79226 152854
rect 79462 152618 79546 152854
rect 79782 152618 115226 152854
rect 115462 152618 115546 152854
rect 115782 152618 151226 152854
rect 151462 152618 151546 152854
rect 151782 152618 187226 152854
rect 187462 152618 187546 152854
rect 187782 152618 223226 152854
rect 223462 152618 223546 152854
rect 223782 152618 259226 152854
rect 259462 152618 259546 152854
rect 259782 152618 295226 152854
rect 295462 152618 295546 152854
rect 295782 152618 331226 152854
rect 331462 152618 331546 152854
rect 331782 152618 367226 152854
rect 367462 152618 367546 152854
rect 367782 152618 403226 152854
rect 403462 152618 403546 152854
rect 403782 152618 439226 152854
rect 439462 152618 439546 152854
rect 439782 152618 475226 152854
rect 475462 152618 475546 152854
rect 475782 152618 511226 152854
rect 511462 152618 511546 152854
rect 511782 152618 547226 152854
rect 547462 152618 547546 152854
rect 547782 152618 590142 152854
rect 590378 152618 590462 152854
rect 590698 152618 592650 152854
rect -8726 152534 592650 152618
rect -8726 152298 -6774 152534
rect -6538 152298 -6454 152534
rect -6218 152298 7226 152534
rect 7462 152298 7546 152534
rect 7782 152298 43226 152534
rect 43462 152298 43546 152534
rect 43782 152298 79226 152534
rect 79462 152298 79546 152534
rect 79782 152298 115226 152534
rect 115462 152298 115546 152534
rect 115782 152298 151226 152534
rect 151462 152298 151546 152534
rect 151782 152298 187226 152534
rect 187462 152298 187546 152534
rect 187782 152298 223226 152534
rect 223462 152298 223546 152534
rect 223782 152298 259226 152534
rect 259462 152298 259546 152534
rect 259782 152298 295226 152534
rect 295462 152298 295546 152534
rect 295782 152298 331226 152534
rect 331462 152298 331546 152534
rect 331782 152298 367226 152534
rect 367462 152298 367546 152534
rect 367782 152298 403226 152534
rect 403462 152298 403546 152534
rect 403782 152298 439226 152534
rect 439462 152298 439546 152534
rect 439782 152298 475226 152534
rect 475462 152298 475546 152534
rect 475782 152298 511226 152534
rect 511462 152298 511546 152534
rect 511782 152298 547226 152534
rect 547462 152298 547546 152534
rect 547782 152298 590142 152534
rect 590378 152298 590462 152534
rect 590698 152298 592650 152534
rect -8726 152266 592650 152298
rect -8726 151614 592650 151646
rect -8726 151378 -5814 151614
rect -5578 151378 -5494 151614
rect -5258 151378 5986 151614
rect 6222 151378 6306 151614
rect 6542 151378 41986 151614
rect 42222 151378 42306 151614
rect 42542 151378 77986 151614
rect 78222 151378 78306 151614
rect 78542 151378 113986 151614
rect 114222 151378 114306 151614
rect 114542 151378 149986 151614
rect 150222 151378 150306 151614
rect 150542 151378 185986 151614
rect 186222 151378 186306 151614
rect 186542 151378 221986 151614
rect 222222 151378 222306 151614
rect 222542 151378 257986 151614
rect 258222 151378 258306 151614
rect 258542 151378 293986 151614
rect 294222 151378 294306 151614
rect 294542 151378 329986 151614
rect 330222 151378 330306 151614
rect 330542 151378 365986 151614
rect 366222 151378 366306 151614
rect 366542 151378 401986 151614
rect 402222 151378 402306 151614
rect 402542 151378 437986 151614
rect 438222 151378 438306 151614
rect 438542 151378 473986 151614
rect 474222 151378 474306 151614
rect 474542 151378 509986 151614
rect 510222 151378 510306 151614
rect 510542 151378 545986 151614
rect 546222 151378 546306 151614
rect 546542 151378 581986 151614
rect 582222 151378 582306 151614
rect 582542 151378 589182 151614
rect 589418 151378 589502 151614
rect 589738 151378 592650 151614
rect -8726 151294 592650 151378
rect -8726 151058 -5814 151294
rect -5578 151058 -5494 151294
rect -5258 151058 5986 151294
rect 6222 151058 6306 151294
rect 6542 151058 41986 151294
rect 42222 151058 42306 151294
rect 42542 151058 77986 151294
rect 78222 151058 78306 151294
rect 78542 151058 113986 151294
rect 114222 151058 114306 151294
rect 114542 151058 149986 151294
rect 150222 151058 150306 151294
rect 150542 151058 185986 151294
rect 186222 151058 186306 151294
rect 186542 151058 221986 151294
rect 222222 151058 222306 151294
rect 222542 151058 257986 151294
rect 258222 151058 258306 151294
rect 258542 151058 293986 151294
rect 294222 151058 294306 151294
rect 294542 151058 329986 151294
rect 330222 151058 330306 151294
rect 330542 151058 365986 151294
rect 366222 151058 366306 151294
rect 366542 151058 401986 151294
rect 402222 151058 402306 151294
rect 402542 151058 437986 151294
rect 438222 151058 438306 151294
rect 438542 151058 473986 151294
rect 474222 151058 474306 151294
rect 474542 151058 509986 151294
rect 510222 151058 510306 151294
rect 510542 151058 545986 151294
rect 546222 151058 546306 151294
rect 546542 151058 581986 151294
rect 582222 151058 582306 151294
rect 582542 151058 589182 151294
rect 589418 151058 589502 151294
rect 589738 151058 592650 151294
rect -8726 151026 592650 151058
rect -8726 150374 592650 150406
rect -8726 150138 -4854 150374
rect -4618 150138 -4534 150374
rect -4298 150138 4746 150374
rect 4982 150138 5066 150374
rect 5302 150138 40746 150374
rect 40982 150138 41066 150374
rect 41302 150138 76746 150374
rect 76982 150138 77066 150374
rect 77302 150138 112746 150374
rect 112982 150138 113066 150374
rect 113302 150138 148746 150374
rect 148982 150138 149066 150374
rect 149302 150138 184746 150374
rect 184982 150138 185066 150374
rect 185302 150138 220746 150374
rect 220982 150138 221066 150374
rect 221302 150138 256746 150374
rect 256982 150138 257066 150374
rect 257302 150138 292746 150374
rect 292982 150138 293066 150374
rect 293302 150138 328746 150374
rect 328982 150138 329066 150374
rect 329302 150138 364746 150374
rect 364982 150138 365066 150374
rect 365302 150138 400746 150374
rect 400982 150138 401066 150374
rect 401302 150138 436746 150374
rect 436982 150138 437066 150374
rect 437302 150138 472746 150374
rect 472982 150138 473066 150374
rect 473302 150138 508746 150374
rect 508982 150138 509066 150374
rect 509302 150138 544746 150374
rect 544982 150138 545066 150374
rect 545302 150138 580746 150374
rect 580982 150138 581066 150374
rect 581302 150138 588222 150374
rect 588458 150138 588542 150374
rect 588778 150138 592650 150374
rect -8726 150054 592650 150138
rect -8726 149818 -4854 150054
rect -4618 149818 -4534 150054
rect -4298 149818 4746 150054
rect 4982 149818 5066 150054
rect 5302 149818 40746 150054
rect 40982 149818 41066 150054
rect 41302 149818 76746 150054
rect 76982 149818 77066 150054
rect 77302 149818 112746 150054
rect 112982 149818 113066 150054
rect 113302 149818 148746 150054
rect 148982 149818 149066 150054
rect 149302 149818 184746 150054
rect 184982 149818 185066 150054
rect 185302 149818 220746 150054
rect 220982 149818 221066 150054
rect 221302 149818 256746 150054
rect 256982 149818 257066 150054
rect 257302 149818 292746 150054
rect 292982 149818 293066 150054
rect 293302 149818 328746 150054
rect 328982 149818 329066 150054
rect 329302 149818 364746 150054
rect 364982 149818 365066 150054
rect 365302 149818 400746 150054
rect 400982 149818 401066 150054
rect 401302 149818 436746 150054
rect 436982 149818 437066 150054
rect 437302 149818 472746 150054
rect 472982 149818 473066 150054
rect 473302 149818 508746 150054
rect 508982 149818 509066 150054
rect 509302 149818 544746 150054
rect 544982 149818 545066 150054
rect 545302 149818 580746 150054
rect 580982 149818 581066 150054
rect 581302 149818 588222 150054
rect 588458 149818 588542 150054
rect 588778 149818 592650 150054
rect -8726 149786 592650 149818
rect -8726 149134 592650 149166
rect -8726 148898 -3894 149134
rect -3658 148898 -3574 149134
rect -3338 148898 3506 149134
rect 3742 148898 3826 149134
rect 4062 148898 39506 149134
rect 39742 148898 39826 149134
rect 40062 148898 75506 149134
rect 75742 148898 75826 149134
rect 76062 148898 111506 149134
rect 111742 148898 111826 149134
rect 112062 148898 147506 149134
rect 147742 148898 147826 149134
rect 148062 148898 183506 149134
rect 183742 148898 183826 149134
rect 184062 148898 219506 149134
rect 219742 148898 219826 149134
rect 220062 148898 255506 149134
rect 255742 148898 255826 149134
rect 256062 148898 291506 149134
rect 291742 148898 291826 149134
rect 292062 148898 327506 149134
rect 327742 148898 327826 149134
rect 328062 148898 363506 149134
rect 363742 148898 363826 149134
rect 364062 148898 399506 149134
rect 399742 148898 399826 149134
rect 400062 148898 435506 149134
rect 435742 148898 435826 149134
rect 436062 148898 471506 149134
rect 471742 148898 471826 149134
rect 472062 148898 507506 149134
rect 507742 148898 507826 149134
rect 508062 148898 543506 149134
rect 543742 148898 543826 149134
rect 544062 148898 579506 149134
rect 579742 148898 579826 149134
rect 580062 148898 587262 149134
rect 587498 148898 587582 149134
rect 587818 148898 592650 149134
rect -8726 148814 592650 148898
rect -8726 148578 -3894 148814
rect -3658 148578 -3574 148814
rect -3338 148578 3506 148814
rect 3742 148578 3826 148814
rect 4062 148578 39506 148814
rect 39742 148578 39826 148814
rect 40062 148578 75506 148814
rect 75742 148578 75826 148814
rect 76062 148578 111506 148814
rect 111742 148578 111826 148814
rect 112062 148578 147506 148814
rect 147742 148578 147826 148814
rect 148062 148578 183506 148814
rect 183742 148578 183826 148814
rect 184062 148578 219506 148814
rect 219742 148578 219826 148814
rect 220062 148578 255506 148814
rect 255742 148578 255826 148814
rect 256062 148578 291506 148814
rect 291742 148578 291826 148814
rect 292062 148578 327506 148814
rect 327742 148578 327826 148814
rect 328062 148578 363506 148814
rect 363742 148578 363826 148814
rect 364062 148578 399506 148814
rect 399742 148578 399826 148814
rect 400062 148578 435506 148814
rect 435742 148578 435826 148814
rect 436062 148578 471506 148814
rect 471742 148578 471826 148814
rect 472062 148578 507506 148814
rect 507742 148578 507826 148814
rect 508062 148578 543506 148814
rect 543742 148578 543826 148814
rect 544062 148578 579506 148814
rect 579742 148578 579826 148814
rect 580062 148578 587262 148814
rect 587498 148578 587582 148814
rect 587818 148578 592650 148814
rect -8726 148546 592650 148578
rect -8726 147894 592650 147926
rect -8726 147658 -2934 147894
rect -2698 147658 -2614 147894
rect -2378 147658 2266 147894
rect 2502 147658 2586 147894
rect 2822 147658 38266 147894
rect 38502 147658 38586 147894
rect 38822 147658 74266 147894
rect 74502 147658 74586 147894
rect 74822 147658 110266 147894
rect 110502 147658 110586 147894
rect 110822 147658 146266 147894
rect 146502 147658 146586 147894
rect 146822 147658 182266 147894
rect 182502 147658 182586 147894
rect 182822 147658 218266 147894
rect 218502 147658 218586 147894
rect 218822 147658 254266 147894
rect 254502 147658 254586 147894
rect 254822 147658 290266 147894
rect 290502 147658 290586 147894
rect 290822 147658 326266 147894
rect 326502 147658 326586 147894
rect 326822 147658 362266 147894
rect 362502 147658 362586 147894
rect 362822 147658 398266 147894
rect 398502 147658 398586 147894
rect 398822 147658 434266 147894
rect 434502 147658 434586 147894
rect 434822 147658 470266 147894
rect 470502 147658 470586 147894
rect 470822 147658 506266 147894
rect 506502 147658 506586 147894
rect 506822 147658 542266 147894
rect 542502 147658 542586 147894
rect 542822 147658 578266 147894
rect 578502 147658 578586 147894
rect 578822 147658 586302 147894
rect 586538 147658 586622 147894
rect 586858 147658 592650 147894
rect -8726 147574 592650 147658
rect -8726 147338 -2934 147574
rect -2698 147338 -2614 147574
rect -2378 147338 2266 147574
rect 2502 147338 2586 147574
rect 2822 147338 38266 147574
rect 38502 147338 38586 147574
rect 38822 147338 74266 147574
rect 74502 147338 74586 147574
rect 74822 147338 110266 147574
rect 110502 147338 110586 147574
rect 110822 147338 146266 147574
rect 146502 147338 146586 147574
rect 146822 147338 182266 147574
rect 182502 147338 182586 147574
rect 182822 147338 218266 147574
rect 218502 147338 218586 147574
rect 218822 147338 254266 147574
rect 254502 147338 254586 147574
rect 254822 147338 290266 147574
rect 290502 147338 290586 147574
rect 290822 147338 326266 147574
rect 326502 147338 326586 147574
rect 326822 147338 362266 147574
rect 362502 147338 362586 147574
rect 362822 147338 398266 147574
rect 398502 147338 398586 147574
rect 398822 147338 434266 147574
rect 434502 147338 434586 147574
rect 434822 147338 470266 147574
rect 470502 147338 470586 147574
rect 470822 147338 506266 147574
rect 506502 147338 506586 147574
rect 506822 147338 542266 147574
rect 542502 147338 542586 147574
rect 542822 147338 578266 147574
rect 578502 147338 578586 147574
rect 578822 147338 586302 147574
rect 586538 147338 586622 147574
rect 586858 147338 592650 147574
rect -8726 147306 592650 147338
rect -8726 146654 592650 146686
rect -8726 146418 -1974 146654
rect -1738 146418 -1654 146654
rect -1418 146418 1026 146654
rect 1262 146418 1346 146654
rect 1582 146418 37026 146654
rect 37262 146418 37346 146654
rect 37582 146418 73026 146654
rect 73262 146418 73346 146654
rect 73582 146418 109026 146654
rect 109262 146418 109346 146654
rect 109582 146418 145026 146654
rect 145262 146418 145346 146654
rect 145582 146418 181026 146654
rect 181262 146418 181346 146654
rect 181582 146418 217026 146654
rect 217262 146418 217346 146654
rect 217582 146418 253026 146654
rect 253262 146418 253346 146654
rect 253582 146418 289026 146654
rect 289262 146418 289346 146654
rect 289582 146418 325026 146654
rect 325262 146418 325346 146654
rect 325582 146418 361026 146654
rect 361262 146418 361346 146654
rect 361582 146418 397026 146654
rect 397262 146418 397346 146654
rect 397582 146418 433026 146654
rect 433262 146418 433346 146654
rect 433582 146418 469026 146654
rect 469262 146418 469346 146654
rect 469582 146418 505026 146654
rect 505262 146418 505346 146654
rect 505582 146418 541026 146654
rect 541262 146418 541346 146654
rect 541582 146418 577026 146654
rect 577262 146418 577346 146654
rect 577582 146418 585342 146654
rect 585578 146418 585662 146654
rect 585898 146418 592650 146654
rect -8726 146334 592650 146418
rect -8726 146098 -1974 146334
rect -1738 146098 -1654 146334
rect -1418 146098 1026 146334
rect 1262 146098 1346 146334
rect 1582 146098 37026 146334
rect 37262 146098 37346 146334
rect 37582 146098 73026 146334
rect 73262 146098 73346 146334
rect 73582 146098 109026 146334
rect 109262 146098 109346 146334
rect 109582 146098 145026 146334
rect 145262 146098 145346 146334
rect 145582 146098 181026 146334
rect 181262 146098 181346 146334
rect 181582 146098 217026 146334
rect 217262 146098 217346 146334
rect 217582 146098 253026 146334
rect 253262 146098 253346 146334
rect 253582 146098 289026 146334
rect 289262 146098 289346 146334
rect 289582 146098 325026 146334
rect 325262 146098 325346 146334
rect 325582 146098 361026 146334
rect 361262 146098 361346 146334
rect 361582 146098 397026 146334
rect 397262 146098 397346 146334
rect 397582 146098 433026 146334
rect 433262 146098 433346 146334
rect 433582 146098 469026 146334
rect 469262 146098 469346 146334
rect 469582 146098 505026 146334
rect 505262 146098 505346 146334
rect 505582 146098 541026 146334
rect 541262 146098 541346 146334
rect 541582 146098 577026 146334
rect 577262 146098 577346 146334
rect 577582 146098 585342 146334
rect 585578 146098 585662 146334
rect 585898 146098 592650 146334
rect -8726 146066 592650 146098
rect -8726 119334 592650 119366
rect -8726 119098 -8694 119334
rect -8458 119098 -8374 119334
rect -8138 119098 9706 119334
rect 9942 119098 10026 119334
rect 10262 119098 45706 119334
rect 45942 119098 46026 119334
rect 46262 119098 81706 119334
rect 81942 119098 82026 119334
rect 82262 119098 117706 119334
rect 117942 119098 118026 119334
rect 118262 119098 153706 119334
rect 153942 119098 154026 119334
rect 154262 119098 189706 119334
rect 189942 119098 190026 119334
rect 190262 119098 225706 119334
rect 225942 119098 226026 119334
rect 226262 119098 261706 119334
rect 261942 119098 262026 119334
rect 262262 119098 297706 119334
rect 297942 119098 298026 119334
rect 298262 119098 333706 119334
rect 333942 119098 334026 119334
rect 334262 119098 369706 119334
rect 369942 119098 370026 119334
rect 370262 119098 405706 119334
rect 405942 119098 406026 119334
rect 406262 119098 441706 119334
rect 441942 119098 442026 119334
rect 442262 119098 477706 119334
rect 477942 119098 478026 119334
rect 478262 119098 513706 119334
rect 513942 119098 514026 119334
rect 514262 119098 549706 119334
rect 549942 119098 550026 119334
rect 550262 119098 592062 119334
rect 592298 119098 592382 119334
rect 592618 119098 592650 119334
rect -8726 119014 592650 119098
rect -8726 118778 -8694 119014
rect -8458 118778 -8374 119014
rect -8138 118778 9706 119014
rect 9942 118778 10026 119014
rect 10262 118778 45706 119014
rect 45942 118778 46026 119014
rect 46262 118778 81706 119014
rect 81942 118778 82026 119014
rect 82262 118778 117706 119014
rect 117942 118778 118026 119014
rect 118262 118778 153706 119014
rect 153942 118778 154026 119014
rect 154262 118778 189706 119014
rect 189942 118778 190026 119014
rect 190262 118778 225706 119014
rect 225942 118778 226026 119014
rect 226262 118778 261706 119014
rect 261942 118778 262026 119014
rect 262262 118778 297706 119014
rect 297942 118778 298026 119014
rect 298262 118778 333706 119014
rect 333942 118778 334026 119014
rect 334262 118778 369706 119014
rect 369942 118778 370026 119014
rect 370262 118778 405706 119014
rect 405942 118778 406026 119014
rect 406262 118778 441706 119014
rect 441942 118778 442026 119014
rect 442262 118778 477706 119014
rect 477942 118778 478026 119014
rect 478262 118778 513706 119014
rect 513942 118778 514026 119014
rect 514262 118778 549706 119014
rect 549942 118778 550026 119014
rect 550262 118778 592062 119014
rect 592298 118778 592382 119014
rect 592618 118778 592650 119014
rect -8726 118746 592650 118778
rect -8726 118094 592650 118126
rect -8726 117858 -7734 118094
rect -7498 117858 -7414 118094
rect -7178 117858 8466 118094
rect 8702 117858 8786 118094
rect 9022 117858 44466 118094
rect 44702 117858 44786 118094
rect 45022 117858 80466 118094
rect 80702 117858 80786 118094
rect 81022 117858 116466 118094
rect 116702 117858 116786 118094
rect 117022 117858 152466 118094
rect 152702 117858 152786 118094
rect 153022 117858 188466 118094
rect 188702 117858 188786 118094
rect 189022 117858 224466 118094
rect 224702 117858 224786 118094
rect 225022 117858 260466 118094
rect 260702 117858 260786 118094
rect 261022 117858 296466 118094
rect 296702 117858 296786 118094
rect 297022 117858 332466 118094
rect 332702 117858 332786 118094
rect 333022 117858 368466 118094
rect 368702 117858 368786 118094
rect 369022 117858 404466 118094
rect 404702 117858 404786 118094
rect 405022 117858 440466 118094
rect 440702 117858 440786 118094
rect 441022 117858 476466 118094
rect 476702 117858 476786 118094
rect 477022 117858 512466 118094
rect 512702 117858 512786 118094
rect 513022 117858 548466 118094
rect 548702 117858 548786 118094
rect 549022 117858 591102 118094
rect 591338 117858 591422 118094
rect 591658 117858 592650 118094
rect -8726 117774 592650 117858
rect -8726 117538 -7734 117774
rect -7498 117538 -7414 117774
rect -7178 117538 8466 117774
rect 8702 117538 8786 117774
rect 9022 117538 44466 117774
rect 44702 117538 44786 117774
rect 45022 117538 80466 117774
rect 80702 117538 80786 117774
rect 81022 117538 116466 117774
rect 116702 117538 116786 117774
rect 117022 117538 152466 117774
rect 152702 117538 152786 117774
rect 153022 117538 188466 117774
rect 188702 117538 188786 117774
rect 189022 117538 224466 117774
rect 224702 117538 224786 117774
rect 225022 117538 260466 117774
rect 260702 117538 260786 117774
rect 261022 117538 296466 117774
rect 296702 117538 296786 117774
rect 297022 117538 332466 117774
rect 332702 117538 332786 117774
rect 333022 117538 368466 117774
rect 368702 117538 368786 117774
rect 369022 117538 404466 117774
rect 404702 117538 404786 117774
rect 405022 117538 440466 117774
rect 440702 117538 440786 117774
rect 441022 117538 476466 117774
rect 476702 117538 476786 117774
rect 477022 117538 512466 117774
rect 512702 117538 512786 117774
rect 513022 117538 548466 117774
rect 548702 117538 548786 117774
rect 549022 117538 591102 117774
rect 591338 117538 591422 117774
rect 591658 117538 592650 117774
rect -8726 117506 592650 117538
rect -8726 116854 592650 116886
rect -8726 116618 -6774 116854
rect -6538 116618 -6454 116854
rect -6218 116618 7226 116854
rect 7462 116618 7546 116854
rect 7782 116618 43226 116854
rect 43462 116618 43546 116854
rect 43782 116618 79226 116854
rect 79462 116618 79546 116854
rect 79782 116618 115226 116854
rect 115462 116618 115546 116854
rect 115782 116618 151226 116854
rect 151462 116618 151546 116854
rect 151782 116618 187226 116854
rect 187462 116618 187546 116854
rect 187782 116618 223226 116854
rect 223462 116618 223546 116854
rect 223782 116618 259226 116854
rect 259462 116618 259546 116854
rect 259782 116618 295226 116854
rect 295462 116618 295546 116854
rect 295782 116618 331226 116854
rect 331462 116618 331546 116854
rect 331782 116618 367226 116854
rect 367462 116618 367546 116854
rect 367782 116618 403226 116854
rect 403462 116618 403546 116854
rect 403782 116618 439226 116854
rect 439462 116618 439546 116854
rect 439782 116618 475226 116854
rect 475462 116618 475546 116854
rect 475782 116618 511226 116854
rect 511462 116618 511546 116854
rect 511782 116618 547226 116854
rect 547462 116618 547546 116854
rect 547782 116618 590142 116854
rect 590378 116618 590462 116854
rect 590698 116618 592650 116854
rect -8726 116534 592650 116618
rect -8726 116298 -6774 116534
rect -6538 116298 -6454 116534
rect -6218 116298 7226 116534
rect 7462 116298 7546 116534
rect 7782 116298 43226 116534
rect 43462 116298 43546 116534
rect 43782 116298 79226 116534
rect 79462 116298 79546 116534
rect 79782 116298 115226 116534
rect 115462 116298 115546 116534
rect 115782 116298 151226 116534
rect 151462 116298 151546 116534
rect 151782 116298 187226 116534
rect 187462 116298 187546 116534
rect 187782 116298 223226 116534
rect 223462 116298 223546 116534
rect 223782 116298 259226 116534
rect 259462 116298 259546 116534
rect 259782 116298 295226 116534
rect 295462 116298 295546 116534
rect 295782 116298 331226 116534
rect 331462 116298 331546 116534
rect 331782 116298 367226 116534
rect 367462 116298 367546 116534
rect 367782 116298 403226 116534
rect 403462 116298 403546 116534
rect 403782 116298 439226 116534
rect 439462 116298 439546 116534
rect 439782 116298 475226 116534
rect 475462 116298 475546 116534
rect 475782 116298 511226 116534
rect 511462 116298 511546 116534
rect 511782 116298 547226 116534
rect 547462 116298 547546 116534
rect 547782 116298 590142 116534
rect 590378 116298 590462 116534
rect 590698 116298 592650 116534
rect -8726 116266 592650 116298
rect -8726 115614 592650 115646
rect -8726 115378 -5814 115614
rect -5578 115378 -5494 115614
rect -5258 115378 5986 115614
rect 6222 115378 6306 115614
rect 6542 115378 41986 115614
rect 42222 115378 42306 115614
rect 42542 115378 77986 115614
rect 78222 115378 78306 115614
rect 78542 115378 113986 115614
rect 114222 115378 114306 115614
rect 114542 115378 149986 115614
rect 150222 115378 150306 115614
rect 150542 115378 185986 115614
rect 186222 115378 186306 115614
rect 186542 115378 221986 115614
rect 222222 115378 222306 115614
rect 222542 115378 257986 115614
rect 258222 115378 258306 115614
rect 258542 115378 293986 115614
rect 294222 115378 294306 115614
rect 294542 115378 329986 115614
rect 330222 115378 330306 115614
rect 330542 115378 365986 115614
rect 366222 115378 366306 115614
rect 366542 115378 401986 115614
rect 402222 115378 402306 115614
rect 402542 115378 437986 115614
rect 438222 115378 438306 115614
rect 438542 115378 473986 115614
rect 474222 115378 474306 115614
rect 474542 115378 509986 115614
rect 510222 115378 510306 115614
rect 510542 115378 545986 115614
rect 546222 115378 546306 115614
rect 546542 115378 581986 115614
rect 582222 115378 582306 115614
rect 582542 115378 589182 115614
rect 589418 115378 589502 115614
rect 589738 115378 592650 115614
rect -8726 115294 592650 115378
rect -8726 115058 -5814 115294
rect -5578 115058 -5494 115294
rect -5258 115058 5986 115294
rect 6222 115058 6306 115294
rect 6542 115058 41986 115294
rect 42222 115058 42306 115294
rect 42542 115058 77986 115294
rect 78222 115058 78306 115294
rect 78542 115058 113986 115294
rect 114222 115058 114306 115294
rect 114542 115058 149986 115294
rect 150222 115058 150306 115294
rect 150542 115058 185986 115294
rect 186222 115058 186306 115294
rect 186542 115058 221986 115294
rect 222222 115058 222306 115294
rect 222542 115058 257986 115294
rect 258222 115058 258306 115294
rect 258542 115058 293986 115294
rect 294222 115058 294306 115294
rect 294542 115058 329986 115294
rect 330222 115058 330306 115294
rect 330542 115058 365986 115294
rect 366222 115058 366306 115294
rect 366542 115058 401986 115294
rect 402222 115058 402306 115294
rect 402542 115058 437986 115294
rect 438222 115058 438306 115294
rect 438542 115058 473986 115294
rect 474222 115058 474306 115294
rect 474542 115058 509986 115294
rect 510222 115058 510306 115294
rect 510542 115058 545986 115294
rect 546222 115058 546306 115294
rect 546542 115058 581986 115294
rect 582222 115058 582306 115294
rect 582542 115058 589182 115294
rect 589418 115058 589502 115294
rect 589738 115058 592650 115294
rect -8726 115026 592650 115058
rect -8726 114374 592650 114406
rect -8726 114138 -4854 114374
rect -4618 114138 -4534 114374
rect -4298 114138 4746 114374
rect 4982 114138 5066 114374
rect 5302 114138 40746 114374
rect 40982 114138 41066 114374
rect 41302 114138 76746 114374
rect 76982 114138 77066 114374
rect 77302 114138 112746 114374
rect 112982 114138 113066 114374
rect 113302 114138 148746 114374
rect 148982 114138 149066 114374
rect 149302 114138 184746 114374
rect 184982 114138 185066 114374
rect 185302 114138 220746 114374
rect 220982 114138 221066 114374
rect 221302 114138 256746 114374
rect 256982 114138 257066 114374
rect 257302 114138 292746 114374
rect 292982 114138 293066 114374
rect 293302 114138 328746 114374
rect 328982 114138 329066 114374
rect 329302 114138 364746 114374
rect 364982 114138 365066 114374
rect 365302 114138 400746 114374
rect 400982 114138 401066 114374
rect 401302 114138 436746 114374
rect 436982 114138 437066 114374
rect 437302 114138 472746 114374
rect 472982 114138 473066 114374
rect 473302 114138 508746 114374
rect 508982 114138 509066 114374
rect 509302 114138 544746 114374
rect 544982 114138 545066 114374
rect 545302 114138 580746 114374
rect 580982 114138 581066 114374
rect 581302 114138 588222 114374
rect 588458 114138 588542 114374
rect 588778 114138 592650 114374
rect -8726 114054 592650 114138
rect -8726 113818 -4854 114054
rect -4618 113818 -4534 114054
rect -4298 113818 4746 114054
rect 4982 113818 5066 114054
rect 5302 113818 40746 114054
rect 40982 113818 41066 114054
rect 41302 113818 76746 114054
rect 76982 113818 77066 114054
rect 77302 113818 112746 114054
rect 112982 113818 113066 114054
rect 113302 113818 148746 114054
rect 148982 113818 149066 114054
rect 149302 113818 184746 114054
rect 184982 113818 185066 114054
rect 185302 113818 220746 114054
rect 220982 113818 221066 114054
rect 221302 113818 256746 114054
rect 256982 113818 257066 114054
rect 257302 113818 292746 114054
rect 292982 113818 293066 114054
rect 293302 113818 328746 114054
rect 328982 113818 329066 114054
rect 329302 113818 364746 114054
rect 364982 113818 365066 114054
rect 365302 113818 400746 114054
rect 400982 113818 401066 114054
rect 401302 113818 436746 114054
rect 436982 113818 437066 114054
rect 437302 113818 472746 114054
rect 472982 113818 473066 114054
rect 473302 113818 508746 114054
rect 508982 113818 509066 114054
rect 509302 113818 544746 114054
rect 544982 113818 545066 114054
rect 545302 113818 580746 114054
rect 580982 113818 581066 114054
rect 581302 113818 588222 114054
rect 588458 113818 588542 114054
rect 588778 113818 592650 114054
rect -8726 113786 592650 113818
rect -8726 113134 592650 113166
rect -8726 112898 -3894 113134
rect -3658 112898 -3574 113134
rect -3338 112898 3506 113134
rect 3742 112898 3826 113134
rect 4062 112898 39506 113134
rect 39742 112898 39826 113134
rect 40062 112898 75506 113134
rect 75742 112898 75826 113134
rect 76062 112898 111506 113134
rect 111742 112898 111826 113134
rect 112062 112898 147506 113134
rect 147742 112898 147826 113134
rect 148062 112898 183506 113134
rect 183742 112898 183826 113134
rect 184062 112898 219506 113134
rect 219742 112898 219826 113134
rect 220062 112898 255506 113134
rect 255742 112898 255826 113134
rect 256062 112898 291506 113134
rect 291742 112898 291826 113134
rect 292062 112898 327506 113134
rect 327742 112898 327826 113134
rect 328062 112898 363506 113134
rect 363742 112898 363826 113134
rect 364062 112898 399506 113134
rect 399742 112898 399826 113134
rect 400062 112898 435506 113134
rect 435742 112898 435826 113134
rect 436062 112898 471506 113134
rect 471742 112898 471826 113134
rect 472062 112898 507506 113134
rect 507742 112898 507826 113134
rect 508062 112898 543506 113134
rect 543742 112898 543826 113134
rect 544062 112898 579506 113134
rect 579742 112898 579826 113134
rect 580062 112898 587262 113134
rect 587498 112898 587582 113134
rect 587818 112898 592650 113134
rect -8726 112814 592650 112898
rect -8726 112578 -3894 112814
rect -3658 112578 -3574 112814
rect -3338 112578 3506 112814
rect 3742 112578 3826 112814
rect 4062 112578 39506 112814
rect 39742 112578 39826 112814
rect 40062 112578 75506 112814
rect 75742 112578 75826 112814
rect 76062 112578 111506 112814
rect 111742 112578 111826 112814
rect 112062 112578 147506 112814
rect 147742 112578 147826 112814
rect 148062 112578 183506 112814
rect 183742 112578 183826 112814
rect 184062 112578 219506 112814
rect 219742 112578 219826 112814
rect 220062 112578 255506 112814
rect 255742 112578 255826 112814
rect 256062 112578 291506 112814
rect 291742 112578 291826 112814
rect 292062 112578 327506 112814
rect 327742 112578 327826 112814
rect 328062 112578 363506 112814
rect 363742 112578 363826 112814
rect 364062 112578 399506 112814
rect 399742 112578 399826 112814
rect 400062 112578 435506 112814
rect 435742 112578 435826 112814
rect 436062 112578 471506 112814
rect 471742 112578 471826 112814
rect 472062 112578 507506 112814
rect 507742 112578 507826 112814
rect 508062 112578 543506 112814
rect 543742 112578 543826 112814
rect 544062 112578 579506 112814
rect 579742 112578 579826 112814
rect 580062 112578 587262 112814
rect 587498 112578 587582 112814
rect 587818 112578 592650 112814
rect -8726 112546 592650 112578
rect -8726 111894 592650 111926
rect -8726 111658 -2934 111894
rect -2698 111658 -2614 111894
rect -2378 111658 2266 111894
rect 2502 111658 2586 111894
rect 2822 111658 38266 111894
rect 38502 111658 38586 111894
rect 38822 111658 74266 111894
rect 74502 111658 74586 111894
rect 74822 111658 110266 111894
rect 110502 111658 110586 111894
rect 110822 111658 146266 111894
rect 146502 111658 146586 111894
rect 146822 111658 182266 111894
rect 182502 111658 182586 111894
rect 182822 111658 218266 111894
rect 218502 111658 218586 111894
rect 218822 111658 254266 111894
rect 254502 111658 254586 111894
rect 254822 111658 290266 111894
rect 290502 111658 290586 111894
rect 290822 111658 326266 111894
rect 326502 111658 326586 111894
rect 326822 111658 362266 111894
rect 362502 111658 362586 111894
rect 362822 111658 398266 111894
rect 398502 111658 398586 111894
rect 398822 111658 434266 111894
rect 434502 111658 434586 111894
rect 434822 111658 470266 111894
rect 470502 111658 470586 111894
rect 470822 111658 506266 111894
rect 506502 111658 506586 111894
rect 506822 111658 542266 111894
rect 542502 111658 542586 111894
rect 542822 111658 578266 111894
rect 578502 111658 578586 111894
rect 578822 111658 586302 111894
rect 586538 111658 586622 111894
rect 586858 111658 592650 111894
rect -8726 111574 592650 111658
rect -8726 111338 -2934 111574
rect -2698 111338 -2614 111574
rect -2378 111338 2266 111574
rect 2502 111338 2586 111574
rect 2822 111338 38266 111574
rect 38502 111338 38586 111574
rect 38822 111338 74266 111574
rect 74502 111338 74586 111574
rect 74822 111338 110266 111574
rect 110502 111338 110586 111574
rect 110822 111338 146266 111574
rect 146502 111338 146586 111574
rect 146822 111338 182266 111574
rect 182502 111338 182586 111574
rect 182822 111338 218266 111574
rect 218502 111338 218586 111574
rect 218822 111338 254266 111574
rect 254502 111338 254586 111574
rect 254822 111338 290266 111574
rect 290502 111338 290586 111574
rect 290822 111338 326266 111574
rect 326502 111338 326586 111574
rect 326822 111338 362266 111574
rect 362502 111338 362586 111574
rect 362822 111338 398266 111574
rect 398502 111338 398586 111574
rect 398822 111338 434266 111574
rect 434502 111338 434586 111574
rect 434822 111338 470266 111574
rect 470502 111338 470586 111574
rect 470822 111338 506266 111574
rect 506502 111338 506586 111574
rect 506822 111338 542266 111574
rect 542502 111338 542586 111574
rect 542822 111338 578266 111574
rect 578502 111338 578586 111574
rect 578822 111338 586302 111574
rect 586538 111338 586622 111574
rect 586858 111338 592650 111574
rect -8726 111306 592650 111338
rect -8726 110654 592650 110686
rect -8726 110418 -1974 110654
rect -1738 110418 -1654 110654
rect -1418 110418 1026 110654
rect 1262 110418 1346 110654
rect 1582 110418 37026 110654
rect 37262 110418 37346 110654
rect 37582 110418 73026 110654
rect 73262 110418 73346 110654
rect 73582 110418 109026 110654
rect 109262 110418 109346 110654
rect 109582 110418 145026 110654
rect 145262 110418 145346 110654
rect 145582 110418 181026 110654
rect 181262 110418 181346 110654
rect 181582 110418 217026 110654
rect 217262 110418 217346 110654
rect 217582 110418 253026 110654
rect 253262 110418 253346 110654
rect 253582 110418 289026 110654
rect 289262 110418 289346 110654
rect 289582 110418 325026 110654
rect 325262 110418 325346 110654
rect 325582 110418 361026 110654
rect 361262 110418 361346 110654
rect 361582 110418 397026 110654
rect 397262 110418 397346 110654
rect 397582 110418 433026 110654
rect 433262 110418 433346 110654
rect 433582 110418 469026 110654
rect 469262 110418 469346 110654
rect 469582 110418 505026 110654
rect 505262 110418 505346 110654
rect 505582 110418 541026 110654
rect 541262 110418 541346 110654
rect 541582 110418 577026 110654
rect 577262 110418 577346 110654
rect 577582 110418 585342 110654
rect 585578 110418 585662 110654
rect 585898 110418 592650 110654
rect -8726 110334 592650 110418
rect -8726 110098 -1974 110334
rect -1738 110098 -1654 110334
rect -1418 110098 1026 110334
rect 1262 110098 1346 110334
rect 1582 110098 37026 110334
rect 37262 110098 37346 110334
rect 37582 110098 73026 110334
rect 73262 110098 73346 110334
rect 73582 110098 109026 110334
rect 109262 110098 109346 110334
rect 109582 110098 145026 110334
rect 145262 110098 145346 110334
rect 145582 110098 181026 110334
rect 181262 110098 181346 110334
rect 181582 110098 217026 110334
rect 217262 110098 217346 110334
rect 217582 110098 253026 110334
rect 253262 110098 253346 110334
rect 253582 110098 289026 110334
rect 289262 110098 289346 110334
rect 289582 110098 325026 110334
rect 325262 110098 325346 110334
rect 325582 110098 361026 110334
rect 361262 110098 361346 110334
rect 361582 110098 397026 110334
rect 397262 110098 397346 110334
rect 397582 110098 433026 110334
rect 433262 110098 433346 110334
rect 433582 110098 469026 110334
rect 469262 110098 469346 110334
rect 469582 110098 505026 110334
rect 505262 110098 505346 110334
rect 505582 110098 541026 110334
rect 541262 110098 541346 110334
rect 541582 110098 577026 110334
rect 577262 110098 577346 110334
rect 577582 110098 585342 110334
rect 585578 110098 585662 110334
rect 585898 110098 592650 110334
rect -8726 110066 592650 110098
rect -8726 83334 592650 83366
rect -8726 83098 -8694 83334
rect -8458 83098 -8374 83334
rect -8138 83098 9706 83334
rect 9942 83098 10026 83334
rect 10262 83098 45706 83334
rect 45942 83098 46026 83334
rect 46262 83098 81706 83334
rect 81942 83098 82026 83334
rect 82262 83098 117706 83334
rect 117942 83098 118026 83334
rect 118262 83098 153706 83334
rect 153942 83098 154026 83334
rect 154262 83098 189706 83334
rect 189942 83098 190026 83334
rect 190262 83098 225706 83334
rect 225942 83098 226026 83334
rect 226262 83098 261706 83334
rect 261942 83098 262026 83334
rect 262262 83098 297706 83334
rect 297942 83098 298026 83334
rect 298262 83098 333706 83334
rect 333942 83098 334026 83334
rect 334262 83098 369706 83334
rect 369942 83098 370026 83334
rect 370262 83098 405706 83334
rect 405942 83098 406026 83334
rect 406262 83098 441706 83334
rect 441942 83098 442026 83334
rect 442262 83098 477706 83334
rect 477942 83098 478026 83334
rect 478262 83098 513706 83334
rect 513942 83098 514026 83334
rect 514262 83098 549706 83334
rect 549942 83098 550026 83334
rect 550262 83098 592062 83334
rect 592298 83098 592382 83334
rect 592618 83098 592650 83334
rect -8726 83014 592650 83098
rect -8726 82778 -8694 83014
rect -8458 82778 -8374 83014
rect -8138 82778 9706 83014
rect 9942 82778 10026 83014
rect 10262 82778 45706 83014
rect 45942 82778 46026 83014
rect 46262 82778 81706 83014
rect 81942 82778 82026 83014
rect 82262 82778 117706 83014
rect 117942 82778 118026 83014
rect 118262 82778 153706 83014
rect 153942 82778 154026 83014
rect 154262 82778 189706 83014
rect 189942 82778 190026 83014
rect 190262 82778 225706 83014
rect 225942 82778 226026 83014
rect 226262 82778 261706 83014
rect 261942 82778 262026 83014
rect 262262 82778 297706 83014
rect 297942 82778 298026 83014
rect 298262 82778 333706 83014
rect 333942 82778 334026 83014
rect 334262 82778 369706 83014
rect 369942 82778 370026 83014
rect 370262 82778 405706 83014
rect 405942 82778 406026 83014
rect 406262 82778 441706 83014
rect 441942 82778 442026 83014
rect 442262 82778 477706 83014
rect 477942 82778 478026 83014
rect 478262 82778 513706 83014
rect 513942 82778 514026 83014
rect 514262 82778 549706 83014
rect 549942 82778 550026 83014
rect 550262 82778 592062 83014
rect 592298 82778 592382 83014
rect 592618 82778 592650 83014
rect -8726 82746 592650 82778
rect -8726 82094 592650 82126
rect -8726 81858 -7734 82094
rect -7498 81858 -7414 82094
rect -7178 81858 8466 82094
rect 8702 81858 8786 82094
rect 9022 81858 44466 82094
rect 44702 81858 44786 82094
rect 45022 81858 80466 82094
rect 80702 81858 80786 82094
rect 81022 81858 116466 82094
rect 116702 81858 116786 82094
rect 117022 81858 152466 82094
rect 152702 81858 152786 82094
rect 153022 81858 188466 82094
rect 188702 81858 188786 82094
rect 189022 81858 224466 82094
rect 224702 81858 224786 82094
rect 225022 81858 260466 82094
rect 260702 81858 260786 82094
rect 261022 81858 296466 82094
rect 296702 81858 296786 82094
rect 297022 81858 332466 82094
rect 332702 81858 332786 82094
rect 333022 81858 368466 82094
rect 368702 81858 368786 82094
rect 369022 81858 404466 82094
rect 404702 81858 404786 82094
rect 405022 81858 440466 82094
rect 440702 81858 440786 82094
rect 441022 81858 476466 82094
rect 476702 81858 476786 82094
rect 477022 81858 512466 82094
rect 512702 81858 512786 82094
rect 513022 81858 548466 82094
rect 548702 81858 548786 82094
rect 549022 81858 591102 82094
rect 591338 81858 591422 82094
rect 591658 81858 592650 82094
rect -8726 81774 592650 81858
rect -8726 81538 -7734 81774
rect -7498 81538 -7414 81774
rect -7178 81538 8466 81774
rect 8702 81538 8786 81774
rect 9022 81538 44466 81774
rect 44702 81538 44786 81774
rect 45022 81538 80466 81774
rect 80702 81538 80786 81774
rect 81022 81538 116466 81774
rect 116702 81538 116786 81774
rect 117022 81538 152466 81774
rect 152702 81538 152786 81774
rect 153022 81538 188466 81774
rect 188702 81538 188786 81774
rect 189022 81538 224466 81774
rect 224702 81538 224786 81774
rect 225022 81538 260466 81774
rect 260702 81538 260786 81774
rect 261022 81538 296466 81774
rect 296702 81538 296786 81774
rect 297022 81538 332466 81774
rect 332702 81538 332786 81774
rect 333022 81538 368466 81774
rect 368702 81538 368786 81774
rect 369022 81538 404466 81774
rect 404702 81538 404786 81774
rect 405022 81538 440466 81774
rect 440702 81538 440786 81774
rect 441022 81538 476466 81774
rect 476702 81538 476786 81774
rect 477022 81538 512466 81774
rect 512702 81538 512786 81774
rect 513022 81538 548466 81774
rect 548702 81538 548786 81774
rect 549022 81538 591102 81774
rect 591338 81538 591422 81774
rect 591658 81538 592650 81774
rect -8726 81506 592650 81538
rect -8726 80854 592650 80886
rect -8726 80618 -6774 80854
rect -6538 80618 -6454 80854
rect -6218 80618 7226 80854
rect 7462 80618 7546 80854
rect 7782 80618 43226 80854
rect 43462 80618 43546 80854
rect 43782 80618 79226 80854
rect 79462 80618 79546 80854
rect 79782 80618 115226 80854
rect 115462 80618 115546 80854
rect 115782 80618 151226 80854
rect 151462 80618 151546 80854
rect 151782 80618 187226 80854
rect 187462 80618 187546 80854
rect 187782 80618 223226 80854
rect 223462 80618 223546 80854
rect 223782 80618 259226 80854
rect 259462 80618 259546 80854
rect 259782 80618 295226 80854
rect 295462 80618 295546 80854
rect 295782 80618 331226 80854
rect 331462 80618 331546 80854
rect 331782 80618 367226 80854
rect 367462 80618 367546 80854
rect 367782 80618 403226 80854
rect 403462 80618 403546 80854
rect 403782 80618 439226 80854
rect 439462 80618 439546 80854
rect 439782 80618 475226 80854
rect 475462 80618 475546 80854
rect 475782 80618 511226 80854
rect 511462 80618 511546 80854
rect 511782 80618 547226 80854
rect 547462 80618 547546 80854
rect 547782 80618 590142 80854
rect 590378 80618 590462 80854
rect 590698 80618 592650 80854
rect -8726 80534 592650 80618
rect -8726 80298 -6774 80534
rect -6538 80298 -6454 80534
rect -6218 80298 7226 80534
rect 7462 80298 7546 80534
rect 7782 80298 43226 80534
rect 43462 80298 43546 80534
rect 43782 80298 79226 80534
rect 79462 80298 79546 80534
rect 79782 80298 115226 80534
rect 115462 80298 115546 80534
rect 115782 80298 151226 80534
rect 151462 80298 151546 80534
rect 151782 80298 187226 80534
rect 187462 80298 187546 80534
rect 187782 80298 223226 80534
rect 223462 80298 223546 80534
rect 223782 80298 259226 80534
rect 259462 80298 259546 80534
rect 259782 80298 295226 80534
rect 295462 80298 295546 80534
rect 295782 80298 331226 80534
rect 331462 80298 331546 80534
rect 331782 80298 367226 80534
rect 367462 80298 367546 80534
rect 367782 80298 403226 80534
rect 403462 80298 403546 80534
rect 403782 80298 439226 80534
rect 439462 80298 439546 80534
rect 439782 80298 475226 80534
rect 475462 80298 475546 80534
rect 475782 80298 511226 80534
rect 511462 80298 511546 80534
rect 511782 80298 547226 80534
rect 547462 80298 547546 80534
rect 547782 80298 590142 80534
rect 590378 80298 590462 80534
rect 590698 80298 592650 80534
rect -8726 80266 592650 80298
rect -8726 79614 592650 79646
rect -8726 79378 -5814 79614
rect -5578 79378 -5494 79614
rect -5258 79378 5986 79614
rect 6222 79378 6306 79614
rect 6542 79378 41986 79614
rect 42222 79378 42306 79614
rect 42542 79378 77986 79614
rect 78222 79378 78306 79614
rect 78542 79378 113986 79614
rect 114222 79378 114306 79614
rect 114542 79378 149986 79614
rect 150222 79378 150306 79614
rect 150542 79378 185986 79614
rect 186222 79378 186306 79614
rect 186542 79378 221986 79614
rect 222222 79378 222306 79614
rect 222542 79378 257986 79614
rect 258222 79378 258306 79614
rect 258542 79378 293986 79614
rect 294222 79378 294306 79614
rect 294542 79378 329986 79614
rect 330222 79378 330306 79614
rect 330542 79378 365986 79614
rect 366222 79378 366306 79614
rect 366542 79378 401986 79614
rect 402222 79378 402306 79614
rect 402542 79378 437986 79614
rect 438222 79378 438306 79614
rect 438542 79378 473986 79614
rect 474222 79378 474306 79614
rect 474542 79378 509986 79614
rect 510222 79378 510306 79614
rect 510542 79378 545986 79614
rect 546222 79378 546306 79614
rect 546542 79378 581986 79614
rect 582222 79378 582306 79614
rect 582542 79378 589182 79614
rect 589418 79378 589502 79614
rect 589738 79378 592650 79614
rect -8726 79294 592650 79378
rect -8726 79058 -5814 79294
rect -5578 79058 -5494 79294
rect -5258 79058 5986 79294
rect 6222 79058 6306 79294
rect 6542 79058 41986 79294
rect 42222 79058 42306 79294
rect 42542 79058 77986 79294
rect 78222 79058 78306 79294
rect 78542 79058 113986 79294
rect 114222 79058 114306 79294
rect 114542 79058 149986 79294
rect 150222 79058 150306 79294
rect 150542 79058 185986 79294
rect 186222 79058 186306 79294
rect 186542 79058 221986 79294
rect 222222 79058 222306 79294
rect 222542 79058 257986 79294
rect 258222 79058 258306 79294
rect 258542 79058 293986 79294
rect 294222 79058 294306 79294
rect 294542 79058 329986 79294
rect 330222 79058 330306 79294
rect 330542 79058 365986 79294
rect 366222 79058 366306 79294
rect 366542 79058 401986 79294
rect 402222 79058 402306 79294
rect 402542 79058 437986 79294
rect 438222 79058 438306 79294
rect 438542 79058 473986 79294
rect 474222 79058 474306 79294
rect 474542 79058 509986 79294
rect 510222 79058 510306 79294
rect 510542 79058 545986 79294
rect 546222 79058 546306 79294
rect 546542 79058 581986 79294
rect 582222 79058 582306 79294
rect 582542 79058 589182 79294
rect 589418 79058 589502 79294
rect 589738 79058 592650 79294
rect -8726 79026 592650 79058
rect -8726 78374 592650 78406
rect -8726 78138 -4854 78374
rect -4618 78138 -4534 78374
rect -4298 78138 4746 78374
rect 4982 78138 5066 78374
rect 5302 78138 40746 78374
rect 40982 78138 41066 78374
rect 41302 78138 76746 78374
rect 76982 78138 77066 78374
rect 77302 78138 112746 78374
rect 112982 78138 113066 78374
rect 113302 78138 148746 78374
rect 148982 78138 149066 78374
rect 149302 78138 184746 78374
rect 184982 78138 185066 78374
rect 185302 78138 220746 78374
rect 220982 78138 221066 78374
rect 221302 78138 256746 78374
rect 256982 78138 257066 78374
rect 257302 78138 292746 78374
rect 292982 78138 293066 78374
rect 293302 78138 328746 78374
rect 328982 78138 329066 78374
rect 329302 78138 364746 78374
rect 364982 78138 365066 78374
rect 365302 78138 400746 78374
rect 400982 78138 401066 78374
rect 401302 78138 436746 78374
rect 436982 78138 437066 78374
rect 437302 78138 472746 78374
rect 472982 78138 473066 78374
rect 473302 78138 508746 78374
rect 508982 78138 509066 78374
rect 509302 78138 544746 78374
rect 544982 78138 545066 78374
rect 545302 78138 580746 78374
rect 580982 78138 581066 78374
rect 581302 78138 588222 78374
rect 588458 78138 588542 78374
rect 588778 78138 592650 78374
rect -8726 78054 592650 78138
rect -8726 77818 -4854 78054
rect -4618 77818 -4534 78054
rect -4298 77818 4746 78054
rect 4982 77818 5066 78054
rect 5302 77818 40746 78054
rect 40982 77818 41066 78054
rect 41302 77818 76746 78054
rect 76982 77818 77066 78054
rect 77302 77818 112746 78054
rect 112982 77818 113066 78054
rect 113302 77818 148746 78054
rect 148982 77818 149066 78054
rect 149302 77818 184746 78054
rect 184982 77818 185066 78054
rect 185302 77818 220746 78054
rect 220982 77818 221066 78054
rect 221302 77818 256746 78054
rect 256982 77818 257066 78054
rect 257302 77818 292746 78054
rect 292982 77818 293066 78054
rect 293302 77818 328746 78054
rect 328982 77818 329066 78054
rect 329302 77818 364746 78054
rect 364982 77818 365066 78054
rect 365302 77818 400746 78054
rect 400982 77818 401066 78054
rect 401302 77818 436746 78054
rect 436982 77818 437066 78054
rect 437302 77818 472746 78054
rect 472982 77818 473066 78054
rect 473302 77818 508746 78054
rect 508982 77818 509066 78054
rect 509302 77818 544746 78054
rect 544982 77818 545066 78054
rect 545302 77818 580746 78054
rect 580982 77818 581066 78054
rect 581302 77818 588222 78054
rect 588458 77818 588542 78054
rect 588778 77818 592650 78054
rect -8726 77786 592650 77818
rect -8726 77134 592650 77166
rect -8726 76898 -3894 77134
rect -3658 76898 -3574 77134
rect -3338 76898 3506 77134
rect 3742 76898 3826 77134
rect 4062 76898 39506 77134
rect 39742 76898 39826 77134
rect 40062 76898 75506 77134
rect 75742 76898 75826 77134
rect 76062 76898 111506 77134
rect 111742 76898 111826 77134
rect 112062 76898 147506 77134
rect 147742 76898 147826 77134
rect 148062 76898 183506 77134
rect 183742 76898 183826 77134
rect 184062 76898 219506 77134
rect 219742 76898 219826 77134
rect 220062 76898 255506 77134
rect 255742 76898 255826 77134
rect 256062 76898 291506 77134
rect 291742 76898 291826 77134
rect 292062 76898 327506 77134
rect 327742 76898 327826 77134
rect 328062 76898 363506 77134
rect 363742 76898 363826 77134
rect 364062 76898 399506 77134
rect 399742 76898 399826 77134
rect 400062 76898 435506 77134
rect 435742 76898 435826 77134
rect 436062 76898 471506 77134
rect 471742 76898 471826 77134
rect 472062 76898 507506 77134
rect 507742 76898 507826 77134
rect 508062 76898 543506 77134
rect 543742 76898 543826 77134
rect 544062 76898 579506 77134
rect 579742 76898 579826 77134
rect 580062 76898 587262 77134
rect 587498 76898 587582 77134
rect 587818 76898 592650 77134
rect -8726 76814 592650 76898
rect -8726 76578 -3894 76814
rect -3658 76578 -3574 76814
rect -3338 76578 3506 76814
rect 3742 76578 3826 76814
rect 4062 76578 39506 76814
rect 39742 76578 39826 76814
rect 40062 76578 75506 76814
rect 75742 76578 75826 76814
rect 76062 76578 111506 76814
rect 111742 76578 111826 76814
rect 112062 76578 147506 76814
rect 147742 76578 147826 76814
rect 148062 76578 183506 76814
rect 183742 76578 183826 76814
rect 184062 76578 219506 76814
rect 219742 76578 219826 76814
rect 220062 76578 255506 76814
rect 255742 76578 255826 76814
rect 256062 76578 291506 76814
rect 291742 76578 291826 76814
rect 292062 76578 327506 76814
rect 327742 76578 327826 76814
rect 328062 76578 363506 76814
rect 363742 76578 363826 76814
rect 364062 76578 399506 76814
rect 399742 76578 399826 76814
rect 400062 76578 435506 76814
rect 435742 76578 435826 76814
rect 436062 76578 471506 76814
rect 471742 76578 471826 76814
rect 472062 76578 507506 76814
rect 507742 76578 507826 76814
rect 508062 76578 543506 76814
rect 543742 76578 543826 76814
rect 544062 76578 579506 76814
rect 579742 76578 579826 76814
rect 580062 76578 587262 76814
rect 587498 76578 587582 76814
rect 587818 76578 592650 76814
rect -8726 76546 592650 76578
rect -8726 75894 592650 75926
rect -8726 75658 -2934 75894
rect -2698 75658 -2614 75894
rect -2378 75658 2266 75894
rect 2502 75658 2586 75894
rect 2822 75658 38266 75894
rect 38502 75658 38586 75894
rect 38822 75658 74266 75894
rect 74502 75658 74586 75894
rect 74822 75658 110266 75894
rect 110502 75658 110586 75894
rect 110822 75658 146266 75894
rect 146502 75658 146586 75894
rect 146822 75658 182266 75894
rect 182502 75658 182586 75894
rect 182822 75658 218266 75894
rect 218502 75658 218586 75894
rect 218822 75658 254266 75894
rect 254502 75658 254586 75894
rect 254822 75658 290266 75894
rect 290502 75658 290586 75894
rect 290822 75658 326266 75894
rect 326502 75658 326586 75894
rect 326822 75658 362266 75894
rect 362502 75658 362586 75894
rect 362822 75658 398266 75894
rect 398502 75658 398586 75894
rect 398822 75658 434266 75894
rect 434502 75658 434586 75894
rect 434822 75658 470266 75894
rect 470502 75658 470586 75894
rect 470822 75658 506266 75894
rect 506502 75658 506586 75894
rect 506822 75658 542266 75894
rect 542502 75658 542586 75894
rect 542822 75658 578266 75894
rect 578502 75658 578586 75894
rect 578822 75658 586302 75894
rect 586538 75658 586622 75894
rect 586858 75658 592650 75894
rect -8726 75574 592650 75658
rect -8726 75338 -2934 75574
rect -2698 75338 -2614 75574
rect -2378 75338 2266 75574
rect 2502 75338 2586 75574
rect 2822 75338 38266 75574
rect 38502 75338 38586 75574
rect 38822 75338 74266 75574
rect 74502 75338 74586 75574
rect 74822 75338 110266 75574
rect 110502 75338 110586 75574
rect 110822 75338 146266 75574
rect 146502 75338 146586 75574
rect 146822 75338 182266 75574
rect 182502 75338 182586 75574
rect 182822 75338 218266 75574
rect 218502 75338 218586 75574
rect 218822 75338 254266 75574
rect 254502 75338 254586 75574
rect 254822 75338 290266 75574
rect 290502 75338 290586 75574
rect 290822 75338 326266 75574
rect 326502 75338 326586 75574
rect 326822 75338 362266 75574
rect 362502 75338 362586 75574
rect 362822 75338 398266 75574
rect 398502 75338 398586 75574
rect 398822 75338 434266 75574
rect 434502 75338 434586 75574
rect 434822 75338 470266 75574
rect 470502 75338 470586 75574
rect 470822 75338 506266 75574
rect 506502 75338 506586 75574
rect 506822 75338 542266 75574
rect 542502 75338 542586 75574
rect 542822 75338 578266 75574
rect 578502 75338 578586 75574
rect 578822 75338 586302 75574
rect 586538 75338 586622 75574
rect 586858 75338 592650 75574
rect -8726 75306 592650 75338
rect -8726 74654 592650 74686
rect -8726 74418 -1974 74654
rect -1738 74418 -1654 74654
rect -1418 74418 1026 74654
rect 1262 74418 1346 74654
rect 1582 74418 37026 74654
rect 37262 74418 37346 74654
rect 37582 74418 73026 74654
rect 73262 74418 73346 74654
rect 73582 74418 109026 74654
rect 109262 74418 109346 74654
rect 109582 74418 145026 74654
rect 145262 74418 145346 74654
rect 145582 74418 181026 74654
rect 181262 74418 181346 74654
rect 181582 74418 217026 74654
rect 217262 74418 217346 74654
rect 217582 74418 253026 74654
rect 253262 74418 253346 74654
rect 253582 74418 289026 74654
rect 289262 74418 289346 74654
rect 289582 74418 325026 74654
rect 325262 74418 325346 74654
rect 325582 74418 361026 74654
rect 361262 74418 361346 74654
rect 361582 74418 397026 74654
rect 397262 74418 397346 74654
rect 397582 74418 433026 74654
rect 433262 74418 433346 74654
rect 433582 74418 469026 74654
rect 469262 74418 469346 74654
rect 469582 74418 505026 74654
rect 505262 74418 505346 74654
rect 505582 74418 541026 74654
rect 541262 74418 541346 74654
rect 541582 74418 577026 74654
rect 577262 74418 577346 74654
rect 577582 74418 585342 74654
rect 585578 74418 585662 74654
rect 585898 74418 592650 74654
rect -8726 74334 592650 74418
rect -8726 74098 -1974 74334
rect -1738 74098 -1654 74334
rect -1418 74098 1026 74334
rect 1262 74098 1346 74334
rect 1582 74098 37026 74334
rect 37262 74098 37346 74334
rect 37582 74098 73026 74334
rect 73262 74098 73346 74334
rect 73582 74098 109026 74334
rect 109262 74098 109346 74334
rect 109582 74098 145026 74334
rect 145262 74098 145346 74334
rect 145582 74098 181026 74334
rect 181262 74098 181346 74334
rect 181582 74098 217026 74334
rect 217262 74098 217346 74334
rect 217582 74098 253026 74334
rect 253262 74098 253346 74334
rect 253582 74098 289026 74334
rect 289262 74098 289346 74334
rect 289582 74098 325026 74334
rect 325262 74098 325346 74334
rect 325582 74098 361026 74334
rect 361262 74098 361346 74334
rect 361582 74098 397026 74334
rect 397262 74098 397346 74334
rect 397582 74098 433026 74334
rect 433262 74098 433346 74334
rect 433582 74098 469026 74334
rect 469262 74098 469346 74334
rect 469582 74098 505026 74334
rect 505262 74098 505346 74334
rect 505582 74098 541026 74334
rect 541262 74098 541346 74334
rect 541582 74098 577026 74334
rect 577262 74098 577346 74334
rect 577582 74098 585342 74334
rect 585578 74098 585662 74334
rect 585898 74098 592650 74334
rect -8726 74066 592650 74098
rect -8726 47334 592650 47366
rect -8726 47098 -8694 47334
rect -8458 47098 -8374 47334
rect -8138 47098 9706 47334
rect 9942 47098 10026 47334
rect 10262 47098 45706 47334
rect 45942 47098 46026 47334
rect 46262 47098 81706 47334
rect 81942 47098 82026 47334
rect 82262 47098 117706 47334
rect 117942 47098 118026 47334
rect 118262 47098 153706 47334
rect 153942 47098 154026 47334
rect 154262 47098 189706 47334
rect 189942 47098 190026 47334
rect 190262 47098 225706 47334
rect 225942 47098 226026 47334
rect 226262 47098 261706 47334
rect 261942 47098 262026 47334
rect 262262 47098 297706 47334
rect 297942 47098 298026 47334
rect 298262 47098 333706 47334
rect 333942 47098 334026 47334
rect 334262 47098 369706 47334
rect 369942 47098 370026 47334
rect 370262 47098 405706 47334
rect 405942 47098 406026 47334
rect 406262 47098 441706 47334
rect 441942 47098 442026 47334
rect 442262 47098 477706 47334
rect 477942 47098 478026 47334
rect 478262 47098 513706 47334
rect 513942 47098 514026 47334
rect 514262 47098 549706 47334
rect 549942 47098 550026 47334
rect 550262 47098 592062 47334
rect 592298 47098 592382 47334
rect 592618 47098 592650 47334
rect -8726 47014 592650 47098
rect -8726 46778 -8694 47014
rect -8458 46778 -8374 47014
rect -8138 46778 9706 47014
rect 9942 46778 10026 47014
rect 10262 46778 45706 47014
rect 45942 46778 46026 47014
rect 46262 46778 81706 47014
rect 81942 46778 82026 47014
rect 82262 46778 117706 47014
rect 117942 46778 118026 47014
rect 118262 46778 153706 47014
rect 153942 46778 154026 47014
rect 154262 46778 189706 47014
rect 189942 46778 190026 47014
rect 190262 46778 225706 47014
rect 225942 46778 226026 47014
rect 226262 46778 261706 47014
rect 261942 46778 262026 47014
rect 262262 46778 297706 47014
rect 297942 46778 298026 47014
rect 298262 46778 333706 47014
rect 333942 46778 334026 47014
rect 334262 46778 369706 47014
rect 369942 46778 370026 47014
rect 370262 46778 405706 47014
rect 405942 46778 406026 47014
rect 406262 46778 441706 47014
rect 441942 46778 442026 47014
rect 442262 46778 477706 47014
rect 477942 46778 478026 47014
rect 478262 46778 513706 47014
rect 513942 46778 514026 47014
rect 514262 46778 549706 47014
rect 549942 46778 550026 47014
rect 550262 46778 592062 47014
rect 592298 46778 592382 47014
rect 592618 46778 592650 47014
rect -8726 46746 592650 46778
rect -8726 46094 592650 46126
rect -8726 45858 -7734 46094
rect -7498 45858 -7414 46094
rect -7178 45858 8466 46094
rect 8702 45858 8786 46094
rect 9022 45858 44466 46094
rect 44702 45858 44786 46094
rect 45022 45858 80466 46094
rect 80702 45858 80786 46094
rect 81022 45858 116466 46094
rect 116702 45858 116786 46094
rect 117022 45858 152466 46094
rect 152702 45858 152786 46094
rect 153022 45858 188466 46094
rect 188702 45858 188786 46094
rect 189022 45858 224466 46094
rect 224702 45858 224786 46094
rect 225022 45858 260466 46094
rect 260702 45858 260786 46094
rect 261022 45858 296466 46094
rect 296702 45858 296786 46094
rect 297022 45858 332466 46094
rect 332702 45858 332786 46094
rect 333022 45858 368466 46094
rect 368702 45858 368786 46094
rect 369022 45858 404466 46094
rect 404702 45858 404786 46094
rect 405022 45858 440466 46094
rect 440702 45858 440786 46094
rect 441022 45858 476466 46094
rect 476702 45858 476786 46094
rect 477022 45858 512466 46094
rect 512702 45858 512786 46094
rect 513022 45858 548466 46094
rect 548702 45858 548786 46094
rect 549022 45858 591102 46094
rect 591338 45858 591422 46094
rect 591658 45858 592650 46094
rect -8726 45774 592650 45858
rect -8726 45538 -7734 45774
rect -7498 45538 -7414 45774
rect -7178 45538 8466 45774
rect 8702 45538 8786 45774
rect 9022 45538 44466 45774
rect 44702 45538 44786 45774
rect 45022 45538 80466 45774
rect 80702 45538 80786 45774
rect 81022 45538 116466 45774
rect 116702 45538 116786 45774
rect 117022 45538 152466 45774
rect 152702 45538 152786 45774
rect 153022 45538 188466 45774
rect 188702 45538 188786 45774
rect 189022 45538 224466 45774
rect 224702 45538 224786 45774
rect 225022 45538 260466 45774
rect 260702 45538 260786 45774
rect 261022 45538 296466 45774
rect 296702 45538 296786 45774
rect 297022 45538 332466 45774
rect 332702 45538 332786 45774
rect 333022 45538 368466 45774
rect 368702 45538 368786 45774
rect 369022 45538 404466 45774
rect 404702 45538 404786 45774
rect 405022 45538 440466 45774
rect 440702 45538 440786 45774
rect 441022 45538 476466 45774
rect 476702 45538 476786 45774
rect 477022 45538 512466 45774
rect 512702 45538 512786 45774
rect 513022 45538 548466 45774
rect 548702 45538 548786 45774
rect 549022 45538 591102 45774
rect 591338 45538 591422 45774
rect 591658 45538 592650 45774
rect -8726 45506 592650 45538
rect -8726 44854 592650 44886
rect -8726 44618 -6774 44854
rect -6538 44618 -6454 44854
rect -6218 44618 7226 44854
rect 7462 44618 7546 44854
rect 7782 44618 43226 44854
rect 43462 44618 43546 44854
rect 43782 44618 79226 44854
rect 79462 44618 79546 44854
rect 79782 44618 115226 44854
rect 115462 44618 115546 44854
rect 115782 44618 151226 44854
rect 151462 44618 151546 44854
rect 151782 44618 187226 44854
rect 187462 44618 187546 44854
rect 187782 44618 223226 44854
rect 223462 44618 223546 44854
rect 223782 44618 259226 44854
rect 259462 44618 259546 44854
rect 259782 44618 295226 44854
rect 295462 44618 295546 44854
rect 295782 44618 331226 44854
rect 331462 44618 331546 44854
rect 331782 44618 367226 44854
rect 367462 44618 367546 44854
rect 367782 44618 403226 44854
rect 403462 44618 403546 44854
rect 403782 44618 439226 44854
rect 439462 44618 439546 44854
rect 439782 44618 475226 44854
rect 475462 44618 475546 44854
rect 475782 44618 511226 44854
rect 511462 44618 511546 44854
rect 511782 44618 547226 44854
rect 547462 44618 547546 44854
rect 547782 44618 590142 44854
rect 590378 44618 590462 44854
rect 590698 44618 592650 44854
rect -8726 44534 592650 44618
rect -8726 44298 -6774 44534
rect -6538 44298 -6454 44534
rect -6218 44298 7226 44534
rect 7462 44298 7546 44534
rect 7782 44298 43226 44534
rect 43462 44298 43546 44534
rect 43782 44298 79226 44534
rect 79462 44298 79546 44534
rect 79782 44298 115226 44534
rect 115462 44298 115546 44534
rect 115782 44298 151226 44534
rect 151462 44298 151546 44534
rect 151782 44298 187226 44534
rect 187462 44298 187546 44534
rect 187782 44298 223226 44534
rect 223462 44298 223546 44534
rect 223782 44298 259226 44534
rect 259462 44298 259546 44534
rect 259782 44298 295226 44534
rect 295462 44298 295546 44534
rect 295782 44298 331226 44534
rect 331462 44298 331546 44534
rect 331782 44298 367226 44534
rect 367462 44298 367546 44534
rect 367782 44298 403226 44534
rect 403462 44298 403546 44534
rect 403782 44298 439226 44534
rect 439462 44298 439546 44534
rect 439782 44298 475226 44534
rect 475462 44298 475546 44534
rect 475782 44298 511226 44534
rect 511462 44298 511546 44534
rect 511782 44298 547226 44534
rect 547462 44298 547546 44534
rect 547782 44298 590142 44534
rect 590378 44298 590462 44534
rect 590698 44298 592650 44534
rect -8726 44266 592650 44298
rect -8726 43614 592650 43646
rect -8726 43378 -5814 43614
rect -5578 43378 -5494 43614
rect -5258 43378 5986 43614
rect 6222 43378 6306 43614
rect 6542 43378 41986 43614
rect 42222 43378 42306 43614
rect 42542 43378 77986 43614
rect 78222 43378 78306 43614
rect 78542 43378 113986 43614
rect 114222 43378 114306 43614
rect 114542 43378 149986 43614
rect 150222 43378 150306 43614
rect 150542 43378 185986 43614
rect 186222 43378 186306 43614
rect 186542 43378 221986 43614
rect 222222 43378 222306 43614
rect 222542 43378 257986 43614
rect 258222 43378 258306 43614
rect 258542 43378 293986 43614
rect 294222 43378 294306 43614
rect 294542 43378 329986 43614
rect 330222 43378 330306 43614
rect 330542 43378 365986 43614
rect 366222 43378 366306 43614
rect 366542 43378 401986 43614
rect 402222 43378 402306 43614
rect 402542 43378 437986 43614
rect 438222 43378 438306 43614
rect 438542 43378 473986 43614
rect 474222 43378 474306 43614
rect 474542 43378 509986 43614
rect 510222 43378 510306 43614
rect 510542 43378 545986 43614
rect 546222 43378 546306 43614
rect 546542 43378 581986 43614
rect 582222 43378 582306 43614
rect 582542 43378 589182 43614
rect 589418 43378 589502 43614
rect 589738 43378 592650 43614
rect -8726 43294 592650 43378
rect -8726 43058 -5814 43294
rect -5578 43058 -5494 43294
rect -5258 43058 5986 43294
rect 6222 43058 6306 43294
rect 6542 43058 41986 43294
rect 42222 43058 42306 43294
rect 42542 43058 77986 43294
rect 78222 43058 78306 43294
rect 78542 43058 113986 43294
rect 114222 43058 114306 43294
rect 114542 43058 149986 43294
rect 150222 43058 150306 43294
rect 150542 43058 185986 43294
rect 186222 43058 186306 43294
rect 186542 43058 221986 43294
rect 222222 43058 222306 43294
rect 222542 43058 257986 43294
rect 258222 43058 258306 43294
rect 258542 43058 293986 43294
rect 294222 43058 294306 43294
rect 294542 43058 329986 43294
rect 330222 43058 330306 43294
rect 330542 43058 365986 43294
rect 366222 43058 366306 43294
rect 366542 43058 401986 43294
rect 402222 43058 402306 43294
rect 402542 43058 437986 43294
rect 438222 43058 438306 43294
rect 438542 43058 473986 43294
rect 474222 43058 474306 43294
rect 474542 43058 509986 43294
rect 510222 43058 510306 43294
rect 510542 43058 545986 43294
rect 546222 43058 546306 43294
rect 546542 43058 581986 43294
rect 582222 43058 582306 43294
rect 582542 43058 589182 43294
rect 589418 43058 589502 43294
rect 589738 43058 592650 43294
rect -8726 43026 592650 43058
rect -8726 42374 592650 42406
rect -8726 42138 -4854 42374
rect -4618 42138 -4534 42374
rect -4298 42138 4746 42374
rect 4982 42138 5066 42374
rect 5302 42138 40746 42374
rect 40982 42138 41066 42374
rect 41302 42138 76746 42374
rect 76982 42138 77066 42374
rect 77302 42138 112746 42374
rect 112982 42138 113066 42374
rect 113302 42138 148746 42374
rect 148982 42138 149066 42374
rect 149302 42138 184746 42374
rect 184982 42138 185066 42374
rect 185302 42138 220746 42374
rect 220982 42138 221066 42374
rect 221302 42138 256746 42374
rect 256982 42138 257066 42374
rect 257302 42138 292746 42374
rect 292982 42138 293066 42374
rect 293302 42138 328746 42374
rect 328982 42138 329066 42374
rect 329302 42138 364746 42374
rect 364982 42138 365066 42374
rect 365302 42138 400746 42374
rect 400982 42138 401066 42374
rect 401302 42138 436746 42374
rect 436982 42138 437066 42374
rect 437302 42138 472746 42374
rect 472982 42138 473066 42374
rect 473302 42138 508746 42374
rect 508982 42138 509066 42374
rect 509302 42138 544746 42374
rect 544982 42138 545066 42374
rect 545302 42138 580746 42374
rect 580982 42138 581066 42374
rect 581302 42138 588222 42374
rect 588458 42138 588542 42374
rect 588778 42138 592650 42374
rect -8726 42054 592650 42138
rect -8726 41818 -4854 42054
rect -4618 41818 -4534 42054
rect -4298 41818 4746 42054
rect 4982 41818 5066 42054
rect 5302 41818 40746 42054
rect 40982 41818 41066 42054
rect 41302 41818 76746 42054
rect 76982 41818 77066 42054
rect 77302 41818 112746 42054
rect 112982 41818 113066 42054
rect 113302 41818 148746 42054
rect 148982 41818 149066 42054
rect 149302 41818 184746 42054
rect 184982 41818 185066 42054
rect 185302 41818 220746 42054
rect 220982 41818 221066 42054
rect 221302 41818 256746 42054
rect 256982 41818 257066 42054
rect 257302 41818 292746 42054
rect 292982 41818 293066 42054
rect 293302 41818 328746 42054
rect 328982 41818 329066 42054
rect 329302 41818 364746 42054
rect 364982 41818 365066 42054
rect 365302 41818 400746 42054
rect 400982 41818 401066 42054
rect 401302 41818 436746 42054
rect 436982 41818 437066 42054
rect 437302 41818 472746 42054
rect 472982 41818 473066 42054
rect 473302 41818 508746 42054
rect 508982 41818 509066 42054
rect 509302 41818 544746 42054
rect 544982 41818 545066 42054
rect 545302 41818 580746 42054
rect 580982 41818 581066 42054
rect 581302 41818 588222 42054
rect 588458 41818 588542 42054
rect 588778 41818 592650 42054
rect -8726 41786 592650 41818
rect -8726 41134 592650 41166
rect -8726 40898 -3894 41134
rect -3658 40898 -3574 41134
rect -3338 40898 3506 41134
rect 3742 40898 3826 41134
rect 4062 40898 39506 41134
rect 39742 40898 39826 41134
rect 40062 40898 75506 41134
rect 75742 40898 75826 41134
rect 76062 40898 111506 41134
rect 111742 40898 111826 41134
rect 112062 40898 147506 41134
rect 147742 40898 147826 41134
rect 148062 40898 183506 41134
rect 183742 40898 183826 41134
rect 184062 40898 219506 41134
rect 219742 40898 219826 41134
rect 220062 40898 255506 41134
rect 255742 40898 255826 41134
rect 256062 40898 291506 41134
rect 291742 40898 291826 41134
rect 292062 40898 327506 41134
rect 327742 40898 327826 41134
rect 328062 40898 363506 41134
rect 363742 40898 363826 41134
rect 364062 40898 399506 41134
rect 399742 40898 399826 41134
rect 400062 40898 435506 41134
rect 435742 40898 435826 41134
rect 436062 40898 471506 41134
rect 471742 40898 471826 41134
rect 472062 40898 507506 41134
rect 507742 40898 507826 41134
rect 508062 40898 543506 41134
rect 543742 40898 543826 41134
rect 544062 40898 579506 41134
rect 579742 40898 579826 41134
rect 580062 40898 587262 41134
rect 587498 40898 587582 41134
rect 587818 40898 592650 41134
rect -8726 40814 592650 40898
rect -8726 40578 -3894 40814
rect -3658 40578 -3574 40814
rect -3338 40578 3506 40814
rect 3742 40578 3826 40814
rect 4062 40578 39506 40814
rect 39742 40578 39826 40814
rect 40062 40578 75506 40814
rect 75742 40578 75826 40814
rect 76062 40578 111506 40814
rect 111742 40578 111826 40814
rect 112062 40578 147506 40814
rect 147742 40578 147826 40814
rect 148062 40578 183506 40814
rect 183742 40578 183826 40814
rect 184062 40578 219506 40814
rect 219742 40578 219826 40814
rect 220062 40578 255506 40814
rect 255742 40578 255826 40814
rect 256062 40578 291506 40814
rect 291742 40578 291826 40814
rect 292062 40578 327506 40814
rect 327742 40578 327826 40814
rect 328062 40578 363506 40814
rect 363742 40578 363826 40814
rect 364062 40578 399506 40814
rect 399742 40578 399826 40814
rect 400062 40578 435506 40814
rect 435742 40578 435826 40814
rect 436062 40578 471506 40814
rect 471742 40578 471826 40814
rect 472062 40578 507506 40814
rect 507742 40578 507826 40814
rect 508062 40578 543506 40814
rect 543742 40578 543826 40814
rect 544062 40578 579506 40814
rect 579742 40578 579826 40814
rect 580062 40578 587262 40814
rect 587498 40578 587582 40814
rect 587818 40578 592650 40814
rect -8726 40546 592650 40578
rect -8726 39894 592650 39926
rect -8726 39658 -2934 39894
rect -2698 39658 -2614 39894
rect -2378 39658 2266 39894
rect 2502 39658 2586 39894
rect 2822 39658 38266 39894
rect 38502 39658 38586 39894
rect 38822 39658 74266 39894
rect 74502 39658 74586 39894
rect 74822 39658 110266 39894
rect 110502 39658 110586 39894
rect 110822 39658 146266 39894
rect 146502 39658 146586 39894
rect 146822 39658 182266 39894
rect 182502 39658 182586 39894
rect 182822 39658 218266 39894
rect 218502 39658 218586 39894
rect 218822 39658 254266 39894
rect 254502 39658 254586 39894
rect 254822 39658 290266 39894
rect 290502 39658 290586 39894
rect 290822 39658 326266 39894
rect 326502 39658 326586 39894
rect 326822 39658 362266 39894
rect 362502 39658 362586 39894
rect 362822 39658 398266 39894
rect 398502 39658 398586 39894
rect 398822 39658 434266 39894
rect 434502 39658 434586 39894
rect 434822 39658 470266 39894
rect 470502 39658 470586 39894
rect 470822 39658 506266 39894
rect 506502 39658 506586 39894
rect 506822 39658 542266 39894
rect 542502 39658 542586 39894
rect 542822 39658 578266 39894
rect 578502 39658 578586 39894
rect 578822 39658 586302 39894
rect 586538 39658 586622 39894
rect 586858 39658 592650 39894
rect -8726 39574 592650 39658
rect -8726 39338 -2934 39574
rect -2698 39338 -2614 39574
rect -2378 39338 2266 39574
rect 2502 39338 2586 39574
rect 2822 39338 38266 39574
rect 38502 39338 38586 39574
rect 38822 39338 74266 39574
rect 74502 39338 74586 39574
rect 74822 39338 110266 39574
rect 110502 39338 110586 39574
rect 110822 39338 146266 39574
rect 146502 39338 146586 39574
rect 146822 39338 182266 39574
rect 182502 39338 182586 39574
rect 182822 39338 218266 39574
rect 218502 39338 218586 39574
rect 218822 39338 254266 39574
rect 254502 39338 254586 39574
rect 254822 39338 290266 39574
rect 290502 39338 290586 39574
rect 290822 39338 326266 39574
rect 326502 39338 326586 39574
rect 326822 39338 362266 39574
rect 362502 39338 362586 39574
rect 362822 39338 398266 39574
rect 398502 39338 398586 39574
rect 398822 39338 434266 39574
rect 434502 39338 434586 39574
rect 434822 39338 470266 39574
rect 470502 39338 470586 39574
rect 470822 39338 506266 39574
rect 506502 39338 506586 39574
rect 506822 39338 542266 39574
rect 542502 39338 542586 39574
rect 542822 39338 578266 39574
rect 578502 39338 578586 39574
rect 578822 39338 586302 39574
rect 586538 39338 586622 39574
rect 586858 39338 592650 39574
rect -8726 39306 592650 39338
rect -8726 38654 592650 38686
rect -8726 38418 -1974 38654
rect -1738 38418 -1654 38654
rect -1418 38418 1026 38654
rect 1262 38418 1346 38654
rect 1582 38418 37026 38654
rect 37262 38418 37346 38654
rect 37582 38418 73026 38654
rect 73262 38418 73346 38654
rect 73582 38418 109026 38654
rect 109262 38418 109346 38654
rect 109582 38418 145026 38654
rect 145262 38418 145346 38654
rect 145582 38418 181026 38654
rect 181262 38418 181346 38654
rect 181582 38418 217026 38654
rect 217262 38418 217346 38654
rect 217582 38418 253026 38654
rect 253262 38418 253346 38654
rect 253582 38418 289026 38654
rect 289262 38418 289346 38654
rect 289582 38418 325026 38654
rect 325262 38418 325346 38654
rect 325582 38418 361026 38654
rect 361262 38418 361346 38654
rect 361582 38418 397026 38654
rect 397262 38418 397346 38654
rect 397582 38418 433026 38654
rect 433262 38418 433346 38654
rect 433582 38418 469026 38654
rect 469262 38418 469346 38654
rect 469582 38418 505026 38654
rect 505262 38418 505346 38654
rect 505582 38418 541026 38654
rect 541262 38418 541346 38654
rect 541582 38418 577026 38654
rect 577262 38418 577346 38654
rect 577582 38418 585342 38654
rect 585578 38418 585662 38654
rect 585898 38418 592650 38654
rect -8726 38334 592650 38418
rect -8726 38098 -1974 38334
rect -1738 38098 -1654 38334
rect -1418 38098 1026 38334
rect 1262 38098 1346 38334
rect 1582 38098 37026 38334
rect 37262 38098 37346 38334
rect 37582 38098 73026 38334
rect 73262 38098 73346 38334
rect 73582 38098 109026 38334
rect 109262 38098 109346 38334
rect 109582 38098 145026 38334
rect 145262 38098 145346 38334
rect 145582 38098 181026 38334
rect 181262 38098 181346 38334
rect 181582 38098 217026 38334
rect 217262 38098 217346 38334
rect 217582 38098 253026 38334
rect 253262 38098 253346 38334
rect 253582 38098 289026 38334
rect 289262 38098 289346 38334
rect 289582 38098 325026 38334
rect 325262 38098 325346 38334
rect 325582 38098 361026 38334
rect 361262 38098 361346 38334
rect 361582 38098 397026 38334
rect 397262 38098 397346 38334
rect 397582 38098 433026 38334
rect 433262 38098 433346 38334
rect 433582 38098 469026 38334
rect 469262 38098 469346 38334
rect 469582 38098 505026 38334
rect 505262 38098 505346 38334
rect 505582 38098 541026 38334
rect 541262 38098 541346 38334
rect 541582 38098 577026 38334
rect 577262 38098 577346 38334
rect 577582 38098 585342 38334
rect 585578 38098 585662 38334
rect 585898 38098 592650 38334
rect -8726 38066 592650 38098
rect -8726 11334 592650 11366
rect -8726 11098 -8694 11334
rect -8458 11098 -8374 11334
rect -8138 11098 9706 11334
rect 9942 11098 10026 11334
rect 10262 11098 45706 11334
rect 45942 11098 46026 11334
rect 46262 11098 81706 11334
rect 81942 11098 82026 11334
rect 82262 11098 117706 11334
rect 117942 11098 118026 11334
rect 118262 11098 153706 11334
rect 153942 11098 154026 11334
rect 154262 11098 189706 11334
rect 189942 11098 190026 11334
rect 190262 11098 225706 11334
rect 225942 11098 226026 11334
rect 226262 11098 261706 11334
rect 261942 11098 262026 11334
rect 262262 11098 297706 11334
rect 297942 11098 298026 11334
rect 298262 11098 333706 11334
rect 333942 11098 334026 11334
rect 334262 11098 369706 11334
rect 369942 11098 370026 11334
rect 370262 11098 405706 11334
rect 405942 11098 406026 11334
rect 406262 11098 441706 11334
rect 441942 11098 442026 11334
rect 442262 11098 477706 11334
rect 477942 11098 478026 11334
rect 478262 11098 513706 11334
rect 513942 11098 514026 11334
rect 514262 11098 549706 11334
rect 549942 11098 550026 11334
rect 550262 11098 592062 11334
rect 592298 11098 592382 11334
rect 592618 11098 592650 11334
rect -8726 11014 592650 11098
rect -8726 10778 -8694 11014
rect -8458 10778 -8374 11014
rect -8138 10778 9706 11014
rect 9942 10778 10026 11014
rect 10262 10778 45706 11014
rect 45942 10778 46026 11014
rect 46262 10778 81706 11014
rect 81942 10778 82026 11014
rect 82262 10778 117706 11014
rect 117942 10778 118026 11014
rect 118262 10778 153706 11014
rect 153942 10778 154026 11014
rect 154262 10778 189706 11014
rect 189942 10778 190026 11014
rect 190262 10778 225706 11014
rect 225942 10778 226026 11014
rect 226262 10778 261706 11014
rect 261942 10778 262026 11014
rect 262262 10778 297706 11014
rect 297942 10778 298026 11014
rect 298262 10778 333706 11014
rect 333942 10778 334026 11014
rect 334262 10778 369706 11014
rect 369942 10778 370026 11014
rect 370262 10778 405706 11014
rect 405942 10778 406026 11014
rect 406262 10778 441706 11014
rect 441942 10778 442026 11014
rect 442262 10778 477706 11014
rect 477942 10778 478026 11014
rect 478262 10778 513706 11014
rect 513942 10778 514026 11014
rect 514262 10778 549706 11014
rect 549942 10778 550026 11014
rect 550262 10778 592062 11014
rect 592298 10778 592382 11014
rect 592618 10778 592650 11014
rect -8726 10746 592650 10778
rect -8726 10094 592650 10126
rect -8726 9858 -7734 10094
rect -7498 9858 -7414 10094
rect -7178 9858 8466 10094
rect 8702 9858 8786 10094
rect 9022 9858 44466 10094
rect 44702 9858 44786 10094
rect 45022 9858 80466 10094
rect 80702 9858 80786 10094
rect 81022 9858 116466 10094
rect 116702 9858 116786 10094
rect 117022 9858 152466 10094
rect 152702 9858 152786 10094
rect 153022 9858 188466 10094
rect 188702 9858 188786 10094
rect 189022 9858 224466 10094
rect 224702 9858 224786 10094
rect 225022 9858 260466 10094
rect 260702 9858 260786 10094
rect 261022 9858 296466 10094
rect 296702 9858 296786 10094
rect 297022 9858 332466 10094
rect 332702 9858 332786 10094
rect 333022 9858 368466 10094
rect 368702 9858 368786 10094
rect 369022 9858 404466 10094
rect 404702 9858 404786 10094
rect 405022 9858 440466 10094
rect 440702 9858 440786 10094
rect 441022 9858 476466 10094
rect 476702 9858 476786 10094
rect 477022 9858 512466 10094
rect 512702 9858 512786 10094
rect 513022 9858 548466 10094
rect 548702 9858 548786 10094
rect 549022 9858 591102 10094
rect 591338 9858 591422 10094
rect 591658 9858 592650 10094
rect -8726 9774 592650 9858
rect -8726 9538 -7734 9774
rect -7498 9538 -7414 9774
rect -7178 9538 8466 9774
rect 8702 9538 8786 9774
rect 9022 9538 44466 9774
rect 44702 9538 44786 9774
rect 45022 9538 80466 9774
rect 80702 9538 80786 9774
rect 81022 9538 116466 9774
rect 116702 9538 116786 9774
rect 117022 9538 152466 9774
rect 152702 9538 152786 9774
rect 153022 9538 188466 9774
rect 188702 9538 188786 9774
rect 189022 9538 224466 9774
rect 224702 9538 224786 9774
rect 225022 9538 260466 9774
rect 260702 9538 260786 9774
rect 261022 9538 296466 9774
rect 296702 9538 296786 9774
rect 297022 9538 332466 9774
rect 332702 9538 332786 9774
rect 333022 9538 368466 9774
rect 368702 9538 368786 9774
rect 369022 9538 404466 9774
rect 404702 9538 404786 9774
rect 405022 9538 440466 9774
rect 440702 9538 440786 9774
rect 441022 9538 476466 9774
rect 476702 9538 476786 9774
rect 477022 9538 512466 9774
rect 512702 9538 512786 9774
rect 513022 9538 548466 9774
rect 548702 9538 548786 9774
rect 549022 9538 591102 9774
rect 591338 9538 591422 9774
rect 591658 9538 592650 9774
rect -8726 9506 592650 9538
rect -8726 8854 592650 8886
rect -8726 8618 -6774 8854
rect -6538 8618 -6454 8854
rect -6218 8618 7226 8854
rect 7462 8618 7546 8854
rect 7782 8618 43226 8854
rect 43462 8618 43546 8854
rect 43782 8618 79226 8854
rect 79462 8618 79546 8854
rect 79782 8618 115226 8854
rect 115462 8618 115546 8854
rect 115782 8618 151226 8854
rect 151462 8618 151546 8854
rect 151782 8618 187226 8854
rect 187462 8618 187546 8854
rect 187782 8618 223226 8854
rect 223462 8618 223546 8854
rect 223782 8618 259226 8854
rect 259462 8618 259546 8854
rect 259782 8618 295226 8854
rect 295462 8618 295546 8854
rect 295782 8618 331226 8854
rect 331462 8618 331546 8854
rect 331782 8618 367226 8854
rect 367462 8618 367546 8854
rect 367782 8618 403226 8854
rect 403462 8618 403546 8854
rect 403782 8618 439226 8854
rect 439462 8618 439546 8854
rect 439782 8618 475226 8854
rect 475462 8618 475546 8854
rect 475782 8618 511226 8854
rect 511462 8618 511546 8854
rect 511782 8618 547226 8854
rect 547462 8618 547546 8854
rect 547782 8618 590142 8854
rect 590378 8618 590462 8854
rect 590698 8618 592650 8854
rect -8726 8534 592650 8618
rect -8726 8298 -6774 8534
rect -6538 8298 -6454 8534
rect -6218 8298 7226 8534
rect 7462 8298 7546 8534
rect 7782 8298 43226 8534
rect 43462 8298 43546 8534
rect 43782 8298 79226 8534
rect 79462 8298 79546 8534
rect 79782 8298 115226 8534
rect 115462 8298 115546 8534
rect 115782 8298 151226 8534
rect 151462 8298 151546 8534
rect 151782 8298 187226 8534
rect 187462 8298 187546 8534
rect 187782 8298 223226 8534
rect 223462 8298 223546 8534
rect 223782 8298 259226 8534
rect 259462 8298 259546 8534
rect 259782 8298 295226 8534
rect 295462 8298 295546 8534
rect 295782 8298 331226 8534
rect 331462 8298 331546 8534
rect 331782 8298 367226 8534
rect 367462 8298 367546 8534
rect 367782 8298 403226 8534
rect 403462 8298 403546 8534
rect 403782 8298 439226 8534
rect 439462 8298 439546 8534
rect 439782 8298 475226 8534
rect 475462 8298 475546 8534
rect 475782 8298 511226 8534
rect 511462 8298 511546 8534
rect 511782 8298 547226 8534
rect 547462 8298 547546 8534
rect 547782 8298 590142 8534
rect 590378 8298 590462 8534
rect 590698 8298 592650 8534
rect -8726 8266 592650 8298
rect -8726 7614 592650 7646
rect -8726 7378 -5814 7614
rect -5578 7378 -5494 7614
rect -5258 7378 5986 7614
rect 6222 7378 6306 7614
rect 6542 7378 41986 7614
rect 42222 7378 42306 7614
rect 42542 7378 77986 7614
rect 78222 7378 78306 7614
rect 78542 7378 113986 7614
rect 114222 7378 114306 7614
rect 114542 7378 149986 7614
rect 150222 7378 150306 7614
rect 150542 7378 185986 7614
rect 186222 7378 186306 7614
rect 186542 7378 221986 7614
rect 222222 7378 222306 7614
rect 222542 7378 257986 7614
rect 258222 7378 258306 7614
rect 258542 7378 293986 7614
rect 294222 7378 294306 7614
rect 294542 7378 329986 7614
rect 330222 7378 330306 7614
rect 330542 7378 365986 7614
rect 366222 7378 366306 7614
rect 366542 7378 401986 7614
rect 402222 7378 402306 7614
rect 402542 7378 437986 7614
rect 438222 7378 438306 7614
rect 438542 7378 473986 7614
rect 474222 7378 474306 7614
rect 474542 7378 509986 7614
rect 510222 7378 510306 7614
rect 510542 7378 545986 7614
rect 546222 7378 546306 7614
rect 546542 7378 581986 7614
rect 582222 7378 582306 7614
rect 582542 7378 589182 7614
rect 589418 7378 589502 7614
rect 589738 7378 592650 7614
rect -8726 7294 592650 7378
rect -8726 7058 -5814 7294
rect -5578 7058 -5494 7294
rect -5258 7058 5986 7294
rect 6222 7058 6306 7294
rect 6542 7058 41986 7294
rect 42222 7058 42306 7294
rect 42542 7058 77986 7294
rect 78222 7058 78306 7294
rect 78542 7058 113986 7294
rect 114222 7058 114306 7294
rect 114542 7058 149986 7294
rect 150222 7058 150306 7294
rect 150542 7058 185986 7294
rect 186222 7058 186306 7294
rect 186542 7058 221986 7294
rect 222222 7058 222306 7294
rect 222542 7058 257986 7294
rect 258222 7058 258306 7294
rect 258542 7058 293986 7294
rect 294222 7058 294306 7294
rect 294542 7058 329986 7294
rect 330222 7058 330306 7294
rect 330542 7058 365986 7294
rect 366222 7058 366306 7294
rect 366542 7058 401986 7294
rect 402222 7058 402306 7294
rect 402542 7058 437986 7294
rect 438222 7058 438306 7294
rect 438542 7058 473986 7294
rect 474222 7058 474306 7294
rect 474542 7058 509986 7294
rect 510222 7058 510306 7294
rect 510542 7058 545986 7294
rect 546222 7058 546306 7294
rect 546542 7058 581986 7294
rect 582222 7058 582306 7294
rect 582542 7058 589182 7294
rect 589418 7058 589502 7294
rect 589738 7058 592650 7294
rect -8726 7026 592650 7058
rect -8726 6374 592650 6406
rect -8726 6138 -4854 6374
rect -4618 6138 -4534 6374
rect -4298 6138 4746 6374
rect 4982 6138 5066 6374
rect 5302 6138 40746 6374
rect 40982 6138 41066 6374
rect 41302 6138 76746 6374
rect 76982 6138 77066 6374
rect 77302 6138 112746 6374
rect 112982 6138 113066 6374
rect 113302 6138 148746 6374
rect 148982 6138 149066 6374
rect 149302 6138 184746 6374
rect 184982 6138 185066 6374
rect 185302 6138 220746 6374
rect 220982 6138 221066 6374
rect 221302 6138 256746 6374
rect 256982 6138 257066 6374
rect 257302 6138 292746 6374
rect 292982 6138 293066 6374
rect 293302 6138 328746 6374
rect 328982 6138 329066 6374
rect 329302 6138 364746 6374
rect 364982 6138 365066 6374
rect 365302 6138 400746 6374
rect 400982 6138 401066 6374
rect 401302 6138 436746 6374
rect 436982 6138 437066 6374
rect 437302 6138 472746 6374
rect 472982 6138 473066 6374
rect 473302 6138 508746 6374
rect 508982 6138 509066 6374
rect 509302 6138 544746 6374
rect 544982 6138 545066 6374
rect 545302 6138 580746 6374
rect 580982 6138 581066 6374
rect 581302 6138 588222 6374
rect 588458 6138 588542 6374
rect 588778 6138 592650 6374
rect -8726 6054 592650 6138
rect -8726 5818 -4854 6054
rect -4618 5818 -4534 6054
rect -4298 5818 4746 6054
rect 4982 5818 5066 6054
rect 5302 5818 40746 6054
rect 40982 5818 41066 6054
rect 41302 5818 76746 6054
rect 76982 5818 77066 6054
rect 77302 5818 112746 6054
rect 112982 5818 113066 6054
rect 113302 5818 148746 6054
rect 148982 5818 149066 6054
rect 149302 5818 184746 6054
rect 184982 5818 185066 6054
rect 185302 5818 220746 6054
rect 220982 5818 221066 6054
rect 221302 5818 256746 6054
rect 256982 5818 257066 6054
rect 257302 5818 292746 6054
rect 292982 5818 293066 6054
rect 293302 5818 328746 6054
rect 328982 5818 329066 6054
rect 329302 5818 364746 6054
rect 364982 5818 365066 6054
rect 365302 5818 400746 6054
rect 400982 5818 401066 6054
rect 401302 5818 436746 6054
rect 436982 5818 437066 6054
rect 437302 5818 472746 6054
rect 472982 5818 473066 6054
rect 473302 5818 508746 6054
rect 508982 5818 509066 6054
rect 509302 5818 544746 6054
rect 544982 5818 545066 6054
rect 545302 5818 580746 6054
rect 580982 5818 581066 6054
rect 581302 5818 588222 6054
rect 588458 5818 588542 6054
rect 588778 5818 592650 6054
rect -8726 5786 592650 5818
rect -8726 5134 592650 5166
rect -8726 4898 -3894 5134
rect -3658 4898 -3574 5134
rect -3338 4898 3506 5134
rect 3742 4898 3826 5134
rect 4062 4898 39506 5134
rect 39742 4898 39826 5134
rect 40062 4898 75506 5134
rect 75742 4898 75826 5134
rect 76062 4898 111506 5134
rect 111742 4898 111826 5134
rect 112062 4898 147506 5134
rect 147742 4898 147826 5134
rect 148062 4898 183506 5134
rect 183742 4898 183826 5134
rect 184062 4898 219506 5134
rect 219742 4898 219826 5134
rect 220062 4898 255506 5134
rect 255742 4898 255826 5134
rect 256062 4898 291506 5134
rect 291742 4898 291826 5134
rect 292062 4898 327506 5134
rect 327742 4898 327826 5134
rect 328062 4898 363506 5134
rect 363742 4898 363826 5134
rect 364062 4898 399506 5134
rect 399742 4898 399826 5134
rect 400062 4898 435506 5134
rect 435742 4898 435826 5134
rect 436062 4898 471506 5134
rect 471742 4898 471826 5134
rect 472062 4898 507506 5134
rect 507742 4898 507826 5134
rect 508062 4898 543506 5134
rect 543742 4898 543826 5134
rect 544062 4898 579506 5134
rect 579742 4898 579826 5134
rect 580062 4898 587262 5134
rect 587498 4898 587582 5134
rect 587818 4898 592650 5134
rect -8726 4814 592650 4898
rect -8726 4578 -3894 4814
rect -3658 4578 -3574 4814
rect -3338 4578 3506 4814
rect 3742 4578 3826 4814
rect 4062 4578 39506 4814
rect 39742 4578 39826 4814
rect 40062 4578 75506 4814
rect 75742 4578 75826 4814
rect 76062 4578 111506 4814
rect 111742 4578 111826 4814
rect 112062 4578 147506 4814
rect 147742 4578 147826 4814
rect 148062 4578 183506 4814
rect 183742 4578 183826 4814
rect 184062 4578 219506 4814
rect 219742 4578 219826 4814
rect 220062 4578 255506 4814
rect 255742 4578 255826 4814
rect 256062 4578 291506 4814
rect 291742 4578 291826 4814
rect 292062 4578 327506 4814
rect 327742 4578 327826 4814
rect 328062 4578 363506 4814
rect 363742 4578 363826 4814
rect 364062 4578 399506 4814
rect 399742 4578 399826 4814
rect 400062 4578 435506 4814
rect 435742 4578 435826 4814
rect 436062 4578 471506 4814
rect 471742 4578 471826 4814
rect 472062 4578 507506 4814
rect 507742 4578 507826 4814
rect 508062 4578 543506 4814
rect 543742 4578 543826 4814
rect 544062 4578 579506 4814
rect 579742 4578 579826 4814
rect 580062 4578 587262 4814
rect 587498 4578 587582 4814
rect 587818 4578 592650 4814
rect -8726 4546 592650 4578
rect -8726 3894 592650 3926
rect -8726 3658 -2934 3894
rect -2698 3658 -2614 3894
rect -2378 3658 2266 3894
rect 2502 3658 2586 3894
rect 2822 3658 38266 3894
rect 38502 3658 38586 3894
rect 38822 3658 74266 3894
rect 74502 3658 74586 3894
rect 74822 3658 110266 3894
rect 110502 3658 110586 3894
rect 110822 3658 146266 3894
rect 146502 3658 146586 3894
rect 146822 3658 182266 3894
rect 182502 3658 182586 3894
rect 182822 3658 218266 3894
rect 218502 3658 218586 3894
rect 218822 3658 254266 3894
rect 254502 3658 254586 3894
rect 254822 3658 290266 3894
rect 290502 3658 290586 3894
rect 290822 3658 326266 3894
rect 326502 3658 326586 3894
rect 326822 3658 362266 3894
rect 362502 3658 362586 3894
rect 362822 3658 398266 3894
rect 398502 3658 398586 3894
rect 398822 3658 434266 3894
rect 434502 3658 434586 3894
rect 434822 3658 470266 3894
rect 470502 3658 470586 3894
rect 470822 3658 506266 3894
rect 506502 3658 506586 3894
rect 506822 3658 542266 3894
rect 542502 3658 542586 3894
rect 542822 3658 578266 3894
rect 578502 3658 578586 3894
rect 578822 3658 586302 3894
rect 586538 3658 586622 3894
rect 586858 3658 592650 3894
rect -8726 3574 592650 3658
rect -8726 3338 -2934 3574
rect -2698 3338 -2614 3574
rect -2378 3338 2266 3574
rect 2502 3338 2586 3574
rect 2822 3338 38266 3574
rect 38502 3338 38586 3574
rect 38822 3338 74266 3574
rect 74502 3338 74586 3574
rect 74822 3338 110266 3574
rect 110502 3338 110586 3574
rect 110822 3338 146266 3574
rect 146502 3338 146586 3574
rect 146822 3338 182266 3574
rect 182502 3338 182586 3574
rect 182822 3338 218266 3574
rect 218502 3338 218586 3574
rect 218822 3338 254266 3574
rect 254502 3338 254586 3574
rect 254822 3338 290266 3574
rect 290502 3338 290586 3574
rect 290822 3338 326266 3574
rect 326502 3338 326586 3574
rect 326822 3338 362266 3574
rect 362502 3338 362586 3574
rect 362822 3338 398266 3574
rect 398502 3338 398586 3574
rect 398822 3338 434266 3574
rect 434502 3338 434586 3574
rect 434822 3338 470266 3574
rect 470502 3338 470586 3574
rect 470822 3338 506266 3574
rect 506502 3338 506586 3574
rect 506822 3338 542266 3574
rect 542502 3338 542586 3574
rect 542822 3338 578266 3574
rect 578502 3338 578586 3574
rect 578822 3338 586302 3574
rect 586538 3338 586622 3574
rect 586858 3338 592650 3574
rect -8726 3306 592650 3338
rect -8726 2654 592650 2686
rect -8726 2418 -1974 2654
rect -1738 2418 -1654 2654
rect -1418 2418 1026 2654
rect 1262 2418 1346 2654
rect 1582 2418 37026 2654
rect 37262 2418 37346 2654
rect 37582 2418 73026 2654
rect 73262 2418 73346 2654
rect 73582 2418 109026 2654
rect 109262 2418 109346 2654
rect 109582 2418 145026 2654
rect 145262 2418 145346 2654
rect 145582 2418 181026 2654
rect 181262 2418 181346 2654
rect 181582 2418 217026 2654
rect 217262 2418 217346 2654
rect 217582 2418 253026 2654
rect 253262 2418 253346 2654
rect 253582 2418 289026 2654
rect 289262 2418 289346 2654
rect 289582 2418 325026 2654
rect 325262 2418 325346 2654
rect 325582 2418 361026 2654
rect 361262 2418 361346 2654
rect 361582 2418 397026 2654
rect 397262 2418 397346 2654
rect 397582 2418 433026 2654
rect 433262 2418 433346 2654
rect 433582 2418 469026 2654
rect 469262 2418 469346 2654
rect 469582 2418 505026 2654
rect 505262 2418 505346 2654
rect 505582 2418 541026 2654
rect 541262 2418 541346 2654
rect 541582 2418 577026 2654
rect 577262 2418 577346 2654
rect 577582 2418 585342 2654
rect 585578 2418 585662 2654
rect 585898 2418 592650 2654
rect -8726 2334 592650 2418
rect -8726 2098 -1974 2334
rect -1738 2098 -1654 2334
rect -1418 2098 1026 2334
rect 1262 2098 1346 2334
rect 1582 2098 37026 2334
rect 37262 2098 37346 2334
rect 37582 2098 73026 2334
rect 73262 2098 73346 2334
rect 73582 2098 109026 2334
rect 109262 2098 109346 2334
rect 109582 2098 145026 2334
rect 145262 2098 145346 2334
rect 145582 2098 181026 2334
rect 181262 2098 181346 2334
rect 181582 2098 217026 2334
rect 217262 2098 217346 2334
rect 217582 2098 253026 2334
rect 253262 2098 253346 2334
rect 253582 2098 289026 2334
rect 289262 2098 289346 2334
rect 289582 2098 325026 2334
rect 325262 2098 325346 2334
rect 325582 2098 361026 2334
rect 361262 2098 361346 2334
rect 361582 2098 397026 2334
rect 397262 2098 397346 2334
rect 397582 2098 433026 2334
rect 433262 2098 433346 2334
rect 433582 2098 469026 2334
rect 469262 2098 469346 2334
rect 469582 2098 505026 2334
rect 505262 2098 505346 2334
rect 505582 2098 541026 2334
rect 541262 2098 541346 2334
rect 541582 2098 577026 2334
rect 577262 2098 577346 2334
rect 577582 2098 585342 2334
rect 585578 2098 585662 2334
rect 585898 2098 592650 2334
rect -8726 2066 592650 2098
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1026 -346
rect 1262 -582 1346 -346
rect 1582 -582 37026 -346
rect 37262 -582 37346 -346
rect 37582 -582 73026 -346
rect 73262 -582 73346 -346
rect 73582 -582 109026 -346
rect 109262 -582 109346 -346
rect 109582 -582 145026 -346
rect 145262 -582 145346 -346
rect 145582 -582 181026 -346
rect 181262 -582 181346 -346
rect 181582 -582 217026 -346
rect 217262 -582 217346 -346
rect 217582 -582 253026 -346
rect 253262 -582 253346 -346
rect 253582 -582 289026 -346
rect 289262 -582 289346 -346
rect 289582 -582 325026 -346
rect 325262 -582 325346 -346
rect 325582 -582 361026 -346
rect 361262 -582 361346 -346
rect 361582 -582 397026 -346
rect 397262 -582 397346 -346
rect 397582 -582 433026 -346
rect 433262 -582 433346 -346
rect 433582 -582 469026 -346
rect 469262 -582 469346 -346
rect 469582 -582 505026 -346
rect 505262 -582 505346 -346
rect 505582 -582 541026 -346
rect 541262 -582 541346 -346
rect 541582 -582 577026 -346
rect 577262 -582 577346 -346
rect 577582 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1026 -666
rect 1262 -902 1346 -666
rect 1582 -902 37026 -666
rect 37262 -902 37346 -666
rect 37582 -902 73026 -666
rect 73262 -902 73346 -666
rect 73582 -902 109026 -666
rect 109262 -902 109346 -666
rect 109582 -902 145026 -666
rect 145262 -902 145346 -666
rect 145582 -902 181026 -666
rect 181262 -902 181346 -666
rect 181582 -902 217026 -666
rect 217262 -902 217346 -666
rect 217582 -902 253026 -666
rect 253262 -902 253346 -666
rect 253582 -902 289026 -666
rect 289262 -902 289346 -666
rect 289582 -902 325026 -666
rect 325262 -902 325346 -666
rect 325582 -902 361026 -666
rect 361262 -902 361346 -666
rect 361582 -902 397026 -666
rect 397262 -902 397346 -666
rect 397582 -902 433026 -666
rect 433262 -902 433346 -666
rect 433582 -902 469026 -666
rect 469262 -902 469346 -666
rect 469582 -902 505026 -666
rect 505262 -902 505346 -666
rect 505582 -902 541026 -666
rect 541262 -902 541346 -666
rect 541582 -902 577026 -666
rect 577262 -902 577346 -666
rect 577582 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 2266 -1306
rect 2502 -1542 2586 -1306
rect 2822 -1542 38266 -1306
rect 38502 -1542 38586 -1306
rect 38822 -1542 74266 -1306
rect 74502 -1542 74586 -1306
rect 74822 -1542 110266 -1306
rect 110502 -1542 110586 -1306
rect 110822 -1542 146266 -1306
rect 146502 -1542 146586 -1306
rect 146822 -1542 182266 -1306
rect 182502 -1542 182586 -1306
rect 182822 -1542 218266 -1306
rect 218502 -1542 218586 -1306
rect 218822 -1542 254266 -1306
rect 254502 -1542 254586 -1306
rect 254822 -1542 290266 -1306
rect 290502 -1542 290586 -1306
rect 290822 -1542 326266 -1306
rect 326502 -1542 326586 -1306
rect 326822 -1542 362266 -1306
rect 362502 -1542 362586 -1306
rect 362822 -1542 398266 -1306
rect 398502 -1542 398586 -1306
rect 398822 -1542 434266 -1306
rect 434502 -1542 434586 -1306
rect 434822 -1542 470266 -1306
rect 470502 -1542 470586 -1306
rect 470822 -1542 506266 -1306
rect 506502 -1542 506586 -1306
rect 506822 -1542 542266 -1306
rect 542502 -1542 542586 -1306
rect 542822 -1542 578266 -1306
rect 578502 -1542 578586 -1306
rect 578822 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 2266 -1626
rect 2502 -1862 2586 -1626
rect 2822 -1862 38266 -1626
rect 38502 -1862 38586 -1626
rect 38822 -1862 74266 -1626
rect 74502 -1862 74586 -1626
rect 74822 -1862 110266 -1626
rect 110502 -1862 110586 -1626
rect 110822 -1862 146266 -1626
rect 146502 -1862 146586 -1626
rect 146822 -1862 182266 -1626
rect 182502 -1862 182586 -1626
rect 182822 -1862 218266 -1626
rect 218502 -1862 218586 -1626
rect 218822 -1862 254266 -1626
rect 254502 -1862 254586 -1626
rect 254822 -1862 290266 -1626
rect 290502 -1862 290586 -1626
rect 290822 -1862 326266 -1626
rect 326502 -1862 326586 -1626
rect 326822 -1862 362266 -1626
rect 362502 -1862 362586 -1626
rect 362822 -1862 398266 -1626
rect 398502 -1862 398586 -1626
rect 398822 -1862 434266 -1626
rect 434502 -1862 434586 -1626
rect 434822 -1862 470266 -1626
rect 470502 -1862 470586 -1626
rect 470822 -1862 506266 -1626
rect 506502 -1862 506586 -1626
rect 506822 -1862 542266 -1626
rect 542502 -1862 542586 -1626
rect 542822 -1862 578266 -1626
rect 578502 -1862 578586 -1626
rect 578822 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 3506 -2266
rect 3742 -2502 3826 -2266
rect 4062 -2502 39506 -2266
rect 39742 -2502 39826 -2266
rect 40062 -2502 75506 -2266
rect 75742 -2502 75826 -2266
rect 76062 -2502 111506 -2266
rect 111742 -2502 111826 -2266
rect 112062 -2502 147506 -2266
rect 147742 -2502 147826 -2266
rect 148062 -2502 183506 -2266
rect 183742 -2502 183826 -2266
rect 184062 -2502 219506 -2266
rect 219742 -2502 219826 -2266
rect 220062 -2502 255506 -2266
rect 255742 -2502 255826 -2266
rect 256062 -2502 291506 -2266
rect 291742 -2502 291826 -2266
rect 292062 -2502 327506 -2266
rect 327742 -2502 327826 -2266
rect 328062 -2502 363506 -2266
rect 363742 -2502 363826 -2266
rect 364062 -2502 399506 -2266
rect 399742 -2502 399826 -2266
rect 400062 -2502 435506 -2266
rect 435742 -2502 435826 -2266
rect 436062 -2502 471506 -2266
rect 471742 -2502 471826 -2266
rect 472062 -2502 507506 -2266
rect 507742 -2502 507826 -2266
rect 508062 -2502 543506 -2266
rect 543742 -2502 543826 -2266
rect 544062 -2502 579506 -2266
rect 579742 -2502 579826 -2266
rect 580062 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 3506 -2586
rect 3742 -2822 3826 -2586
rect 4062 -2822 39506 -2586
rect 39742 -2822 39826 -2586
rect 40062 -2822 75506 -2586
rect 75742 -2822 75826 -2586
rect 76062 -2822 111506 -2586
rect 111742 -2822 111826 -2586
rect 112062 -2822 147506 -2586
rect 147742 -2822 147826 -2586
rect 148062 -2822 183506 -2586
rect 183742 -2822 183826 -2586
rect 184062 -2822 219506 -2586
rect 219742 -2822 219826 -2586
rect 220062 -2822 255506 -2586
rect 255742 -2822 255826 -2586
rect 256062 -2822 291506 -2586
rect 291742 -2822 291826 -2586
rect 292062 -2822 327506 -2586
rect 327742 -2822 327826 -2586
rect 328062 -2822 363506 -2586
rect 363742 -2822 363826 -2586
rect 364062 -2822 399506 -2586
rect 399742 -2822 399826 -2586
rect 400062 -2822 435506 -2586
rect 435742 -2822 435826 -2586
rect 436062 -2822 471506 -2586
rect 471742 -2822 471826 -2586
rect 472062 -2822 507506 -2586
rect 507742 -2822 507826 -2586
rect 508062 -2822 543506 -2586
rect 543742 -2822 543826 -2586
rect 544062 -2822 579506 -2586
rect 579742 -2822 579826 -2586
rect 580062 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 4746 -3226
rect 4982 -3462 5066 -3226
rect 5302 -3462 40746 -3226
rect 40982 -3462 41066 -3226
rect 41302 -3462 76746 -3226
rect 76982 -3462 77066 -3226
rect 77302 -3462 112746 -3226
rect 112982 -3462 113066 -3226
rect 113302 -3462 148746 -3226
rect 148982 -3462 149066 -3226
rect 149302 -3462 184746 -3226
rect 184982 -3462 185066 -3226
rect 185302 -3462 220746 -3226
rect 220982 -3462 221066 -3226
rect 221302 -3462 256746 -3226
rect 256982 -3462 257066 -3226
rect 257302 -3462 292746 -3226
rect 292982 -3462 293066 -3226
rect 293302 -3462 328746 -3226
rect 328982 -3462 329066 -3226
rect 329302 -3462 364746 -3226
rect 364982 -3462 365066 -3226
rect 365302 -3462 400746 -3226
rect 400982 -3462 401066 -3226
rect 401302 -3462 436746 -3226
rect 436982 -3462 437066 -3226
rect 437302 -3462 472746 -3226
rect 472982 -3462 473066 -3226
rect 473302 -3462 508746 -3226
rect 508982 -3462 509066 -3226
rect 509302 -3462 544746 -3226
rect 544982 -3462 545066 -3226
rect 545302 -3462 580746 -3226
rect 580982 -3462 581066 -3226
rect 581302 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 4746 -3546
rect 4982 -3782 5066 -3546
rect 5302 -3782 40746 -3546
rect 40982 -3782 41066 -3546
rect 41302 -3782 76746 -3546
rect 76982 -3782 77066 -3546
rect 77302 -3782 112746 -3546
rect 112982 -3782 113066 -3546
rect 113302 -3782 148746 -3546
rect 148982 -3782 149066 -3546
rect 149302 -3782 184746 -3546
rect 184982 -3782 185066 -3546
rect 185302 -3782 220746 -3546
rect 220982 -3782 221066 -3546
rect 221302 -3782 256746 -3546
rect 256982 -3782 257066 -3546
rect 257302 -3782 292746 -3546
rect 292982 -3782 293066 -3546
rect 293302 -3782 328746 -3546
rect 328982 -3782 329066 -3546
rect 329302 -3782 364746 -3546
rect 364982 -3782 365066 -3546
rect 365302 -3782 400746 -3546
rect 400982 -3782 401066 -3546
rect 401302 -3782 436746 -3546
rect 436982 -3782 437066 -3546
rect 437302 -3782 472746 -3546
rect 472982 -3782 473066 -3546
rect 473302 -3782 508746 -3546
rect 508982 -3782 509066 -3546
rect 509302 -3782 544746 -3546
rect 544982 -3782 545066 -3546
rect 545302 -3782 580746 -3546
rect 580982 -3782 581066 -3546
rect 581302 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 5986 -4186
rect 6222 -4422 6306 -4186
rect 6542 -4422 41986 -4186
rect 42222 -4422 42306 -4186
rect 42542 -4422 77986 -4186
rect 78222 -4422 78306 -4186
rect 78542 -4422 113986 -4186
rect 114222 -4422 114306 -4186
rect 114542 -4422 149986 -4186
rect 150222 -4422 150306 -4186
rect 150542 -4422 185986 -4186
rect 186222 -4422 186306 -4186
rect 186542 -4422 221986 -4186
rect 222222 -4422 222306 -4186
rect 222542 -4422 257986 -4186
rect 258222 -4422 258306 -4186
rect 258542 -4422 293986 -4186
rect 294222 -4422 294306 -4186
rect 294542 -4422 329986 -4186
rect 330222 -4422 330306 -4186
rect 330542 -4422 365986 -4186
rect 366222 -4422 366306 -4186
rect 366542 -4422 401986 -4186
rect 402222 -4422 402306 -4186
rect 402542 -4422 437986 -4186
rect 438222 -4422 438306 -4186
rect 438542 -4422 473986 -4186
rect 474222 -4422 474306 -4186
rect 474542 -4422 509986 -4186
rect 510222 -4422 510306 -4186
rect 510542 -4422 545986 -4186
rect 546222 -4422 546306 -4186
rect 546542 -4422 581986 -4186
rect 582222 -4422 582306 -4186
rect 582542 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 5986 -4506
rect 6222 -4742 6306 -4506
rect 6542 -4742 41986 -4506
rect 42222 -4742 42306 -4506
rect 42542 -4742 77986 -4506
rect 78222 -4742 78306 -4506
rect 78542 -4742 113986 -4506
rect 114222 -4742 114306 -4506
rect 114542 -4742 149986 -4506
rect 150222 -4742 150306 -4506
rect 150542 -4742 185986 -4506
rect 186222 -4742 186306 -4506
rect 186542 -4742 221986 -4506
rect 222222 -4742 222306 -4506
rect 222542 -4742 257986 -4506
rect 258222 -4742 258306 -4506
rect 258542 -4742 293986 -4506
rect 294222 -4742 294306 -4506
rect 294542 -4742 329986 -4506
rect 330222 -4742 330306 -4506
rect 330542 -4742 365986 -4506
rect 366222 -4742 366306 -4506
rect 366542 -4742 401986 -4506
rect 402222 -4742 402306 -4506
rect 402542 -4742 437986 -4506
rect 438222 -4742 438306 -4506
rect 438542 -4742 473986 -4506
rect 474222 -4742 474306 -4506
rect 474542 -4742 509986 -4506
rect 510222 -4742 510306 -4506
rect 510542 -4742 545986 -4506
rect 546222 -4742 546306 -4506
rect 546542 -4742 581986 -4506
rect 582222 -4742 582306 -4506
rect 582542 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 7226 -5146
rect 7462 -5382 7546 -5146
rect 7782 -5382 43226 -5146
rect 43462 -5382 43546 -5146
rect 43782 -5382 79226 -5146
rect 79462 -5382 79546 -5146
rect 79782 -5382 115226 -5146
rect 115462 -5382 115546 -5146
rect 115782 -5382 151226 -5146
rect 151462 -5382 151546 -5146
rect 151782 -5382 187226 -5146
rect 187462 -5382 187546 -5146
rect 187782 -5382 223226 -5146
rect 223462 -5382 223546 -5146
rect 223782 -5382 259226 -5146
rect 259462 -5382 259546 -5146
rect 259782 -5382 295226 -5146
rect 295462 -5382 295546 -5146
rect 295782 -5382 331226 -5146
rect 331462 -5382 331546 -5146
rect 331782 -5382 367226 -5146
rect 367462 -5382 367546 -5146
rect 367782 -5382 403226 -5146
rect 403462 -5382 403546 -5146
rect 403782 -5382 439226 -5146
rect 439462 -5382 439546 -5146
rect 439782 -5382 475226 -5146
rect 475462 -5382 475546 -5146
rect 475782 -5382 511226 -5146
rect 511462 -5382 511546 -5146
rect 511782 -5382 547226 -5146
rect 547462 -5382 547546 -5146
rect 547782 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 7226 -5466
rect 7462 -5702 7546 -5466
rect 7782 -5702 43226 -5466
rect 43462 -5702 43546 -5466
rect 43782 -5702 79226 -5466
rect 79462 -5702 79546 -5466
rect 79782 -5702 115226 -5466
rect 115462 -5702 115546 -5466
rect 115782 -5702 151226 -5466
rect 151462 -5702 151546 -5466
rect 151782 -5702 187226 -5466
rect 187462 -5702 187546 -5466
rect 187782 -5702 223226 -5466
rect 223462 -5702 223546 -5466
rect 223782 -5702 259226 -5466
rect 259462 -5702 259546 -5466
rect 259782 -5702 295226 -5466
rect 295462 -5702 295546 -5466
rect 295782 -5702 331226 -5466
rect 331462 -5702 331546 -5466
rect 331782 -5702 367226 -5466
rect 367462 -5702 367546 -5466
rect 367782 -5702 403226 -5466
rect 403462 -5702 403546 -5466
rect 403782 -5702 439226 -5466
rect 439462 -5702 439546 -5466
rect 439782 -5702 475226 -5466
rect 475462 -5702 475546 -5466
rect 475782 -5702 511226 -5466
rect 511462 -5702 511546 -5466
rect 511782 -5702 547226 -5466
rect 547462 -5702 547546 -5466
rect 547782 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 8466 -6106
rect 8702 -6342 8786 -6106
rect 9022 -6342 44466 -6106
rect 44702 -6342 44786 -6106
rect 45022 -6342 80466 -6106
rect 80702 -6342 80786 -6106
rect 81022 -6342 116466 -6106
rect 116702 -6342 116786 -6106
rect 117022 -6342 152466 -6106
rect 152702 -6342 152786 -6106
rect 153022 -6342 188466 -6106
rect 188702 -6342 188786 -6106
rect 189022 -6342 224466 -6106
rect 224702 -6342 224786 -6106
rect 225022 -6342 260466 -6106
rect 260702 -6342 260786 -6106
rect 261022 -6342 296466 -6106
rect 296702 -6342 296786 -6106
rect 297022 -6342 332466 -6106
rect 332702 -6342 332786 -6106
rect 333022 -6342 368466 -6106
rect 368702 -6342 368786 -6106
rect 369022 -6342 404466 -6106
rect 404702 -6342 404786 -6106
rect 405022 -6342 440466 -6106
rect 440702 -6342 440786 -6106
rect 441022 -6342 476466 -6106
rect 476702 -6342 476786 -6106
rect 477022 -6342 512466 -6106
rect 512702 -6342 512786 -6106
rect 513022 -6342 548466 -6106
rect 548702 -6342 548786 -6106
rect 549022 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 8466 -6426
rect 8702 -6662 8786 -6426
rect 9022 -6662 44466 -6426
rect 44702 -6662 44786 -6426
rect 45022 -6662 80466 -6426
rect 80702 -6662 80786 -6426
rect 81022 -6662 116466 -6426
rect 116702 -6662 116786 -6426
rect 117022 -6662 152466 -6426
rect 152702 -6662 152786 -6426
rect 153022 -6662 188466 -6426
rect 188702 -6662 188786 -6426
rect 189022 -6662 224466 -6426
rect 224702 -6662 224786 -6426
rect 225022 -6662 260466 -6426
rect 260702 -6662 260786 -6426
rect 261022 -6662 296466 -6426
rect 296702 -6662 296786 -6426
rect 297022 -6662 332466 -6426
rect 332702 -6662 332786 -6426
rect 333022 -6662 368466 -6426
rect 368702 -6662 368786 -6426
rect 369022 -6662 404466 -6426
rect 404702 -6662 404786 -6426
rect 405022 -6662 440466 -6426
rect 440702 -6662 440786 -6426
rect 441022 -6662 476466 -6426
rect 476702 -6662 476786 -6426
rect 477022 -6662 512466 -6426
rect 512702 -6662 512786 -6426
rect 513022 -6662 548466 -6426
rect 548702 -6662 548786 -6426
rect 549022 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 9706 -7066
rect 9942 -7302 10026 -7066
rect 10262 -7302 45706 -7066
rect 45942 -7302 46026 -7066
rect 46262 -7302 81706 -7066
rect 81942 -7302 82026 -7066
rect 82262 -7302 117706 -7066
rect 117942 -7302 118026 -7066
rect 118262 -7302 153706 -7066
rect 153942 -7302 154026 -7066
rect 154262 -7302 189706 -7066
rect 189942 -7302 190026 -7066
rect 190262 -7302 225706 -7066
rect 225942 -7302 226026 -7066
rect 226262 -7302 261706 -7066
rect 261942 -7302 262026 -7066
rect 262262 -7302 297706 -7066
rect 297942 -7302 298026 -7066
rect 298262 -7302 333706 -7066
rect 333942 -7302 334026 -7066
rect 334262 -7302 369706 -7066
rect 369942 -7302 370026 -7066
rect 370262 -7302 405706 -7066
rect 405942 -7302 406026 -7066
rect 406262 -7302 441706 -7066
rect 441942 -7302 442026 -7066
rect 442262 -7302 477706 -7066
rect 477942 -7302 478026 -7066
rect 478262 -7302 513706 -7066
rect 513942 -7302 514026 -7066
rect 514262 -7302 549706 -7066
rect 549942 -7302 550026 -7066
rect 550262 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 9706 -7386
rect 9942 -7622 10026 -7386
rect 10262 -7622 45706 -7386
rect 45942 -7622 46026 -7386
rect 46262 -7622 81706 -7386
rect 81942 -7622 82026 -7386
rect 82262 -7622 117706 -7386
rect 117942 -7622 118026 -7386
rect 118262 -7622 153706 -7386
rect 153942 -7622 154026 -7386
rect 154262 -7622 189706 -7386
rect 189942 -7622 190026 -7386
rect 190262 -7622 225706 -7386
rect 225942 -7622 226026 -7386
rect 226262 -7622 261706 -7386
rect 261942 -7622 262026 -7386
rect 262262 -7622 297706 -7386
rect 297942 -7622 298026 -7386
rect 298262 -7622 333706 -7386
rect 333942 -7622 334026 -7386
rect 334262 -7622 369706 -7386
rect 369942 -7622 370026 -7386
rect 370262 -7622 405706 -7386
rect 405942 -7622 406026 -7386
rect 406262 -7622 441706 -7386
rect 441942 -7622 442026 -7386
rect 442262 -7622 477706 -7386
rect 477942 -7622 478026 -7386
rect 478262 -7622 513706 -7386
rect 513942 -7622 514026 -7386
rect 514262 -7622 549706 -7386
rect 549942 -7622 550026 -7386
rect 550262 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use mux16x1_project  mprj1
timestamp 0
transform 1 0 538000 0 1 423800
box 0 552 10000 22000
use mux16x1_project  mprj2
timestamp 0
transform 1 0 538000 0 1 387800
box 0 552 10000 22000
use mux16x1_project  mprj3
timestamp 0
transform 1 0 538000 0 1 351800
box 0 552 10000 22000
use mux16x1_project  mprj4
timestamp 0
transform 1 0 538000 0 1 315800
box 0 552 10000 22000
use mux16x1_project  mprj5
timestamp 0
transform 1 0 538000 0 1 279800
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro1
timestamp 0
transform 1 0 468600 0 1 449000
box 0 0 20145 2491
use sky130_osu_ring_oscillator_mpr2ct_8_b0r1  ro2
timestamp 0
transform 1 0 468600 0 1 430600
box 0 0 20785 2492
use sky130_osu_ring_oscillator_mpr2ea_8_b0r1  ro3
timestamp 0
transform 1 0 468600 0 1 409600
box 0 0 19886 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r1  ro4
timestamp 0
transform 1 0 468600 0 1 388600
box 0 0 22123 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r1  ro5
timestamp 0
transform 1 0 468600 0 1 356000
box 0 0 20809 2493
use sky130_osu_ring_oscillator_mpr2ca_8_b0r2  ro6
timestamp 0
transform 1 0 468600 0 1 340000
box 0 0 20217 2494
use sky130_osu_ring_oscillator_mpr2ct_8_b0r2  ro7
timestamp 0
transform 1 0 468600 0 1 320000
box 0 0 20783 2493
use sky130_osu_ring_oscillator_mpr2ea_8_b0r2  ro8
timestamp 0
transform 1 0 468600 0 1 304600
box 0 0 19885 2492
use sky130_osu_ring_oscillator_mpr2et_8_b0r2  ro9
timestamp 0
transform 1 0 468600 0 1 285000
box 0 0 22120 2493
use sky130_osu_ring_oscillator_mpr2xa_8_b0r2  ro10
timestamp 0
transform 1 0 468600 0 1 265000
box 0 0 20819 2493
use sky130_fd_sc_hd__conb_1  TIE_ZERO_zero_ pdk/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1689802698
transform 1 0 426328 0 1 373184
box -38 -48 314 592
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 994 -7654 1614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 36994 -7654 37614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 72994 -7654 73614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 108994 -7654 109614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 144994 -7654 145614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 180994 -7654 181614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 216994 -7654 217614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 252994 -7654 253614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 288994 -7654 289614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 324994 -7654 325614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 360994 -7654 361614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 396994 -7654 397614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 432994 -7654 433614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 468994 -7654 469614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 504994 -7654 505614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 540994 -7654 541614 279788 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 540994 445572 541614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 576994 -7654 577614 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2066 592650 2686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38066 592650 38686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74066 592650 74686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110066 592650 110686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146066 592650 146686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182066 592650 182686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218066 592650 218686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254066 592650 254686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290066 592650 290686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326066 592650 326686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362066 592650 362686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398066 592650 398686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434066 592650 434686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470066 592650 470686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506066 592650 506686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542066 592650 542686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578066 592650 578686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614066 592650 614686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650066 592650 650686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686066 592650 686686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 3474 -7654 4094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 39474 -7654 40094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 75474 -7654 76094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 111474 -7654 112094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 147474 -7654 148094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 183474 -7654 184094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 219474 -7654 220094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 255474 -7654 256094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 291474 -7654 292094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 327474 -7654 328094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 363474 -7654 364094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 399474 -7654 400094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 435474 -7654 436094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 471474 -7654 472094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 507474 -7654 508094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 543474 -7654 544094 279788 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 543474 445572 544094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 579474 -7654 580094 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 4546 592650 5166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 40546 592650 41166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 76546 592650 77166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 112546 592650 113166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 148546 592650 149166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 184546 592650 185166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 220546 592650 221166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 256546 592650 257166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 292546 592650 293166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 328546 592650 329166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 364546 592650 365166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 400546 592650 401166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 436546 592650 437166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 472546 592650 473166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 508546 592650 509166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 544546 592650 545166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 580546 592650 581166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 616546 592650 617166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 652546 592650 653166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 688546 592650 689166 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 5954 -7654 6574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 41954 -7654 42574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 77954 -7654 78574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 113954 -7654 114574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 149954 -7654 150574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 185954 -7654 186574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 221954 -7654 222574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 257954 -7654 258574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 293954 -7654 294574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 329954 -7654 330574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 365954 -7654 366574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 401954 -7654 402574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 437954 -7654 438574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 -7654 474574 263615 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 268060 474574 354615 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 473954 359060 474574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 509954 -7654 510574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 545954 -7654 546574 279788 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 545954 445572 546574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 581954 -7654 582574 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 7026 592650 7646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 43026 592650 43646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 79026 592650 79646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 115026 592650 115646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 151026 592650 151646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 187026 592650 187646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 223026 592650 223646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 259026 592650 259646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 295026 592650 295646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 331026 592650 331646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 367026 592650 367646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 403026 592650 403646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 439026 592650 439646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 475026 592650 475646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 511026 592650 511646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 547026 592650 547646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 583026 592650 583646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 619026 592650 619646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 655026 592650 655646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 691026 592650 691646 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 8434 -7654 9054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 44434 -7654 45054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 80434 -7654 81054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 116434 -7654 117054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 152434 -7654 153054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 188434 -7654 189054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 224434 -7654 225054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 260434 -7654 261054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 296434 -7654 297054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 332434 -7654 333054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 368434 -7654 369054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 404434 -7654 405054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 440434 -7654 441054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 -7654 477054 263615 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 268060 477054 354615 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 476434 359060 477054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 512434 -7654 513054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 548434 -7654 549054 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 9506 592650 10126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 45506 592650 46126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 81506 592650 82126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 117506 592650 118126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 153506 592650 154126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 189506 592650 190126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 225506 592650 226126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 261506 592650 262126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 297506 592650 298126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 333506 592650 334126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 369506 592650 370126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 405506 592650 406126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 441506 592650 442126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 477506 592650 478126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 513506 592650 514126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 549506 592650 550126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 585506 592650 586126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 621506 592650 622126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 657506 592650 658126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 693506 592650 694126 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 7194 -7654 7814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 43194 -7654 43814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 79194 -7654 79814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 115194 -7654 115814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 151194 -7654 151814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 187194 -7654 187814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 223194 -7654 223814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 259194 -7654 259814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 295194 -7654 295814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 331194 -7654 331814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 367194 -7654 367814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 403194 -7654 403814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 439194 -7654 439814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 -7654 475814 263615 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 268060 475814 354615 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 475194 359060 475814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 511194 -7654 511814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 547194 -7654 547814 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 8266 592650 8886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 44266 592650 44886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 80266 592650 80886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 116266 592650 116886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 152266 592650 152886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 188266 592650 188886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 224266 592650 224886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 260266 592650 260886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 296266 592650 296886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 332266 592650 332886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 368266 592650 368886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 404266 592650 404886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 440266 592650 440886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 476266 592650 476886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 512266 592650 512886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 548266 592650 548886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 584266 592650 584886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 620266 592650 620886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 656266 592650 656886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 692266 592650 692886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 9674 -7654 10294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 45674 -7654 46294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 81674 -7654 82294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 117674 -7654 118294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 153674 -7654 154294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 189674 -7654 190294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 225674 -7654 226294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 261674 -7654 262294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 297674 -7654 298294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 333674 -7654 334294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 369674 -7654 370294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 405674 -7654 406294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 441674 -7654 442294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 -7654 478294 263615 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 268060 478294 354615 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 477674 359060 478294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 513674 -7654 514294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 549674 -7654 550294 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 10746 592650 11366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 46746 592650 47366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 82746 592650 83366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 118746 592650 119366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 154746 592650 155366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 190746 592650 191366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 226746 592650 227366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 262746 592650 263366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 298746 592650 299366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 334746 592650 335366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 370746 592650 371366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 406746 592650 407366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 442746 592650 443366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 478746 592650 479366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 514746 592650 515366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 550746 592650 551366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 586746 592650 587366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 622746 592650 623366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 658746 592650 659366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 694746 592650 695366 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 2234 -7654 2854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 38234 -7654 38854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 74234 -7654 74854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 110234 -7654 110854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 146234 -7654 146854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 182234 -7654 182854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 218234 -7654 218854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 254234 -7654 254854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 290234 -7654 290854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 326234 -7654 326854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 362234 -7654 362854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 398234 -7654 398854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 434234 -7654 434854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 470234 -7654 470854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 506234 -7654 506854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 542234 -7654 542854 279788 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 542234 445572 542854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 578234 -7654 578854 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 3306 592650 3926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 39306 592650 39926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 75306 592650 75926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 111306 592650 111926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 147306 592650 147926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 183306 592650 183926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 219306 592650 219926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 255306 592650 255926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 291306 592650 291926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 327306 592650 327926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 363306 592650 363926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 399306 592650 399926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 435306 592650 435926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 471306 592650 471926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 507306 592650 507926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 543306 592650 543926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 579306 592650 579926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 615306 592650 615926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 651306 592650 651926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 687306 592650 687926 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 4714 -7654 5334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 40714 -7654 41334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 76714 -7654 77334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 112714 -7654 113334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 148714 -7654 149334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 184714 -7654 185334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 220714 -7654 221334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 256714 -7654 257334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 292714 -7654 293334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 328714 -7654 329334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 364714 -7654 365334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 400714 -7654 401334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 436714 -7654 437334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 -7654 473334 263615 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 268060 473334 354615 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 472714 359060 473334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 508714 -7654 509334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 544714 -7654 545334 279788 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 544714 445572 545334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 580714 -7654 581334 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 5786 592650 6406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 41786 592650 42406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 77786 592650 78406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 113786 592650 114406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 149786 592650 150406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 185786 592650 186406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 221786 592650 222406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 257786 592650 258406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 293786 592650 294406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 329786 592650 330406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 365786 592650 366406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 401786 592650 402406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 437786 592650 438406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 473786 592650 474406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 509786 592650 510406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 545786 592650 546406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 581786 592650 582406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 617786 592650 618406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 653786 592650 654406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 689786 592650 690406 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
